* NGSPICE file created from housekeeping.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufbuf_16 abstract view
.subckt sky130_fd_sc_hd__bufbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtn_1 abstract view
.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

.subckt housekeeping VGND VPWR debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oeb
+ pad_flash_csb pad_flash_csb_oeb pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ieb
+ pad_flash_io0_oeb pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ieb pad_flash_io1_oeb
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out[0] pwr_ctrl_out[1]
+ pwr_ctrl_out[2] pwr_ctrl_out[3] qspi_enabled reset ser_rx ser_tx serial_clock serial_data_1
+ serial_data_2 serial_load serial_resetn spi_csb spi_enabled spi_sck spi_sdi spi_sdo
+ spi_sdoenb spimemio_flash_clk spimemio_flash_csb spimemio_flash_io0_di spimemio_flash_io0_do
+ spimemio_flash_io0_oeb spimemio_flash_io1_di spimemio_flash_io1_do spimemio_flash_io1_oeb
+ spimemio_flash_io2_di spimemio_flash_io2_do spimemio_flash_io2_oeb spimemio_flash_io3_di
+ spimemio_flash_io3_do spimemio_flash_io3_oeb trap uart_enabled user_clock usr1_vcc_pwrgood
+ usr1_vdd_pwrgood usr2_vcc_pwrgood usr2_vdd_pwrgood wb_ack_o wb_adr_i[0] wb_adr_i[10]
+ wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17]
+ wb_adr_i[18] wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23]
+ wb_adr_i[24] wb_adr_i[25] wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2]
+ wb_adr_i[30] wb_adr_i[31] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7]
+ wb_adr_i[8] wb_adr_i[9] wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11]
+ wb_dat_i[12] wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18]
+ wb_dat_i[19] wb_dat_i[1] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24]
+ wb_dat_i[25] wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30]
+ wb_dat_i[31] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8]
+ wb_dat_i[9] wb_dat_o[0] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14]
+ wb_dat_o[15] wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20]
+ wb_dat_o[21] wb_dat_o[22] wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27]
+ wb_dat_o[28] wb_dat_o[29] wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4]
+ wb_dat_o[5] wb_dat_o[6] wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0]
+ wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] wb_stb_i wb_we_i
XFILLER_39_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6914_ _7154_/CLK _6914_/D fanout451/X VGND VGND VPWR VPWR _6914_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_70_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6845_ _6845_/CLK _6845_/D _6455_/A VGND VGND VPWR VPWR _6845_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3988_ hold470/X _6411_/A0 _3994_/S VGND VGND VPWR VPWR _3988_/X sky130_fd_sc_hd__mux2_1
X_6776_ _6851_/CLK _6776_/D fanout418/X VGND VGND VPWR VPWR _6776_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_109_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5727_ _7038_/Q _5683_/X _5704_/X _6934_/Q _5724_/X VGND VGND VPWR VPWR _5734_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5658_ _5665_/A _7173_/Q _5658_/S VGND VGND VPWR VPWR _7173_/D sky130_fd_sc_hd__mux2_1
XFILLER_190_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5589_ hold71/X _7144_/Q _5593_/S VGND VGND VPWR VPWR _5589_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4609_ _4987_/A _4992_/B _4586_/B VGND VGND VPWR VPWR _4619_/A sky130_fd_sc_hd__o21ai_1
XFILLER_2_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold340 _6872_/Q VGND VGND VPWR VPWR hold340/X sky130_fd_sc_hd__bufbuf_16
Xhold351 _6998_/Q VGND VGND VPWR VPWR hold351/X sky130_fd_sc_hd__bufbuf_16
Xhold362 _7134_/Q VGND VGND VPWR VPWR hold362/X sky130_fd_sc_hd__bufbuf_16
Xhold384 _6519_/Q VGND VGND VPWR VPWR hold384/X sky130_fd_sc_hd__bufbuf_16
Xhold373 _7030_/Q VGND VGND VPWR VPWR hold373/X sky130_fd_sc_hd__bufbuf_16
Xhold395 _6854_/Q VGND VGND VPWR VPWR hold395/X sky130_fd_sc_hd__bufbuf_16
XFILLER_132_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1040 _4102_/X VGND VGND VPWR VPWR _6580_/D sky130_fd_sc_hd__bufbuf_16
Xhold1051 _4134_/X VGND VGND VPWR VPWR _6607_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1084 _6819_/Q VGND VGND VPWR VPWR _5217_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1073 _6820_/Q VGND VGND VPWR VPWR _5219_/A0 sky130_fd_sc_hd__bufbuf_16
Xhold1062 _7021_/Q VGND VGND VPWR VPWR _5451_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_45_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_202 _7016_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_213 _6787_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1095 _6989_/Q VGND VGND VPWR VPWR _5415_/A1 sky130_fd_sc_hd__bufbuf_16
XANTENNA_224 _6480_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_268 wb_adr_i[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_257 _7174_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_235 mask_rev_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_246 mask_rev_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_279 wb_dat_i[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4960_ _4949_/A _4949_/C _4959_/X _4907_/A VGND VGND VPWR VPWR _4974_/A sky130_fd_sc_hd__a31o_4
XFILLER_91_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4891_ _4986_/A _4617_/A _5005_/C _4757_/B VGND VGND VPWR VPWR _5174_/C sky130_fd_sc_hd__o22ai_4
X_3911_ _7157_/Q _7159_/Q _7160_/Q _7158_/Q VGND VGND VPWR VPWR _3918_/B sky130_fd_sc_hd__or4b_2
X_6630_ _6746_/CLK _6630_/D fanout427/X VGND VGND VPWR VPWR _6630_/Q sky130_fd_sc_hd__dfrtp_2
X_3842_ _6487_/Q _6485_/Q _6664_/Q VGND VGND VPWR VPWR _3876_/S sky130_fd_sc_hd__and3_1
X_6561_ _7209_/CLK _6561_/D VGND VGND VPWR VPWR _6561_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_20_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5512_ _5584_/A0 hold486/X hold93/X VGND VGND VPWR VPWR _5512_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3773_ _7045_/Q _5477_/A _3344_/Y _6496_/Q _3772_/X VGND VGND VPWR VPWR _3773_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_145_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6492_ _6825_/CLK _6492_/D fanout421/X VGND VGND VPWR VPWR _6492_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_172_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5443_ _5578_/A0 hold361/X _5449_/S VGND VGND VPWR VPWR _7014_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5374_ _5599_/A0 hold849/X _5377_/S VGND VGND VPWR VPWR _5374_/X sky130_fd_sc_hd__mux2_1
X_7113_ _7150_/CLK _7113_/D fanout446/X VGND VGND VPWR VPWR _7113_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_114_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4325_ _6409_/A0 _4325_/A1 _4327_/S VGND VGND VPWR VPWR _6770_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4256_ _4256_/A hold47/X VGND VGND VPWR VPWR _4261_/S sky130_fd_sc_hd__and2_4
X_7044_ _7132_/CLK _7044_/D fanout428/X VGND VGND VPWR VPWR _7044_/Q sky130_fd_sc_hd__dfrtp_2
X_3207_ _7120_/Q VGND VGND VPWR VPWR _3207_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4187_ hold689/X _5561_/A0 _4189_/S VGND VGND VPWR VPWR _6651_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6828_ _7035_/CLK _6828_/D fanout432/X VGND VGND VPWR VPWR _6828_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6759_ _6759_/CLK _6759_/D fanout420/X VGND VGND VPWR VPWR _6759_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold170 _5228_/X VGND VGND VPWR VPWR _6826_/D sky130_fd_sc_hd__bufbuf_16
Xhold181 hold181/A VGND VGND VPWR VPWR hold181/X sky130_fd_sc_hd__bufbuf_16
XFILLER_120_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold192 _3257_/X VGND VGND VPWR VPWR hold192/X sky130_fd_sc_hd__bufbuf_16
XFILLER_144_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5090_ _5121_/C _5121_/D _5140_/C _5118_/D VGND VGND VPWR VPWR _5091_/C sky130_fd_sc_hd__or4_1
XFILLER_111_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4110_ _6587_/Q _3415_/X _4111_/S VGND VGND VPWR VPWR _6587_/D sky130_fd_sc_hd__mux2_1
X_4041_ hold209/A _4041_/A1 _4042_/S VGND VGND VPWR VPWR _4041_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5992_ _6014_/A _6036_/B VGND VGND VPWR VPWR _6020_/A sky130_fd_sc_hd__nor2_8
XFILLER_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4943_ _4745_/A _4697_/A _4756_/B VGND VGND VPWR VPWR _4943_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6613_ _6725_/CLK _6613_/D fanout440/X VGND VGND VPWR VPWR _6613_/Q sky130_fd_sc_hd__dfrtp_2
X_4874_ _5003_/A _4874_/B VGND VGND VPWR VPWR _5060_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3825_ _6482_/Q _3825_/B VGND VGND VPWR VPWR _3826_/B sky130_fd_sc_hd__nand2_1
X_3756_ _6589_/Q _4112_/A _3739_/X VGND VGND VPWR VPWR _3759_/B sky130_fd_sc_hd__a21o_1
X_6544_ _6777_/CLK _6544_/D fanout424/X VGND VGND VPWR VPWR _6544_/Q sky130_fd_sc_hd__dfrtp_2
Xclkbuf_3_5_0_csclk clkbuf_3_5_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_5_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_145_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6475_ _6668_/CLK _6475_/D _6430_/X VGND VGND VPWR VPWR _6475_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_106_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5426_ hold43/X _5426_/A1 hold48/X VGND VGND VPWR VPWR hold49/A sky130_fd_sc_hd__mux2_1
X_3687_ _3687_/A _3687_/B _3687_/C VGND VGND VPWR VPWR _3727_/A sky130_fd_sc_hd__or3_1
Xoutput231 _6516_/Q VGND VGND VPWR VPWR mgmt_gpio_out[26] sky130_fd_sc_hd__buf_8
Xoutput242 _3930_/X VGND VGND VPWR VPWR mgmt_gpio_out[36] sky130_fd_sc_hd__buf_8
Xoutput220 _6669_/Q VGND VGND VPWR VPWR mgmt_gpio_out[16] sky130_fd_sc_hd__buf_8
Xoutput253 _3955_/X VGND VGND VPWR VPWR pad_flash_csb sky130_fd_sc_hd__buf_8
XFILLER_160_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5357_ _5600_/A0 hold442/X _5359_/S VGND VGND VPWR VPWR _5357_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput275 _6496_/Q VGND VGND VPWR VPWR pll_trim[0] sky130_fd_sc_hd__buf_8
Xoutput264 _6819_/Q VGND VGND VPWR VPWR pll_bypass sky130_fd_sc_hd__buf_8
Xoutput286 _6497_/Q VGND VGND VPWR VPWR pll_trim[1] sky130_fd_sc_hd__buf_8
X_5288_ _5288_/A _5594_/B VGND VGND VPWR VPWR _5296_/S sky130_fd_sc_hd__nand2_8
XFILLER_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput297 _6502_/Q VGND VGND VPWR VPWR pll_trim[6] sky130_fd_sc_hd__buf_8
X_4308_ _4308_/A0 _6410_/A0 _4309_/S VGND VGND VPWR VPWR _4308_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4239_ _6703_/Q _6706_/Q _6705_/Q _6707_/Q VGND VGND VPWR VPWR _4239_/X sky130_fd_sc_hd__or4_4
XFILLER_75_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7027_ _7104_/CLK _7027_/D fanout435/X VGND VGND VPWR VPWR _7027_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_101_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4590_ _4590_/A _4590_/B VGND VGND VPWR VPWR _4591_/B sky130_fd_sc_hd__or2_4
X_3610_ _3970_/A _5245_/A _4124_/A _6601_/Q VGND VGND VPWR VPWR _3610_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3541_ _6712_/Q _4250_/A _4268_/A _6727_/Q VGND VGND VPWR VPWR _3541_/X sky130_fd_sc_hd__a22o_1
Xhold906 _4281_/X VGND VGND VPWR VPWR _6733_/D sky130_fd_sc_hd__bufbuf_16
Xhold917 _4210_/X VGND VGND VPWR VPWR _6672_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_127_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold928 _6774_/Q VGND VGND VPWR VPWR hold928/X sky130_fd_sc_hd__bufbuf_16
Xhold939 _5489_/X VGND VGND VPWR VPWR _7055_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_142_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3472_ _3472_/A _3472_/B _3472_/C _3472_/D VGND VGND VPWR VPWR _3548_/A sky130_fd_sc_hd__or4_1
X_6260_ _7197_/Q _6309_/S _6258_/X _6259_/X VGND VGND VPWR VPWR _7197_/D sky130_fd_sc_hd__o22a_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5211_ hold903/X _6410_/A0 _5215_/S VGND VGND VPWR VPWR _5211_/X sky130_fd_sc_hd__mux2_1
X_6191_ _7003_/Q _5987_/Y _6022_/D _6923_/Q _6190_/X VGND VGND VPWR VPWR _6194_/C
+ sky130_fd_sc_hd__a221o_1
X_5142_ _5142_/A _5142_/B _5124_/C VGND VGND VPWR VPWR _5143_/C sky130_fd_sc_hd__or3b_2
XFILLER_97_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5073_ _5079_/B _5073_/B _5073_/C _5073_/D VGND VGND VPWR VPWR _5145_/C sky130_fd_sc_hd__or4_2
XFILLER_96_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4024_ hold281/X _4023_/X _4024_/S VGND VGND VPWR VPWR _4024_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5975_ _6717_/Q _5676_/X _5702_/X _6554_/Q _5974_/X VGND VGND VPWR VPWR _5976_/D
+ sky130_fd_sc_hd__a221o_2
X_4926_ _4988_/A _4398_/Y _4660_/X _4746_/X VGND VGND VPWR VPWR _4926_/X sky130_fd_sc_hd__o22a_2
XFILLER_178_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4857_ _4622_/B _4845_/B _5071_/A _4849_/A VGND VGND VPWR VPWR _4857_/X sky130_fd_sc_hd__a211o_1
XFILLER_20_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3808_ _6485_/Q _3841_/B VGND VGND VPWR VPWR _3898_/A sky130_fd_sc_hd__nand2_4
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6527_ _7141_/CLK _6527_/D fanout447/X VGND VGND VPWR VPWR _6527_/Q sky130_fd_sc_hd__dfrtp_1
X_4788_ _4758_/B _4652_/B _4758_/C _5136_/A VGND VGND VPWR VPWR _4802_/C sky130_fd_sc_hd__a31o_1
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3739_ _6925_/Q _5342_/A _5405_/A _6981_/Q VGND VGND VPWR VPWR _3739_/X sky130_fd_sc_hd__a22o_2
XFILLER_4_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6458_ _6458_/CLK _6458_/D _3878_/X VGND VGND VPWR VPWR _6458_/Q sky130_fd_sc_hd__dfstp_4
X_6389_ _6705_/Q _6389_/A2 _6389_/B1 _4238_/B VGND VGND VPWR VPWR _6389_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5409_ hold617/X _5571_/A0 _5413_/S VGND VGND VPWR VPWR _5409_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5760_ _7007_/Q _5678_/X _5699_/X _6927_/Q _5759_/X VGND VGND VPWR VPWR _5763_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_98_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4711_ _4711_/A _4758_/A _4711_/C VGND VGND VPWR VPWR _4936_/A sky130_fd_sc_hd__and3_1
X_5691_ _5864_/B _5704_/B _5701_/C VGND VGND VPWR VPWR _5691_/X sky130_fd_sc_hd__and3_4
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4642_ _4642_/A _5069_/A _4922_/A _4641_/X VGND VGND VPWR VPWR _4642_/X sky130_fd_sc_hd__or4b_2
XFILLER_135_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4573_ _4947_/B _4875_/A VGND VGND VPWR VPWR _5128_/A sky130_fd_sc_hd__nor2_2
XFILLER_128_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold703 _5480_/X VGND VGND VPWR VPWR _7047_/D sky130_fd_sc_hd__bufbuf_16
Xhold736 _5329_/X VGND VGND VPWR VPWR _6913_/D sky130_fd_sc_hd__bufbuf_16
Xhold725 _6834_/Q VGND VGND VPWR VPWR hold725/X sky130_fd_sc_hd__bufbuf_16
XFILLER_116_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3524_ _4241_/A _3543_/B VGND VGND VPWR VPWR _4292_/A sky130_fd_sc_hd__nor2_8
Xhold714 _5520_/X VGND VGND VPWR VPWR _7083_/D sky130_fd_sc_hd__bufbuf_16
X_6312_ _6736_/Q _6020_/B _6011_/X _6788_/Q VGND VGND VPWR VPWR _6312_/X sky130_fd_sc_hd__a22o_1
Xhold758 hold882/X VGND VGND VPWR VPWR hold883/A sky130_fd_sc_hd__bufbuf_16
XFILLER_170_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold747 _5394_/X VGND VGND VPWR VPWR _6971_/D sky130_fd_sc_hd__bufbuf_16
X_6243_ _6604_/Q _6025_/A _6022_/A _6614_/Q VGND VGND VPWR VPWR _6243_/X sky130_fd_sc_hd__a22o_1
X_3455_ _3457_/A _3543_/B VGND VGND VPWR VPWR _4130_/A sky130_fd_sc_hd__nor2_8
Xhold769 _6500_/Q VGND VGND VPWR VPWR hold769/X sky130_fd_sc_hd__bufbuf_16
XFILLER_103_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6174_ _6954_/Q _6022_/A _6025_/C _6930_/Q VGND VGND VPWR VPWR _6174_/X sky130_fd_sc_hd__a22o_1
X_3386_ _3476_/A _3386_/B VGND VGND VPWR VPWR _3726_/A sky130_fd_sc_hd__nor2_8
XFILLER_97_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5125_ _4748_/A _4719_/X _4907_/C _4974_/A _5114_/B VGND VGND VPWR VPWR _5126_/B
+ sky130_fd_sc_hd__a2111o_1
X_5056_ _5056_/A _5056_/B _5157_/A _5056_/D VGND VGND VPWR VPWR _5057_/B sky130_fd_sc_hd__or4_1
XFILLER_111_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4007_ _6421_/B _4025_/A VGND VGND VPWR VPWR _4007_/X sky130_fd_sc_hd__and2b_4
XFILLER_65_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_1_wb_clk_i clkbuf_1_0_1_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_25_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5958_ _6612_/Q _5705_/X _5707_/X _6761_/Q _5957_/X VGND VGND VPWR VPWR _5959_/D
+ sky130_fd_sc_hd__a221o_1
X_4909_ _5145_/A _4909_/B _5075_/A _4909_/D VGND VGND VPWR VPWR _4910_/C sky130_fd_sc_hd__or4_1
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5889_ _6708_/Q _5691_/X _5701_/X _6614_/Q VGND VGND VPWR VPWR _5889_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_csclk clkbuf_2_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_5_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_20_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold41 hold41/A VGND VGND VPWR VPWR hold41/X sky130_fd_sc_hd__bufbuf_16
XFILLER_130_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold30 hold30/A VGND VGND VPWR VPWR hold30/X sky130_fd_sc_hd__bufbuf_16
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold74 hold5/X VGND VGND VPWR VPWR hold74/X sky130_fd_sc_hd__bufbuf_16
XFILLER_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold52 hold52/A VGND VGND VPWR VPWR hold52/X sky130_fd_sc_hd__bufbuf_16
Xhold63 hold63/A VGND VGND VPWR VPWR hold63/X sky130_fd_sc_hd__bufbuf_16
Xhold96 hold96/A VGND VGND VPWR VPWR hold96/X sky130_fd_sc_hd__bufbuf_16
Xhold85 hold85/A VGND VGND VPWR VPWR hold85/X sky130_fd_sc_hd__bufbuf_16
XFILLER_91_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_749 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_5 _6498_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6930_ _7130_/CLK _6930_/D fanout452/X VGND VGND VPWR VPWR _6930_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_81_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6861_ _7141_/CLK _6861_/D fanout448/X VGND VGND VPWR VPWR _6861_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_35_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5812_ _6898_/Q _5694_/X _5706_/X _7058_/Q VGND VGND VPWR VPWR _5812_/X sky130_fd_sc_hd__a22o_2
XFILLER_34_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6792_ _3545_/A1 _6792_/D _6450_/X VGND VGND VPWR VPWR _6792_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_179_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR clkbuf_2_1_0_mgmt_gpio_in[4]/A
+ sky130_fd_sc_hd__clkbuf_8
X_5743_ _5663_/A _7176_/Q _6358_/B1 VGND VGND VPWR VPWR _5743_/X sky130_fd_sc_hd__a21o_1
XFILLER_22_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5674_ _5864_/B _5705_/B _5703_/B VGND VGND VPWR VPWR _5674_/X sky130_fd_sc_hd__and3_4
XFILLER_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4625_ _4995_/A _4749_/C VGND VGND VPWR VPWR _5114_/B sky130_fd_sc_hd__nor2_4
Xhold511 _6911_/Q VGND VGND VPWR VPWR hold511/X sky130_fd_sc_hd__bufbuf_16
XFILLER_163_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4556_ _5118_/A _4840_/A _4805_/A _4556_/D VGND VGND VPWR VPWR _4557_/D sky130_fd_sc_hd__or4_1
Xhold500 _5377_/X VGND VGND VPWR VPWR _6956_/D sky130_fd_sc_hd__bufbuf_16
Xhold522 _4248_/X VGND VGND VPWR VPWR _6696_/D sky130_fd_sc_hd__bufbuf_16
Xhold533 _7151_/Q VGND VGND VPWR VPWR hold533/X sky130_fd_sc_hd__bufbuf_16
Xhold544 _5552_/X VGND VGND VPWR VPWR _7111_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_150_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3507_ _6643_/Q _4172_/A _4286_/A _6742_/Q VGND VGND VPWR VPWR _3507_/X sky130_fd_sc_hd__a22o_1
Xhold588 _5290_/X VGND VGND VPWR VPWR _6878_/D sky130_fd_sc_hd__bufbuf_16
X_4487_ _4655_/A _5050_/A VGND VGND VPWR VPWR _4746_/A sky130_fd_sc_hd__or2_4
Xhold555 _4244_/X VGND VGND VPWR VPWR _6692_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_104_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold577 _7042_/Q VGND VGND VPWR VPWR hold577/X sky130_fd_sc_hd__bufbuf_16
Xhold566 _6734_/Q VGND VGND VPWR VPWR hold566/X sky130_fd_sc_hd__bufbuf_16
Xhold599 _6883_/Q VGND VGND VPWR VPWR hold599/X sky130_fd_sc_hd__bufbuf_16
X_6226_ _6876_/Q _6023_/C _6025_/B _6900_/Q _6225_/X VGND VGND VPWR VPWR _6231_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_104_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3438_ _6994_/Q _3299_/Y hold21/A _7106_/Q _3437_/X VGND VGND VPWR VPWR _3452_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6157_ _6356_/A _6157_/B _6157_/C VGND VGND VPWR VPWR _6157_/X sky130_fd_sc_hd__or3_2
XFILLER_103_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1200 _6824_/Q VGND VGND VPWR VPWR _5224_/A1 sky130_fd_sc_hd__bufbuf_16
X_3369_ _3457_/A hold20/X VGND VGND VPWR VPWR _5396_/A sky130_fd_sc_hd__nor2_8
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _5108_/A _5108_/B _5108_/C VGND VGND VPWR VPWR _5155_/A sky130_fd_sc_hd__or3_2
Xhold1222 _6644_/Q VGND VGND VPWR VPWR _4179_/A0 sky130_fd_sc_hd__bufbuf_16
XFILLER_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1211 _6758_/Q VGND VGND VPWR VPWR _4311_/A0 sky130_fd_sc_hd__bufbuf_16
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1233 _4317_/X VGND VGND VPWR VPWR _6763_/D sky130_fd_sc_hd__bufbuf_16
Xhold1255 _6866_/Q VGND VGND VPWR VPWR _5276_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1266 _6691_/Q VGND VGND VPWR VPWR hold317/A sky130_fd_sc_hd__bufbuf_16
Xhold1244 _6615_/Q VGND VGND VPWR VPWR _4144_/A1 sky130_fd_sc_hd__bufbuf_16
X_6088_ _7135_/Q _6020_/B _6011_/X _7095_/Q VGND VGND VPWR VPWR _6088_/X sky130_fd_sc_hd__a22o_1
XFILLER_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5039_ _4832_/C _5050_/C _4689_/Y _4453_/Y VGND VGND VPWR VPWR _5039_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA_406 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_417 _3969_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_439 hold254/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_428 _5581_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput120 wb_adr_i[29] VGND VGND VPWR VPWR input120/X sky130_fd_sc_hd__clkbuf_4
XFILLER_122_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput153 wb_dat_i[29] VGND VGND VPWR VPWR _6393_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput131 wb_cyc_i VGND VGND VPWR VPWR input131/X sky130_fd_sc_hd__clkbuf_4
Xinput142 wb_dat_i[19] VGND VGND VPWR VPWR _6387_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_76_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput164 wb_rstn_i VGND VGND VPWR VPWR input164/X sky130_fd_sc_hd__buf_6
XFILLER_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4410_ _4707_/B _4478_/C _4410_/C _4410_/D VGND VGND VPWR VPWR _4997_/A sky130_fd_sc_hd__or4_4
X_5390_ _5597_/A0 hold550/X _5395_/S VGND VGND VPWR VPWR _5390_/X sky130_fd_sc_hd__mux2_1
X_4341_ _4654_/A _4696_/A _4413_/C _4654_/B VGND VGND VPWR VPWR _4341_/X sky130_fd_sc_hd__a31o_2
XFILLER_125_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7060_ _7152_/CLK _7060_/D fanout454/X VGND VGND VPWR VPWR _7060_/Q sky130_fd_sc_hd__dfrtp_2
X_4272_ hold870/X _4326_/A0 _4273_/S VGND VGND VPWR VPWR _4272_/X sky130_fd_sc_hd__mux2_1
X_3223_ _6992_/Q VGND VGND VPWR VPWR _3223_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6011_ _6012_/A _6035_/A _6037_/C VGND VGND VPWR VPWR _6011_/X sky130_fd_sc_hd__and3_4
XFILLER_101_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6913_ _7151_/CLK _6913_/D fanout446/X VGND VGND VPWR VPWR _6913_/Q sky130_fd_sc_hd__dfrtp_2
X_6844_ _7121_/CLK hold96/X _6421_/A VGND VGND VPWR VPWR hold95/A sky130_fd_sc_hd__dfrtp_2
XFILLER_50_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3987_ hold181/X hold200/X _6689_/Q VGND VGND VPWR VPWR _3987_/X sky130_fd_sc_hd__mux2_8
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6775_ _6840_/CLK _6775_/D fanout424/X VGND VGND VPWR VPWR _6775_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_167_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5726_ _7086_/Q _5685_/X _5699_/X _6926_/Q VGND VGND VPWR VPWR _5726_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5657_ _5612_/B _5620_/Y _5656_/X _6680_/Q VGND VGND VPWR VPWR _5658_/S sky130_fd_sc_hd__a22o_1
XFILLER_190_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5588_ _5588_/A0 _5588_/A1 _5593_/S VGND VGND VPWR VPWR _5588_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4608_ _4986_/B _4694_/A _4874_/B VGND VGND VPWR VPWR _4712_/B sky130_fd_sc_hd__o21ai_1
XFILLER_190_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4539_ _4818_/A _4672_/A _4740_/A _4539_/D VGND VGND VPWR VPWR _4542_/B sky130_fd_sc_hd__and4_1
XFILLER_104_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold330 _3511_/Y VGND VGND VPWR VPWR _4142_/A sky130_fd_sc_hd__bufbuf_16
Xhold341 _7126_/Q VGND VGND VPWR VPWR hold341/X sky130_fd_sc_hd__bufbuf_16
Xhold352 _5425_/X VGND VGND VPWR VPWR _6998_/D sky130_fd_sc_hd__bufbuf_16
Xhold363 _7060_/Q VGND VGND VPWR VPWR hold363/X sky130_fd_sc_hd__bufbuf_16
Xhold385 _4031_/X VGND VGND VPWR VPWR _6519_/D sky130_fd_sc_hd__bufbuf_16
Xhold374 _6930_/Q VGND VGND VPWR VPWR hold374/X sky130_fd_sc_hd__bufbuf_16
XFILLER_132_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold396 _5263_/X VGND VGND VPWR VPWR _6854_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_104_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6209_ _5663_/A _7194_/Q _5664_/X _6208_/X VGND VGND VPWR VPWR _6209_/X sky130_fd_sc_hd__a211o_1
X_7189_ _7197_/CLK _7189_/D fanout431/X VGND VGND VPWR VPWR _7189_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1030 _6598_/Q VGND VGND VPWR VPWR _4123_/A0 sky130_fd_sc_hd__bufbuf_16
Xhold1041 _6813_/Q VGND VGND VPWR VPWR _5210_/A0 sky130_fd_sc_hd__bufbuf_16
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1085 _6863_/Q VGND VGND VPWR VPWR _5273_/A1 sky130_fd_sc_hd__bufbuf_16
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1063 _6618_/Q VGND VGND VPWR VPWR _4147_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_85_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1052 _6608_/Q VGND VGND VPWR VPWR _4135_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1074 _5219_/X VGND VGND VPWR VPWR _6820_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_46_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_203 _7016_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_225 _6487_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1096 _6770_/Q VGND VGND VPWR VPWR _4325_/A1 sky130_fd_sc_hd__bufbuf_16
XANTENNA_214 _7096_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_258 spi_csb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_236 mask_rev_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_247 mask_rev_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_269 wb_adr_i[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_71_csclk clkbuf_opt_1_0_csclk/X VGND VGND VPWR VPWR _6825_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_36_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4890_ _4443_/X _4537_/X _4956_/C _5136_/B VGND VGND VPWR VPWR _5075_/A sky130_fd_sc_hd__a31o_1
X_3910_ _5663_/A _3905_/X _3921_/B _6832_/Q _6677_/Q VGND VGND VPWR VPWR _6679_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_17_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3841_ _6664_/Q _3841_/B VGND VGND VPWR VPWR _3847_/B sky130_fd_sc_hd__nand2_1
XFILLER_149_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6560_ _7208_/CLK _6560_/D VGND VGND VPWR VPWR _6560_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3772_ _6773_/Q _4328_/A _4172_/A _6639_/Q VGND VGND VPWR VPWR _3772_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5511_ hold209/X hold307/X hold93/X VGND VGND VPWR VPWR _5511_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6491_ _6759_/CLK _6491_/D fanout421/X VGND VGND VPWR VPWR _6491_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_8_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5442_ _5541_/A0 _5442_/A1 _5449_/S VGND VGND VPWR VPWR _7013_/D sky130_fd_sc_hd__mux2_1
X_5373_ _5571_/A0 hold796/X _5377_/S VGND VGND VPWR VPWR _5373_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7112_ _7130_/CLK _7112_/D fanout454/X VGND VGND VPWR VPWR _7112_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_172_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_24_csclk _7137_/CLK VGND VGND VPWR VPWR _6975_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_114_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4324_ _6408_/A0 hold501/X _4327_/S VGND VGND VPWR VPWR _4324_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7043_ _7131_/CLK _7043_/D fanout432/X VGND VGND VPWR VPWR _7043_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_101_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4255_ _5545_/A0 _4255_/A1 _4255_/S VGND VGND VPWR VPWR _4255_/X sky130_fd_sc_hd__mux2_1
X_3206_ _7128_/Q VGND VGND VPWR VPWR _3206_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_39_csclk _7137_/CLK VGND VGND VPWR VPWR _6971_/CLK sky130_fd_sc_hd__clkbuf_8
X_4186_ hold342/X _5587_/A0 _4189_/S VGND VGND VPWR VPWR _4186_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_1_0_csclk clkbuf_3_1_0_csclk/A VGND VGND VPWR VPWR _6722_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_55_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6827_ _7035_/CLK _6827_/D fanout433/X VGND VGND VPWR VPWR _6827_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6758_ _7222_/CLK _6758_/D fanout420/X VGND VGND VPWR VPWR _6758_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_109_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5709_ _7045_/Q _5687_/X _5701_/X _6949_/Q _5708_/X VGND VGND VPWR VPWR _5709_/X
+ sky130_fd_sc_hd__a221o_2
X_6689_ _7220_/CLK _6689_/D _6362_/B VGND VGND VPWR VPWR _6689_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_128_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold171 _6864_/Q VGND VGND VPWR VPWR hold171/X sky130_fd_sc_hd__bufbuf_16
Xhold160 _3981_/X VGND VGND VPWR VPWR hold66/A sky130_fd_sc_hd__bufbuf_16
XFILLER_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold182 hold201/X VGND VGND VPWR VPWR hold202/A sky130_fd_sc_hd__bufbuf_16
XFILLER_104_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold193 _3258_/X VGND VGND VPWR VPWR hold193/X sky130_fd_sc_hd__bufbuf_16
XFILLER_132_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4040_ _5600_/A0 hold411/X _4042_/S VGND VGND VPWR VPWR _4040_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5991_ _6037_/A _6035_/C VGND VGND VPWR VPWR _6036_/B sky130_fd_sc_hd__nand2_8
XFILLER_64_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4942_ _4395_/D _4469_/Y _4689_/Y _4798_/C _4847_/A VGND VGND VPWR VPWR _5180_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6612_ _6725_/CLK _6612_/D fanout440/X VGND VGND VPWR VPWR _6612_/Q sky130_fd_sc_hd__dfrtp_2
X_4873_ _4947_/B _4898_/B _4591_/B VGND VGND VPWR VPWR _5128_/B sky130_fd_sc_hd__a21oi_1
XFILLER_177_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3824_ _3840_/S _3824_/B _6481_/Q VGND VGND VPWR VPWR _3826_/A sky130_fd_sc_hd__or3b_2
XFILLER_165_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3755_ _6594_/Q _4118_/A _4262_/A _6718_/Q _3734_/X VGND VGND VPWR VPWR _3759_/A
+ sky130_fd_sc_hd__a221o_1
X_6543_ _6777_/CLK _6543_/D fanout418/X VGND VGND VPWR VPWR _6543_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_145_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3686_ _6564_/Q _4082_/A _3511_/Y _6615_/Q _3685_/X VGND VGND VPWR VPWR _3687_/C
+ sky130_fd_sc_hd__a221o_4
X_6474_ _6668_/CLK _6474_/D _6429_/X VGND VGND VPWR VPWR _6474_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_146_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput210 _3233_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[7] sky130_fd_sc_hd__buf_8
X_5425_ _5578_/A0 hold351/X hold48/X VGND VGND VPWR VPWR _5425_/X sky130_fd_sc_hd__mux2_1
Xoutput232 _6517_/Q VGND VGND VPWR VPWR mgmt_gpio_out[27] sky130_fd_sc_hd__buf_8
Xoutput243 _3929_/X VGND VGND VPWR VPWR mgmt_gpio_out[37] sky130_fd_sc_hd__buf_8
Xoutput221 _6670_/Q VGND VGND VPWR VPWR mgmt_gpio_out[17] sky130_fd_sc_hd__buf_8
XFILLER_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5356_ _5599_/A0 hold845/X _5359_/S VGND VGND VPWR VPWR _5356_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput276 _6490_/Q VGND VGND VPWR VPWR pll_trim[10] sky130_fd_sc_hd__buf_8
Xoutput265 _6799_/Q VGND VGND VPWR VPWR pll_dco_ena sky130_fd_sc_hd__buf_8
Xoutput254 _3956_/Y VGND VGND VPWR VPWR pad_flash_csb_oeb sky130_fd_sc_hd__buf_8
X_5287_ _5602_/A0 hold519/X _5287_/S VGND VGND VPWR VPWR _5287_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput287 _6815_/Q VGND VGND VPWR VPWR pll_trim[20] sky130_fd_sc_hd__buf_8
Xoutput298 _6503_/Q VGND VGND VPWR VPWR pll_trim[7] sky130_fd_sc_hd__buf_8
X_4307_ _4307_/A0 _6409_/A0 _4309_/S VGND VGND VPWR VPWR _4307_/X sky130_fd_sc_hd__mux2_1
X_4238_ _6703_/Q _4238_/B VGND VGND VPWR VPWR _6376_/A sky130_fd_sc_hd__and2b_4
XFILLER_102_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7026_ _7090_/CLK _7026_/D fanout438/X VGND VGND VPWR VPWR _7026_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_68_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4169_ _6409_/A0 _4169_/A1 _4171_/S VGND VGND VPWR VPWR _6636_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3540_ _3540_/A _3733_/B VGND VGND VPWR VPWR _4268_/A sky130_fd_sc_hd__nor2_8
XFILLER_128_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold918 _6973_/Q VGND VGND VPWR VPWR hold918/X sky130_fd_sc_hd__bufbuf_16
Xhold907 _6749_/Q VGND VGND VPWR VPWR hold907/X sky130_fd_sc_hd__bufbuf_16
XFILLER_170_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5210_ _5210_/A0 _6409_/A0 _5215_/S VGND VGND VPWR VPWR _6813_/D sky130_fd_sc_hd__mux2_1
Xhold929 _4330_/X VGND VGND VPWR VPWR _6774_/D sky130_fd_sc_hd__bufbuf_16
X_3471_ _7105_/Q hold21/A _4310_/A _6762_/Q _3469_/X VGND VGND VPWR VPWR _3472_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6190_ _7123_/Q _6023_/D _6030_/Y _7035_/Q VGND VGND VPWR VPWR _6190_/X sky130_fd_sc_hd__a22o_1
X_5141_ _5172_/B _5171_/C _5172_/A VGND VGND VPWR VPWR _5169_/A sky130_fd_sc_hd__o21ba_1
X_5072_ _4748_/A _4689_/Y _4905_/C _4973_/C _4850_/B VGND VGND VPWR VPWR _5175_/A
+ sky130_fd_sc_hd__a2111o_1
X_4023_ hold355/X hold14/X _4023_/S VGND VGND VPWR VPWR _4023_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5974_ _6663_/Q _5669_/X _5698_/B _5963_/X VGND VGND VPWR VPWR _5974_/X sky130_fd_sc_hd__a22o_1
X_4925_ _4930_/D _4586_/B _4933_/B _4748_/B VGND VGND VPWR VPWR _5022_/D sky130_fd_sc_hd__a22o_1
XFILLER_100_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4856_ _4586_/B _4845_/B _4850_/X _4855_/X _5116_/B VGND VGND VPWR VPWR _4856_/X
+ sky130_fd_sc_hd__a2111o_1
X_3807_ _6487_/Q _6486_/Q _6485_/Q VGND VGND VPWR VPWR _3843_/B sky130_fd_sc_hd__and3_4
XFILLER_193_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4787_ _4808_/A _4787_/B VGND VGND VPWR VPWR _5132_/A sky130_fd_sc_hd__or2_4
X_6526_ _6987_/CLK _6526_/D fanout450/X VGND VGND VPWR VPWR _6526_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3738_ _6563_/Q _4082_/A _4124_/A _6599_/Q VGND VGND VPWR VPWR _3738_/X sky130_fd_sc_hd__a22o_2
XFILLER_118_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3669_ _6729_/Q _4274_/A _4004_/A _6505_/Q VGND VGND VPWR VPWR _3669_/X sky130_fd_sc_hd__a22o_2
X_6457_ _3957_/A1 _6457_/D _6413_/X VGND VGND VPWR VPWR _6457_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6388_ _6387_/X _7214_/Q _6400_/S VGND VGND VPWR VPWR _7214_/D sky130_fd_sc_hd__mux2_1
X_5408_ hold515/X _5597_/A0 _5413_/S VGND VGND VPWR VPWR _5408_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5339_ hold404/X _5600_/A0 _5341_/S VGND VGND VPWR VPWR _5339_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7009_ _7118_/CLK _7009_/D fanout436/X VGND VGND VPWR VPWR _7009_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4710_ _5023_/A _4671_/A _5031_/B VGND VGND VPWR VPWR _4713_/C sky130_fd_sc_hd__a21oi_1
X_5690_ _7165_/Q _5704_/B _5701_/C VGND VGND VPWR VPWR _5690_/X sky130_fd_sc_hd__and3_4
XFILLER_91_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4641_ _4965_/A _5005_/C _4639_/X _4640_/X VGND VGND VPWR VPWR _4641_/X sky130_fd_sc_hd__o211a_1
XFILLER_175_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4572_ _4572_/A _4572_/B _5147_/A VGND VGND VPWR VPWR _4875_/A sky130_fd_sc_hd__or3_4
XFILLER_162_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold737 _6907_/Q VGND VGND VPWR VPWR hold737/X sky130_fd_sc_hd__bufbuf_16
Xhold726 _5239_/X VGND VGND VPWR VPWR _6834_/D sky130_fd_sc_hd__bufbuf_16
Xhold715 _6525_/Q VGND VGND VPWR VPWR hold715/X sky130_fd_sc_hd__bufbuf_16
XFILLER_116_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3523_ _6857_/Q _3315_/Y _3334_/Y _7041_/Q VGND VGND VPWR VPWR _3523_/X sky130_fd_sc_hd__a22o_1
Xhold704 _6828_/Q VGND VGND VPWR VPWR hold704/X sky130_fd_sc_hd__bufbuf_16
X_6311_ _6657_/Q _6311_/B VGND VGND VPWR VPWR _6311_/X sky130_fd_sc_hd__and2_1
Xhold759 hold884/X VGND VGND VPWR VPWR hold885/A sky130_fd_sc_hd__bufbuf_16
X_6242_ _6576_/Q _6021_/A _6011_/X _6785_/Q _6241_/X VGND VGND VPWR VPWR _6247_/B
+ sky130_fd_sc_hd__a221o_1
Xhold748 _6752_/Q VGND VGND VPWR VPWR hold748/X sky130_fd_sc_hd__bufbuf_16
X_3454_ _3453_/X _6795_/Q _3928_/A VGND VGND VPWR VPWR _6795_/D sky130_fd_sc_hd__mux2_1
XFILLER_103_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6173_ _7130_/Q _6023_/A _6033_/X _7010_/Q _6172_/X VGND VGND VPWR VPWR _6182_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3385_ _7201_/Q _6830_/Q _6831_/Q VGND VGND VPWR VPWR _3385_/X sky130_fd_sc_hd__mux2_8
X_5124_ _5142_/A _5124_/B _5124_/C _5124_/D VGND VGND VPWR VPWR _5131_/A sky130_fd_sc_hd__nand4b_4
XFILLER_97_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5055_ _5156_/B _5105_/C VGND VGND VPWR VPWR _5056_/D sky130_fd_sc_hd__or2_1
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4006_ _5578_/A0 _6505_/Q _4006_/S VGND VGND VPWR VPWR _4006_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5957_ _6741_/Q _5678_/X _5692_/X _7224_/Q VGND VGND VPWR VPWR _5957_/X sky130_fd_sc_hd__a22o_1
X_4908_ _4956_/C _4719_/X _5073_/C _4907_/X _4628_/Y VGND VGND VPWR VPWR _4909_/D
+ sky130_fd_sc_hd__a2111o_2
XFILLER_178_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5888_ _6599_/Q _5699_/X _5706_/X _6649_/Q _5887_/X VGND VGND VPWR VPWR _5893_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_138_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4839_ _5087_/B _5087_/C _4719_/C VGND VGND VPWR VPWR _4839_/X sky130_fd_sc_hd__o21a_4
XFILLER_193_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6509_ _6672_/CLK _6509_/D fanout453/X VGND VGND VPWR VPWR _6509_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_146_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold31 hold38/X VGND VGND VPWR VPWR hold39/A sky130_fd_sc_hd__bufbuf_16
Xhold20 hold20/A VGND VGND VPWR VPWR hold20/X sky130_fd_sc_hd__bufbuf_16
XFILLER_29_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold64 hold64/A VGND VGND VPWR VPWR hold64/X sky130_fd_sc_hd__bufbuf_16
Xhold42 hold42/A VGND VGND VPWR VPWR hold42/X sky130_fd_sc_hd__bufbuf_16
Xhold53 hold53/A VGND VGND VPWR VPWR hold53/X sky130_fd_sc_hd__bufbuf_16
Xhold75 hold75/A VGND VGND VPWR VPWR hold6/A sky130_fd_sc_hd__bufbuf_16
Xhold86 hold86/A VGND VGND VPWR VPWR hold86/X sky130_fd_sc_hd__bufbuf_16
XFILLER_152_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold97 hold97/A VGND VGND VPWR VPWR hold97/X sky130_fd_sc_hd__bufbuf_16
XFILLER_56_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_6 _6499_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6860_ _7088_/CLK _6860_/D fanout438/X VGND VGND VPWR VPWR _6860_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_179_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5811_ _7090_/Q _5685_/X _5699_/X _6930_/Q VGND VGND VPWR VPWR _5811_/X sky130_fd_sc_hd__a22o_1
X_6791_ _3957_/A1 _6791_/D _6449_/X VGND VGND VPWR VPWR _6791_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_15_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5742_ _6854_/Q _5722_/B _5734_/X _5741_/X _3197_/Y VGND VGND VPWR VPWR _5742_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_50_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5673_ _5864_/B _5707_/B _5701_/C VGND VGND VPWR VPWR _5673_/X sky130_fd_sc_hd__and3_4
XFILLER_163_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4624_ _4987_/A _4624_/B VGND VGND VPWR VPWR _4624_/Y sky130_fd_sc_hd__nand2_1
XFILLER_135_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4555_ _4987_/B _4845_/A _4552_/X _4554_/X VGND VGND VPWR VPWR _4556_/D sky130_fd_sc_hd__a211o_1
XFILLER_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold501 _6769_/Q VGND VGND VPWR VPWR hold501/X sky130_fd_sc_hd__bufbuf_16
Xhold534 _5597_/X VGND VGND VPWR VPWR _7151_/D sky130_fd_sc_hd__bufbuf_16
Xhold512 _5327_/X VGND VGND VPWR VPWR _6911_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_144_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold545 _6931_/Q VGND VGND VPWR VPWR hold545/X sky130_fd_sc_hd__bufbuf_16
X_3506_ _3506_/A _5234_/B VGND VGND VPWR VPWR _4286_/A sky130_fd_sc_hd__nor2_8
Xhold523 _6687_/Q VGND VGND VPWR VPWR hold523/X sky130_fd_sc_hd__bufbuf_16
Xhold556 _6870_/Q VGND VGND VPWR VPWR hold556/X sky130_fd_sc_hd__bufbuf_16
X_4486_ _4735_/B _4486_/B _4507_/A VGND VGND VPWR VPWR _5118_/A sky130_fd_sc_hd__and3_2
Xhold578 _5474_/X VGND VGND VPWR VPWR _7042_/D sky130_fd_sc_hd__bufbuf_16
Xhold567 _4282_/X VGND VGND VPWR VPWR _6734_/D sky130_fd_sc_hd__bufbuf_16
Xhold589 _6923_/Q VGND VGND VPWR VPWR hold589/X sky130_fd_sc_hd__bufbuf_16
X_6225_ _6964_/Q _6022_/C _6032_/X _7060_/Q VGND VGND VPWR VPWR _6225_/X sky130_fd_sc_hd__a22o_1
XFILLER_106_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3437_ _7074_/Q hold92/A _5227_/A _3423_/X VGND VGND VPWR VPWR _3437_/X sky130_fd_sc_hd__a22o_1
X_6156_ _6156_/A _6156_/B _6156_/C _6156_/D VGND VGND VPWR VPWR _6157_/C sky130_fd_sc_hd__or4_2
X_3368_ _5225_/A _3473_/B VGND VGND VPWR VPWR _3368_/Y sky130_fd_sc_hd__nor2_8
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _4756_/B _5050_/C _4823_/X VGND VGND VPWR VPWR _5108_/C sky130_fd_sc_hd__o21ai_2
Xhold1234 _6528_/Q VGND VGND VPWR VPWR _4041_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_112_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1223 _4179_/X VGND VGND VPWR VPWR _6644_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1201 _5224_/X VGND VGND VPWR VPWR _6824_/D sky130_fd_sc_hd__bufbuf_16
Xhold1212 _4311_/X VGND VGND VPWR VPWR _6758_/D sky130_fd_sc_hd__bufbuf_16
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6087_ _7063_/Q _5996_/X _6020_/C _6911_/Q VGND VGND VPWR VPWR _6087_/X sky130_fd_sc_hd__a22o_1
XFILLER_111_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1256 _6826_/Q VGND VGND VPWR VPWR _5228_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1245 _6827_/Q VGND VGND VPWR VPWR _5229_/A1 sky130_fd_sc_hd__bufbuf_16
X_3299_ _3514_/A _3668_/A VGND VGND VPWR VPWR _3299_/Y sky130_fd_sc_hd__nor2_8
Xhold1267 _7118_/Q VGND VGND VPWR VPWR _5560_/A1 sky130_fd_sc_hd__bufbuf_16
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_407 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5038_ _6376_/A _5158_/A VGND VGND VPWR VPWR _5038_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_418 _3202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_429 _5561_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_750 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6989_ _7101_/CLK _6989_/D fanout430/X VGND VGND VPWR VPWR _6989_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_178_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput110 wb_adr_i[1] VGND VGND VPWR VPWR _4818_/A sky130_fd_sc_hd__buf_8
XFILLER_163_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput121 wb_adr_i[2] VGND VGND VPWR VPWR _4395_/D sky130_fd_sc_hd__buf_8
Xinput132 wb_dat_i[0] VGND VGND VPWR VPWR _6378_/B1 sky130_fd_sc_hd__clkbuf_4
Xinput154 wb_dat_i[2] VGND VGND VPWR VPWR _6383_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_163_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput143 wb_dat_i[1] VGND VGND VPWR VPWR _6381_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput165 wb_sel_i[0] VGND VGND VPWR VPWR _6374_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4340_ _4654_/A _4340_/B VGND VGND VPWR VPWR _4408_/A sky130_fd_sc_hd__xor2_4
XFILLER_125_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4271_ hold942/X _5300_/A0 _4273_/S VGND VGND VPWR VPWR _6725_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3222_ _7000_/Q VGND VGND VPWR VPWR _3222_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_140_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6010_ _6036_/A _6010_/B VGND VGND VPWR VPWR _6010_/Y sky130_fd_sc_hd__nor2_8
XFILLER_67_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6912_ _6987_/CLK _6912_/D fanout450/X VGND VGND VPWR VPWR _6912_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_82_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6843_ _6843_/CLK _6843_/D _6421_/A VGND VGND VPWR VPWR _6843_/Q sky130_fd_sc_hd__dfrtp_2
X_3986_ _3986_/A0 _6410_/A0 _3994_/S VGND VGND VPWR VPWR _6491_/D sky130_fd_sc_hd__mux2_1
X_6774_ _6851_/CLK _6774_/D fanout418/X VGND VGND VPWR VPWR _6774_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_148_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5725_ _6894_/Q _5694_/X _5706_/X _7054_/Q VGND VGND VPWR VPWR _5725_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5656_ _7159_/Q _7160_/Q _5610_/Y VGND VGND VPWR VPWR _5656_/X sky130_fd_sc_hd__or3b_1
X_4607_ _4917_/A VGND VGND VPWR VPWR _4980_/C sky130_fd_sc_hd__inv_2
XFILLER_191_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold320 _4033_/X VGND VGND VPWR VPWR _6521_/D sky130_fd_sc_hd__bufbuf_16
X_5587_ _5587_/A0 hold461/X _5593_/S VGND VGND VPWR VPWR _7142_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4538_ _4538_/A _4949_/B VGND VGND VPWR VPWR _4970_/B sky130_fd_sc_hd__nand2_1
Xhold342 _6650_/Q VGND VGND VPWR VPWR hold342/X sky130_fd_sc_hd__bufbuf_16
XFILLER_104_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold331 _4144_/X VGND VGND VPWR VPWR _6615_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold353 _6821_/Q VGND VGND VPWR VPWR hold353/X sky130_fd_sc_hd__bufbuf_16
Xhold364 _5494_/X VGND VGND VPWR VPWR _7060_/D sky130_fd_sc_hd__bufbuf_16
X_4469_ _4469_/A _4663_/B VGND VGND VPWR VPWR _4469_/Y sky130_fd_sc_hd__nor2_8
Xhold386 _6900_/Q VGND VGND VPWR VPWR hold386/X sky130_fd_sc_hd__bufbuf_16
Xhold375 _5348_/X VGND VGND VPWR VPWR _6930_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_117_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6208_ _6859_/Q _6060_/B _6207_/X _6308_/S VGND VGND VPWR VPWR _6208_/X sky130_fd_sc_hd__o211a_1
Xhold397 _6990_/Q VGND VGND VPWR VPWR hold397/X sky130_fd_sc_hd__bufbuf_16
XFILLER_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7188_ _7201_/CLK _7188_/D fanout419/X VGND VGND VPWR VPWR _7188_/Q sky130_fd_sc_hd__dfrtp_2
Xhold1042 _6933_/Q VGND VGND VPWR VPWR _5352_/A1 sky130_fd_sc_hd__bufbuf_16
X_6139_ _7017_/Q _6036_/Y _6335_/B _7041_/Q _6136_/X VGND VGND VPWR VPWR _6144_/B
+ sky130_fd_sc_hd__a221o_1
Xhold1031 _4123_/X VGND VGND VPWR VPWR _6598_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_58_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1020 _4176_/X VGND VGND VPWR VPWR _6642_/D sky130_fd_sc_hd__bufbuf_16
Xhold1075 _6901_/Q VGND VGND VPWR VPWR _5316_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1064 _4147_/X VGND VGND VPWR VPWR _6618_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1053 _4135_/X VGND VGND VPWR VPWR _6608_/D sky130_fd_sc_hd__bufbuf_16
Xhold1086 _5273_/X VGND VGND VPWR VPWR _6863_/D sky130_fd_sc_hd__bufbuf_16
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_215 _6766_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1097 _6633_/Q VGND VGND VPWR VPWR _4165_/A1 sky130_fd_sc_hd__bufbuf_16
XANTENNA_204 _7024_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_259 spi_sck VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_226 _6473_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_237 mask_rev_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_248 mask_rev_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_5_csclk _6722_/CLK VGND VGND VPWR VPWR _6713_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_174_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3840_ _3839_/X hold80/A _3840_/S VGND VGND VPWR VPWR _6477_/D sky130_fd_sc_hd__mux2_1
XFILLER_60_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3771_ _6763_/Q _4316_/A _4196_/A _6659_/Q VGND VGND VPWR VPWR _3771_/X sky130_fd_sc_hd__a22o_1
XFILLER_157_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5510_ _5582_/A0 hold765/X hold93/X VGND VGND VPWR VPWR _5510_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6490_ _6759_/CLK _6490_/D fanout421/X VGND VGND VPWR VPWR _6490_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_8_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5441_ _5441_/A _5576_/B VGND VGND VPWR VPWR _5441_/Y sky130_fd_sc_hd__nand2_8
X_5372_ _5588_/A0 _5372_/A1 _5377_/S VGND VGND VPWR VPWR _5372_/X sky130_fd_sc_hd__mux2_1
X_7111_ _7111_/CLK _7111_/D fanout444/X VGND VGND VPWR VPWR _7111_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_160_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4323_ _6407_/A0 _4323_/A1 _4327_/S VGND VGND VPWR VPWR _4323_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7042_ _7131_/CLK _7042_/D fanout432/X VGND VGND VPWR VPWR _7042_/Q sky130_fd_sc_hd__dfrtp_2
X_4254_ _4326_/A0 hold772/X _4255_/S VGND VGND VPWR VPWR _4254_/X sky130_fd_sc_hd__mux2_1
X_4185_ _4185_/A0 _5289_/A0 _4189_/S VGND VGND VPWR VPWR _4185_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3205_ _7136_/Q VGND VGND VPWR VPWR _3205_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6826_ _7035_/CLK _6826_/D fanout433/X VGND VGND VPWR VPWR _6826_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_51_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6757_ _7222_/CLK _6757_/D fanout423/X VGND VGND VPWR VPWR _6757_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_109_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5708_ _7029_/Q _5688_/X _5707_/X _7021_/Q _5670_/X VGND VGND VPWR VPWR _5708_/X
+ sky130_fd_sc_hd__a221o_1
X_3969_ _3969_/A _3969_/B VGND VGND VPWR VPWR _3969_/X sky130_fd_sc_hd__and2_2
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6688_ _7107_/CLK _6688_/D fanout434/X VGND VGND VPWR VPWR _6688_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5639_ _7167_/Q _7166_/Q _6679_/Q VGND VGND VPWR VPWR _5648_/B sky130_fd_sc_hd__and3_2
XFILLER_163_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold161 hold66/X VGND VGND VPWR VPWR hold36/A sky130_fd_sc_hd__bufbuf_16
XFILLER_105_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold150 _5445_/X VGND VGND VPWR VPWR _7016_/D sky130_fd_sc_hd__bufbuf_16
Xhold172 _5274_/X VGND VGND VPWR VPWR _6864_/D sky130_fd_sc_hd__bufbuf_16
Xhold183 hold183/A VGND VGND VPWR VPWR hold183/X sky130_fd_sc_hd__bufbuf_16
Xhold194 _3259_/Y VGND VGND VPWR VPWR hold52/A sky130_fd_sc_hd__bufbuf_16
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5990_ _7167_/Q _7166_/Q VGND VGND VPWR VPWR _6035_/C sky130_fd_sc_hd__nor2_8
X_4941_ _5163_/A _4941_/B _4941_/C _4941_/D VGND VGND VPWR VPWR _4946_/A sky130_fd_sc_hd__or4_1
X_4872_ _4953_/A _4899_/B VGND VGND VPWR VPWR _5099_/C sky130_fd_sc_hd__nor2_2
XFILLER_60_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6611_ _6725_/CLK _6611_/D fanout440/X VGND VGND VPWR VPWR _6611_/Q sky130_fd_sc_hd__dfstp_4
X_3823_ _3845_/A _3828_/S VGND VGND VPWR VPWR _3824_/B sky130_fd_sc_hd__nor2_1
XFILLER_20_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6542_ _6616_/CLK _6542_/D fanout440/X VGND VGND VPWR VPWR _6542_/Q sky130_fd_sc_hd__dfstp_4
X_3754_ _3754_/A _3754_/B _3754_/C _3754_/D VGND VGND VPWR VPWR _3794_/A sky130_fd_sc_hd__or4_2
XFILLER_145_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3685_ _6918_/Q _5333_/A _4112_/A _6590_/Q VGND VGND VPWR VPWR _3685_/X sky130_fd_sc_hd__a22o_1
X_6473_ _6668_/CLK _6473_/D _6428_/X VGND VGND VPWR VPWR _6473_/Q sky130_fd_sc_hd__dfrtp_2
Xoutput200 _3208_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[32] sky130_fd_sc_hd__buf_8
XFILLER_161_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5424_ _5541_/A0 _5424_/A1 hold48/X VGND VGND VPWR VPWR _6997_/D sky130_fd_sc_hd__mux2_1
Xoutput233 _6518_/Q VGND VGND VPWR VPWR mgmt_gpio_out[28] sky130_fd_sc_hd__buf_8
Xoutput222 _6671_/Q VGND VGND VPWR VPWR mgmt_gpio_out[18] sky130_fd_sc_hd__buf_8
Xoutput211 _3232_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[8] sky130_fd_sc_hd__buf_8
Xoutput244 _6684_/Q VGND VGND VPWR VPWR mgmt_gpio_out[3] sky130_fd_sc_hd__buf_8
XFILLER_161_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5355_ _5571_/A0 hold793/X _5359_/S VGND VGND VPWR VPWR _6936_/D sky130_fd_sc_hd__mux2_1
Xoutput266 _6800_/Q VGND VGND VPWR VPWR pll_div[0] sky130_fd_sc_hd__buf_8
Xoutput255 _3963_/X VGND VGND VPWR VPWR pad_flash_io0_do sky130_fd_sc_hd__buf_8
Xoutput277 _6491_/Q VGND VGND VPWR VPWR pll_trim[11] sky130_fd_sc_hd__buf_8
X_5286_ _5601_/A0 hold767/X _5287_/S VGND VGND VPWR VPWR _5286_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput299 _6488_/Q VGND VGND VPWR VPWR pll_trim[8] sky130_fd_sc_hd__buf_8
Xoutput288 _6816_/Q VGND VGND VPWR VPWR pll_trim[21] sky130_fd_sc_hd__buf_8
X_4306_ hold497/X _6408_/A0 _4309_/S VGND VGND VPWR VPWR _4306_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7025_ _7081_/CLK _7025_/D fanout437/X VGND VGND VPWR VPWR _7025_/Q sky130_fd_sc_hd__dfrtp_2
X_4237_ _6700_/Q _6704_/D _6701_/Q _6702_/Q VGND VGND VPWR VPWR _4237_/X sky130_fd_sc_hd__or4_2
XFILLER_67_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4168_ _5254_/A0 hold895/X _4171_/S VGND VGND VPWR VPWR _4168_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4099_ _6408_/A0 hold495/X _4102_/S VGND VGND VPWR VPWR _4099_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6809_ _6810_/CLK _6809_/D fanout419/X VGND VGND VPWR VPWR _6809_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_70_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6770_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_164_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_23_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7133_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_38_csclk _7137_/CLK VGND VGND VPWR VPWR _6976_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_128_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold919 _6806_/Q VGND VGND VPWR VPWR hold919/X sky130_fd_sc_hd__bufbuf_16
Xhold908 _4300_/X VGND VGND VPWR VPWR _6749_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_170_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3470_ _3506_/A _3534_/A VGND VGND VPWR VPWR _4310_/A sky130_fd_sc_hd__nor2_8
XFILLER_170_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5140_ _5140_/A _5140_/B _5140_/C _5139_/X VGND VGND VPWR VPWR _5171_/C sky130_fd_sc_hd__or4b_4
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5071_ _5071_/A _5071_/B _5071_/C _5071_/D VGND VGND VPWR VPWR _5126_/A sky130_fd_sc_hd__or4_4
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4022_ hold889/X _4021_/X _4024_/S VGND VGND VPWR VPWR _4022_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5973_ _6638_/Q _5675_/X _5684_/X _6727_/Q _5972_/X VGND VGND VPWR VPWR _5976_/C
+ sky130_fd_sc_hd__a221o_1
X_4924_ _4756_/B _4660_/X _4624_/B _4930_/D VGND VGND VPWR VPWR _5098_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_80_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4855_ _4539_/D _4845_/B _4853_/X _4854_/X VGND VGND VPWR VPWR _4855_/X sky130_fd_sc_hd__a211o_1
X_4786_ _4772_/A _4399_/Y _4453_/Y _4689_/Y VGND VGND VPWR VPWR _4798_/C sky130_fd_sc_hd__a22o_1
X_3806_ _6487_/Q _6486_/Q VGND VGND VPWR VPWR _3841_/B sky130_fd_sc_hd__and2_2
XFILLER_193_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6525_ _6672_/CLK _6525_/D fanout453/X VGND VGND VPWR VPWR _6525_/Q sky130_fd_sc_hd__dfrtp_1
X_3737_ _6877_/Q _5288_/A _4055_/A _6540_/Q VGND VGND VPWR VPWR _3737_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3668_ _3668_/A _5234_/A VGND VGND VPWR VPWR _4004_/A sky130_fd_sc_hd__nor2_2
X_6456_ _6668_/CLK _6456_/D _6412_/X VGND VGND VPWR VPWR _6456_/Q sky130_fd_sc_hd__dfrtn_1
X_6387_ _6705_/Q _6387_/A2 _6387_/B1 _4238_/B _6386_/X VGND VGND VPWR VPWR _6387_/X
+ sky130_fd_sc_hd__a221o_1
X_5407_ hold314/X _5596_/A0 _5413_/S VGND VGND VPWR VPWR _6982_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3599_ _7072_/Q hold92/A _4166_/A _6637_/Q _3563_/X VGND VGND VPWR VPWR _3605_/A
+ sky130_fd_sc_hd__a221o_1
X_5338_ hold837/X _5599_/A0 _5341_/S VGND VGND VPWR VPWR _5338_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7008_ _7139_/CLK _7008_/D fanout434/X VGND VGND VPWR VPWR _7008_/Q sky130_fd_sc_hd__dfrtp_2
X_5269_ _5269_/A0 hold14/X _5269_/S VGND VGND VPWR VPWR _5269_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4640_ _4603_/B _5005_/C _5135_/A VGND VGND VPWR VPWR _4640_/X sky130_fd_sc_hd__o21ba_1
XFILLER_147_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4571_ _4572_/B _5147_/A VGND VGND VPWR VPWR _4571_/Y sky130_fd_sc_hd__nor2_4
XFILLER_128_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6310_ _6622_/Q _6022_/C _6032_/X _6652_/Q VGND VGND VPWR VPWR _6310_/X sky130_fd_sc_hd__a22o_1
Xhold727 _6670_/Q VGND VGND VPWR VPWR hold727/X sky130_fd_sc_hd__bufbuf_16
Xhold716 _4038_/X VGND VGND VPWR VPWR _6525_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3522_ _3522_/A _3522_/B _3522_/C _3522_/D VGND VGND VPWR VPWR _3547_/B sky130_fd_sc_hd__or4_1
Xhold705 _5230_/X VGND VGND VPWR VPWR _6828_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_171_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold738 _5322_/X VGND VGND VPWR VPWR _6907_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_116_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6241_ _6634_/Q _5653_/X _6311_/B _6654_/Q VGND VGND VPWR VPWR _6241_/X sky130_fd_sc_hd__a22o_1
XFILLER_89_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3453_ _3452_/X _6794_/Q _3857_/C VGND VGND VPWR VPWR _3453_/X sky130_fd_sc_hd__mux2_1
Xhold749 _4303_/X VGND VGND VPWR VPWR _6752_/D sky130_fd_sc_hd__bufbuf_16
X_6172_ _6890_/Q _6020_/A _6021_/D _7146_/Q _6171_/X VGND VGND VPWR VPWR _6172_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_131_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5123_ _5129_/B _5123_/B _5123_/C _5123_/D VGND VGND VPWR VPWR _5124_/D sky130_fd_sc_hd__and4b_4
XFILLER_97_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3384_ _5234_/A _5234_/B VGND VGND VPWR VPWR _5227_/A sky130_fd_sc_hd__nor2_8
XFILLER_57_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5054_ _4505_/X _4812_/C _5144_/B _4812_/X _4836_/X VGND VGND VPWR VPWR _5105_/C
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_97_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4005_ _6407_/A0 _4005_/A1 _4006_/S VGND VGND VPWR VPWR _6504_/D sky130_fd_sc_hd__mux2_1
XFILLER_38_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5956_ _6788_/Q _5690_/X _5693_/X _6657_/Q _5955_/X VGND VGND VPWR VPWR _5959_/C
+ sky130_fd_sc_hd__a221o_1
X_5887_ _6576_/Q _5689_/X _5698_/B _5886_/X VGND VGND VPWR VPWR _5887_/X sky130_fd_sc_hd__a22o_1
X_4907_ _4907_/A _5071_/C _4907_/C _4907_/D VGND VGND VPWR VPWR _4907_/X sky130_fd_sc_hd__or4_2
X_4838_ _5037_/A _4838_/B VGND VGND VPWR VPWR _4838_/X sky130_fd_sc_hd__or2_1
XFILLER_193_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4769_ _5013_/A _5135_/A VGND VGND VPWR VPWR _5142_/A sky130_fd_sc_hd__or2_4
X_6508_ _6987_/CLK _6508_/D fanout450/X VGND VGND VPWR VPWR _6508_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_134_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6439_ _6439_/A _6446_/B VGND VGND VPWR VPWR _6439_/X sky130_fd_sc_hd__and2_1
XFILLER_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold10 hold1/X VGND VGND VPWR VPWR hold10/X sky130_fd_sc_hd__bufbuf_16
Xhold32 hold40/X VGND VGND VPWR VPWR hold41/A sky130_fd_sc_hd__bufbuf_16
XFILLER_88_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold21 hold21/A VGND VGND VPWR VPWR hold21/X sky130_fd_sc_hd__bufbuf_16
XFILLER_48_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold65 hold65/A VGND VGND VPWR VPWR hold65/X sky130_fd_sc_hd__bufbuf_16
XFILLER_152_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold54 hold54/A VGND VGND VPWR VPWR hold54/X sky130_fd_sc_hd__bufbuf_16
XFILLER_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold43 hold43/A VGND VGND VPWR VPWR hold43/X sky130_fd_sc_hd__bufbuf_16
Xhold76 hold6/X VGND VGND VPWR VPWR hold76/X sky130_fd_sc_hd__bufbuf_16
XFILLER_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold87 hold87/A VGND VGND VPWR VPWR hold87/X sky130_fd_sc_hd__bufbuf_16
XFILLER_75_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold98 hold98/A VGND VGND VPWR VPWR hold98/X sky130_fd_sc_hd__bufbuf_16
XFILLER_152_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3240__1 _3545_/A1 VGND VGND VPWR VPWR _6458_/CLK sky130_fd_sc_hd__inv_2
XFILLER_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_7 _4002_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5810_ _7002_/Q _5667_/X _5687_/X _7050_/Q VGND VGND VPWR VPWR _5810_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6790_ _3545_/A1 _6790_/D _6448_/X VGND VGND VPWR VPWR _6790_/Q sky130_fd_sc_hd__dfrtn_1
X_5741_ _5741_/A _5741_/B _5741_/C VGND VGND VPWR VPWR _5741_/X sky130_fd_sc_hd__or3_1
XFILLER_50_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5672_ _7164_/Q _7163_/Q VGND VGND VPWR VPWR _5701_/C sky130_fd_sc_hd__and2_4
XFILLER_30_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4623_ _4623_/A _4623_/B _4623_/C _4623_/D VGND VGND VPWR VPWR _4623_/X sky130_fd_sc_hd__and4_1
XFILLER_175_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4554_ _4554_/A _4554_/B VGND VGND VPWR VPWR _4554_/X sky130_fd_sc_hd__and2_2
XFILLER_135_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold502 _4324_/X VGND VGND VPWR VPWR _6769_/D sky130_fd_sc_hd__bufbuf_16
Xhold535 _6625_/Q VGND VGND VPWR VPWR hold535/X sky130_fd_sc_hd__bufbuf_16
XFILLER_116_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold513 _6595_/Q VGND VGND VPWR VPWR hold513/X sky130_fd_sc_hd__bufbuf_16
X_3505_ _3514_/A _5252_/B VGND VGND VPWR VPWR _4172_/A sky130_fd_sc_hd__nor2_8
Xhold524 _4233_/X VGND VGND VPWR VPWR _6687_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_171_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4485_ _4485_/A VGND VGND VPWR VPWR _4554_/A sky130_fd_sc_hd__clkinv_2
Xhold579 _6962_/Q VGND VGND VPWR VPWR hold579/X sky130_fd_sc_hd__bufbuf_16
Xhold546 _5349_/X VGND VGND VPWR VPWR _6931_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_144_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6224_ _6908_/Q _6021_/A _6025_/A _6940_/Q _6223_/X VGND VGND VPWR VPWR _6231_/A
+ sky130_fd_sc_hd__a221o_1
Xhold557 _6590_/Q VGND VGND VPWR VPWR hold557/X sky130_fd_sc_hd__bufbuf_16
Xhold568 _6744_/Q VGND VGND VPWR VPWR hold568/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3436_ _3436_/A _3436_/B _3436_/C _3436_/D VGND VGND VPWR VPWR _3452_/A sky130_fd_sc_hd__or4_4
X_6155_ _6977_/Q _6023_/B _6021_/C _6881_/Q _6154_/X VGND VGND VPWR VPWR _6156_/D
+ sky130_fd_sc_hd__a221o_1
X_3367_ hold90/X _3421_/C VGND VGND VPWR VPWR _3473_/B sky130_fd_sc_hd__or2_4
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _4745_/A _4947_/B _5017_/A VGND VGND VPWR VPWR _5108_/B sky130_fd_sc_hd__a21oi_1
Xhold1202 _6722_/Q VGND VGND VPWR VPWR _4267_/A0 sky130_fd_sc_hd__bufbuf_16
Xhold1213 _6535_/Q VGND VGND VPWR VPWR _4050_/A0 sky130_fd_sc_hd__bufbuf_16
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6086_ _7190_/Q _6309_/S _6084_/X _6085_/X VGND VGND VPWR VPWR _7190_/D sky130_fd_sc_hd__o22a_1
Xhold1224 _6837_/Q VGND VGND VPWR VPWR _5243_/A1 sky130_fd_sc_hd__bufbuf_16
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1235 _4041_/X VGND VGND VPWR VPWR hold131/A sky130_fd_sc_hd__bufbuf_16
Xhold1246 _7114_/Q VGND VGND VPWR VPWR _5555_/A0 sky130_fd_sc_hd__bufbuf_16
X_5037_ _5037_/A _5037_/B _5003_/X VGND VGND VPWR VPWR _5158_/A sky130_fd_sc_hd__or3b_4
XFILLER_57_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1257 _7087_/Q VGND VGND VPWR VPWR _5525_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_45_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3298_ _3501_/A _3668_/A VGND VGND VPWR VPWR _5486_/A sky130_fd_sc_hd__nor2_8
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_408 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_419 _3971_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6988_ _7156_/CLK _6988_/D fanout452/X VGND VGND VPWR VPWR _6988_/Q sky130_fd_sc_hd__dfrtp_2
X_5939_ _5611_/A _7185_/Q _6358_/B1 VGND VGND VPWR VPWR _5939_/X sky130_fd_sc_hd__a21o_1
XFILLER_193_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput111 wb_adr_i[20] VGND VGND VPWR VPWR _4722_/A sky130_fd_sc_hd__buf_8
Xinput100 wb_adr_i[10] VGND VGND VPWR VPWR _4351_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_163_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput133 wb_dat_i[10] VGND VGND VPWR VPWR _6384_/B1 sky130_fd_sc_hd__clkbuf_4
Xinput144 wb_dat_i[20] VGND VGND VPWR VPWR _6389_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput122 wb_adr_i[30] VGND VGND VPWR VPWR _3892_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_163_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput166 wb_sel_i[1] VGND VGND VPWR VPWR _6371_/B sky130_fd_sc_hd__clkbuf_4
Xinput155 wb_dat_i[30] VGND VGND VPWR VPWR _6396_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_76_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4270_ hold609/X _6408_/A0 _4273_/S VGND VGND VPWR VPWR _4270_/X sky130_fd_sc_hd__mux2_1
X_3221_ _7008_/Q VGND VGND VPWR VPWR _3221_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6911_ _7151_/CLK _6911_/D fanout446/X VGND VGND VPWR VPWR _6911_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_62_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6842_ _6851_/CLK _6842_/D _6454_/A VGND VGND VPWR VPWR _6842_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3985_ hold133/X hold151/X _6689_/Q VGND VGND VPWR VPWR _3985_/X sky130_fd_sc_hd__mux2_8
X_6773_ _6851_/CLK _6773_/D fanout418/X VGND VGND VPWR VPWR _6773_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_176_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5724_ _6998_/Q _5667_/X _5687_/X _7046_/Q VGND VGND VPWR VPWR _5724_/X sky130_fd_sc_hd__a22o_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5655_ _6679_/Q _5653_/X _5654_/Y _7171_/Q VGND VGND VPWR VPWR _7171_/D sky130_fd_sc_hd__a22o_1
XFILLER_190_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4606_ _4775_/A _4694_/A VGND VGND VPWR VPWR _4917_/A sky130_fd_sc_hd__or2_2
XFILLER_136_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold310 _4027_/X VGND VGND VPWR VPWR _6515_/D sky130_fd_sc_hd__bufbuf_16
X_5586_ _5595_/A0 hold988/X _5593_/S VGND VGND VPWR VPWR _7141_/D sky130_fd_sc_hd__mux2_1
XFILLER_190_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4537_ _4533_/A _4533_/B _4537_/C _4538_/A VGND VGND VPWR VPWR _4537_/X sky130_fd_sc_hd__and4bb_4
Xhold332 _6934_/Q VGND VGND VPWR VPWR hold332/X sky130_fd_sc_hd__bufbuf_16
Xhold321 _6523_/Q VGND VGND VPWR VPWR hold321/X sky130_fd_sc_hd__bufbuf_16
XFILLER_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold343 _4186_/X VGND VGND VPWR VPWR _6650_/D sky130_fd_sc_hd__bufbuf_16
X_4468_ _4758_/A _5004_/A VGND VGND VPWR VPWR _4818_/C sky130_fd_sc_hd__nand2_4
Xhold387 _5314_/X VGND VGND VPWR VPWR _6900_/D sky130_fd_sc_hd__bufbuf_16
Xhold365 _7054_/Q VGND VGND VPWR VPWR hold365/X sky130_fd_sc_hd__bufbuf_16
Xhold376 _6632_/Q VGND VGND VPWR VPWR hold376/X sky130_fd_sc_hd__bufbuf_16
Xhold354 _5220_/X VGND VGND VPWR VPWR _6821_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_131_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6207_ _6232_/A _6207_/B _6207_/C _6207_/D VGND VGND VPWR VPWR _6207_/X sky130_fd_sc_hd__or4_4
X_7187_ _7201_/CLK _7187_/D fanout419/X VGND VGND VPWR VPWR _7187_/Q sky130_fd_sc_hd__dfrtp_4
X_3419_ _3419_/A _3421_/C VGND VGND VPWR VPWR _3732_/B sky130_fd_sc_hd__or2_4
Xhold398 _6948_/Q VGND VGND VPWR VPWR hold398/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4399_ _4400_/A _4513_/A VGND VGND VPWR VPWR _4399_/Y sky130_fd_sc_hd__nor2_4
X_6138_ _7025_/Q _6010_/Y _6031_/X _7089_/Q _6137_/X VGND VGND VPWR VPWR _6144_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_98_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1021 _6965_/Q VGND VGND VPWR VPWR _5388_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_133_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1032 _6661_/Q VGND VGND VPWR VPWR _4199_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1010 _6842_/Q VGND VGND VPWR VPWR _5249_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_93_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1065 _6593_/Q VGND VGND VPWR VPWR _4117_/A1 sky130_fd_sc_hd__bufbuf_16
X_6069_ _7070_/Q _6009_/X _6020_/D _6966_/Q VGND VGND VPWR VPWR _6069_/X sky130_fd_sc_hd__a22o_1
Xhold1043 _6549_/Q VGND VGND VPWR VPWR _4066_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_58_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1076 _6853_/Q VGND VGND VPWR VPWR _5262_/A0 sky130_fd_sc_hd__bufbuf_16
Xhold1054 _6777_/Q VGND VGND VPWR VPWR _4333_/A1 sky130_fd_sc_hd__bufbuf_16
XANTENNA_216 _6735_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_205 _7033_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1098 _7045_/Q VGND VGND VPWR VPWR _5478_/A0 sky130_fd_sc_hd__bufbuf_16
Xhold1087 _7093_/Q VGND VGND VPWR VPWR _5532_/A1 sky130_fd_sc_hd__bufbuf_16
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_227 _6475_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_238 mask_rev_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_249 mask_rev_in[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3770_ _7109_/Q hold85/A _5185_/A _6785_/Q _3745_/X VGND VGND VPWR VPWR _3793_/A
+ sky130_fd_sc_hd__a221o_4
XFILLER_13_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5440_ _5584_/A0 hold474/X _5440_/S VGND VGND VPWR VPWR _5440_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5371_ _5587_/A0 hold695/X _5377_/S VGND VGND VPWR VPWR _6950_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7110_ _7150_/CLK _7110_/D fanout446/X VGND VGND VPWR VPWR _7110_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_153_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4322_ _4322_/A _6406_/B VGND VGND VPWR VPWR _4327_/S sky130_fd_sc_hd__nand2_4
XFILLER_141_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4253_ _5561_/A0 hold690/X _4255_/S VGND VGND VPWR VPWR _6710_/D sky130_fd_sc_hd__mux2_1
X_7041_ _7129_/CLK _7041_/D fanout429/X VGND VGND VPWR VPWR _7041_/Q sky130_fd_sc_hd__dfrtp_2
X_3204_ _7144_/Q VGND VGND VPWR VPWR _3204_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4184_ _4184_/A _5558_/B VGND VGND VPWR VPWR _4189_/S sky130_fd_sc_hd__and2_4
XFILLER_79_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A VGND VGND VPWR VPWR _3949_/A1 sky130_fd_sc_hd__clkbuf_8
X_6825_ _6825_/CLK _6825_/D fanout429/X VGND VGND VPWR VPWR _6825_/Q sky130_fd_sc_hd__dfrtp_2
X_3968_ _6706_/Q _3974_/B VGND VGND VPWR VPWR _6700_/D sky130_fd_sc_hd__and2_1
X_6756_ _6770_/CLK _6756_/D fanout423/X VGND VGND VPWR VPWR _6756_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5707_ _7165_/Q _5707_/B _5707_/C VGND VGND VPWR VPWR _5707_/X sky130_fd_sc_hd__and3_4
XFILLER_176_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3899_ _6664_/Q _3898_/A _3898_/Y _6666_/Q VGND VGND VPWR VPWR _6664_/D sky130_fd_sc_hd__a22o_1
X_6687_ _6851_/CLK _6687_/D _6455_/A VGND VGND VPWR VPWR _6687_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5638_ _7167_/Q _7166_/Q VGND VGND VPWR VPWR _6037_/B sky130_fd_sc_hd__and2_4
XFILLER_163_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5569_ _5578_/A0 hold341/X _5575_/S VGND VGND VPWR VPWR _7126_/D sky130_fd_sc_hd__mux2_1
Xhold151 _7214_/Q VGND VGND VPWR VPWR hold151/X sky130_fd_sc_hd__bufbuf_16
Xhold140 _7152_/Q VGND VGND VPWR VPWR hold140/X sky130_fd_sc_hd__bufbuf_16
XFILLER_163_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold162 _4006_/X VGND VGND VPWR VPWR _6505_/D sky130_fd_sc_hd__bufbuf_16
Xhold184 hold184/A VGND VGND VPWR VPWR hold184/X sky130_fd_sc_hd__bufbuf_16
Xhold173 _6782_/Q VGND VGND VPWR VPWR hold173/X sky130_fd_sc_hd__bufbuf_16
XFILLER_2_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold195 hold52/X VGND VGND VPWR VPWR _3275_/C sky130_fd_sc_hd__bufbuf_16
XFILLER_120_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4940_ _5034_/A _4940_/B _4940_/C _4940_/D VGND VGND VPWR VPWR _4941_/D sky130_fd_sc_hd__or4_1
XFILLER_91_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4871_ _4871_/A _5164_/B VGND VGND VPWR VPWR _4899_/B sky130_fd_sc_hd__and2_4
XFILLER_32_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6610_ _6843_/CLK _6610_/D fanout440/X VGND VGND VPWR VPWR _6610_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3822_ _3821_/X hold50/A _3840_/S VGND VGND VPWR VPWR _6483_/D sky130_fd_sc_hd__mux2_1
XFILLER_60_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6541_ _6786_/CLK _6541_/D fanout417/X VGND VGND VPWR VPWR _6541_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_193_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3753_ _6973_/Q _5396_/A _4130_/A _6604_/Q _3752_/X VGND VGND VPWR VPWR _3754_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6472_ _3957_/A1 _6472_/D _6427_/X VGND VGND VPWR VPWR _6472_/Q sky130_fd_sc_hd__dfrtp_2
X_3684_ _7086_/Q hold54/A _5513_/A _7078_/Q _3683_/X VGND VGND VPWR VPWR _3687_/B
+ sky130_fd_sc_hd__a221o_1
Xoutput201 _3207_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[33] sky130_fd_sc_hd__buf_8
XFILLER_173_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5423_ _5423_/A hold47/X VGND VGND VPWR VPWR hold48/A sky130_fd_sc_hd__nand2_8
Xoutput234 _6519_/Q VGND VGND VPWR VPWR mgmt_gpio_out[29] sky130_fd_sc_hd__buf_8
X_5354_ _5588_/A0 _5354_/A1 _5359_/S VGND VGND VPWR VPWR _5354_/X sky130_fd_sc_hd__mux2_1
Xoutput223 _6672_/Q VGND VGND VPWR VPWR mgmt_gpio_out[19] sky130_fd_sc_hd__buf_8
XFILLER_133_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput212 _3231_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[9] sky130_fd_sc_hd__buf_8
XFILLER_99_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput245 _6685_/Q VGND VGND VPWR VPWR mgmt_gpio_out[4] sky130_fd_sc_hd__buf_8
Xoutput256 _3960_/A VGND VGND VPWR VPWR pad_flash_io0_ieb sky130_fd_sc_hd__buf_8
Xoutput267 _6801_/Q VGND VGND VPWR VPWR pll_div[1] sky130_fd_sc_hd__buf_8
X_4305_ _4305_/A0 _6407_/A0 _4309_/S VGND VGND VPWR VPWR _4305_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5285_ hold78/X hold264/X _5287_/S VGND VGND VPWR VPWR _5285_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput278 _6492_/Q VGND VGND VPWR VPWR pll_trim[12] sky130_fd_sc_hd__buf_8
Xoutput289 _6817_/Q VGND VGND VPWR VPWR pll_trim[22] sky130_fd_sc_hd__buf_8
X_4236_ _6706_/Q _6705_/Q _6707_/Q VGND VGND VPWR VPWR _4238_/B sky130_fd_sc_hd__nor3_4
XFILLER_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7024_ _7101_/CLK _7024_/D fanout430/X VGND VGND VPWR VPWR _7024_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_101_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4167_ _5234_/C _4167_/A1 _4171_/S VGND VGND VPWR VPWR _4167_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4098_ _6407_/A0 _4098_/A1 _4102_/S VGND VGND VPWR VPWR _4098_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_4_csclk _6722_/CLK VGND VGND VPWR VPWR _6717_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_82_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6808_ _6810_/CLK _6808_/D fanout419/X VGND VGND VPWR VPWR _6808_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_51_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6739_ _6759_/CLK _6739_/D fanout421/X VGND VGND VPWR VPWR _6739_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout450 fanout451/X VGND VGND VPWR VPWR fanout450/X sky130_fd_sc_hd__buf_8
XFILLER_171_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold909 _6497_/Q VGND VGND VPWR VPWR hold909/X sky130_fd_sc_hd__bufbuf_16
XFILLER_115_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5070_ _4749_/C _5005_/C _4965_/A VGND VGND VPWR VPWR _5076_/C sky130_fd_sc_hd__a21oi_1
XFILLER_97_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4021_ _4041_/A1 _5601_/A0 _4023_/S VGND VGND VPWR VPWR _4021_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5972_ _6549_/Q _5674_/X _5688_/X _6772_/Q VGND VGND VPWR VPWR _5972_/X sky130_fd_sc_hd__a22o_1
XFILLER_64_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4923_ _4672_/A _4672_/B _4711_/C _4936_/B _4936_/C VGND VGND VPWR VPWR _5024_/C
+ sky130_fd_sc_hd__a311o_1
XFILLER_80_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4854_ _4409_/Y _4845_/B _4846_/X VGND VGND VPWR VPWR _4854_/X sky130_fd_sc_hd__a21o_1
XFILLER_178_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4785_ _4500_/A _4622_/B _4758_/C _4689_/Y VGND VGND VPWR VPWR _5180_/A sky130_fd_sc_hd__a22o_1
X_3805_ _6664_/Q _3845_/A VGND VGND VPWR VPWR _3825_/B sky130_fd_sc_hd__nand2b_2
X_6524_ _6987_/CLK _6524_/D fanout450/X VGND VGND VPWR VPWR _6524_/Q sky130_fd_sc_hd__dfrtp_1
X_3736_ input43/X _4217_/S _3552_/Y _6820_/Q VGND VGND VPWR VPWR _3736_/X sky130_fd_sc_hd__a22o_2
XFILLER_119_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6455_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6455_/X sky130_fd_sc_hd__and2_1
X_3667_ _3666_/X _6792_/Q _3928_/A VGND VGND VPWR VPWR _6792_/D sky130_fd_sc_hd__mux2_1
X_6386_ _6707_/Q _6386_/A2 _6386_/B1 _6706_/Q VGND VGND VPWR VPWR _6386_/X sky130_fd_sc_hd__a22o_1
X_5406_ hold975/X _5595_/A0 _5413_/S VGND VGND VPWR VPWR _6981_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3598_ _3598_/A _3598_/B _3598_/C _3598_/D VGND VGND VPWR VPWR _3606_/C sky130_fd_sc_hd__or4_4
X_5337_ hold663/X _5571_/A0 _5341_/S VGND VGND VPWR VPWR _5337_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5268_ hold706/X _5583_/A0 _5269_/S VGND VGND VPWR VPWR _5268_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4219_ _5252_/B _6454_/B _4007_/X _4234_/S hold47/X VGND VGND VPWR VPWR _4235_/S
+ sky130_fd_sc_hd__o221a_4
X_7007_ _7135_/CLK _7007_/D fanout431/X VGND VGND VPWR VPWR _7007_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_75_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5199_ _6411_/A0 hold823/X _5199_/S VGND VGND VPWR VPWR _5199_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4570_ _5071_/A VGND VGND VPWR VPWR _4623_/B sky130_fd_sc_hd__inv_2
X_3521_ _6937_/Q _5351_/A _4280_/A _6737_/Q _3519_/X VGND VGND VPWR VPWR _3522_/D
+ sky130_fd_sc_hd__a221o_4
XFILLER_128_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold728 _4206_/X VGND VGND VPWR VPWR _6670_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_116_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold706 _6859_/Q VGND VGND VPWR VPWR hold706/X sky130_fd_sc_hd__bufbuf_16
Xhold717 _7007_/Q VGND VGND VPWR VPWR hold717/X sky130_fd_sc_hd__bufbuf_16
X_6240_ _6535_/Q _6025_/D _6029_/X _6639_/Q _6239_/X VGND VGND VPWR VPWR _6247_/A
+ sky130_fd_sc_hd__a221o_2
X_3452_ _3452_/A _3452_/B _3452_/C _3452_/D VGND VGND VPWR VPWR _3452_/X sky130_fd_sc_hd__or4_4
Xhold739 _6742_/Q VGND VGND VPWR VPWR hold739/X sky130_fd_sc_hd__bufbuf_16
XFILLER_170_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6171_ _7114_/Q _6027_/B _6021_/B _7154_/Q VGND VGND VPWR VPWR _6171_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3383_ _3421_/A _3421_/B _3383_/C VGND VGND VPWR VPWR _5234_/B sky130_fd_sc_hd__or3_4
X_5122_ _4749_/C _5005_/C _4898_/B _4953_/A VGND VGND VPWR VPWR _5124_/C sky130_fd_sc_hd__a31o_2
XFILLER_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5053_ _4745_/A _4648_/B _5164_/B _4818_/C _5052_/X VGND VGND VPWR VPWR _5157_/A
+ sky130_fd_sc_hd__o221ai_2
XFILLER_84_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4004_ _4004_/A _5576_/B VGND VGND VPWR VPWR _4006_/S sky130_fd_sc_hd__nand2_1
XFILLER_38_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5955_ _6751_/Q _5682_/X _5703_/X _6543_/Q VGND VGND VPWR VPWR _5955_/X sky130_fd_sc_hd__a22o_1
X_5886_ _6624_/Q _5963_/B VGND VGND VPWR VPWR _5886_/X sky130_fd_sc_hd__or2_1
X_4906_ _5174_/C _4906_/B _4906_/C _4906_/D VGND VGND VPWR VPWR _4907_/D sky130_fd_sc_hd__or4_1
X_4837_ _4588_/X _4717_/B _4757_/B _5164_/B VGND VGND VPWR VPWR _4837_/X sky130_fd_sc_hd__o22a_1
XFILLER_139_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4768_ _4772_/A _4409_/Y _4453_/Y _4656_/X VGND VGND VPWR VPWR _4796_/B sky130_fd_sc_hd__a22o_1
X_6507_ _6672_/CLK _6507_/D fanout453/X VGND VGND VPWR VPWR _6507_/Q sky130_fd_sc_hd__dfrtp_2
X_4699_ _4595_/B _4697_/Y _4698_/Y _5165_/A VGND VGND VPWR VPWR _4713_/A sky130_fd_sc_hd__o31a_1
XFILLER_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3719_ input72/X _4023_/S _4178_/A _6645_/Q _3718_/X VGND VGND VPWR VPWR _3725_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6438_ _6439_/A _6446_/B VGND VGND VPWR VPWR _6438_/X sky130_fd_sc_hd__and2_1
XFILLER_115_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_22_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _6833_/CLK sky130_fd_sc_hd__clkbuf_8
X_6369_ _7209_/Q _3415_/X _6370_/S VGND VGND VPWR VPWR _7209_/D sky130_fd_sc_hd__mux2_1
Xhold11 hold11/A VGND VGND VPWR VPWR hold2/A sky130_fd_sc_hd__bufbuf_16
Xhold22 hold22/A VGND VGND VPWR VPWR hold22/X sky130_fd_sc_hd__bufbuf_16
Xhold33 hold42/X VGND VGND VPWR VPWR hold43/A sky130_fd_sc_hd__bufbuf_16
XFILLER_75_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold44 hold44/A VGND VGND VPWR VPWR hold44/X sky130_fd_sc_hd__bufbuf_16
Xhold55 hold55/A VGND VGND VPWR VPWR hold55/X sky130_fd_sc_hd__bufbuf_16
Xhold77 hold77/A VGND VGND VPWR VPWR hold7/A sky130_fd_sc_hd__bufbuf_16
XFILLER_152_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold66 hold66/A VGND VGND VPWR VPWR hold66/X sky130_fd_sc_hd__bufbuf_16
Xhold88 hold88/A VGND VGND VPWR VPWR hold88/X sky130_fd_sc_hd__bufbuf_16
Xhold99 hold99/A VGND VGND VPWR VPWR hold99/X sky130_fd_sc_hd__bufbuf_16
XFILLER_29_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_37_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _6987_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_90_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] VGND VGND VPWR VPWR clkbuf_0_mgmt_gpio_in[4]/X
+ sky130_fd_sc_hd__clkbuf_8
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_8 _4016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5740_ _6942_/Q _5705_/X _5707_/X _7022_/Q _5739_/X VGND VGND VPWR VPWR _5741_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_188_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5671_ _7162_/Q _7161_/Q VGND VGND VPWR VPWR _5707_/B sky130_fd_sc_hd__and2b_4
XFILLER_30_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4622_ _4987_/A _4622_/B VGND VGND VPWR VPWR _4623_/D sky130_fd_sc_hd__nand2_1
X_4553_ _4553_/A _4553_/B _4986_/C VGND VGND VPWR VPWR _4554_/B sky130_fd_sc_hd__nor3_2
XFILLER_116_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4484_ _4533_/A _4484_/B _4484_/C VGND VGND VPWR VPWR _4485_/A sky130_fd_sc_hd__or3_2
Xhold536 _4156_/X VGND VGND VPWR VPWR _6625_/D sky130_fd_sc_hd__bufbuf_16
Xhold525 _6524_/Q VGND VGND VPWR VPWR hold525/X sky130_fd_sc_hd__bufbuf_16
Xhold503 _6605_/Q VGND VGND VPWR VPWR hold503/X sky130_fd_sc_hd__bufbuf_16
Xhold514 _4120_/X VGND VGND VPWR VPWR _6595_/D sky130_fd_sc_hd__bufbuf_16
X_3504_ _3504_/A _3504_/B _3504_/C _3504_/D VGND VGND VPWR VPWR _3547_/A sky130_fd_sc_hd__or4_4
Xhold547 _7110_/Q VGND VGND VPWR VPWR hold547/X sky130_fd_sc_hd__bufbuf_16
X_3435_ input57/X _4025_/A _5594_/A _7154_/Q _3424_/X VGND VGND VPWR VPWR _3436_/D
+ sky130_fd_sc_hd__a221o_4
XFILLER_116_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6223_ _6956_/Q _6022_/A _6025_/C _6932_/Q VGND VGND VPWR VPWR _6223_/X sky130_fd_sc_hd__a22o_1
Xhold558 _4114_/X VGND VGND VPWR VPWR _6590_/D sky130_fd_sc_hd__bufbuf_16
Xhold569 _4294_/X VGND VGND VPWR VPWR _6744_/D sky130_fd_sc_hd__bufbuf_16
X_6154_ _7065_/Q _5996_/X _6020_/C _6913_/Q VGND VGND VPWR VPWR _6154_/X sky130_fd_sc_hd__a22o_1
XFILLER_106_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3366_ _7084_/Q _5513_/A hold61/A _7140_/Q VGND VGND VPWR VPWR _3366_/X sky130_fd_sc_hd__a22o_1
X_5105_ _5105_/A _5105_/B _5105_/C VGND VGND VPWR VPWR _5157_/B sky130_fd_sc_hd__or3_2
X_3297_ _7012_/Q _5432_/A hold92/A _7076_/Q _3296_/X VGND VGND VPWR VPWR _3379_/A
+ sky130_fd_sc_hd__a221o_1
Xhold1214 _4050_/X VGND VGND VPWR VPWR _6535_/D sky130_fd_sc_hd__bufbuf_16
Xhold1203 _6488_/Q VGND VGND VPWR VPWR _3980_/A0 sky130_fd_sc_hd__bufbuf_16
X_6085_ _5663_/A _7189_/Q _6358_/B1 VGND VGND VPWR VPWR _6085_/X sky130_fd_sc_hd__a21o_1
Xhold1225 _5243_/X VGND VGND VPWR VPWR _6837_/D sky130_fd_sc_hd__bufbuf_16
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1236 _6695_/Q VGND VGND VPWR VPWR _4247_/A1 sky130_fd_sc_hd__bufbuf_16
X_5036_ _5036_/A _5101_/A _5036_/C VGND VGND VPWR VPWR _5036_/X sky130_fd_sc_hd__or3_1
XFILLER_57_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1258 _7041_/Q VGND VGND VPWR VPWR _5473_/A1 sky130_fd_sc_hd__bufbuf_16
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1247 _6860_/Q VGND VGND VPWR VPWR _5269_/A0 sky130_fd_sc_hd__bufbuf_16
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_409 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6987_ _6987_/CLK _6987_/D fanout453/X VGND VGND VPWR VPWR _6987_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5938_ _6532_/Q _5722_/B _5927_/X _5937_/X _6308_/S VGND VGND VPWR VPWR _5938_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5869_ _7092_/Q _5685_/X _5701_/X _6956_/Q VGND VGND VPWR VPWR _5869_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput101 wb_adr_i[11] VGND VGND VPWR VPWR _4351_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_163_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput145 wb_dat_i[21] VGND VGND VPWR VPWR _6392_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput134 wb_dat_i[11] VGND VGND VPWR VPWR _6386_/B1 sky130_fd_sc_hd__clkbuf_4
Xinput123 wb_adr_i[31] VGND VGND VPWR VPWR _3892_/A sky130_fd_sc_hd__clkbuf_4
Xinput112 wb_adr_i[21] VGND VGND VPWR VPWR _4368_/A sky130_fd_sc_hd__buf_4
XFILLER_103_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput167 wb_sel_i[2] VGND VGND VPWR VPWR _6372_/B sky130_fd_sc_hd__clkbuf_4
Xinput156 wb_dat_i[31] VGND VGND VPWR VPWR _6398_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_102_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3220_ _7016_/Q VGND VGND VPWR VPWR _3220_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6910_ _7151_/CLK _6910_/D fanout446/X VGND VGND VPWR VPWR _6910_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_63_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6841_ _6939_/CLK _6841_/D fanout453/X VGND VGND VPWR VPWR _6841_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_62_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3984_ hold997/X _6409_/A0 _3994_/S VGND VGND VPWR VPWR _6490_/D sky130_fd_sc_hd__mux2_1
X_6772_ _7222_/CLK _6772_/D fanout422/X VGND VGND VPWR VPWR _6772_/Q sky130_fd_sc_hd__dfrtp_2
X_5723_ _5663_/Y _5721_/X _5722_/X _6358_/B1 _7176_/Q VGND VGND VPWR VPWR _7176_/D
+ sky130_fd_sc_hd__a32o_1
X_5654_ _5654_/A _5654_/B VGND VGND VPWR VPWR _5654_/Y sky130_fd_sc_hd__nor2_1
XFILLER_176_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4605_ _5023_/A _4694_/A VGND VGND VPWR VPWR _4787_/B sky130_fd_sc_hd__nor2_1
XFILLER_117_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold311 _6926_/Q VGND VGND VPWR VPWR hold311/X sky130_fd_sc_hd__bufbuf_16
X_5585_ _5585_/A _5594_/B VGND VGND VPWR VPWR _5593_/S sky130_fd_sc_hd__nand2_8
XFILLER_163_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold300 _5518_/X VGND VGND VPWR VPWR _7081_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_7_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4536_ _4949_/B _4536_/B VGND VGND VPWR VPWR _4536_/X sky130_fd_sc_hd__and2_4
Xhold333 _6966_/Q VGND VGND VPWR VPWR hold333/X sky130_fd_sc_hd__bufbuf_16
Xhold322 _4036_/X VGND VGND VPWR VPWR _6523_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_144_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold344 _6564_/Q VGND VGND VPWR VPWR hold344/X sky130_fd_sc_hd__bufbuf_16
X_4467_ _4722_/A _4467_/B VGND VGND VPWR VPWR _4819_/B sky130_fd_sc_hd__nand2_8
Xhold355 _6529_/Q VGND VGND VPWR VPWR hold355/X sky130_fd_sc_hd__bufbuf_16
Xhold377 _6884_/Q VGND VGND VPWR VPWR hold377/X sky130_fd_sc_hd__bufbuf_16
XFILLER_171_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold366 _6892_/Q VGND VGND VPWR VPWR hold366/X sky130_fd_sc_hd__bufbuf_16
XFILLER_132_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold388 _7130_/Q VGND VGND VPWR VPWR hold388/X sky130_fd_sc_hd__bufbuf_16
XFILLER_132_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4398_ _4930_/D VGND VGND VPWR VPWR _4398_/Y sky130_fd_sc_hd__inv_2
X_3418_ _7130_/Q _5567_/A _5558_/A _7122_/Q VGND VGND VPWR VPWR _3418_/X sky130_fd_sc_hd__a22o_1
X_6206_ _6206_/A _6206_/B _6206_/C _6206_/D VGND VGND VPWR VPWR _6207_/D sky130_fd_sc_hd__or4_2
X_7186_ _7201_/CLK _7186_/D fanout420/X VGND VGND VPWR VPWR _7186_/Q sky130_fd_sc_hd__dfrtp_4
Xhold399 _5368_/X VGND VGND VPWR VPWR _6948_/D sky130_fd_sc_hd__bufbuf_16
X_6137_ _7137_/Q _6020_/B _6011_/X _7097_/Q VGND VGND VPWR VPWR _6137_/X sky130_fd_sc_hd__a22o_1
XFILLER_58_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3349_ _3506_/A _3386_/B VGND VGND VPWR VPWR _5423_/A sky130_fd_sc_hd__nor2_8
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1000 _6776_/Q VGND VGND VPWR VPWR _4332_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_112_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1033 _6662_/Q VGND VGND VPWR VPWR _4200_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1011 _5249_/X VGND VGND VPWR VPWR _6842_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_46_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1022 _6767_/Q VGND VGND VPWR VPWR _4321_/A0 sky130_fd_sc_hd__bufbuf_16
XFILLER_133_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1066 _4117_/X VGND VGND VPWR VPWR _6593_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_73_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1044 _4066_/X VGND VGND VPWR VPWR _6549_/D sky130_fd_sc_hd__bufbuf_16
Xhold1055 _4333_/X VGND VGND VPWR VPWR _6777_/D sky130_fd_sc_hd__bufbuf_16
X_6068_ _6998_/Q _5987_/Y _6022_/D _6918_/Q _6067_/X VGND VGND VPWR VPWR _6071_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1099 _6540_/Q VGND VGND VPWR VPWR _4056_/A1 sky130_fd_sc_hd__bufbuf_16
X_5019_ _5003_/X _5018_/X _6376_/A VGND VGND VPWR VPWR _5019_/X sky130_fd_sc_hd__a21o_1
XFILLER_100_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1077 _7061_/Q VGND VGND VPWR VPWR _5496_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1088 _6756_/Q VGND VGND VPWR VPWR _4308_/A0 sky130_fd_sc_hd__bufbuf_16
XANTENNA_206 _7055_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_217 _7141_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_228 _6475_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_239 mask_rev_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5370_ _5595_/A0 _5370_/A1 _5377_/S VGND VGND VPWR VPWR _6949_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4321_ _4321_/A0 _5545_/A0 _4321_/S VGND VGND VPWR VPWR _4321_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4252_ _6408_/A0 hold489/X _4255_/S VGND VGND VPWR VPWR _4252_/X sky130_fd_sc_hd__mux2_1
X_7040_ _7140_/CLK _7040_/D fanout432/X VGND VGND VPWR VPWR _7040_/Q sky130_fd_sc_hd__dfrtp_2
X_3203_ _7152_/Q VGND VGND VPWR VPWR _3203_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_67_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4183_ _4183_/A0 _5545_/A0 _4183_/S VGND VGND VPWR VPWR _4183_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6824_ _6824_/CLK _6824_/D _6446_/A VGND VGND VPWR VPWR _6824_/Q sky130_fd_sc_hd__dfrtp_4
X_3967_ _6703_/Q _3974_/B VGND VGND VPWR VPWR _6701_/D sky130_fd_sc_hd__and2_1
X_6755_ _6770_/CLK _6755_/D fanout423/X VGND VGND VPWR VPWR _6755_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_50_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5706_ _7165_/Q _5706_/B _5707_/B VGND VGND VPWR VPWR _5706_/X sky130_fd_sc_hd__and3_4
XFILLER_50_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6686_ _7138_/CLK _6686_/D fanout438/X VGND VGND VPWR VPWR _6686_/Q sky130_fd_sc_hd__dfrtp_2
X_3898_ _3898_/A _3898_/B VGND VGND VPWR VPWR _3898_/Y sky130_fd_sc_hd__nor2_1
XFILLER_148_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5637_ _5621_/X _5663_/B _7166_/Q VGND VGND VPWR VPWR _7166_/D sky130_fd_sc_hd__mux2_1
X_5568_ _5595_/A0 hold961/X _5575_/S VGND VGND VPWR VPWR _7125_/D sky130_fd_sc_hd__mux2_1
XFILLER_151_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold130 hold208/X VGND VGND VPWR VPWR hold209/A sky130_fd_sc_hd__bufbuf_16
Xhold141 _5598_/X VGND VGND VPWR VPWR _7152_/D sky130_fd_sc_hd__bufbuf_16
Xhold152 _3985_/X VGND VGND VPWR VPWR hold152/X sky130_fd_sc_hd__bufbuf_16
X_4519_ _4871_/A _4995_/A VGND VGND VPWR VPWR _4519_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5499_ hold71/X hold163/X _5503_/S VGND VGND VPWR VPWR _5499_/X sky130_fd_sc_hd__mux2_1
Xhold163 _7064_/Q VGND VGND VPWR VPWR hold163/X sky130_fd_sc_hd__bufbuf_16
Xhold174 _3251_/X VGND VGND VPWR VPWR hold59/A sky130_fd_sc_hd__bufbuf_16
Xhold185 hold185/A VGND VGND VPWR VPWR hold185/X sky130_fd_sc_hd__bufbuf_16
XFILLER_132_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold196 _3334_/Y VGND VGND VPWR VPWR _5468_/A sky130_fd_sc_hd__bufbuf_16
X_7169_ _7193_/CLK _7169_/D fanout455/X VGND VGND VPWR VPWR _7169_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_86_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4870_ _4870_/A VGND VGND VPWR VPWR _4903_/A sky130_fd_sc_hd__inv_2
XFILLER_60_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3821_ _6482_/Q _3845_/A _3820_/X VGND VGND VPWR VPWR _3821_/X sky130_fd_sc_hd__a21o_1
XFILLER_177_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6540_ _6725_/CLK _6540_/D fanout440/X VGND VGND VPWR VPWR _6540_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_60_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3752_ _7125_/Q _5567_/A _4097_/A _6576_/Q VGND VGND VPWR VPWR _3752_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6471_ _3957_/A1 _6471_/D _6426_/X VGND VGND VPWR VPWR _6471_/Q sky130_fd_sc_hd__dfrtp_4
X_3683_ _6854_/Q _3315_/Y _5351_/A _6934_/Q VGND VGND VPWR VPWR _3683_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5422_ _5584_/A0 hold482/X _5422_/S VGND VGND VPWR VPWR _5422_/X sky130_fd_sc_hd__mux2_1
Xoutput202 _3206_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[34] sky130_fd_sc_hd__buf_8
X_5353_ _5596_/A0 hold332/X _5359_/S VGND VGND VPWR VPWR _6934_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput213 _3945_/X VGND VGND VPWR VPWR mgmt_gpio_out[0] sky130_fd_sc_hd__buf_8
Xoutput224 _3944_/X VGND VGND VPWR VPWR mgmt_gpio_out[1] sky130_fd_sc_hd__buf_8
Xoutput235 _6683_/Q VGND VGND VPWR VPWR mgmt_gpio_out[2] sky130_fd_sc_hd__buf_8
XFILLER_160_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput246 _6686_/Q VGND VGND VPWR VPWR mgmt_gpio_out[5] sky130_fd_sc_hd__buf_8
Xoutput268 _6802_/Q VGND VGND VPWR VPWR pll_div[2] sky130_fd_sc_hd__buf_8
Xoutput257 _3960_/Y VGND VGND VPWR VPWR pad_flash_io0_oeb sky130_fd_sc_hd__buf_8
X_4304_ _4304_/A _6406_/B VGND VGND VPWR VPWR _4309_/S sky130_fd_sc_hd__and2_4
X_5284_ _5599_/A0 hold855/X _5287_/S VGND VGND VPWR VPWR _5284_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput279 _6493_/Q VGND VGND VPWR VPWR pll_trim[13] sky130_fd_sc_hd__buf_8
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7023_ _7140_/CLK hold34/X fanout430/X VGND VGND VPWR VPWR _7023_/Q sky130_fd_sc_hd__dfrtp_2
X_4235_ hold847/X _4234_/X _4235_/S VGND VGND VPWR VPWR _4235_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4166_ _4166_/A _6406_/B VGND VGND VPWR VPWR _4171_/S sky130_fd_sc_hd__nand2_4
XFILLER_55_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4097_ _4097_/A hold47/X VGND VGND VPWR VPWR _4102_/S sky130_fd_sc_hd__nand2_4
XFILLER_82_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6807_ _6810_/CLK _6807_/D fanout419/X VGND VGND VPWR VPWR _6807_/Q sky130_fd_sc_hd__dfrtp_2
X_4999_ _5121_/C _5118_/C _5078_/C _4985_/Y VGND VGND VPWR VPWR _5001_/C sky130_fd_sc_hd__or4b_1
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6738_ _6810_/CLK _6738_/D fanout419/X VGND VGND VPWR VPWR _6738_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6669_ _6672_/CLK _6669_/D fanout453/X VGND VGND VPWR VPWR _6669_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout440 fanout442/X VGND VGND VPWR VPWR fanout440/X sky130_fd_sc_hd__buf_8
XFILLER_120_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout451 fanout455/X VGND VGND VPWR VPWR fanout451/X sky130_fd_sc_hd__buf_8
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4020_ hold802/X _4019_/X _4024_/S VGND VGND VPWR VPWR _4020_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5971_ _6623_/Q _5673_/X _5681_/X _6598_/Q _5970_/X VGND VGND VPWR VPWR _5976_/B
+ sky130_fd_sc_hd__a221o_2
X_4922_ _4922_/A _5142_/A VGND VGND VPWR VPWR _5034_/A sky130_fd_sc_hd__or2_2
XFILLER_92_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4853_ _4581_/B _4634_/B _4839_/X _4842_/X _5140_/A VGND VGND VPWR VPWR _4853_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_100_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4784_ _4724_/B _4756_/B _4519_/Y VGND VGND VPWR VPWR _4800_/C sky130_fd_sc_hd__o21bai_1
X_3804_ _3797_/X _3803_/X _3801_/B VGND VGND VPWR VPWR _6485_/D sky130_fd_sc_hd__o21ba_1
X_6523_ _6672_/CLK _6523_/D fanout453/X VGND VGND VPWR VPWR _6523_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_opt_2_0_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR clkbuf_opt_2_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
X_3735_ _5225_/A _5225_/B VGND VGND VPWR VPWR _3735_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6454_ _6454_/A _6454_/B VGND VGND VPWR VPWR _6454_/X sky130_fd_sc_hd__and2_1
X_5405_ _5405_/A _5594_/B VGND VGND VPWR VPWR _5413_/S sky130_fd_sc_hd__and2_4
X_3666_ _3665_/X _6791_/Q _3857_/C VGND VGND VPWR VPWR _3666_/X sky130_fd_sc_hd__mux2_1
X_6385_ _6384_/X _7213_/Q _6400_/S VGND VGND VPWR VPWR _7213_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3597_ input29/X _3283_/Y _3320_/Y input6/X _3562_/X VGND VGND VPWR VPWR _3598_/D
+ sky130_fd_sc_hd__a221o_2
X_5336_ _5336_/A0 _5588_/A0 _5341_/S VGND VGND VPWR VPWR _5336_/X sky130_fd_sc_hd__mux2_1
X_5267_ hold649/X _5582_/A0 _5269_/S VGND VGND VPWR VPWR _5267_/X sky130_fd_sc_hd__mux2_1
X_4218_ hold254/X _4217_/X _4218_/S VGND VGND VPWR VPWR _4218_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7006_ _7078_/CLK _7006_/D fanout430/X VGND VGND VPWR VPWR _7006_/Q sky130_fd_sc_hd__dfstp_2
X_5198_ _6410_/A0 _5198_/A1 _5199_/S VGND VGND VPWR VPWR _5198_/X sky130_fd_sc_hd__mux2_1
X_4149_ _4149_/A0 _5289_/A0 _4153_/S VGND VGND VPWR VPWR _4149_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3520_ _4241_/A _5234_/B VGND VGND VPWR VPWR _4280_/A sky130_fd_sc_hd__nor2_8
XFILLER_183_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold707 _5268_/X VGND VGND VPWR VPWR _6859_/D sky130_fd_sc_hd__bufbuf_16
Xhold718 _5435_/X VGND VGND VPWR VPWR _7007_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_143_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3451_ _3451_/A _3451_/B _3451_/C _3451_/D VGND VGND VPWR VPWR _3452_/D sky130_fd_sc_hd__or4_1
Xhold729 _7027_/Q VGND VGND VPWR VPWR hold729/X sky130_fd_sc_hd__bufbuf_16
XFILLER_170_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6170_ _6170_/A _6170_/B _6170_/C _6170_/D VGND VGND VPWR VPWR _6170_/X sky130_fd_sc_hd__or4_1
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3382_ _3381_/X _6797_/Q _3928_/A VGND VGND VPWR VPWR _6797_/D sky130_fd_sc_hd__mux2_1
X_5121_ _5121_/A _5121_/B _5121_/C _5121_/D VGND VGND VPWR VPWR _5135_/D sky130_fd_sc_hd__or4_1
XFILLER_130_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_3_csclk _6722_/CLK VGND VGND VPWR VPWR _6840_/CLK sky130_fd_sc_hd__clkbuf_8
X_5052_ _4660_/X _4724_/B _4819_/B _4724_/A VGND VGND VPWR VPWR _5052_/X sky130_fd_sc_hd__a211o_1
XFILLER_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4003_ hold488/X _5584_/A0 _4003_/S VGND VGND VPWR VPWR _6503_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5954_ _6579_/Q _5689_/X _5941_/X _5944_/X VGND VGND VPWR VPWR _5959_/B sky130_fd_sc_hd__a211o_2
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4905_ _4950_/B _4905_/B _4905_/C _4905_/D VGND VGND VPWR VPWR _4906_/D sky130_fd_sc_hd__or4_4
X_5885_ _6563_/Q _5694_/X _5703_/X _6540_/Q _5884_/X VGND VGND VPWR VPWR _5893_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4836_ _4697_/A _5005_/C _4832_/B VGND VGND VPWR VPWR _4836_/X sky130_fd_sc_hd__a21o_1
XFILLER_166_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6506_ _6987_/CLK _6506_/D fanout450/X VGND VGND VPWR VPWR _6506_/Q sky130_fd_sc_hd__dfrtp_2
X_4767_ _4871_/A _4997_/A _4724_/B _4886_/B VGND VGND VPWR VPWR _4767_/X sky130_fd_sc_hd__o22a_1
X_4698_ _4745_/A _5147_/B VGND VGND VPWR VPWR _4698_/Y sky130_fd_sc_hd__nor2_2
X_3718_ _7102_/Q hold21/A _4328_/A _6774_/Q VGND VGND VPWR VPWR _3718_/X sky130_fd_sc_hd__a22o_1
X_6437_ _6446_/A _6446_/B VGND VGND VPWR VPWR _6437_/X sky130_fd_sc_hd__and2_1
X_3649_ _7047_/Q _5477_/A _5207_/A _6813_/Q _3648_/X VGND VGND VPWR VPWR _3654_/B
+ sky130_fd_sc_hd__a221o_1
X_6368_ _7208_/Q _3452_/X _6370_/S VGND VGND VPWR VPWR _7208_/D sky130_fd_sc_hd__mux2_1
X_5319_ _5571_/A0 hold778/X _5323_/S VGND VGND VPWR VPWR _5319_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold12 hold2/X VGND VGND VPWR VPWR hold12/X sky130_fd_sc_hd__bufbuf_16
X_6299_ _6621_/Q _6022_/C _6032_/X _6651_/Q VGND VGND VPWR VPWR _6299_/X sky130_fd_sc_hd__a22o_1
XFILLER_76_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold23 hold23/A VGND VGND VPWR VPWR hold23/X sky130_fd_sc_hd__bufbuf_16
XFILLER_130_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold56 hold56/A VGND VGND VPWR VPWR hold56/X sky130_fd_sc_hd__bufbuf_16
Xhold34 hold34/A VGND VGND VPWR VPWR hold34/X sky130_fd_sc_hd__bufbuf_16
Xhold45 hold45/A VGND VGND VPWR VPWR hold98/A sky130_fd_sc_hd__bufbuf_16
Xhold78 hold7/X VGND VGND VPWR VPWR hold78/X sky130_fd_sc_hd__bufbuf_16
Xhold67 hold67/A VGND VGND VPWR VPWR hold67/X sky130_fd_sc_hd__bufbuf_16
XFILLER_75_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold89 hold89/A VGND VGND VPWR VPWR hold89/X sky130_fd_sc_hd__bufbuf_16
XFILLER_16_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_9 _4018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5670_ _6997_/Q _5667_/X _5669_/X _7061_/Q VGND VGND VPWR VPWR _5670_/X sky130_fd_sc_hd__a22o_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4621_ _4988_/A _4986_/C _4619_/X _4620_/X VGND VGND VPWR VPWR _4623_/C sky130_fd_sc_hd__o211a_1
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4552_ _4376_/Y _4987_/B _4920_/A _5136_/A _4551_/X VGND VGND VPWR VPWR _4552_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_116_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold515 _6983_/Q VGND VGND VPWR VPWR hold515/X sky130_fd_sc_hd__bufbuf_16
X_4483_ _4533_/A _4484_/C VGND VGND VPWR VPWR _4693_/B sky130_fd_sc_hd__nor2_2
Xhold526 _4037_/X VGND VGND VPWR VPWR _6524_/D sky130_fd_sc_hd__bufbuf_16
Xhold504 _4132_/X VGND VGND VPWR VPWR _6605_/D sky130_fd_sc_hd__bufbuf_16
X_3503_ _7017_/Q _3359_/Y _4166_/A _6638_/Q _3502_/X VGND VGND VPWR VPWR _3504_/D
+ sky130_fd_sc_hd__a221o_1
Xhold537 _6520_/Q VGND VGND VPWR VPWR hold537/X sky130_fd_sc_hd__bufbuf_16
Xhold559 _6918_/Q VGND VGND VPWR VPWR hold559/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3434_ input40/X _4023_/S _5333_/A _6922_/Q _3418_/X VGND VGND VPWR VPWR _3436_/C
+ sky130_fd_sc_hd__a221o_1
X_6222_ _7132_/Q _6023_/A _6033_/X _7012_/Q _6221_/X VGND VGND VPWR VPWR _6232_/B
+ sky130_fd_sc_hd__a221o_1
Xhold548 _6685_/Q VGND VGND VPWR VPWR hold548/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6153_ _6865_/Q _6025_/D _6029_/X _7049_/Q _6152_/X VGND VGND VPWR VPWR _6156_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3365_ hold91/A hold60/X VGND VGND VPWR VPWR hold61/A sky130_fd_sc_hd__nor2_8
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5104_ _4898_/B _5050_/C _4754_/B VGND VGND VPWR VPWR _5104_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3296_ _7052_/Q _5477_/A hold28/A _6868_/Q _3287_/X VGND VGND VPWR VPWR _3296_/X
+ sky130_fd_sc_hd__a221o_1
Xhold1204 _3980_/X VGND VGND VPWR VPWR _6488_/D sky130_fd_sc_hd__bufbuf_16
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1215 _6768_/Q VGND VGND VPWR VPWR _4323_/A1 sky130_fd_sc_hd__bufbuf_16
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ _6854_/Q _6060_/B _6071_/X _6083_/X _3197_/Y VGND VGND VPWR VPWR _6084_/X
+ sky130_fd_sc_hd__o221a_2
X_5035_ _5035_/A _5035_/B _5035_/C _5035_/D VGND VGND VPWR VPWR _5166_/C sky130_fd_sc_hd__or4_1
Xhold1237 _6522_/Q VGND VGND VPWR VPWR _4035_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1248 _6566_/Q VGND VGND VPWR VPWR _4086_/A0 sky130_fd_sc_hd__bufbuf_16
XFILLER_85_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1226 _6681_/Q VGND VGND VPWR VPWR _4221_/A0 sky130_fd_sc_hd__bufbuf_16
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1259 _7147_/Q VGND VGND VPWR VPWR _5592_/A1 sky130_fd_sc_hd__bufbuf_16
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6986_ _7130_/CLK _6986_/D fanout452/X VGND VGND VPWR VPWR _6986_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_81_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5937_ _5937_/A _5937_/B _5937_/C _5937_/D VGND VGND VPWR VPWR _5937_/X sky130_fd_sc_hd__or4_1
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5868_ _7084_/Q _5693_/X _5694_/X _6900_/Q _5867_/X VGND VGND VPWR VPWR _5871_/C
+ sky130_fd_sc_hd__a221o_1
X_4819_ _4819_/A _4819_/B _5005_/A _4819_/D VGND VGND VPWR VPWR _4820_/B sky130_fd_sc_hd__or4_1
X_5799_ _6985_/Q _5963_/B VGND VGND VPWR VPWR _5799_/X sky130_fd_sc_hd__or2_1
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput102 wb_adr_i[12] VGND VGND VPWR VPWR _4350_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_163_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput124 wb_adr_i[3] VGND VGND VPWR VPWR _4469_/A sky130_fd_sc_hd__buf_8
XFILLER_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput135 wb_dat_i[12] VGND VGND VPWR VPWR _6390_/B1 sky130_fd_sc_hd__clkbuf_4
Xinput113 wb_adr_i[22] VGND VGND VPWR VPWR _4345_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_103_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput146 wb_dat_i[22] VGND VGND VPWR VPWR _6395_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput168 wb_sel_i[3] VGND VGND VPWR VPWR _6402_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput157 wb_dat_i[3] VGND VGND VPWR VPWR _6387_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6840_ _6840_/CLK _6840_/D _6454_/A VGND VGND VPWR VPWR _6840_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6771_ _7222_/CLK _6771_/D fanout422/X VGND VGND VPWR VPWR _6771_/Q sky130_fd_sc_hd__dfrtp_2
X_3983_ hold39/X _7213_/Q _6689_/Q VGND VGND VPWR VPWR hold40/A sky130_fd_sc_hd__mux2_4
X_5722_ _6853_/Q _5722_/B VGND VGND VPWR VPWR _5722_/X sky130_fd_sc_hd__or2_1
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_21_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _6951_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_31_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5653_ _6037_/B _6035_/A _6037_/C VGND VGND VPWR VPWR _5653_/X sky130_fd_sc_hd__and3_4
XFILLER_191_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4604_ _4694_/A _4898_/B VGND VGND VPWR VPWR _4887_/B sky130_fd_sc_hd__nor2_1
X_5584_ _5584_/A0 hold427/X hold62/X VGND VGND VPWR VPWR _5584_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4535_ _4533_/A _4533_/B _4537_/C _4956_/B VGND VGND VPWR VPWR _4536_/B sky130_fd_sc_hd__and4bb_4
Xhold301 _6929_/Q VGND VGND VPWR VPWR hold301/X sky130_fd_sc_hd__bufbuf_16
Xclkbuf_leaf_36_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _6672_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_144_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold334 _5389_/X VGND VGND VPWR VPWR _6966_/D sky130_fd_sc_hd__bufbuf_16
Xhold312 _6627_/Q VGND VGND VPWR VPWR hold312/X sky130_fd_sc_hd__bufbuf_16
Xhold323 _6546_/Q VGND VGND VPWR VPWR hold323/X sky130_fd_sc_hd__bufbuf_16
X_4466_ _4722_/A _4467_/B VGND VGND VPWR VPWR _5004_/A sky130_fd_sc_hd__and2_4
Xhold356 _4042_/X VGND VGND VPWR VPWR _6529_/D sky130_fd_sc_hd__bufbuf_16
Xhold378 _5296_/X VGND VGND VPWR VPWR _6884_/D sky130_fd_sc_hd__bufbuf_16
Xhold367 _5305_/X VGND VGND VPWR VPWR _6892_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_117_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold345 _4084_/X VGND VGND VPWR VPWR _6564_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_171_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold389 _5573_/X VGND VGND VPWR VPWR _7130_/D sky130_fd_sc_hd__bufbuf_16
X_4397_ _4775_/A _4671_/A VGND VGND VPWR VPWR _4930_/D sky130_fd_sc_hd__nand2_4
X_6205_ _6979_/Q _6023_/B _6021_/C _6883_/Q _6204_/X VGND VGND VPWR VPWR _6206_/D
+ sky130_fd_sc_hd__a221o_1
X_7185_ _7201_/CLK _7185_/D _6446_/A VGND VGND VPWR VPWR _7185_/Q sky130_fd_sc_hd__dfrtp_4
X_3417_ _3416_/X _6796_/Q _3928_/A VGND VGND VPWR VPWR _6796_/D sky130_fd_sc_hd__mux2_1
X_3348_ _7148_/Q _5585_/A _5297_/A _6892_/Q VGND VGND VPWR VPWR _3348_/X sky130_fd_sc_hd__a22o_1
X_6136_ _7081_/Q _6311_/B VGND VGND VPWR VPWR _6136_/X sky130_fd_sc_hd__and2_1
XFILLER_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1012 _6766_/Q VGND VGND VPWR VPWR _4320_/A0 sky130_fd_sc_hd__bufbuf_16
Xhold1001 _4332_/X VGND VGND VPWR VPWR _6776_/D sky130_fd_sc_hd__bufbuf_16
Xhold1023 _4321_/X VGND VGND VPWR VPWR _6767_/D sky130_fd_sc_hd__bufbuf_16
Xhold1067 _6836_/Q VGND VGND VPWR VPWR _5241_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_100_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1056 _6539_/Q VGND VGND VPWR VPWR _4054_/A0 sky130_fd_sc_hd__bufbuf_16
X_3279_ _3309_/A _3314_/B VGND VGND VPWR VPWR _3476_/A sky130_fd_sc_hd__or2_4
Xhold1045 _6760_/Q VGND VGND VPWR VPWR _4313_/A0 sky130_fd_sc_hd__bufbuf_16
Xhold1034 _4200_/X VGND VGND VPWR VPWR _6662_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_39_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6067_ _7118_/Q _6023_/D _6030_/Y _7030_/Q VGND VGND VPWR VPWR _6067_/X sky130_fd_sc_hd__a22o_1
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5018_ _5037_/A _5037_/B _5018_/C VGND VGND VPWR VPWR _5018_/X sky130_fd_sc_hd__or3_1
XANTENNA_207 _7060_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1078 _7037_/Q VGND VGND VPWR VPWR _5469_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1089 _4308_/X VGND VGND VPWR VPWR _6756_/D sky130_fd_sc_hd__bufbuf_16
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_218 _6914_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_229 _6476_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6969_ _7111_/CLK _6969_/D fanout444/X VGND VGND VPWR VPWR _6969_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_139_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold890 _4022_/X VGND VGND VPWR VPWR _6512_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4320_ _4320_/A0 _6410_/A0 _4321_/S VGND VGND VPWR VPWR _4320_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4251_ _6407_/A0 _4251_/A1 _4255_/S VGND VGND VPWR VPWR _4251_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3202_ _3202_/A VGND VGND VPWR VPWR _3202_/Y sky130_fd_sc_hd__clkinv_2
X_4182_ hold861/X _4326_/A0 _4183_/S VGND VGND VPWR VPWR _4182_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6823_ _7035_/CLK _6823_/D fanout433/X VGND VGND VPWR VPWR _6823_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3966_ _6705_/Q _3974_/B VGND VGND VPWR VPWR _6702_/D sky130_fd_sc_hd__and2_1
X_6754_ _7222_/CLK _6754_/D fanout422/X VGND VGND VPWR VPWR _6754_/Q sky130_fd_sc_hd__dfrtp_2
X_5705_ _5864_/B _5705_/B _5706_/B VGND VGND VPWR VPWR _5705_/X sky130_fd_sc_hd__and3_4
X_6685_ _7138_/CLK _6685_/D fanout438/X VGND VGND VPWR VPWR _6685_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_10_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5636_ _5635_/Y _5963_/B _5636_/S VGND VGND VPWR VPWR _7165_/D sky130_fd_sc_hd__mux2_1
X_3897_ _6703_/Q _3883_/X _3915_/B _6698_/Q VGND VGND VPWR VPWR _6703_/D sky130_fd_sc_hd__a22o_1
XFILLER_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5567_ _5567_/A hold47/X VGND VGND VPWR VPWR _5575_/S sky130_fd_sc_hd__nand2_8
X_5498_ _5597_/A0 hold431/X _5503_/S VGND VGND VPWR VPWR _5498_/X sky130_fd_sc_hd__mux2_1
Xhold153 _5589_/X VGND VGND VPWR VPWR _7144_/D sky130_fd_sc_hd__bufbuf_16
Xhold131 hold131/A VGND VGND VPWR VPWR _6528_/D sky130_fd_sc_hd__bufbuf_16
Xhold142 _7122_/Q VGND VGND VPWR VPWR hold142/X sky130_fd_sc_hd__bufbuf_16
X_4518_ _4871_/A _4990_/A VGND VGND VPWR VPWR _5081_/A sky130_fd_sc_hd__nor2_2
Xhold120 _5546_/X VGND VGND VPWR VPWR _7106_/D sky130_fd_sc_hd__bufbuf_16
Xhold164 _5499_/X VGND VGND VPWR VPWR _7064_/D sky130_fd_sc_hd__bufbuf_16
X_4449_ _4534_/B _4449_/B VGND VGND VPWR VPWR _4572_/B sky130_fd_sc_hd__nand2_2
XFILLER_132_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold186 _5473_/X VGND VGND VPWR VPWR _7041_/D sky130_fd_sc_hd__bufbuf_16
Xhold175 hold59/X VGND VGND VPWR VPWR _3309_/A sky130_fd_sc_hd__bufbuf_16
XFILLER_144_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold197 _5472_/X VGND VGND VPWR VPWR _7040_/D sky130_fd_sc_hd__bufbuf_16
X_7168_ _7193_/CLK _7168_/D fanout455/X VGND VGND VPWR VPWR _7168_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6119_ _7072_/Q _6009_/X _6020_/D _6968_/Q VGND VGND VPWR VPWR _6119_/X sky130_fd_sc_hd__a22o_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7099_ _7139_/CLK _7099_/D fanout435/X VGND VGND VPWR VPWR _7099_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3820_ _3845_/A _3820_/B _3820_/C VGND VGND VPWR VPWR _3820_/X sky130_fd_sc_hd__and3b_1
X_3751_ _6949_/Q _5369_/A _4067_/A _6550_/Q _3750_/X VGND VGND VPWR VPWR _3754_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6470_ _6668_/CLK _6470_/D _6425_/X VGND VGND VPWR VPWR _6470_/Q sky130_fd_sc_hd__dfrtp_2
X_3682_ input15/X _3283_/Y _4280_/A _6734_/Q _3681_/X VGND VGND VPWR VPWR _3687_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5421_ _5583_/A0 hold774/X _5422_/S VGND VGND VPWR VPWR _5421_/X sky130_fd_sc_hd__mux2_1
Xoutput225 _6673_/Q VGND VGND VPWR VPWR mgmt_gpio_out[20] sky130_fd_sc_hd__buf_8
Xoutput203 _3933_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[35] sky130_fd_sc_hd__buf_8
XFILLER_161_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5352_ _5595_/A0 _5352_/A1 _5359_/S VGND VGND VPWR VPWR _6933_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput214 _3937_/X VGND VGND VPWR VPWR mgmt_gpio_out[10] sky130_fd_sc_hd__buf_8
Xoutput236 _6520_/Q VGND VGND VPWR VPWR mgmt_gpio_out[30] sky130_fd_sc_hd__buf_8
XFILLER_126_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput247 _3940_/X VGND VGND VPWR VPWR mgmt_gpio_out[6] sky130_fd_sc_hd__buf_8
Xoutput258 _7227_/X VGND VGND VPWR VPWR pad_flash_io1_do sky130_fd_sc_hd__buf_8
X_4303_ _6411_/A0 hold748/X _4303_/S VGND VGND VPWR VPWR _4303_/X sky130_fd_sc_hd__mux2_1
X_5283_ hold71/X hold340/X _5287_/S VGND VGND VPWR VPWR _6872_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput269 _6803_/Q VGND VGND VPWR VPWR pll_div[3] sky130_fd_sc_hd__buf_8
X_7022_ _7078_/CLK _7022_/D fanout430/X VGND VGND VPWR VPWR _7022_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_141_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4234_ hold429/X _5584_/A0 _4234_/S VGND VGND VPWR VPWR _4234_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4165_ _5545_/A0 _4165_/A1 _4165_/S VGND VGND VPWR VPWR _6633_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_634 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4096_ _6575_/Q _3379_/X _4096_/S VGND VGND VPWR VPWR _6575_/D sky130_fd_sc_hd__mux2_1
XFILLER_70_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6806_ _6810_/CLK _6806_/D _6439_/A VGND VGND VPWR VPWR _6806_/Q sky130_fd_sc_hd__dfstp_4
X_4998_ _5114_/C _5116_/C VGND VGND VPWR VPWR _5001_/B sky130_fd_sc_hd__or2_2
XFILLER_23_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3949_ _6512_/Q _3949_/A1 _6834_/Q VGND VGND VPWR VPWR _3949_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6737_ _6744_/CLK _6737_/D fanout427/X VGND VGND VPWR VPWR _6737_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6668_ _6668_/CLK _6668_/D _6447_/X VGND VGND VPWR VPWR _6668_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6599_ _6951_/CLK _6599_/D fanout440/X VGND VGND VPWR VPWR _6599_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_109_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5619_ _7160_/Q _5616_/A _5618_/Y VGND VGND VPWR VPWR _7160_/D sky130_fd_sc_hd__o21a_1
XFILLER_164_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout441 fanout442/X VGND VGND VPWR VPWR _6421_/A sky130_fd_sc_hd__buf_8
Xfanout430 fanout431/X VGND VGND VPWR VPWR fanout430/X sky130_fd_sc_hd__buf_8
Xfanout452 fanout454/X VGND VGND VPWR VPWR fanout452/X sky130_fd_sc_hd__buf_8
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5970_ _6712_/Q _5691_/X _5701_/X _6618_/Q VGND VGND VPWR VPWR _5970_/X sky130_fd_sc_hd__a22o_1
XFILLER_18_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4921_ _4930_/D _4575_/B _4933_/B _4684_/Y VGND VGND VPWR VPWR _4941_/B sky130_fd_sc_hd__a22o_1
XFILLER_33_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4852_ _4986_/C _4989_/B VGND VGND VPWR VPWR _5118_/B sky130_fd_sc_hd__nor2_1
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_390 _5694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3803_ _6485_/Q _6664_/Q VGND VGND VPWR VPWR _3803_/X sky130_fd_sc_hd__or2_1
X_4783_ _4920_/B _5047_/A VGND VGND VPWR VPWR _4802_/B sky130_fd_sc_hd__or2_1
X_6522_ _6987_/CLK _6522_/D fanout450/X VGND VGND VPWR VPWR _6522_/Q sky130_fd_sc_hd__dfrtp_1
X_3734_ input71/X _4023_/S _4234_/S _3971_/A VGND VGND VPWR VPWR _3734_/X sky130_fd_sc_hd__a22o_4
XFILLER_146_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6453_ _6454_/A _6454_/B VGND VGND VPWR VPWR _6453_/X sky130_fd_sc_hd__and2_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3665_ _3665_/A _3665_/B _3665_/C VGND VGND VPWR VPWR _3665_/X sky130_fd_sc_hd__or3_4
XFILLER_161_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5404_ hold493/X _5602_/A0 _5404_/S VGND VGND VPWR VPWR _5404_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6384_ _6707_/Q _6384_/A2 _6384_/B1 _6706_/Q _6383_/X VGND VGND VPWR VPWR _6384_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3596_ _6814_/Q _5207_/A _3344_/Y _6499_/Q _3564_/X VGND VGND VPWR VPWR _3598_/C
+ sky130_fd_sc_hd__a221o_1
X_5335_ hold559/X _5587_/A0 _5341_/S VGND VGND VPWR VPWR _6918_/D sky130_fd_sc_hd__mux2_1
XFILLER_125_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5266_ hold277/X hold185/A _5269_/S VGND VGND VPWR VPWR _5266_/X sky130_fd_sc_hd__mux2_1
X_4217_ _4249_/A1 hold14/X _4217_/S VGND VGND VPWR VPWR _4217_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7005_ _7140_/CLK _7005_/D fanout430/X VGND VGND VPWR VPWR _7005_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_28_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5197_ _6409_/A0 _5197_/A1 _5199_/S VGND VGND VPWR VPWR _6802_/D sky130_fd_sc_hd__mux2_1
X_4148_ _4148_/A _5558_/B VGND VGND VPWR VPWR _4153_/S sky130_fd_sc_hd__and2_4
XFILLER_83_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4079_ _6560_/Q _3452_/X _4081_/S VGND VGND VPWR VPWR _6560_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold719 _6507_/Q VGND VGND VPWR VPWR hold719/X sky130_fd_sc_hd__bufbuf_16
XFILLER_128_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold708 _7099_/Q VGND VGND VPWR VPWR hold708/X sky130_fd_sc_hd__bufbuf_16
XFILLER_171_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3450_ _3450_/A _3450_/B _3450_/C _3450_/D VGND VGND VPWR VPWR _3451_/D sky130_fd_sc_hd__or4_2
XFILLER_130_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3381_ _3379_/X _6796_/Q _3857_/C VGND VGND VPWR VPWR _3381_/X sky130_fd_sc_hd__mux2_1
X_5120_ _5135_/A _5137_/B _5120_/C _5135_/C VGND VGND VPWR VPWR _5120_/X sky130_fd_sc_hd__or4_2
XFILLER_69_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5051_ _4758_/B _5049_/X _5050_/X VGND VGND VPWR VPWR _5056_/B sky130_fd_sc_hd__a21bo_1
XFILLER_85_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4002_ _6502_/Q hold209/X _4003_/S VGND VGND VPWR VPWR _4002_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5953_ _5953_/A _5953_/B _5953_/C _5953_/D VGND VGND VPWR VPWR _5953_/X sky130_fd_sc_hd__or4_2
XFILLER_18_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4904_ _4950_/A _5129_/A _4904_/C _4904_/D VGND VGND VPWR VPWR _4905_/D sky130_fd_sc_hd__or4_1
X_5884_ _6589_/Q _5680_/X _5685_/X _6644_/Q VGND VGND VPWR VPWR _5884_/X sky130_fd_sc_hd__a22o_1
XFILLER_33_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4835_ _4898_/B _4832_/A _4832_/B _5164_/B VGND VGND VPWR VPWR _4835_/X sky130_fd_sc_hd__o22a_1
X_4766_ _4766_/A _5151_/A VGND VGND VPWR VPWR _4802_/A sky130_fd_sc_hd__or2_4
XFILLER_119_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6505_ _6825_/CLK _6505_/D fanout429/X VGND VGND VPWR VPWR _6505_/Q sky130_fd_sc_hd__dfstp_4
X_3717_ _3717_/A _3717_/B _3717_/C _3717_/D VGND VGND VPWR VPWR _3726_/C sky130_fd_sc_hd__or4_1
X_4697_ _4697_/A _5062_/C VGND VGND VPWR VPWR _4697_/Y sky130_fd_sc_hd__nor2_1
XFILLER_162_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6436_ _6439_/A _6446_/B VGND VGND VPWR VPWR _6436_/X sky130_fd_sc_hd__and2_1
XFILLER_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3648_ _7039_/Q _3334_/Y _4196_/A _6661_/Q VGND VGND VPWR VPWR _3648_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3579_ _6617_/Q _3511_/Y _4250_/A _6711_/Q VGND VGND VPWR VPWR _3579_/X sky130_fd_sc_hd__a22o_2
X_6367_ _7207_/Q _6367_/A1 _6370_/S VGND VGND VPWR VPWR _7207_/D sky130_fd_sc_hd__mux2_1
X_5318_ _5588_/A0 _5318_/A1 _5323_/S VGND VGND VPWR VPWR _5318_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold13 hold13/A VGND VGND VPWR VPWR hold3/A sky130_fd_sc_hd__bufbuf_16
XFILLER_130_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6298_ _6578_/Q _6021_/A _6025_/A _6606_/Q _6286_/X VGND VGND VPWR VPWR _6305_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_102_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold35 hold64/X VGND VGND VPWR VPWR hold65/A sky130_fd_sc_hd__bufbuf_16
XFILLER_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold46 hold99/X VGND VGND VPWR VPWR hold46/X sky130_fd_sc_hd__bufbuf_16
Xhold24 hold24/A VGND VGND VPWR VPWR hold24/X sky130_fd_sc_hd__bufbuf_16
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5249_ _6410_/A0 _5249_/A1 _5251_/S VGND VGND VPWR VPWR _5249_/X sky130_fd_sc_hd__mux2_1
Xhold79 hold79/A VGND VGND VPWR VPWR hold79/X sky130_fd_sc_hd__bufbuf_16
XFILLER_152_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold68 hold68/A VGND VGND VPWR VPWR hold68/X sky130_fd_sc_hd__bufbuf_16
Xhold57 hold57/A VGND VGND VPWR VPWR hold57/X sky130_fd_sc_hd__bufbuf_16
XFILLER_29_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4620_ _4986_/A _4617_/A _4749_/C _4988_/A _4893_/A VGND VGND VPWR VPWR _4620_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_175_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4551_ _5079_/A _5078_/A _4551_/C VGND VGND VPWR VPWR _4551_/X sky130_fd_sc_hd__or3_1
Xhold516 _5408_/X VGND VGND VPWR VPWR _6983_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_171_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4482_ _4694_/A _4986_/C VGND VGND VPWR VPWR _4980_/A sky130_fd_sc_hd__nor2_2
XFILLER_143_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold527 _6714_/Q VGND VGND VPWR VPWR hold527/X sky130_fd_sc_hd__bufbuf_16
Xhold505 _7052_/Q VGND VGND VPWR VPWR hold505/X sky130_fd_sc_hd__bufbuf_16
X_3502_ _7073_/Q hold92/A _4178_/A _6648_/Q VGND VGND VPWR VPWR _3502_/X sky130_fd_sc_hd__a22o_2
XFILLER_7_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold538 _4032_/X VGND VGND VPWR VPWR _6520_/D sky130_fd_sc_hd__bufbuf_16
X_6221_ _6892_/Q _6020_/A _6021_/D _7148_/Q _6220_/X VGND VGND VPWR VPWR _6221_/X
+ sky130_fd_sc_hd__a221o_4
X_3433_ _7090_/Q hold54/A _5450_/A _7026_/Q _3425_/X VGND VGND VPWR VPWR _3436_/B
+ sky130_fd_sc_hd__a221o_2
Xhold549 _4229_/X VGND VGND VPWR VPWR _6685_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_131_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6152_ _7105_/Q _5653_/X _6022_/B _6945_/Q VGND VGND VPWR VPWR _6152_/X sky130_fd_sc_hd__a22o_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _5095_/X _5101_/X _5161_/C _4928_/Y VGND VGND VPWR VPWR _5103_/X sky130_fd_sc_hd__o211a_1
XFILLER_106_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _3501_/A _3375_/B VGND VGND VPWR VPWR _5513_/A sky130_fd_sc_hd__nor2_8
Xhold1205 _6594_/Q VGND VGND VPWR VPWR _4119_/A0 sky130_fd_sc_hd__bufbuf_16
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1216 _4323_/X VGND VGND VPWR VPWR _6768_/D sky130_fd_sc_hd__bufbuf_16
X_3295_ hold27/X _3473_/A VGND VGND VPWR VPWR hold28/A sky130_fd_sc_hd__nor2_8
X_6083_ _6232_/A _6083_/B _6083_/C VGND VGND VPWR VPWR _6083_/X sky130_fd_sc_hd__or3_1
X_5034_ _5034_/A _5034_/B _5095_/C _5102_/B VGND VGND VPWR VPWR _5036_/C sky130_fd_sc_hd__or4b_1
Xhold1249 _6623_/Q VGND VGND VPWR VPWR _4153_/A0 sky130_fd_sc_hd__bufbuf_16
XFILLER_85_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1227 _4221_/X VGND VGND VPWR VPWR _6681_/D sky130_fd_sc_hd__bufbuf_16
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1238 _6848_/Q VGND VGND VPWR VPWR _5256_/A1 sky130_fd_sc_hd__bufbuf_16
X_6985_ _7111_/CLK _6985_/D fanout446/X VGND VGND VPWR VPWR _6985_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_25_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5936_ _6730_/Q _5667_/X _5692_/X _7223_/Q _5935_/X VGND VGND VPWR VPWR _5937_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5867_ _6884_/Q _5674_/X _5687_/X _7052_/Q VGND VGND VPWR VPWR _5867_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4818_ _4818_/A _4818_/B _4818_/C VGND VGND VPWR VPWR _5003_/C sky130_fd_sc_hd__or3_4
X_5798_ _7097_/Q _5690_/X _5692_/X _7073_/Q _5797_/X VGND VGND VPWR VPWR _5806_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4749_ _4812_/A _4819_/B _4749_/C VGND VGND VPWR VPWR _4935_/D sky130_fd_sc_hd__or3_4
XFILLER_147_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6419_ _6421_/A _6421_/B VGND VGND VPWR VPWR _6419_/X sky130_fd_sc_hd__and2_1
XFILLER_134_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput125 wb_adr_i[4] VGND VGND VPWR VPWR _5050_/A sky130_fd_sc_hd__buf_8
Xinput114 wb_adr_i[23] VGND VGND VPWR VPWR _4345_/A sky130_fd_sc_hd__clkbuf_4
Xinput103 wb_adr_i[13] VGND VGND VPWR VPWR _4350_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_163_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput136 wb_dat_i[13] VGND VGND VPWR VPWR _6392_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_102_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput147 wb_dat_i[23] VGND VGND VPWR VPWR _6399_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput158 wb_dat_i[4] VGND VGND VPWR VPWR _6389_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_103_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput169 wb_stb_i VGND VGND VPWR VPWR input169/X sky130_fd_sc_hd__buf_6
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_2_csclk _6722_/CLK VGND VGND VPWR VPWR _6777_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_40_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3982_ hold920/X _5254_/A0 _3994_/S VGND VGND VPWR VPWR _6489_/D sky130_fd_sc_hd__mux2_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6770_ _6770_/CLK _6770_/D fanout423/X VGND VGND VPWR VPWR _6770_/Q sky130_fd_sc_hd__dfstp_4
X_5721_ _7069_/Q _5692_/X _5709_/X _5713_/X _5720_/X VGND VGND VPWR VPWR _5721_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_188_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5652_ _7171_/Q _7170_/Q VGND VGND VPWR VPWR _6036_/A sky130_fd_sc_hd__nand2b_4
XFILLER_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4603_ _4871_/A _4603_/B VGND VGND VPWR VPWR _4922_/A sky130_fd_sc_hd__nor2_4
XFILLER_129_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5583_ _5583_/A0 hold723/X hold62/X VGND VGND VPWR VPWR _5583_/X sky130_fd_sc_hd__mux2_1
X_4534_ _4655_/A _4534_/B VGND VGND VPWR VPWR _4956_/B sky130_fd_sc_hd__nor2_2
Xhold302 _5347_/X VGND VGND VPWR VPWR _6929_/D sky130_fd_sc_hd__bufbuf_16
Xhold335 _6932_/Q VGND VGND VPWR VPWR hold335/X sky130_fd_sc_hd__bufbuf_16
Xhold313 _4158_/X VGND VGND VPWR VPWR _6627_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_117_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold324 _4063_/X VGND VGND VPWR VPWR _6546_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4465_ _4685_/A _4651_/B VGND VGND VPWR VPWR _4812_/A sky130_fd_sc_hd__or2_4
Xhold368 _6972_/Q VGND VGND VPWR VPWR hold368/X sky130_fd_sc_hd__bufbuf_16
XFILLER_144_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold346 _7038_/Q VGND VGND VPWR VPWR hold346/X sky130_fd_sc_hd__bufbuf_16
Xhold357 _6778_/Q VGND VGND VPWR VPWR hold357/X sky130_fd_sc_hd__bufbuf_16
X_4396_ _4672_/A _4413_/C VGND VGND VPWR VPWR _4671_/A sky130_fd_sc_hd__nand2_8
XFILLER_131_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6204_ _7067_/Q _5996_/X _6020_/C _6915_/Q VGND VGND VPWR VPWR _6204_/X sky130_fd_sc_hd__a22o_1
Xhold379 _6942_/Q VGND VGND VPWR VPWR hold379/X sky130_fd_sc_hd__bufbuf_16
X_7184_ _7197_/CLK _7184_/D fanout420/X VGND VGND VPWR VPWR _7184_/Q sky130_fd_sc_hd__dfrtp_4
X_3416_ _3415_/X _6795_/Q _3857_/C VGND VGND VPWR VPWR _3416_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3347_ _3543_/A _3375_/B VGND VGND VPWR VPWR _5297_/A sky130_fd_sc_hd__nor2_8
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6135_ _7192_/Q _6309_/S _6134_/X VGND VGND VPWR VPWR _7192_/D sky130_fd_sc_hd__o21a_1
Xhold1024 _6949_/Q VGND VGND VPWR VPWR _5370_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_133_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1002 _6656_/Q VGND VGND VPWR VPWR _4193_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1013 _4320_/X VGND VGND VPWR VPWR _6766_/D sky130_fd_sc_hd__bufbuf_16
X_6066_ _7014_/Q _6036_/Y _6335_/B _7038_/Q _6063_/X VGND VGND VPWR VPWR _6071_/B
+ sky130_fd_sc_hd__a221o_1
X_5017_ _5017_/A _5050_/C VGND VGND VPWR VPWR _5047_/D sky130_fd_sc_hd__nor2_1
XFILLER_100_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1046 _6712_/Q VGND VGND VPWR VPWR _4255_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1035 _6730_/Q VGND VGND VPWR VPWR _4277_/A1 sky130_fd_sc_hd__bufbuf_16
X_3278_ _3293_/B _3278_/B VGND VGND VPWR VPWR _3278_/X sky130_fd_sc_hd__or2_1
Xhold1057 _6534_/Q VGND VGND VPWR VPWR _4048_/A0 sky130_fd_sc_hd__bufbuf_16
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1068 _5241_/X VGND VGND VPWR VPWR _6836_/D sky130_fd_sc_hd__bufbuf_16
Xhold1079 _7085_/Q VGND VGND VPWR VPWR _5523_/A1 sky130_fd_sc_hd__bufbuf_16
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_208 _7062_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_219 _6917_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6968_ _7154_/CLK _6968_/D fanout451/X VGND VGND VPWR VPWR _6968_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_158_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6899_ _6939_/CLK _6899_/D fanout453/X VGND VGND VPWR VPWR _6899_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_167_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5919_ _6552_/Q _5702_/X _5705_/X _6611_/Q VGND VGND VPWR VPWR _5919_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold880 _6843_/Q VGND VGND VPWR VPWR hold880/X sky130_fd_sc_hd__bufbuf_16
XFILLER_150_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold891 _6536_/Q VGND VGND VPWR VPWR hold891/X sky130_fd_sc_hd__bufbuf_16
XFILLER_150_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4250_ _4250_/A _5558_/B VGND VGND VPWR VPWR _4255_/S sky130_fd_sc_hd__nand2_4
X_4181_ _4181_/A0 _6409_/A0 _4183_/S VGND VGND VPWR VPWR _6646_/D sky130_fd_sc_hd__mux2_1
X_3201_ _6668_/Q VGND VGND VPWR VPWR _3201_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6822_ _7035_/CLK _6822_/D fanout433/X VGND VGND VPWR VPWR _6822_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_51_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6753_ _6770_/CLK _6753_/D fanout422/X VGND VGND VPWR VPWR _6753_/Q sky130_fd_sc_hd__dfrtp_2
X_3965_ _6473_/Q _3965_/B VGND VGND VPWR VPWR _3965_/X sky130_fd_sc_hd__and2b_4
X_5704_ _5864_/B _5704_/B _5706_/B VGND VGND VPWR VPWR _5704_/X sky130_fd_sc_hd__and3_4
X_3896_ _6698_/Q _3915_/B VGND VGND VPWR VPWR _3896_/Y sky130_fd_sc_hd__nand2_1
X_6684_ _7107_/CLK _6684_/D fanout434/X VGND VGND VPWR VPWR _6684_/Q sky130_fd_sc_hd__dfrtp_2
X_5635_ _5864_/B _5635_/B VGND VGND VPWR VPWR _5635_/Y sky130_fd_sc_hd__nand2_1
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5566_ _5584_/A0 hold480/X _5566_/S VGND VGND VPWR VPWR _5566_/X sky130_fd_sc_hd__mux2_1
Xhold110 _6480_/Q VGND VGND VPWR VPWR hold57/A sky130_fd_sc_hd__bufbuf_16
X_5497_ _5596_/A0 _7062_/Q _5503_/S VGND VGND VPWR VPWR _5497_/X sky130_fd_sc_hd__mux2_1
Xhold132 _6462_/Q VGND VGND VPWR VPWR hold69/A sky130_fd_sc_hd__bufbuf_16
XFILLER_163_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4517_ _4711_/A _4586_/B VGND VGND VPWR VPWR _4850_/A sky130_fd_sc_hd__and2_1
Xhold143 _5564_/X VGND VGND VPWR VPWR _7122_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_105_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold121 _6780_/Q VGND VGND VPWR VPWR hold121/X sky130_fd_sc_hd__bufbuf_16
Xhold165 _6517_/Q VGND VGND VPWR VPWR hold165/X sky130_fd_sc_hd__bufbuf_16
X_4448_ _4707_/B _4445_/X _4440_/B VGND VGND VPWR VPWR _4449_/B sky130_fd_sc_hd__o21ai_2
XFILLER_171_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold154 _7220_/Q VGND VGND VPWR VPWR hold154/X sky130_fd_sc_hd__bufbuf_16
Xhold176 _3309_/X VGND VGND VPWR VPWR hold60/A sky130_fd_sc_hd__bufbuf_16
Xhold187 _6978_/Q VGND VGND VPWR VPWR hold187/X sky130_fd_sc_hd__bufbuf_16
XFILLER_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold198 _6856_/Q VGND VGND VPWR VPWR hold198/X sky130_fd_sc_hd__bufbuf_16
XFILLER_144_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4379_ _4469_/A _5031_/A VGND VGND VPWR VPWR _4986_/B sky130_fd_sc_hd__or2_4
X_7167_ _3949_/A1 _7167_/D fanout455/X VGND VGND VPWR VPWR _7167_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6118_ _7120_/Q _6023_/D _6030_/Y _7032_/Q _6117_/X VGND VGND VPWR VPWR _6121_/C
+ sky130_fd_sc_hd__a221o_4
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7098_ _7139_/CLK _7098_/D fanout435/X VGND VGND VPWR VPWR _7098_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6049_ _7061_/Q _5996_/X _6029_/X _7045_/Q VGND VGND VPWR VPWR _6049_/X sky130_fd_sc_hd__a22o_2
XFILLER_85_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_20_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _6959_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_49_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_35_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _6939_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3750_ _6619_/Q _4148_/A _4250_/A _6708_/Q VGND VGND VPWR VPWR _3750_/X sky130_fd_sc_hd__a22o_1
XFILLER_60_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3681_ _7038_/Q _3334_/Y _5238_/A _6835_/Q VGND VGND VPWR VPWR _3681_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5420_ hold78/X _5420_/A1 _5422_/S VGND VGND VPWR VPWR _5420_/X sky130_fd_sc_hd__mux2_1
Xoutput226 _6674_/Q VGND VGND VPWR VPWR mgmt_gpio_out[21] sky130_fd_sc_hd__buf_8
Xoutput204 _3932_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[36] sky130_fd_sc_hd__buf_8
XFILLER_160_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5351_ _5351_/A _5594_/B VGND VGND VPWR VPWR _5359_/S sky130_fd_sc_hd__nand2_8
Xoutput215 _6509_/Q VGND VGND VPWR VPWR mgmt_gpio_out[11] sky130_fd_sc_hd__buf_8
Xoutput237 _6521_/Q VGND VGND VPWR VPWR mgmt_gpio_out[31] sky130_fd_sc_hd__buf_8
X_5282_ _5588_/A0 _5282_/A1 _5287_/S VGND VGND VPWR VPWR _5282_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput248 _6688_/Q VGND VGND VPWR VPWR mgmt_gpio_out[7] sky130_fd_sc_hd__buf_8
X_4302_ _6410_/A0 hold993/X _4303_/S VGND VGND VPWR VPWR _4302_/X sky130_fd_sc_hd__mux2_1
Xoutput259 _3962_/Y VGND VGND VPWR VPWR pad_flash_io1_ieb sky130_fd_sc_hd__buf_8
XFILLER_141_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7021_ _7129_/CLK _7021_/D fanout428/X VGND VGND VPWR VPWR _7021_/Q sky130_fd_sc_hd__dfstp_4
X_4233_ hold523/X _4232_/X _4235_/S VGND VGND VPWR VPWR _4233_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4164_ hold71/X hold376/X _4165_/S VGND VGND VPWR VPWR _6632_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4095_ _6574_/Q _3415_/X _4096_/S VGND VGND VPWR VPWR _6574_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_646 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6805_ _6810_/CLK _6805_/D _6439_/A VGND VGND VPWR VPWR _6805_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4997_ _4997_/A _4997_/B VGND VGND VPWR VPWR _5116_/C sky130_fd_sc_hd__nor2_1
XFILLER_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6736_ _6744_/CLK _6736_/D fanout427/X VGND VGND VPWR VPWR _6736_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_177_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3948_ _6513_/Q user_clock _6835_/Q VGND VGND VPWR VPWR _3948_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6667_ _6668_/CLK _6667_/D _6446_/X VGND VGND VPWR VPWR _6667_/Q sky130_fd_sc_hd__dfrtp_2
X_3879_ _6485_/Q _6459_/Q _3847_/B VGND VGND VPWR VPWR _3879_/X sky130_fd_sc_hd__a21o_1
XFILLER_191_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6598_ _6840_/CLK _6598_/D fanout424/X VGND VGND VPWR VPWR _6598_/Q sky130_fd_sc_hd__dfrtp_2
X_5618_ _7160_/Q _5616_/A _5617_/A VGND VGND VPWR VPWR _5618_/Y sky130_fd_sc_hd__a21boi_1
X_5549_ hold85/X _5594_/B VGND VGND VPWR VPWR hold86/A sky130_fd_sc_hd__and2_4
XFILLER_145_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7219_ _7220_/CLK _7219_/D _6362_/B VGND VGND VPWR VPWR _7219_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout431 fanout456/X VGND VGND VPWR VPWR fanout431/X sky130_fd_sc_hd__buf_8
Xfanout420 fanout421/X VGND VGND VPWR VPWR fanout420/X sky130_fd_sc_hd__buf_8
Xfanout453 fanout454/X VGND VGND VPWR VPWR fanout453/X sky130_fd_sc_hd__buf_8
Xfanout442 fanout456/X VGND VGND VPWR VPWR fanout442/X sky130_fd_sc_hd__buf_8
XFILLER_171_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A VGND VGND VPWR VPWR _7208_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4920_ _4920_/A _4920_/B _4920_/C _5047_/A VGND VGND VPWR VPWR _5163_/A sky130_fd_sc_hd__or4_1
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4851_ _4478_/B _4851_/B VGND VGND VPWR VPWR _4989_/B sky130_fd_sc_hd__nand2b_1
XANTENNA_391 _5706_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_380 _3452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3802_ _3802_/A _3802_/B VGND VGND VPWR VPWR _6486_/D sky130_fd_sc_hd__and2_1
XFILLER_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4782_ _4775_/A _4990_/A _4756_/B _4745_/A VGND VGND VPWR VPWR _4800_/B sky130_fd_sc_hd__o22ai_2
XFILLER_193_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6521_ _7130_/CLK _6521_/D fanout452/X VGND VGND VPWR VPWR _6521_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_158_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3733_ _4241_/A _3733_/B VGND VGND VPWR VPWR _5236_/A sky130_fd_sc_hd__nor2_1
XFILLER_119_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6452_ _6454_/A _6454_/B VGND VGND VPWR VPWR _6452_/X sky130_fd_sc_hd__and2_1
X_3664_ _3664_/A _3664_/B _3664_/C _3664_/D VGND VGND VPWR VPWR _3665_/C sky130_fd_sc_hd__or4_1
XFILLER_134_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5403_ hold260/X hold209/X _5404_/S VGND VGND VPWR VPWR _5403_/X sky130_fd_sc_hd__mux2_1
X_6383_ _6705_/Q _6383_/A2 _6383_/B1 _4238_/B VGND VGND VPWR VPWR _6383_/X sky130_fd_sc_hd__a22o_1
XFILLER_127_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3595_ _7064_/Q _3317_/Y _4178_/A _6647_/Q _3558_/X VGND VGND VPWR VPWR _3598_/B
+ sky130_fd_sc_hd__a221o_4
X_5334_ hold960/X _5595_/A0 _5341_/S VGND VGND VPWR VPWR _6917_/D sky130_fd_sc_hd__mux2_1
XFILLER_125_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5265_ hold198/X hold136/X _5269_/S VGND VGND VPWR VPWR _5265_/X sky130_fd_sc_hd__mux2_1
X_4216_ hold874/X _4215_/X _4218_/S VGND VGND VPWR VPWR _4216_/X sky130_fd_sc_hd__mux2_1
X_7004_ _7156_/CLK _7004_/D fanout445/X VGND VGND VPWR VPWR _7004_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_87_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5196_ _5254_/A0 hold932/X _5199_/S VGND VGND VPWR VPWR _5196_/X sky130_fd_sc_hd__mux2_1
X_4147_ _5545_/A0 _4147_/A1 _4147_/S VGND VGND VPWR VPWR _4147_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4078_ _6559_/Q _6367_/A1 _4081_/S VGND VGND VPWR VPWR _6559_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6719_ _6747_/CLK _6719_/D fanout427/X VGND VGND VPWR VPWR _6719_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_109_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold709 _5538_/X VGND VGND VPWR VPWR _7099_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_170_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3380_ _6470_/Q _6666_/Q VGND VGND VPWR VPWR _3928_/A sky130_fd_sc_hd__nand2_8
XFILLER_69_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5050_ _5050_/A _5050_/B _5050_/C VGND VGND VPWR VPWR _5050_/X sky130_fd_sc_hd__or3_1
XFILLER_69_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4001_ hold619/X _5582_/A0 _4003_/S VGND VGND VPWR VPWR _6501_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5952_ _6716_/Q _5676_/X _5702_/X _6553_/Q _5951_/X VGND VGND VPWR VPWR _5953_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4903_ _4903_/A _4936_/C _4903_/C _4878_/A VGND VGND VPWR VPWR _4904_/D sky130_fd_sc_hd__or4b_1
XFILLER_80_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5883_ _5883_/A _5883_/B _5883_/C _5883_/D VGND VGND VPWR VPWR _5883_/X sky130_fd_sc_hd__or4_1
XFILLER_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4834_ _4834_/A _4834_/B _4834_/C _4834_/D VGND VGND VPWR VPWR _4838_/B sky130_fd_sc_hd__or4_4
XFILLER_21_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4765_ _4563_/X _4645_/X _4764_/X _4239_/X _6778_/Q VGND VGND VPWR VPWR _6778_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_193_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6504_ _6825_/CLK _6504_/D fanout429/X VGND VGND VPWR VPWR _6504_/Q sky130_fd_sc_hd__dfstp_4
X_3716_ _7006_/Q _5432_/A _5450_/A _7022_/Q _3715_/X VGND VGND VPWR VPWR _3717_/D
+ sky130_fd_sc_hd__a221o_1
X_4696_ _4696_/A _4696_/B VGND VGND VPWR VPWR _5062_/C sky130_fd_sc_hd__nand2_8
XFILLER_146_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6435_ _6439_/A _6446_/B VGND VGND VPWR VPWR _6435_/X sky130_fd_sc_hd__and2_1
X_3647_ _6807_/Q _5200_/A _5185_/A _6787_/Q _3646_/X VGND VGND VPWR VPWR _3654_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_115_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3578_ _3578_/A _3578_/B _3578_/C _3578_/D VGND VGND VPWR VPWR _3588_/C sky130_fd_sc_hd__or4_1
X_6366_ _7206_/Q _3606_/X _6370_/S VGND VGND VPWR VPWR _7206_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5317_ _5587_/A0 hold741/X _5323_/S VGND VGND VPWR VPWR _6902_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold14 hold3/X VGND VGND VPWR VPWR hold14/X sky130_fd_sc_hd__bufbuf_16
X_6297_ _6745_/Q _6023_/A _6033_/X _6740_/Q _6296_/X VGND VGND VPWR VPWR _6306_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_102_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5248_ _5597_/A0 hold541/X _5251_/S VGND VGND VPWR VPWR _5248_/X sky130_fd_sc_hd__mux2_1
Xhold36 hold36/A VGND VGND VPWR VPWR hold67/A sky130_fd_sc_hd__bufbuf_16
XFILLER_102_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold25 hold25/A VGND VGND VPWR VPWR hold25/X sky130_fd_sc_hd__bufbuf_16
Xhold47 hold47/A VGND VGND VPWR VPWR hold47/X sky130_fd_sc_hd__bufbuf_16
Xhold69 hold69/A VGND VGND VPWR VPWR hold69/X sky130_fd_sc_hd__bufbuf_16
XFILLER_130_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5179_ _5023_/A _4988_/A _5164_/B _4757_/B VGND VGND VPWR VPWR _5179_/X sky130_fd_sc_hd__o22a_1
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold58 hold58/A VGND VGND VPWR VPWR hold58/X sky130_fd_sc_hd__bufbuf_16
XFILLER_56_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4550_ _4987_/B _4575_/B _4519_/Y _4549_/X VGND VGND VPWR VPWR _4551_/C sky130_fd_sc_hd__a211o_1
XFILLER_7_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4481_ _4558_/B _4663_/A VGND VGND VPWR VPWR _4986_/C sky130_fd_sc_hd__or2_4
XFILLER_128_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold506 _5485_/X VGND VGND VPWR VPWR _7052_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold517 _7222_/Q VGND VGND VPWR VPWR hold517/X sky130_fd_sc_hd__bufbuf_16
X_3501_ _3501_/A _3534_/A VGND VGND VPWR VPWR _4178_/A sky130_fd_sc_hd__nor2_8
Xhold539 _6891_/Q VGND VGND VPWR VPWR hold539/X sky130_fd_sc_hd__bufbuf_16
X_6220_ _7116_/Q _6027_/B _6021_/B _7156_/Q VGND VGND VPWR VPWR _6220_/X sky130_fd_sc_hd__a22o_1
XFILLER_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3432_ _6858_/Q _3315_/Y _3317_/Y _7066_/Q _3431_/X VGND VGND VPWR VPWR _3436_/A
+ sky130_fd_sc_hd__a221o_1
Xhold528 _4258_/X VGND VGND VPWR VPWR _6714_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_143_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6151_ _6873_/Q _6023_/C _6025_/B _6897_/Q _6150_/X VGND VGND VPWR VPWR _6156_/B
+ sky130_fd_sc_hd__a221o_1
X_3363_ _3972_/B _4234_/S _5360_/A _6948_/Q _3360_/X VGND VGND VPWR VPWR _3377_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _5037_/B _5102_/B _5102_/C _5102_/D VGND VGND VPWR VPWR _5161_/C sky130_fd_sc_hd__and4b_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _6082_/A _6082_/B _6082_/C _6082_/D VGND VGND VPWR VPWR _6083_/C sky130_fd_sc_hd__or4_4
XFILLER_85_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1206 _4119_/X VGND VGND VPWR VPWR _6594_/D sky130_fd_sc_hd__bufbuf_16
X_3294_ hold59/X _3304_/B VGND VGND VPWR VPWR _3473_/A sky130_fd_sc_hd__or2_4
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1239 _6697_/Q VGND VGND VPWR VPWR _4249_/A1 sky130_fd_sc_hd__bufbuf_16
X_5033_ _5033_/A _5033_/B _5033_/C _5032_/X VGND VGND VPWR VPWR _5095_/C sky130_fd_sc_hd__or4b_2
Xhold1217 _6713_/Q VGND VGND VPWR VPWR _4257_/A0 sky130_fd_sc_hd__bufbuf_16
XFILLER_57_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1228 _6639_/Q VGND VGND VPWR VPWR _4173_/A0 sky130_fd_sc_hd__bufbuf_16
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6984_ _6987_/CLK _6984_/D fanout451/X VGND VGND VPWR VPWR _6984_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_80_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5935_ _6740_/Q _5678_/X _5688_/X _6770_/Q VGND VGND VPWR VPWR _5935_/X sky130_fd_sc_hd__a22o_1
X_5866_ _7012_/Q _5678_/X _5683_/X _7044_/Q _5865_/X VGND VGND VPWR VPWR _5871_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_166_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4817_ _4817_/A _4817_/B _4817_/C _4817_/D VGND VGND VPWR VPWR _4834_/A sky130_fd_sc_hd__or4_1
XFILLER_139_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5797_ _6961_/Q _5673_/X _5681_/X _6921_/Q VGND VGND VPWR VPWR _5797_/X sky130_fd_sc_hd__a22o_2
X_4748_ _4748_/A _4748_/B VGND VGND VPWR VPWR _5123_/B sky130_fd_sc_hd__nand2_2
X_4679_ _4920_/C _5047_/A _4679_/C VGND VGND VPWR VPWR _4680_/C sky130_fd_sc_hd__or3_1
XFILLER_134_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6418_ _6421_/A _6421_/B VGND VGND VPWR VPWR _6418_/X sky130_fd_sc_hd__and2_1
XFILLER_1_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6349_ _6623_/Q _6022_/C _6032_/X _6653_/Q VGND VGND VPWR VPWR _6349_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput115 wb_adr_i[24] VGND VGND VPWR VPWR _3887_/C sky130_fd_sc_hd__clkbuf_4
Xinput126 wb_adr_i[5] VGND VGND VPWR VPWR _5007_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput104 wb_adr_i[14] VGND VGND VPWR VPWR _4350_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_102_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput148 wb_dat_i[24] VGND VGND VPWR VPWR _6378_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput137 wb_dat_i[14] VGND VGND VPWR VPWR _6395_/B1 sky130_fd_sc_hd__clkbuf_4
Xinput159 wb_dat_i[5] VGND VGND VPWR VPWR _6393_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_130_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3981_ hold65/X hold159/X _3991_/S VGND VGND VPWR VPWR _3981_/X sky130_fd_sc_hd__mux2_8
XFILLER_62_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5720_ _5720_/A _5720_/B _5720_/C _5720_/D VGND VGND VPWR VPWR _5720_/X sky130_fd_sc_hd__or4_4
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5651_ _7171_/Q _7170_/Q VGND VGND VPWR VPWR _6037_/C sky130_fd_sc_hd__and2b_4
X_4602_ _4603_/B _4947_/B VGND VGND VPWR VPWR _5069_/A sky130_fd_sc_hd__nor2_1
X_5582_ _5582_/A0 hold661/X hold62/X VGND VGND VPWR VPWR _5582_/X sky130_fd_sc_hd__mux2_1
X_4533_ _4533_/A _4533_/B _4533_/C VGND VGND VPWR VPWR _5147_/A sky130_fd_sc_hd__or3_4
XFILLER_156_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold303 _7001_/Q VGND VGND VPWR VPWR hold303/X sky130_fd_sc_hd__bufbuf_16
Xhold314 _6982_/Q VGND VGND VPWR VPWR hold314/X sky130_fd_sc_hd__bufbuf_16
XFILLER_144_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold325 _6779_/Q VGND VGND VPWR VPWR hold325/X sky130_fd_sc_hd__bufbuf_16
Xhold336 _5350_/X VGND VGND VPWR VPWR _6932_/D sky130_fd_sc_hd__bufbuf_16
X_4464_ _4685_/A _4651_/B VGND VGND VPWR VPWR _4758_/A sky130_fd_sc_hd__nor2_8
Xhold347 _6916_/Q VGND VGND VPWR VPWR hold347/X sky130_fd_sc_hd__bufbuf_16
XFILLER_171_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold369 _5395_/X VGND VGND VPWR VPWR _6972_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_117_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6203_ _6867_/Q _6025_/D _6029_/X _7051_/Q _6202_/X VGND VGND VPWR VPWR _6206_/C
+ sky130_fd_sc_hd__a221o_1
Xhold358 _3271_/X VGND VGND VPWR VPWR hold82/A sky130_fd_sc_hd__bufbuf_16
X_4395_ _4818_/A _4672_/A _4469_/A _4395_/D VGND VGND VPWR VPWR _4711_/A sky130_fd_sc_hd__and4_4
X_7183_ _7197_/CLK _7183_/D fanout432/X VGND VGND VPWR VPWR _7183_/Q sky130_fd_sc_hd__dfrtp_2
X_3415_ _3415_/A _3415_/B _3415_/C _3415_/D VGND VGND VPWR VPWR _3415_/X sky130_fd_sc_hd__or4_4
XFILLER_131_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6134_ _5611_/A _7191_/Q _6358_/B1 _6133_/X VGND VGND VPWR VPWR _6134_/X sky130_fd_sc_hd__a211o_1
X_3346_ _5252_/A _3375_/B VGND VGND VPWR VPWR _5585_/A sky130_fd_sc_hd__nor2_8
Xhold1003 _7149_/Q VGND VGND VPWR VPWR _5595_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_100_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1014 _6803_/Q VGND VGND VPWR VPWR _5198_/A1 sky130_fd_sc_hd__bufbuf_16
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _7022_/Q _6010_/Y _6031_/X _7086_/Q _6064_/X VGND VGND VPWR VPWR _6071_/A
+ sky130_fd_sc_hd__a221o_1
X_5016_ _5016_/A _5156_/B _5016_/C _5015_/X VGND VGND VPWR VPWR _5018_/C sky130_fd_sc_hd__or4b_2
Xhold1025 _6909_/Q VGND VGND VPWR VPWR _5325_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1047 _4255_/X VGND VGND VPWR VPWR _6712_/D sky130_fd_sc_hd__bufbuf_16
Xhold1036 _6717_/Q VGND VGND VPWR VPWR _4261_/A0 sky130_fd_sc_hd__bufbuf_16
Xhold1058 _6653_/Q VGND VGND VPWR VPWR _4189_/A0 sky130_fd_sc_hd__bufbuf_16
X_3277_ _3991_/S hold51/X hold193/X VGND VGND VPWR VPWR _3277_/Y sky130_fd_sc_hd__o21bai_4
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1069 _6723_/Q VGND VGND VPWR VPWR _4269_/A0 sky130_fd_sc_hd__bufbuf_16
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_209 _7062_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6967_ _7111_/CLK _6967_/D fanout444/X VGND VGND VPWR VPWR _6967_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5918_ _7185_/Q _6309_/S _5917_/X VGND VGND VPWR VPWR _7185_/D sky130_fd_sc_hd__o21a_1
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6898_ _6976_/CLK _6898_/D fanout451/X VGND VGND VPWR VPWR _6898_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_139_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5849_ _5849_/A _5849_/B _5849_/C _5849_/D VGND VGND VPWR VPWR _5849_/X sky130_fd_sc_hd__or4_1
XFILLER_167_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold881 _5250_/X VGND VGND VPWR VPWR _6843_/D sky130_fd_sc_hd__bufbuf_16
Xhold870 _6726_/Q VGND VGND VPWR VPWR hold870/X sky130_fd_sc_hd__bufbuf_16
XFILLER_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold892 _4051_/X VGND VGND VPWR VPWR _6536_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4180_ hold607/X _6408_/A0 _4183_/S VGND VGND VPWR VPWR _4180_/X sky130_fd_sc_hd__mux2_1
X_3200_ _6679_/Q VGND VGND VPWR VPWR _5663_/B sky130_fd_sc_hd__clkinv_8
XFILLER_164_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6821_ _7035_/CLK _6821_/D fanout433/X VGND VGND VPWR VPWR _6821_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3964_ _6474_/Q _3964_/B VGND VGND VPWR VPWR _3964_/X sky130_fd_sc_hd__and2b_4
X_6752_ _7225_/CLK _6752_/D fanout420/X VGND VGND VPWR VPWR _6752_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3895_ _3895_/A _3895_/B _3895_/C _3895_/D VGND VGND VPWR VPWR _3915_/B sky130_fd_sc_hd__nor4_4
XFILLER_176_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5703_ _5864_/B _5703_/B _5704_/B VGND VGND VPWR VPWR _5703_/X sky130_fd_sc_hd__and3_4
X_6683_ _7107_/CLK _6683_/D fanout434/X VGND VGND VPWR VPWR _6683_/Q sky130_fd_sc_hd__dfrtp_2
X_5634_ _7164_/Q _5635_/B _5633_/B _5636_/S VGND VGND VPWR VPWR _7164_/D sky130_fd_sc_hd__a31o_1
XFILLER_12_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold100 hold46/X VGND VGND VPWR VPWR _5486_/B sky130_fd_sc_hd__bufbuf_16
X_5565_ _5583_/A0 hold698/X _5566_/S VGND VGND VPWR VPWR _5565_/X sky130_fd_sc_hd__mux2_1
Xhold133 hold69/X VGND VGND VPWR VPWR hold133/X sky130_fd_sc_hd__bufbuf_16
XFILLER_132_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4516_ _4871_/A _4636_/A VGND VGND VPWR VPWR _5136_/A sky130_fd_sc_hd__nor2_2
Xhold144 _6783_/Q VGND VGND VPWR VPWR hold144/X sky130_fd_sc_hd__bufbuf_16
Xhold122 _3262_/X VGND VGND VPWR VPWR hold26/A sky130_fd_sc_hd__bufbuf_16
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5496_ _5541_/A0 _5496_/A1 _5503_/S VGND VGND VPWR VPWR _7061_/D sky130_fd_sc_hd__mux2_1
Xhold111 hold57/X VGND VGND VPWR VPWR hold111/X sky130_fd_sc_hd__bufbuf_16
Xhold166 _4029_/X VGND VGND VPWR VPWR _6517_/D sky130_fd_sc_hd__bufbuf_16
X_4447_ _4696_/A _4446_/B _4445_/X _4707_/B VGND VGND VPWR VPWR _4510_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_104_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold155 _3975_/Y VGND VGND VPWR VPWR hold155/X sky130_fd_sc_hd__bufbuf_16
Xhold177 hold60/X VGND VGND VPWR VPWR _3552_/B sky130_fd_sc_hd__bufbuf_16
Xhold188 _5402_/X VGND VGND VPWR VPWR _6978_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_132_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7166_ _3949_/A1 _7166_/D fanout455/X VGND VGND VPWR VPWR _7166_/Q sky130_fd_sc_hd__dfstp_4
Xhold199 _5265_/X VGND VGND VPWR VPWR _6856_/D sky130_fd_sc_hd__bufbuf_16
X_6117_ _7000_/Q _5987_/Y _6022_/D _6920_/Q VGND VGND VPWR VPWR _6117_/X sky130_fd_sc_hd__a22o_1
X_4378_ _4469_/A _5031_/A VGND VGND VPWR VPWR _4987_/B sky130_fd_sc_hd__nor2_8
XFILLER_86_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_1_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6786_/CLK sky130_fd_sc_hd__clkbuf_8
X_3329_ _4241_/A _4241_/B VGND VGND VPWR VPWR _4217_/S sky130_fd_sc_hd__nor2_8
XFILLER_100_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7097_ _7097_/CLK _7097_/D fanout437/X VGND VGND VPWR VPWR _7097_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6048_ _6885_/Q _6020_/A _6021_/D _7141_/Q _6047_/X VGND VGND VPWR VPWR _6058_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_86_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_0_0_mgmt_gpio_in[4] clkbuf_2_1_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _3957_/A1
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_150_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3680_ _6958_/Q _5378_/A _5405_/A _6982_/Q VGND VGND VPWR VPWR _3680_/X sky130_fd_sc_hd__a22o_4
XFILLER_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5350_ _5602_/A0 hold335/X _5350_/S VGND VGND VPWR VPWR _5350_/X sky130_fd_sc_hd__mux2_1
Xoutput205 _3931_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[37] sky130_fd_sc_hd__buf_8
Xoutput216 _6510_/Q VGND VGND VPWR VPWR mgmt_gpio_out[12] sky130_fd_sc_hd__buf_8
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput227 _6675_/Q VGND VGND VPWR VPWR mgmt_gpio_out[22] sky130_fd_sc_hd__buf_8
Xoutput238 _3934_/X VGND VGND VPWR VPWR mgmt_gpio_out[32] sky130_fd_sc_hd__buf_8
X_5281_ _5587_/A0 hold556/X _5287_/S VGND VGND VPWR VPWR _6870_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput249 _3939_/X VGND VGND VPWR VPWR mgmt_gpio_out[8] sky130_fd_sc_hd__buf_8
XFILLER_5_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4301_ _6409_/A0 _4301_/A1 _4303_/S VGND VGND VPWR VPWR _6750_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7020_ _7140_/CLK _7020_/D fanout430/X VGND VGND VPWR VPWR _7020_/Q sky130_fd_sc_hd__dfrtp_2
X_4232_ hold246/X hold209/A _4234_/S VGND VGND VPWR VPWR _4232_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4163_ _5300_/A0 hold968/X _4165_/S VGND VGND VPWR VPWR _4163_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4094_ _6573_/Q _3452_/X _4096_/S VGND VGND VPWR VPWR _6573_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4996_ _4996_/A _4997_/B VGND VGND VPWR VPWR _5136_/D sky130_fd_sc_hd__nor2_1
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6804_ _6804_/CLK _6804_/D _6439_/A VGND VGND VPWR VPWR _6804_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_51_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6735_ _6745_/CLK _6735_/D _6421_/A VGND VGND VPWR VPWR _6735_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_11_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3947_ _3239_/Y input2/X input1/X VGND VGND VPWR VPWR _3947_/X sky130_fd_sc_hd__mux2_8
XFILLER_51_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3878_ _6455_/A _6455_/B VGND VGND VPWR VPWR _3878_/X sky130_fd_sc_hd__and2_1
X_6666_ _6668_/CLK _6666_/D _6445_/X VGND VGND VPWR VPWR _6666_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_136_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6597_ _6840_/CLK _6597_/D fanout424/X VGND VGND VPWR VPWR _6597_/Q sky130_fd_sc_hd__dfrtp_2
X_5617_ _5617_/A _5617_/B _5617_/C VGND VGND VPWR VPWR _7159_/D sky130_fd_sc_hd__and3_1
XFILLER_155_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5548_ hold14/X _5548_/A1 hold22/X VGND VGND VPWR VPWR hold23/A sky130_fd_sc_hd__mux2_1
XFILLER_117_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7218_ _3949_/A1 _7218_/D fanout458/X VGND VGND VPWR VPWR _7218_/Q sky130_fd_sc_hd__dfrtp_2
X_5479_ hold455/X _5578_/A0 _5485_/S VGND VGND VPWR VPWR _7046_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout421 fanout423/X VGND VGND VPWR VPWR fanout421/X sky130_fd_sc_hd__buf_8
Xfanout432 fanout435/X VGND VGND VPWR VPWR fanout432/X sky130_fd_sc_hd__buf_8
Xfanout410 _6454_/B VGND VGND VPWR VPWR _6446_/B sky130_fd_sc_hd__buf_8
XFILLER_48_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout454 fanout455/X VGND VGND VPWR VPWR fanout454/X sky130_fd_sc_hd__buf_8
X_7149_ _7151_/CLK _7149_/D fanout445/X VGND VGND VPWR VPWR _7149_/Q sky130_fd_sc_hd__dfstp_4
Xfanout443 fanout455/X VGND VGND VPWR VPWR fanout443/X sky130_fd_sc_hd__buf_8
XFILLER_101_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_370 _6690_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4850_ _4850_/A _4850_/B VGND VGND VPWR VPWR _4850_/X sky130_fd_sc_hd__or2_1
XFILLER_33_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_392 _5826_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_381 _4256_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3801_ _6486_/Q _3801_/B VGND VGND VPWR VPWR _3802_/B sky130_fd_sc_hd__or2_1
XFILLER_193_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6520_ _7130_/CLK _6520_/D fanout452/X VGND VGND VPWR VPWR _6520_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4781_ _4622_/B _4772_/A _5178_/A VGND VGND VPWR VPWR _4800_/A sky130_fd_sc_hd__a21o_1
XFILLER_146_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3732_ _5225_/A _3732_/B VGND VGND VPWR VPWR _5216_/A sky130_fd_sc_hd__nor2_2
XFILLER_173_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6451_ _6454_/A _6454_/B VGND VGND VPWR VPWR _6451_/X sky130_fd_sc_hd__and2_1
X_3663_ _3726_/A _3663_/B _3663_/C _3663_/D VGND VGND VPWR VPWR _3664_/D sky130_fd_sc_hd__or4_1
X_6382_ _6381_/X _7212_/Q _6400_/S VGND VGND VPWR VPWR _7212_/D sky130_fd_sc_hd__mux2_1
X_5402_ hold187/X hold78/X _5404_/S VGND VGND VPWR VPWR _5402_/X sky130_fd_sc_hd__mux2_1
X_5333_ _5333_/A _5594_/B VGND VGND VPWR VPWR _5341_/S sky130_fd_sc_hd__and2_4
XFILLER_161_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3594_ _6491_/Q _3978_/A _4298_/A _6751_/Q _3557_/X VGND VGND VPWR VPWR _3598_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_114_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5264_ hold756/X _5561_/A0 _5269_/S VGND VGND VPWR VPWR _5264_/X sky130_fd_sc_hd__mux2_1
X_4215_ hold521/X _5601_/A0 _4217_/S VGND VGND VPWR VPWR _4215_/X sky130_fd_sc_hd__mux2_1
X_7003_ _7154_/CLK _7003_/D fanout452/X VGND VGND VPWR VPWR _7003_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_87_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5195_ _5234_/C _5195_/A1 _5199_/S VGND VGND VPWR VPWR _5195_/X sky130_fd_sc_hd__mux2_1
X_4146_ _4326_/A0 hold808/X _4147_/S VGND VGND VPWR VPWR _4146_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4077_ _6558_/Q _3606_/X _4081_/S VGND VGND VPWR VPWR _6558_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4979_ _4913_/B _4977_/X _5060_/B VGND VGND VPWR VPWR _4979_/X sky130_fd_sc_hd__o21ba_4
X_6718_ _6951_/CLK _6718_/D fanout442/X VGND VGND VPWR VPWR _6718_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_137_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6649_ _6649_/CLK _6649_/D fanout456/X VGND VGND VPWR VPWR _6649_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_125_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_34_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7130_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_164_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_49_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7075_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_74_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4000_ hold769/X _6411_/A0 _4003_/S VGND VGND VPWR VPWR _6500_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5951_ _6662_/Q _5669_/X _5698_/B _5942_/X VGND VGND VPWR VPWR _5951_/X sky130_fd_sc_hd__a22o_1
XFILLER_65_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4902_ _4987_/A _4536_/X _4962_/A _4886_/Y VGND VGND VPWR VPWR _4904_/C sky130_fd_sc_hd__a211o_1
XFILLER_80_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5882_ _6594_/Q _5681_/X _5687_/X _6639_/Q _5881_/X VGND VGND VPWR VPWR _5883_/D
+ sky130_fd_sc_hd__a221o_1
X_4833_ _4697_/A _5005_/C _4832_/X VGND VGND VPWR VPWR _4834_/D sky130_fd_sc_hd__a21oi_1
X_4764_ _5003_/B _4763_/X _6376_/A _4720_/X VGND VGND VPWR VPWR _4764_/X sky130_fd_sc_hd__a211o_4
XFILLER_119_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6503_ _6759_/CLK _6503_/D fanout421/X VGND VGND VPWR VPWR _6503_/Q sky130_fd_sc_hd__dfstp_4
X_3715_ _7054_/Q _5486_/A _3552_/Y _6821_/Q VGND VGND VPWR VPWR _3715_/X sky130_fd_sc_hd__a22o_1
X_4695_ _4696_/A _4696_/B VGND VGND VPWR VPWR _4695_/X sky130_fd_sc_hd__and2_4
X_6434_ _6446_/A _6446_/B VGND VGND VPWR VPWR _6434_/X sky130_fd_sc_hd__and2_1
XFILLER_20_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3646_ _7223_/Q _6406_/A _5194_/A _6802_/Q VGND VGND VPWR VPWR _3646_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3577_ _6872_/Q _5279_/A _4061_/A _6548_/Q _3576_/X VGND VGND VPWR VPWR _3578_/D
+ sky130_fd_sc_hd__a221o_2
X_6365_ _7205_/Q _3665_/X _6370_/S VGND VGND VPWR VPWR _7205_/D sky130_fd_sc_hd__mux2_1
X_5316_ _5595_/A0 _5316_/A1 _5323_/S VGND VGND VPWR VPWR _6901_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6296_ _6552_/Q _6020_/A _6021_/D _6631_/Q _6295_/X VGND VGND VPWR VPWR _6296_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5247_ _6408_/A0 hold491/X _5251_/S VGND VGND VPWR VPWR _5247_/X sky130_fd_sc_hd__mux2_1
Xhold15 hold15/A VGND VGND VPWR VPWR hold15/X sky130_fd_sc_hd__bufbuf_16
XFILLER_88_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold26 hold26/A VGND VGND VPWR VPWR hold26/X sky130_fd_sc_hd__bufbuf_16
Xhold37 hold37/A VGND VGND VPWR VPWR hold37/X sky130_fd_sc_hd__bufbuf_16
X_5178_ _5178_/A _5178_/B _5178_/C _5178_/D VGND VGND VPWR VPWR _5178_/X sky130_fd_sc_hd__or4_4
Xhold59 hold59/A VGND VGND VPWR VPWR hold59/X sky130_fd_sc_hd__bufbuf_16
Xhold48 hold48/A VGND VGND VPWR VPWR hold48/X sky130_fd_sc_hd__bufbuf_16
XFILLER_29_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4129_ hold806/X _5599_/A0 _4129_/S VGND VGND VPWR VPWR _4129_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3500_ hold53/X _4241_/B VGND VGND VPWR VPWR _4166_/A sky130_fd_sc_hd__nor2_8
XFILLER_183_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold507 _6886_/Q VGND VGND VPWR VPWR hold507/X sky130_fd_sc_hd__bufbuf_16
XFILLER_156_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4480_ _4558_/B _4663_/A VGND VGND VPWR VPWR _4992_/B sky130_fd_sc_hd__nor2_4
XFILLER_128_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold518 _6408_/X VGND VGND VPWR VPWR _7222_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_183_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold529 _6908_/Q VGND VGND VPWR VPWR hold529/X sky130_fd_sc_hd__bufbuf_16
XFILLER_143_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3431_ _6866_/Q hold28/A _5245_/A _7229_/A VGND VGND VPWR VPWR _3431_/X sky130_fd_sc_hd__a22o_2
X_6150_ _6961_/Q _6022_/C _6032_/X _7057_/Q VGND VGND VPWR VPWR _6150_/X sky130_fd_sc_hd__a22o_1
X_3362_ hold91/X _3457_/A VGND VGND VPWR VPWR _5360_/A sky130_fd_sc_hd__nor2_8
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _5101_/A _5101_/B _5101_/C _5101_/D VGND VGND VPWR VPWR _5101_/X sky130_fd_sc_hd__or4_1
XFILLER_111_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _7062_/Q _5996_/X _6020_/C _6910_/Q _6080_/X VGND VGND VPWR VPWR _6082_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1207 _6798_/Q VGND VGND VPWR VPWR _5192_/A1 sky130_fd_sc_hd__bufbuf_16
X_3293_ _3278_/B _3293_/B VGND VGND VPWR VPWR _3304_/B sky130_fd_sc_hd__nand2b_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _5023_/A _4997_/A _5164_/B _4754_/B _4767_/X VGND VGND VPWR VPWR _5032_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1218 _4257_/X VGND VGND VPWR VPWR _6713_/D sky130_fd_sc_hd__bufbuf_16
Xhold1229 _4173_/X VGND VGND VPWR VPWR _6639_/D sky130_fd_sc_hd__bufbuf_16
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6983_ _7151_/CLK _6983_/D fanout446/X VGND VGND VPWR VPWR _6983_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_80_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5934_ _6621_/Q _5673_/X _5674_/X _6547_/Q _5933_/X VGND VGND VPWR VPWR _5937_/C
+ sky130_fd_sc_hd__a221o_4
XFILLER_15_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5865_ _6948_/Q _5705_/X _5864_/X _5698_/B VGND VGND VPWR VPWR _5865_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4816_ _4687_/A _4832_/B _4729_/X VGND VGND VPWR VPWR _4817_/D sky130_fd_sc_hd__o21bai_1
XFILLER_193_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5796_ _5796_/A _5796_/B _5796_/C _5796_/D VGND VGND VPWR VPWR _5796_/X sky130_fd_sc_hd__or4_2
XFILLER_21_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4747_ _4728_/X _4735_/X _4746_/X _4740_/B _4745_/X VGND VGND VPWR VPWR _4753_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4678_ _4832_/C _4746_/B _4663_/B VGND VGND VPWR VPWR _4679_/C sky130_fd_sc_hd__a21oi_2
XFILLER_107_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6417_ _6421_/A _6421_/B VGND VGND VPWR VPWR _6417_/X sky130_fd_sc_hd__and2_1
XFILLER_162_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3629_ _3629_/A _3629_/B _3629_/C _3629_/D VGND VGND VPWR VPWR _3636_/C sky130_fd_sc_hd__or4_1
XFILLER_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6348_ _6580_/Q _6021_/A _6025_/A _6608_/Q _6347_/X VGND VGND VPWR VPWR _6355_/A
+ sky130_fd_sc_hd__a221o_1
Xinput127 wb_adr_i[6] VGND VGND VPWR VPWR _4654_/A sky130_fd_sc_hd__buf_8
Xinput116 wb_adr_i[25] VGND VGND VPWR VPWR input116/X sky130_fd_sc_hd__clkbuf_4
Xinput105 wb_adr_i[15] VGND VGND VPWR VPWR _4350_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_102_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6279_ _6660_/Q _5996_/X _6020_/C _6590_/Q VGND VGND VPWR VPWR _6279_/X sky130_fd_sc_hd__a22o_1
Xinput138 wb_dat_i[15] VGND VGND VPWR VPWR _6398_/B1 sky130_fd_sc_hd__clkbuf_4
Xinput149 wb_dat_i[25] VGND VGND VPWR VPWR _6380_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_76_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3980_ _3980_/A0 _6407_/A0 _3994_/S VGND VGND VPWR VPWR _3980_/X sky130_fd_sc_hd__mux2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5650_ _5645_/Y _5649_/Y _5654_/B VGND VGND VPWR VPWR _7170_/D sky130_fd_sc_hd__a21oi_1
XFILLER_175_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4601_ _4603_/B _5062_/A VGND VGND VPWR VPWR _4642_/A sky130_fd_sc_hd__nor2_1
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5581_ _5581_/A0 hold868/X hold62/X VGND VGND VPWR VPWR _5581_/X sky130_fd_sc_hd__mux2_1
X_4532_ _4533_/A _4533_/B _4533_/C VGND VGND VPWR VPWR _4949_/C sky130_fd_sc_hd__nor3_4
XFILLER_156_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4463_ _4654_/A _4958_/A VGND VGND VPWR VPWR _4651_/B sky130_fd_sc_hd__or2_4
Xhold315 _6910_/Q VGND VGND VPWR VPWR hold315/X sky130_fd_sc_hd__bufbuf_16
Xhold304 _5428_/X VGND VGND VPWR VPWR _7001_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_171_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold326 _3269_/X VGND VGND VPWR VPWR hold18/A sky130_fd_sc_hd__bufbuf_16
Xhold337 _6924_/Q VGND VGND VPWR VPWR hold337/X sky130_fd_sc_hd__bufbuf_16
Xhold348 _5332_/X VGND VGND VPWR VPWR _6916_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_131_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6202_ _7107_/Q _5653_/X _6022_/B _6947_/Q VGND VGND VPWR VPWR _6202_/X sky130_fd_sc_hd__a22o_1
Xhold359 _5233_/X VGND VGND VPWR VPWR _6831_/D sky130_fd_sc_hd__bufbuf_16
X_3414_ _3414_/A _3414_/B _3414_/C _3414_/D VGND VGND VPWR VPWR _3415_/D sky130_fd_sc_hd__or4_1
X_4394_ _5031_/A _4663_/A VGND VGND VPWR VPWR _4775_/A sky130_fd_sc_hd__or2_4
X_7182_ _7193_/CLK _7182_/D fanout435/X VGND VGND VPWR VPWR _7182_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6133_ _6856_/Q _6060_/B _6121_/X _6132_/X _3197_/Y VGND VGND VPWR VPWR _6133_/X
+ sky130_fd_sc_hd__o221a_1
X_3345_ _7100_/Q _3341_/Y _3344_/Y _6503_/Q _3340_/X VGND VGND VPWR VPWR _3378_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1004 _6740_/Q VGND VGND VPWR VPWR _4289_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1015 _5198_/X VGND VGND VPWR VPWR _6803_/D sky130_fd_sc_hd__bufbuf_16
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3276_ hold91/X _3501_/A VGND VGND VPWR VPWR hold92/A sky130_fd_sc_hd__nor2_8
X_6064_ _7134_/Q _6020_/B _6011_/X _7094_/Q VGND VGND VPWR VPWR _6064_/X sky130_fd_sc_hd__a22o_1
X_5015_ _4754_/B _4832_/C _5050_/B _4746_/X _5050_/C VGND VGND VPWR VPWR _5015_/X
+ sky130_fd_sc_hd__a41o_1
Xhold1037 _4261_/X VGND VGND VPWR VPWR _6717_/D sky130_fd_sc_hd__bufbuf_16
Xhold1026 _6807_/Q VGND VGND VPWR VPWR _5203_/A1 sky130_fd_sc_hd__bufbuf_16
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1048 _6544_/Q VGND VGND VPWR VPWR _4060_/A1 sky130_fd_sc_hd__bufbuf_16
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1059 _4189_/X VGND VGND VPWR VPWR _6653_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_54_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6966_ _7111_/CLK _6966_/D fanout444/X VGND VGND VPWR VPWR _6966_/Q sky130_fd_sc_hd__dfstp_4
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5917_ _5611_/A _7184_/Q _6358_/B1 _5916_/X VGND VGND VPWR VPWR _5917_/X sky130_fd_sc_hd__a211o_1
XFILLER_41_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6897_ _7121_/CLK _6897_/D _6421_/A VGND VGND VPWR VPWR _6897_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_139_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5848_ _6979_/Q _5676_/X _5684_/X _6995_/Q _5847_/X VGND VGND VPWR VPWR _5849_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_42_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5779_ _6904_/Q _5689_/X _5767_/X _5778_/X VGND VGND VPWR VPWR _5784_/A sky130_fd_sc_hd__a211o_2
XFILLER_108_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold882 _7211_/Q VGND VGND VPWR VPWR hold882/X sky130_fd_sc_hd__bufbuf_16
XFILLER_135_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold871 _4272_/X VGND VGND VPWR VPWR _6726_/D sky130_fd_sc_hd__bufbuf_16
Xhold860 _5543_/X VGND VGND VPWR VPWR _7103_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_103_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold893 _6541_/Q VGND VGND VPWR VPWR hold893/X sky130_fd_sc_hd__bufbuf_16
XFILLER_191_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_728 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6820_ _7035_/CLK _6820_/D fanout433/X VGND VGND VPWR VPWR _6820_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6751_ _6810_/CLK _6751_/D fanout419/X VGND VGND VPWR VPWR _6751_/Q sky130_fd_sc_hd__dfrtp_2
X_3963_ input85/X _3875_/B _6474_/Q VGND VGND VPWR VPWR _3963_/X sky130_fd_sc_hd__mux2_8
X_3894_ _4346_/S _4722_/B _3894_/C _3894_/D VGND VGND VPWR VPWR _3895_/D sky130_fd_sc_hd__or4_4
XFILLER_176_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5702_ _5864_/B _5702_/B _5707_/C VGND VGND VPWR VPWR _5702_/X sky130_fd_sc_hd__and3_4
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_1_1_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
X_6682_ _6851_/CLK _6682_/D _6455_/A VGND VGND VPWR VPWR _6682_/Q sky130_fd_sc_hd__dfrtp_1
X_5633_ _7164_/Q _5633_/B VGND VGND VPWR VPWR _5636_/S sky130_fd_sc_hd__nor2_1
XFILLER_31_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5564_ hold78/X hold142/X _5566_/S VGND VGND VPWR VPWR _5564_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold101 _5378_/Y VGND VGND VPWR VPWR _5386_/S sky130_fd_sc_hd__bufbuf_16
XFILLER_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4515_ _4996_/A _4871_/A VGND VGND VPWR VPWR _5078_/A sky130_fd_sc_hd__nor2_2
Xhold134 hold152/X VGND VGND VPWR VPWR hold70/A sky130_fd_sc_hd__bufbuf_16
XFILLER_144_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5495_ _5495_/A _5594_/B VGND VGND VPWR VPWR _5503_/S sky130_fd_sc_hd__nand2_8
Xhold123 hold26/X VGND VGND VPWR VPWR _3421_/A sky130_fd_sc_hd__bufbuf_16
Xhold112 _3263_/X VGND VGND VPWR VPWR _3264_/B sky130_fd_sc_hd__bufbuf_16
X_4446_ _5050_/A _4446_/B VGND VGND VPWR VPWR _4534_/B sky130_fd_sc_hd__xnor2_4
Xhold156 _5490_/X VGND VGND VPWR VPWR _7056_/D sky130_fd_sc_hd__bufbuf_16
Xhold167 hold180/X VGND VGND VPWR VPWR hold181/A sky130_fd_sc_hd__bufbuf_16
XFILLER_132_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold145 _3254_/X VGND VGND VPWR VPWR hold145/X sky130_fd_sc_hd__bufbuf_16
XFILLER_144_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4377_ _4818_/A _4672_/A VGND VGND VPWR VPWR _5031_/A sky130_fd_sc_hd__nand2_8
X_7165_ _3949_/A1 _7165_/D fanout455/X VGND VGND VPWR VPWR _7165_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_132_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold178 _3552_/Y VGND VGND VPWR VPWR _5218_/A sky130_fd_sc_hd__bufbuf_16
Xhold189 _7017_/Q VGND VGND VPWR VPWR hold189/X sky130_fd_sc_hd__bufbuf_16
XFILLER_98_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6116_ _7016_/Q _6036_/Y _6335_/B _7040_/Q _6111_/X VGND VGND VPWR VPWR _6121_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_86_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3328_ _3383_/C _3419_/A VGND VGND VPWR VPWR _4241_/B sky130_fd_sc_hd__or2_4
XFILLER_100_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7096_ _7104_/CLK _7096_/D fanout434/X VGND VGND VPWR VPWR _7096_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6047_ _7077_/Q _6311_/B _6335_/B _7037_/Q _6046_/X VGND VGND VPWR VPWR _6047_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_100_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3259_ _3991_/S hold51/X hold193/X VGND VGND VPWR VPWR _3259_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_27_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6949_ _7111_/CLK _6949_/D fanout445/X VGND VGND VPWR VPWR _6949_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold690 _6710_/Q VGND VGND VPWR VPWR hold690/X sky130_fd_sc_hd__bufbuf_16
XFILLER_150_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput217 _3950_/X VGND VGND VPWR VPWR mgmt_gpio_out[13] sky130_fd_sc_hd__buf_8
Xoutput206 _3194_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[3] sky130_fd_sc_hd__buf_8
Xoutput228 _6676_/Q VGND VGND VPWR VPWR mgmt_gpio_out[23] sky130_fd_sc_hd__buf_8
Xoutput239 _3935_/X VGND VGND VPWR VPWR mgmt_gpio_out[33] sky130_fd_sc_hd__buf_8
X_5280_ _5595_/A0 hold974/X _5287_/S VGND VGND VPWR VPWR _6869_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4300_ _5254_/A0 hold907/X _4303_/S VGND VGND VPWR VPWR _4300_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4231_ hold930/X _4230_/X _4235_/S VGND VGND VPWR VPWR _4231_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4162_ _6408_/A0 hold595/X _4165_/S VGND VGND VPWR VPWR _4162_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4093_ _6572_/Q _6367_/A1 _4096_/S VGND VGND VPWR VPWR _6572_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4995_ _4995_/A _4997_/B VGND VGND VPWR VPWR _5078_/C sky130_fd_sc_hd__nor2_2
X_6803_ _6804_/CLK _6803_/D _6439_/A VGND VGND VPWR VPWR _6803_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3946_ _3238_/Y _6458_/Q _6454_/B VGND VGND VPWR VPWR _3946_/X sky130_fd_sc_hd__mux2_8
X_6734_ _6744_/CLK _6734_/D fanout427/X VGND VGND VPWR VPWR _6734_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_51_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3877_ _6833_/Q _6880_/Q _3877_/C VGND VGND VPWR VPWR _3877_/Y sky130_fd_sc_hd__nor3_4
X_6665_ _6668_/CLK _6665_/D _6444_/X VGND VGND VPWR VPWR _6665_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_191_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6596_ _6840_/CLK _6596_/D fanout424/X VGND VGND VPWR VPWR _6596_/Q sky130_fd_sc_hd__dfstp_4
X_5616_ _5616_/A VGND VGND VPWR VPWR _5617_/C sky130_fd_sc_hd__inv_2
X_5547_ _5583_/A0 hold639/X hold22/X VGND VGND VPWR VPWR _5547_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5478_ _5478_/A0 _5541_/A0 _5485_/S VGND VGND VPWR VPWR _7045_/D sky130_fd_sc_hd__mux2_1
X_7217_ _3949_/A1 _7217_/D fanout458/X VGND VGND VPWR VPWR _7217_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_160_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4429_ _4507_/A _4851_/B _4499_/C VGND VGND VPWR VPWR _4581_/B sky130_fd_sc_hd__and3_4
XFILLER_160_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout400 _5541_/A0 VGND VGND VPWR VPWR _6407_/A0 sky130_fd_sc_hd__buf_8
Xfanout422 fanout423/X VGND VGND VPWR VPWR fanout422/X sky130_fd_sc_hd__buf_8
Xfanout411 _6454_/B VGND VGND VPWR VPWR _6455_/B sky130_fd_sc_hd__buf_8
X_7148_ _7156_/CLK _7148_/D fanout447/X VGND VGND VPWR VPWR _7148_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout444 fanout455/X VGND VGND VPWR VPWR fanout444/X sky130_fd_sc_hd__buf_8
Xfanout455 fanout456/X VGND VGND VPWR VPWR fanout455/X sky130_fd_sc_hd__buf_8
Xfanout433 fanout435/X VGND VGND VPWR VPWR fanout433/X sky130_fd_sc_hd__buf_8
XFILLER_171_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7079_ _7081_/CLK _7079_/D fanout437/X VGND VGND VPWR VPWR _7079_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_59_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_360 hold335/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4780_ _4772_/A _4586_/B _4748_/B _4453_/Y VGND VGND VPWR VPWR _4799_/B sky130_fd_sc_hd__a22o_1
X_3800_ _6487_/Q _3802_/A VGND VGND VPWR VPWR _6487_/D sky130_fd_sc_hd__xnor2_1
XANTENNA_393 _5937_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_382 _4049_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_371 _5219_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3731_ _5225_/A _4241_/B VGND VGND VPWR VPWR _5223_/A sky130_fd_sc_hd__nor2_4
XFILLER_186_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_0_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6851_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_173_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6450_ _6454_/A _6455_/B VGND VGND VPWR VPWR _6450_/X sky130_fd_sc_hd__and2_1
X_3662_ _6999_/Q _5423_/A _4322_/A _6770_/Q VGND VGND VPWR VPWR _3663_/D sky130_fd_sc_hd__a22o_1
X_6381_ _6705_/Q _6381_/A2 _6381_/B1 _4238_/B _6380_/X VGND VGND VPWR VPWR _6381_/X
+ sky130_fd_sc_hd__a221o_1
X_5401_ hold478/X _5581_/A0 _5404_/S VGND VGND VPWR VPWR _5401_/X sky130_fd_sc_hd__mux2_1
X_3593_ _3593_/A _3593_/B _3593_/C _3593_/D VGND VGND VPWR VPWR _3606_/B sky130_fd_sc_hd__or4_1
X_5332_ _5602_/A0 hold347/X _5332_/S VGND VGND VPWR VPWR _5332_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5263_ hold395/X _5578_/A0 _5269_/S VGND VGND VPWR VPWR _5263_/X sky130_fd_sc_hd__mux2_1
X_4214_ hold273/X _4213_/X _4218_/S VGND VGND VPWR VPWR _4214_/X sky130_fd_sc_hd__mux2_1
X_7002_ _7131_/CLK _7002_/D fanout432/X VGND VGND VPWR VPWR _7002_/Q sky130_fd_sc_hd__dfrtp_2
X_5194_ _5194_/A _6406_/B VGND VGND VPWR VPWR _5199_/S sky130_fd_sc_hd__nand2_4
X_4145_ _5300_/A0 hold979/X _4147_/S VGND VGND VPWR VPWR _6616_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4076_ _6557_/Q _3665_/X _4081_/S VGND VGND VPWR VPWR _6557_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4978_ _4980_/C _4978_/B _4567_/X VGND VGND VPWR VPWR _5060_/B sky130_fd_sc_hd__or3b_2
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3929_ hold95/A input91/X _3932_/S VGND VGND VPWR VPWR _3929_/X sky130_fd_sc_hd__mux2_8
XFILLER_177_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6717_ _6717_/CLK _6717_/D fanout426/X VGND VGND VPWR VPWR _6717_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6648_ _7105_/CLK _6648_/D fanout427/X VGND VGND VPWR VPWR _6648_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6579_ _6717_/CLK _6579_/D fanout426/X VGND VGND VPWR VPWR _6579_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5950_ _6637_/Q _5675_/X _5684_/X _6726_/Q _5949_/X VGND VGND VPWR VPWR _5953_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4901_ _4987_/A _4624_/B _4736_/B _4719_/X VGND VGND VPWR VPWR _4907_/C sky130_fd_sc_hd__a22o_2
XFILLER_80_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5881_ _6723_/Q _5684_/X _5704_/X _6604_/Q VGND VGND VPWR VPWR _5881_/X sky130_fd_sc_hd__a22o_2
XFILLER_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4832_ _4832_/A _4832_/B _4832_/C _4832_/D VGND VGND VPWR VPWR _4832_/X sky130_fd_sc_hd__and4_1
XANTENNA_190 _6259_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4763_ _4808_/A _4763_/B _4980_/B _4763_/D VGND VGND VPWR VPWR _4763_/X sky130_fd_sc_hd__or4_2
XFILLER_174_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4694_ _4694_/A _5005_/C VGND VGND VPWR VPWR _5069_/B sky130_fd_sc_hd__nor2_8
X_6502_ _6759_/CLK _6502_/D fanout421/X VGND VGND VPWR VPWR _6502_/Q sky130_fd_sc_hd__dfstp_4
X_3714_ _7142_/Q _5585_/A _4316_/A _6764_/Q _3713_/X VGND VGND VPWR VPWR _3717_/C
+ sky130_fd_sc_hd__a221o_1
X_6433_ _6446_/A _6446_/B VGND VGND VPWR VPWR _6433_/X sky130_fd_sc_hd__and2_1
XFILLER_174_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3645_ _3645_/A _3645_/B _3645_/C _3645_/D VGND VGND VPWR VPWR _3665_/B sky130_fd_sc_hd__or4_1
XFILLER_161_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3576_ _6880_/Q _5288_/A _4082_/A _6566_/Q VGND VGND VPWR VPWR _3576_/X sky130_fd_sc_hd__a22o_1
X_6364_ _7204_/Q _3727_/X _6370_/S VGND VGND VPWR VPWR _7204_/D sky130_fd_sc_hd__mux2_1
X_5315_ _5315_/A _5558_/B VGND VGND VPWR VPWR _5323_/S sky130_fd_sc_hd__nand2_8
X_6295_ _6765_/Q _6027_/B _6021_/B _6720_/Q VGND VGND VPWR VPWR _6295_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5246_ _6407_/A0 _5246_/A1 _5251_/S VGND VGND VPWR VPWR _5246_/X sky130_fd_sc_hd__mux2_1
Xhold38 hold38/A VGND VGND VPWR VPWR hold38/X sky130_fd_sc_hd__bufbuf_16
XFILLER_102_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold16 hold16/A VGND VGND VPWR VPWR hold16/X sky130_fd_sc_hd__bufbuf_16
Xhold27 hold27/A VGND VGND VPWR VPWR hold27/X sky130_fd_sc_hd__bufbuf_16
X_5177_ _5048_/A _5177_/B VGND VGND VPWR VPWR _5178_/D sky130_fd_sc_hd__nand2b_1
Xhold49 hold49/A VGND VGND VPWR VPWR hold49/X sky130_fd_sc_hd__bufbuf_16
XFILLER_188_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4128_ hold232/X hold71/X _4129_/S VGND VGND VPWR VPWR _4128_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4059_ _6410_/A0 _4059_/A1 _4060_/S VGND VGND VPWR VPWR _4059_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold508 _6974_/Q VGND VGND VPWR VPWR hold508/X sky130_fd_sc_hd__bufbuf_16
XFILLER_143_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold519 _6876_/Q VGND VGND VPWR VPWR hold519/X sky130_fd_sc_hd__bufbuf_16
XFILLER_109_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3430_ _6501_/Q _3344_/Y _3368_/Y input17/X VGND VGND VPWR VPWR _3430_/X sky130_fd_sc_hd__a22o_2
XFILLER_171_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3361_ _5252_/A _5252_/B VGND VGND VPWR VPWR _4234_/S sky130_fd_sc_hd__nor2_8
X_5100_ _4414_/B _5165_/A _5119_/A _4932_/C VGND VGND VPWR VPWR _5101_/D sky130_fd_sc_hd__a211o_1
X_6080_ _6974_/Q _6023_/B _6021_/C _6878_/Q VGND VGND VPWR VPWR _6080_/X sky130_fd_sc_hd__a22o_1
XFILLER_97_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _5031_/A _5031_/B _4584_/A VGND VGND VPWR VPWR _5102_/B sky130_fd_sc_hd__or3b_1
XFILLER_112_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3292_ hold26/X _3421_/B hold19/X VGND VGND VPWR VPWR _3292_/X sky130_fd_sc_hd__or3_4
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1219 _6496_/Q VGND VGND VPWR VPWR _3996_/A0 sky130_fd_sc_hd__bufbuf_16
Xhold1208 _5192_/X VGND VGND VPWR VPWR _6798_/D sky130_fd_sc_hd__bufbuf_16
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6982_ _7151_/CLK _6982_/D fanout447/X VGND VGND VPWR VPWR _6982_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_19_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_33_csclk _7137_/CLK VGND VGND VPWR VPWR _7154_/CLK sky130_fd_sc_hd__clkbuf_8
X_5933_ _6710_/Q _5691_/X _5704_/X _6606_/Q VGND VGND VPWR VPWR _5933_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5864_ _6988_/Q _5864_/B VGND VGND VPWR VPWR _5864_/X sky130_fd_sc_hd__or2_1
XFILLER_21_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4815_ _4687_/A _4728_/X _4881_/B VGND VGND VPWR VPWR _4817_/C sky130_fd_sc_hd__o21ai_4
XFILLER_178_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5795_ _6929_/Q _5699_/X _5707_/X _7025_/Q _5794_/X VGND VGND VPWR VPWR _5796_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_193_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4746_ _4746_/A _4746_/B VGND VGND VPWR VPWR _4746_/X sky130_fd_sc_hd__or2_4
XFILLER_147_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_48_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7106_/CLK sky130_fd_sc_hd__clkbuf_8
X_4677_ _4690_/A _5062_/B VGND VGND VPWR VPWR _4746_/B sky130_fd_sc_hd__or2_4
XFILLER_135_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6416_ _6421_/A _6421_/B VGND VGND VPWR VPWR _6416_/X sky130_fd_sc_hd__and2_1
XFILLER_162_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3628_ input54/X _4025_/A _4292_/A _6745_/Q _3617_/X VGND VGND VPWR VPWR _3629_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6347_ _6618_/Q _6022_/A _6025_/C _6603_/Q VGND VGND VPWR VPWR _6347_/X sky130_fd_sc_hd__a22o_1
X_3559_ _7112_/Q hold85/A _5227_/A _6827_/Q VGND VGND VPWR VPWR _3559_/X sky130_fd_sc_hd__a22o_2
Xinput106 wb_adr_i[16] VGND VGND VPWR VPWR _4349_/B sky130_fd_sc_hd__clkbuf_4
Xinput117 wb_adr_i[26] VGND VGND VPWR VPWR input117/X sky130_fd_sc_hd__clkbuf_4
X_6278_ _6536_/Q _6025_/D _6029_/X _6640_/Q _6277_/X VGND VGND VPWR VPWR _6281_/C
+ sky130_fd_sc_hd__a221o_1
Xinput128 wb_adr_i[7] VGND VGND VPWR VPWR _4958_/A sky130_fd_sc_hd__buf_8
Xinput139 wb_dat_i[16] VGND VGND VPWR VPWR _6377_/A2 sky130_fd_sc_hd__clkbuf_4
X_5229_ hold136/X _5229_/A1 _5233_/S VGND VGND VPWR VPWR _5229_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_90 _3606_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_97_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4600_ _4617_/A _4749_/C VGND VGND VPWR VPWR _4850_/B sky130_fd_sc_hd__nor2_2
XFILLER_30_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5580_ hold136/X hold244/X hold62/X VGND VGND VPWR VPWR _5580_/X sky130_fd_sc_hd__mux2_1
X_4531_ _4529_/B _4529_/C _4650_/B VGND VGND VPWR VPWR _4537_/C sky130_fd_sc_hd__a21bo_1
XFILLER_184_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4462_ _4707_/B _5050_/A VGND VGND VPWR VPWR _4685_/A sky130_fd_sc_hd__or2_4
Xhold316 _5326_/X VGND VGND VPWR VPWR _6910_/D sky130_fd_sc_hd__bufbuf_16
Xhold305 _6553_/Q VGND VGND VPWR VPWR hold305/X sky130_fd_sc_hd__bufbuf_16
XFILLER_129_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold349 _7148_/Q VGND VGND VPWR VPWR hold349/X sky130_fd_sc_hd__bufbuf_16
Xhold338 _5341_/X VGND VGND VPWR VPWR _6924_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_144_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6201_ _6875_/Q _6023_/C _6025_/B _6899_/Q _6200_/X VGND VGND VPWR VPWR _6206_/B
+ sky130_fd_sc_hd__a221o_1
Xhold327 hold18/X VGND VGND VPWR VPWR hold327/X sky130_fd_sc_hd__bufbuf_16
X_3413_ input59/X _4025_/A _3368_/Y input18/X _3412_/X VGND VGND VPWR VPWR _3414_/D
+ sky130_fd_sc_hd__a221o_1
X_4393_ _5031_/A _4663_/A VGND VGND VPWR VPWR _4772_/A sky130_fd_sc_hd__nor2_8
XFILLER_131_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7181_ _7193_/CLK _7181_/D fanout435/X VGND VGND VPWR VPWR _7181_/Q sky130_fd_sc_hd__dfrtp_4
X_6132_ _6306_/A _6132_/B _6132_/C _6132_/D VGND VGND VPWR VPWR _6132_/X sky130_fd_sc_hd__or4_4
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3344_ _3476_/A _5252_/B VGND VGND VPWR VPWR _3344_/Y sky130_fd_sc_hd__nor2_8
XFILLER_98_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1005 _6491_/Q VGND VGND VPWR VPWR _3986_/A0 sky130_fd_sc_hd__bufbuf_16
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ _3314_/A _3275_/B _3275_/C VGND VGND VPWR VPWR hold53/A sky130_fd_sc_hd__or3_4
X_6063_ _7078_/Q _6311_/B VGND VGND VPWR VPWR _6063_/X sky130_fd_sc_hd__and2_1
X_5014_ _4561_/Y _4758_/B _4725_/A _4839_/X VGND VGND VPWR VPWR _5016_/C sky130_fd_sc_hd__a211o_2
XFILLER_100_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1038 _6498_/Q VGND VGND VPWR VPWR _3998_/A0 sky130_fd_sc_hd__bufbuf_16
Xhold1027 _5203_/X VGND VGND VPWR VPWR _6807_/D sky130_fd_sc_hd__bufbuf_16
Xhold1016 _6499_/Q VGND VGND VPWR VPWR _3999_/A0 sky130_fd_sc_hd__bufbuf_16
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1049 _4060_/X VGND VGND VPWR VPWR _6544_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_26_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6965_ _7054_/CLK _6965_/D fanout445/X VGND VGND VPWR VPWR _6965_/Q sky130_fd_sc_hd__dfstp_4
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5916_ _6531_/Q _5722_/B _5915_/X _6308_/S VGND VGND VPWR VPWR _5916_/X sky130_fd_sc_hd__o211a_1
XFILLER_179_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6896_ _6987_/CLK _6896_/D fanout450/X VGND VGND VPWR VPWR _6896_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5847_ _7043_/Q _5683_/X _5702_/X _6891_/Q VGND VGND VPWR VPWR _5847_/X sky130_fd_sc_hd__a22o_1
X_5778_ _6912_/Q _5680_/X _5700_/X _6864_/Q _5768_/X VGND VGND VPWR VPWR _5778_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4729_ _4740_/A _4819_/A _4729_/C VGND VGND VPWR VPWR _4729_/X sky130_fd_sc_hd__and3_1
XFILLER_175_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold850 _5374_/X VGND VGND VPWR VPWR _6953_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_89_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold872 _6727_/Q VGND VGND VPWR VPWR hold872/X sky130_fd_sc_hd__bufbuf_16
Xhold861 _6647_/Q VGND VGND VPWR VPWR hold861/X sky130_fd_sc_hd__bufbuf_16
Xhold883 hold883/A VGND VGND VPWR VPWR hold883/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold894 _4057_/X VGND VGND VPWR VPWR _6541_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_88_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6750_ _7225_/CLK _6750_/D fanout419/X VGND VGND VPWR VPWR _6750_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_35_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5701_ _5864_/B _5702_/B _5701_/C VGND VGND VPWR VPWR _5701_/X sky130_fd_sc_hd__and3_4
X_3962_ _3962_/A VGND VGND VPWR VPWR _3962_/Y sky130_fd_sc_hd__inv_2
X_3893_ _3893_/A _3893_/B input120/X input117/X VGND VGND VPWR VPWR _3894_/D sky130_fd_sc_hd__or4bb_1
X_6681_ _6845_/CLK _6681_/D _6455_/A VGND VGND VPWR VPWR _6681_/Q sky130_fd_sc_hd__dfrtp_2
X_5632_ _7164_/Q _7163_/Q VGND VGND VPWR VPWR _5703_/B sky130_fd_sc_hd__nor2_8
X_5563_ _5599_/A0 hold833/X _5566_/S VGND VGND VPWR VPWR _5563_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4514_ _4671_/A _4995_/A VGND VGND VPWR VPWR _5079_/A sky130_fd_sc_hd__nor2_1
XFILLER_8_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5494_ _5602_/A0 hold363/X _5494_/S VGND VGND VPWR VPWR _5494_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold102 _5386_/X VGND VGND VPWR VPWR _6964_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_144_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold135 hold70/X VGND VGND VPWR VPWR hold135/X sky130_fd_sc_hd__bufbuf_16
Xhold124 _3284_/X VGND VGND VPWR VPWR _3419_/A sky130_fd_sc_hd__bufbuf_16
Xhold113 _3264_/X VGND VGND VPWR VPWR hold113/X sky130_fd_sc_hd__bufbuf_16
X_4445_ _4818_/A _4672_/A _4469_/A _4395_/D _5050_/A VGND VGND VPWR VPWR _4445_/X
+ sky130_fd_sc_hd__o2111a_2
Xhold168 hold202/X VGND VGND VPWR VPWR hold183/A sky130_fd_sc_hd__bufbuf_16
XFILLER_105_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold157 _7079_/Q VGND VGND VPWR VPWR hold157/X sky130_fd_sc_hd__bufbuf_16
Xhold146 _3293_/B VGND VGND VPWR VPWR _3275_/B sky130_fd_sc_hd__bufbuf_16
XFILLER_144_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7164_ _3949_/A1 _7164_/D fanout455/X VGND VGND VPWR VPWR _7164_/Q sky130_fd_sc_hd__dfrtp_2
X_4376_ _4996_/A VGND VGND VPWR VPWR _4376_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold179 _5222_/X VGND VGND VPWR VPWR _6823_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_112_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6115_ _7024_/Q _6010_/Y _6031_/X _7088_/Q _6112_/X VGND VGND VPWR VPWR _6121_/A
+ sky130_fd_sc_hd__a221o_1
X_3327_ _3457_/A _5225_/B VGND VGND VPWR VPWR _5387_/A sky130_fd_sc_hd__nor2_8
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7095_ _7097_/CLK _7095_/D fanout437/X VGND VGND VPWR VPWR _7095_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_58_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ _6941_/Q _6022_/B _6033_/X _7005_/Q VGND VGND VPWR VPWR _6046_/X sky130_fd_sc_hd__a22o_1
XFILLER_100_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ hold192/X _6784_/Q _3991_/S VGND VGND VPWR VPWR _3258_/X sky130_fd_sc_hd__mux2_4
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6948_ _7140_/CLK _6948_/D fanout430/X VGND VGND VPWR VPWR _6948_/Q sky130_fd_sc_hd__dfrtp_2
X_6879_ _7150_/CLK _6879_/D fanout449/X VGND VGND VPWR VPWR _6879_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold680 _6822_/Q VGND VGND VPWR VPWR hold680/X sky130_fd_sc_hd__bufbuf_16
XFILLER_103_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold691 _7026_/Q VGND VGND VPWR VPWR hold691/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput207 _3236_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[4] sky130_fd_sc_hd__buf_8
Xoutput229 _6514_/Q VGND VGND VPWR VPWR mgmt_gpio_out[24] sky130_fd_sc_hd__buf_8
Xoutput218 _3949_/X VGND VGND VPWR VPWR mgmt_gpio_out[14] sky130_fd_sc_hd__clkbuf_4
XFILLER_141_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4230_ hold700/X _5582_/A0 _4234_/S VGND VGND VPWR VPWR _4230_/X sky130_fd_sc_hd__mux2_1
X_4161_ _5289_/A0 _4161_/A1 _4165_/S VGND VGND VPWR VPWR _4161_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4092_ _6571_/Q _3606_/X _4096_/S VGND VGND VPWR VPWR _6571_/D sky130_fd_sc_hd__mux2_1
XFILLER_36_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6802_ _6804_/CLK _6802_/D _6439_/A VGND VGND VPWR VPWR _6802_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_168_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4994_ _4399_/Y _4539_/D _4586_/B _4987_/X VGND VGND VPWR VPWR _5000_/C sky130_fd_sc_hd__o31a_1
X_6733_ _7121_/CLK _6733_/D _6421_/A VGND VGND VPWR VPWR _6733_/Q sky130_fd_sc_hd__dfrtp_2
X_3945_ _6681_/Q input3/X input1/X VGND VGND VPWR VPWR _3945_/X sky130_fd_sc_hd__mux2_8
XFILLER_51_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6664_ _3545_/A1 _6664_/D _6443_/X VGND VGND VPWR VPWR _6664_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_176_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3876_ _6459_/Q _3875_/X _3876_/S VGND VGND VPWR VPWR _6459_/D sky130_fd_sc_hd__mux2_1
X_5615_ _7157_/Q _7158_/Q _7159_/Q _5615_/D VGND VGND VPWR VPWR _5616_/A sky130_fd_sc_hd__and4_2
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6595_ _6840_/CLK _6595_/D fanout424/X VGND VGND VPWR VPWR _6595_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5546_ hold78/X hold119/X hold22/X VGND VGND VPWR VPWR _5546_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5477_ _5477_/A _5576_/B VGND VGND VPWR VPWR _5485_/S sky130_fd_sc_hd__and2_4
X_7216_ _3949_/A1 _7216_/D fanout458/X VGND VGND VPWR VPWR _7216_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_160_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4428_ _4711_/A _5165_/A _4428_/C VGND VGND VPWR VPWR _5140_/A sky130_fd_sc_hd__and3_2
XFILLER_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout401 hold885/X VGND VGND VPWR VPWR _5541_/A0 sky130_fd_sc_hd__buf_8
Xfanout412 _6421_/B VGND VGND VPWR VPWR _6454_/B sky130_fd_sc_hd__buf_8
Xfanout423 fanout456/X VGND VGND VPWR VPWR fanout423/X sky130_fd_sc_hd__buf_8
X_4359_ _4672_/A _4818_/A VGND VGND VPWR VPWR _4558_/B sky130_fd_sc_hd__nand2b_4
X_7147_ _7154_/CLK _7147_/D fanout451/X VGND VGND VPWR VPWR _7147_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout445 fanout455/X VGND VGND VPWR VPWR fanout445/X sky130_fd_sc_hd__buf_8
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout456 input75/X VGND VGND VPWR VPWR fanout456/X sky130_fd_sc_hd__buf_8
Xfanout434 fanout435/X VGND VGND VPWR VPWR fanout434/X sky130_fd_sc_hd__buf_8
XFILLER_48_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7078_ _7078_/CLK _7078_/D fanout430/X VGND VGND VPWR VPWR _7078_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6029_ _6037_/C _6035_/C _6032_/C VGND VGND VPWR VPWR _6029_/X sky130_fd_sc_hd__and3_4
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_361 hold335/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_350 hold209/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_383 _5251_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_394 _6022_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_372 _3980_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3730_ _6474_/Q _6459_/Q _6824_/Q VGND VGND VPWR VPWR _3730_/X sky130_fd_sc_hd__or3_4
XFILLER_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3661_ _3476_/A _3543_/B _4049_/A _6537_/Q VGND VGND VPWR VPWR _3663_/C sky130_fd_sc_hd__a2bb2o_1
X_6380_ _6707_/Q _6380_/A2 _6380_/B1 _6706_/Q VGND VGND VPWR VPWR _6380_/X sky130_fd_sc_hd__a22o_1
X_5400_ hold782/X _5571_/A0 _5404_/S VGND VGND VPWR VPWR _5400_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3592_ _6788_/Q _5185_/A _5194_/A _6803_/Q _3556_/X VGND VGND VPWR VPWR _3593_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_173_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5331_ _5601_/A0 hold585/X _5332_/S VGND VGND VPWR VPWR _5331_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7001_ _7150_/CLK _7001_/D fanout446/X VGND VGND VPWR VPWR _7001_/Q sky130_fd_sc_hd__dfrtp_2
X_5262_ _5262_/A0 _5541_/A0 _5269_/S VGND VGND VPWR VPWR _6853_/D sky130_fd_sc_hd__mux2_1
X_4213_ _4247_/A1 hold78/X _4217_/S VGND VGND VPWR VPWR _4213_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5193_ _5254_/A0 hold927/X _5193_/S VGND VGND VPWR VPWR _6799_/D sky130_fd_sc_hd__mux2_1
X_4144_ _5587_/A0 _4144_/A1 _4147_/S VGND VGND VPWR VPWR _4144_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4075_ _6556_/Q _3727_/X _4081_/S VGND VGND VPWR VPWR _6556_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_3_4_0_csclk clkbuf_3_5_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_4_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_83_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4977_ _5132_/A _5142_/B _5069_/D _4977_/D VGND VGND VPWR VPWR _4977_/X sky130_fd_sc_hd__or4_2
X_6716_ _6717_/CLK _6716_/D fanout426/X VGND VGND VPWR VPWR _6716_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3928_ _3928_/A _3928_/B VGND VGND VPWR VPWR _6458_/D sky130_fd_sc_hd__and2_1
XFILLER_192_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6647_ _6744_/CLK _6647_/D fanout427/X VGND VGND VPWR VPWR _6647_/Q sky130_fd_sc_hd__dfrtp_2
X_3859_ _6666_/Q _3859_/B VGND VGND VPWR VPWR _3874_/S sky130_fd_sc_hd__nand2_8
XFILLER_165_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6578_ _6717_/CLK _6578_/D fanout426/X VGND VGND VPWR VPWR _6578_/Q sky130_fd_sc_hd__dfstp_4
X_5529_ _5583_/A0 hold647/X hold55/X VGND VGND VPWR VPWR _5529_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4900_ _4947_/B _4898_/B _4591_/B VGND VGND VPWR VPWR _5075_/B sky130_fd_sc_hd__a21oi_1
X_5880_ _6728_/Q _5667_/X _5879_/X VGND VGND VPWR VPWR _5883_/C sky130_fd_sc_hd__a21o_1
XFILLER_92_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4831_ _4707_/B _4746_/B _4728_/X _4886_/B VGND VGND VPWR VPWR _4832_/D sky130_fd_sc_hd__o211a_1
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_180 _6030_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_191 _6404_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4762_ _4949_/B _4537_/X _4565_/Y _4759_/Y VGND VGND VPWR VPWR _4763_/D sky130_fd_sc_hd__a31o_2
X_4693_ _4774_/C _4693_/B VGND VGND VPWR VPWR _4711_/C sky130_fd_sc_hd__and2_4
X_6501_ _6759_/CLK _6501_/D fanout419/X VGND VGND VPWR VPWR _6501_/Q sky130_fd_sc_hd__dfstp_4
X_3713_ _6759_/Q _4310_/A _5191_/A _6799_/Q VGND VGND VPWR VPWR _3713_/X sky130_fd_sc_hd__a22o_4
XFILLER_174_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6432_ _6446_/A _6446_/B VGND VGND VPWR VPWR _6432_/X sky130_fd_sc_hd__and2_1
X_3644_ _7023_/Q _5450_/A _4274_/A _6730_/Q _3643_/X VGND VGND VPWR VPWR _3645_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3575_ _6888_/Q _5297_/A _5405_/A _6984_/Q _3574_/X VGND VGND VPWR VPWR _3578_/C
+ sky130_fd_sc_hd__a221o_4
XFILLER_136_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6363_ _7203_/Q _3794_/X _6370_/S VGND VGND VPWR VPWR _7203_/D sky130_fd_sc_hd__mux2_1
X_5314_ _5602_/A0 hold386/X _5314_/S VGND VGND VPWR VPWR _5314_/X sky130_fd_sc_hd__mux2_1
X_6294_ _6656_/Q _6311_/B _6289_/X _6291_/X _6293_/X VGND VGND VPWR VPWR _6294_/X
+ sky130_fd_sc_hd__a2111o_1
X_5245_ _5245_/A _5594_/B VGND VGND VPWR VPWR _5251_/S sky130_fd_sc_hd__nand2_8
XFILLER_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold28 hold28/A VGND VGND VPWR VPWR hold28/X sky130_fd_sc_hd__bufbuf_16
Xhold17 hold17/A VGND VGND VPWR VPWR hold17/X sky130_fd_sc_hd__bufbuf_16
Xhold39 hold39/A VGND VGND VPWR VPWR hold39/X sky130_fd_sc_hd__bufbuf_16
X_5176_ _4947_/B _4757_/B _5050_/C _4717_/B _4837_/X VGND VGND VPWR VPWR _5177_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4127_ _4127_/A0 _5588_/A0 _4129_/S VGND VGND VPWR VPWR _6601_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4058_ _5588_/A0 _4058_/A1 _4060_/S VGND VGND VPWR VPWR _6542_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A VGND VGND VPWR VPWR _7209_/CLK sky130_fd_sc_hd__clkbuf_8
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold509 _6516_/Q VGND VGND VPWR VPWR hold509/X sky130_fd_sc_hd__bufbuf_16
XFILLER_171_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3360_ _7132_/Q _5567_/A _3359_/Y _7020_/Q VGND VGND VPWR VPWR _3360_/X sky130_fd_sc_hd__a22o_1
XFILLER_124_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5030_ _4500_/A _4758_/A _5004_/A _5099_/C _4932_/A VGND VGND VPWR VPWR _5034_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_112_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3291_ _3514_/A hold84/X VGND VGND VPWR VPWR _5477_/A sky130_fd_sc_hd__nor2_8
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1209 _6839_/Q VGND VGND VPWR VPWR _5246_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_66_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6981_ _7141_/CLK _6981_/D fanout447/X VGND VGND VPWR VPWR _6981_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_93_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5932_ _6656_/Q _5693_/X _5707_/X _6760_/Q _5931_/X VGND VGND VPWR VPWR _5937_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_15_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5863_ _6996_/Q _5684_/X _5703_/X _6876_/Q _5862_/X VGND VGND VPWR VPWR _5871_/A
+ sky130_fd_sc_hd__a221o_1
X_4814_ _5095_/A _4950_/B _4814_/C _4812_/X VGND VGND VPWR VPWR _4817_/B sky130_fd_sc_hd__or4b_1
X_5794_ _7081_/Q _5693_/X _5703_/X _6873_/Q VGND VGND VPWR VPWR _5794_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4745_ _4745_/A _4745_/B VGND VGND VPWR VPWR _4745_/X sky130_fd_sc_hd__or2_1
XFILLER_147_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4676_ _4685_/A _5062_/B _4696_/B VGND VGND VPWR VPWR _4832_/C sky130_fd_sc_hd__or3b_4
XFILLER_174_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6415_ _6421_/A _6421_/B VGND VGND VPWR VPWR _6415_/X sky130_fd_sc_hd__and2_1
X_3627_ _6983_/Q _5405_/A _4256_/A _6715_/Q _3616_/X VGND VGND VPWR VPWR _3629_/C
+ sky130_fd_sc_hd__a221o_1
X_6346_ _6747_/Q _6023_/A _6033_/X _6742_/Q _6345_/X VGND VGND VPWR VPWR _6356_/C
+ sky130_fd_sc_hd__a221o_2
X_3558_ _7088_/Q hold54/A _4043_/A _6533_/Q VGND VGND VPWR VPWR _3558_/X sky130_fd_sc_hd__a22o_1
XFILLER_163_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput118 wb_adr_i[27] VGND VGND VPWR VPWR _3893_/A sky130_fd_sc_hd__clkbuf_4
Xinput107 wb_adr_i[17] VGND VGND VPWR VPWR _4349_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_142_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3489_ _3540_/A _5234_/B VGND VGND VPWR VPWR _4136_/A sky130_fd_sc_hd__nor2_8
X_6277_ _6635_/Q _5653_/X _6022_/B _6610_/Q VGND VGND VPWR VPWR _6277_/X sky130_fd_sc_hd__a22o_1
Xinput129 wb_adr_i[8] VGND VGND VPWR VPWR _4351_/B sky130_fd_sc_hd__clkbuf_4
X_5228_ hold185/A _5228_/A1 _5233_/S VGND VGND VPWR VPWR _5228_/X sky130_fd_sc_hd__mux2_1
X_5159_ _4414_/B _5165_/A _4922_/A _4704_/X _5156_/B VGND VGND VPWR VPWR _5159_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_29_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_1_0_csclk clkbuf_2_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_3_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_91 _3606_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_80 _3439_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4530_ _4529_/B _4529_/C _4650_/B VGND VGND VPWR VPWR _4533_/C sky130_fd_sc_hd__a21boi_4
XFILLER_156_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold306 _4071_/X VGND VGND VPWR VPWR _6553_/D sky130_fd_sc_hd__bufbuf_16
X_4461_ _4707_/B _5050_/A VGND VGND VPWR VPWR _4719_/B sky130_fd_sc_hd__nor2_1
Xhold317 hold317/A VGND VGND VPWR VPWR hold317/X sky130_fd_sc_hd__bufbuf_16
XFILLER_116_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6200_ _6963_/Q _6022_/C _6032_/X _7059_/Q VGND VGND VPWR VPWR _6200_/X sky130_fd_sc_hd__a22o_1
Xhold328 _3342_/Y VGND VGND VPWR VPWR _3421_/C sky130_fd_sc_hd__bufbuf_16
Xhold339 _7086_/Q VGND VGND VPWR VPWR hold339/X sky130_fd_sc_hd__bufbuf_16
X_7180_ _7193_/CLK _7180_/D fanout433/X VGND VGND VPWR VPWR _7180_/Q sky130_fd_sc_hd__dfrtp_4
X_3412_ input27/X _3302_/Y _5558_/A _7123_/Q VGND VGND VPWR VPWR _3412_/X sky130_fd_sc_hd__a22o_1
X_4392_ _4469_/A _4395_/D VGND VGND VPWR VPWR _4663_/A sky130_fd_sc_hd__or2_4
X_6131_ _6131_/A _6131_/B _6131_/C _6131_/D VGND VGND VPWR VPWR _6132_/D sky130_fd_sc_hd__or4_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _3343_/A _3421_/C VGND VGND VPWR VPWR _5252_/B sky130_fd_sc_hd__or2_4
X_6062_ _7110_/Q _6027_/B _6021_/B _7150_/Q VGND VGND VPWR VPWR _6062_/X sky130_fd_sc_hd__a22o_1
XFILLER_98_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _3514_/A hold91/X VGND VGND VPWR VPWR _5432_/A sky130_fd_sc_hd__nor2_8
Xhold1006 _6543_/Q VGND VGND VPWR VPWR _4059_/A1 sky130_fd_sc_hd__bufbuf_16
X_5013_ _5013_/A _5013_/B VGND VGND VPWR VPWR _5156_/B sky130_fd_sc_hd__or2_4
XFILLER_85_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1039 _6580_/Q VGND VGND VPWR VPWR _4102_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1017 _6731_/Q VGND VGND VPWR VPWR _4278_/A1 sky130_fd_sc_hd__bufbuf_16
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1028 _6765_/Q VGND VGND VPWR VPWR _4319_/A0 sky130_fd_sc_hd__bufbuf_16
XFILLER_39_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6964_ _6964_/CLK _6964_/D fanout451/X VGND VGND VPWR VPWR _6964_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6895_ _7150_/CLK _6895_/D fanout449/X VGND VGND VPWR VPWR _6895_/Q sky130_fd_sc_hd__dfrtp_2
X_5915_ _5915_/A _5915_/B _5915_/C _5915_/D VGND VGND VPWR VPWR _5915_/X sky130_fd_sc_hd__or4_2
XFILLER_22_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5846_ _6939_/Q _5704_/X _5705_/X _6947_/Q _5845_/X VGND VGND VPWR VPWR _5849_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5777_ _5777_/A _5777_/B _5777_/C _5777_/D VGND VGND VPWR VPWR _5777_/X sky130_fd_sc_hd__or4_4
X_4728_ _4728_/A _4746_/B VGND VGND VPWR VPWR _4728_/X sky130_fd_sc_hd__or2_4
XFILLER_135_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4659_ _4659_/A _4758_/B VGND VGND VPWR VPWR _4832_/B sky130_fd_sc_hd__nand2_8
XFILLER_174_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold840 _5590_/X VGND VGND VPWR VPWR _7145_/D sky130_fd_sc_hd__bufbuf_16
Xhold851 _6889_/Q VGND VGND VPWR VPWR hold851/X sky130_fd_sc_hd__bufbuf_16
XFILLER_150_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold873 _4273_/X VGND VGND VPWR VPWR _6727_/D sky130_fd_sc_hd__bufbuf_16
Xhold862 _4182_/X VGND VGND VPWR VPWR _6647_/D sky130_fd_sc_hd__bufbuf_16
Xhold884 _3979_/X VGND VGND VPWR VPWR hold884/X sky130_fd_sc_hd__bufbuf_16
XFILLER_115_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6329_ _6538_/Q _6025_/D _6029_/X _6642_/Q _6328_/X VGND VGND VPWR VPWR _6330_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_1_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold895 _6635_/Q VGND VGND VPWR VPWR hold895/X sky130_fd_sc_hd__bufbuf_16
XFILLER_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_32_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7156_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_79_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_47_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7138_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_57_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3961_ _6473_/Q _3961_/B VGND VGND VPWR VPWR _3962_/A sky130_fd_sc_hd__or2_4
XFILLER_51_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5700_ _5864_/B _5703_/B _5707_/B VGND VGND VPWR VPWR _5700_/X sky130_fd_sc_hd__and3_4
X_3892_ _3892_/A _3892_/B input131/X input169/X VGND VGND VPWR VPWR _3894_/C sky130_fd_sc_hd__or4bb_1
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6680_ _7196_/CLK _6680_/D fanout433/X VGND VGND VPWR VPWR _6680_/Q sky130_fd_sc_hd__dfrtp_2
X_5631_ _7163_/Q _5629_/B _5635_/B _5630_/Y VGND VGND VPWR VPWR _7163_/D sky130_fd_sc_hd__a31o_1
X_5562_ _5571_/A0 hold564/X _5566_/S VGND VGND VPWR VPWR _5562_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4513_ _4513_/A _4513_/B VGND VGND VPWR VPWR _4990_/A sky130_fd_sc_hd__or2_4
X_5493_ _5601_/A0 hold597/X _5494_/S VGND VGND VPWR VPWR _5493_/X sky130_fd_sc_hd__mux2_1
Xhold103 _6481_/Q VGND VGND VPWR VPWR _3249_/B sky130_fd_sc_hd__bufbuf_16
Xhold114 _3265_/X VGND VGND VPWR VPWR _3421_/B sky130_fd_sc_hd__bufbuf_16
Xhold125 _3551_/B VGND VGND VPWR VPWR _5225_/B sky130_fd_sc_hd__bufbuf_16
X_4444_ _4958_/B _4444_/B VGND VGND VPWR VPWR _4572_/A sky130_fd_sc_hd__nand2_8
XFILLER_171_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold158 _5516_/X VGND VGND VPWR VPWR _7079_/D sky130_fd_sc_hd__bufbuf_16
Xhold147 _3260_/X VGND VGND VPWR VPWR _3506_/A sky130_fd_sc_hd__bufbuf_16
Xhold136 hold136/A VGND VGND VPWR VPWR hold136/X sky130_fd_sc_hd__bufbuf_16
X_7163_ _3949_/A1 _7163_/D fanout455/X VGND VGND VPWR VPWR _7163_/Q sky130_fd_sc_hd__dfrtp_2
X_4375_ _4553_/A _4400_/A VGND VGND VPWR VPWR _4996_/A sky130_fd_sc_hd__or2_4
Xhold169 hold184/X VGND VGND VPWR VPWR hold185/A sky130_fd_sc_hd__bufbuf_16
X_3326_ _6924_/Q _5333_/A _5324_/A _6916_/Q VGND VGND VPWR VPWR _3326_/X sky130_fd_sc_hd__a22o_1
X_6114_ _6976_/Q _6023_/B _6020_/C _6912_/Q VGND VGND VPWR VPWR _6131_/B sky130_fd_sc_hd__a22o_1
XFILLER_113_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7094_ _7135_/CLK _7094_/D fanout430/X VGND VGND VPWR VPWR _7094_/Q sky130_fd_sc_hd__dfstp_2
X_6045_ _7117_/Q _6023_/D _6034_/Y _6989_/Q _6044_/X VGND VGND VPWR VPWR _6059_/C
+ sky130_fd_sc_hd__a221o_4
XFILLER_140_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ hold191/X _3845_/A hold50/X VGND VGND VPWR VPWR _3257_/X sky130_fd_sc_hd__a21o_1
XFILLER_37_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6947_ _7107_/CLK _6947_/D fanout434/X VGND VGND VPWR VPWR _6947_/Q sky130_fd_sc_hd__dfrtp_2
X_6878_ _7121_/CLK _6878_/D _6421_/A VGND VGND VPWR VPWR _6878_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_167_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5829_ _5663_/A _7180_/Q _6358_/B1 VGND VGND VPWR VPWR _5829_/X sky130_fd_sc_hd__a21o_1
XFILLER_182_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold681 _6610_/Q VGND VGND VPWR VPWR hold681/X sky130_fd_sc_hd__bufbuf_16
XFILLER_1_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold670 _7082_/Q VGND VGND VPWR VPWR hold670/X sky130_fd_sc_hd__bufbuf_16
Xhold692 _5456_/X VGND VGND VPWR VPWR _7026_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_134_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput208 _3235_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[5] sky130_fd_sc_hd__buf_8
Xoutput219 _3948_/X VGND VGND VPWR VPWR mgmt_gpio_out[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_126_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4160_ _4160_/A _5558_/B VGND VGND VPWR VPWR _4165_/S sky130_fd_sc_hd__nand2_8
XFILLER_67_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4091_ _6570_/Q _3665_/X _4096_/S VGND VGND VPWR VPWR _6570_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6801_ _6804_/CLK _6801_/D _6439_/A VGND VGND VPWR VPWR _6801_/Q sky130_fd_sc_hd__dfrtp_2
X_4993_ _4478_/B _4992_/Y _4991_/X VGND VGND VPWR VPWR _5118_/C sky130_fd_sc_hd__o21ai_2
XFILLER_90_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6732_ _6804_/CLK _6732_/D _6439_/A VGND VGND VPWR VPWR _6732_/Q sky130_fd_sc_hd__dfrtp_2
X_3944_ _6473_/Q _3965_/B _3942_/X _3943_/Y VGND VGND VPWR VPWR _3944_/X sky130_fd_sc_hd__a22o_4
X_3875_ _6486_/Q _3875_/B VGND VGND VPWR VPWR _3875_/X sky130_fd_sc_hd__and2b_1
X_6663_ _6845_/CLK _6663_/D _6439_/A VGND VGND VPWR VPWR _6663_/Q sky130_fd_sc_hd__dfrtp_2
X_5614_ _7157_/Q _7158_/Q _5615_/D _7159_/Q VGND VGND VPWR VPWR _5617_/B sky130_fd_sc_hd__a31o_1
XFILLER_176_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6594_ _6840_/CLK _6594_/D fanout424/X VGND VGND VPWR VPWR _6594_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_117_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5545_ _5545_/A0 _5545_/A1 hold22/X VGND VGND VPWR VPWR _5545_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5476_ _5584_/A0 hold423/X _5476_/S VGND VGND VPWR VPWR _5476_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_0_0_csclk clkbuf_3_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_0_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
X_7215_ _3949_/A1 _7215_/D fanout458/X VGND VGND VPWR VPWR _7215_/Q sky130_fd_sc_hd__dfrtp_2
X_4427_ _5165_/A _4428_/C VGND VGND VPWR VPWR _5023_/B sky130_fd_sc_hd__nand2_2
Xfanout402 hold885/X VGND VGND VPWR VPWR _5595_/A0 sky130_fd_sc_hd__buf_8
X_7146_ _7154_/CLK _7146_/D fanout452/X VGND VGND VPWR VPWR _7146_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout413 _3877_/Y VGND VGND VPWR VPWR _6421_/B sky130_fd_sc_hd__buf_8
XFILLER_171_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout446 fanout449/X VGND VGND VPWR VPWR fanout446/X sky130_fd_sc_hd__buf_8
X_4358_ _4553_/A _4774_/A _4484_/B VGND VGND VPWR VPWR _4478_/B sky130_fd_sc_hd__or3b_4
XFILLER_101_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout457 fanout458/X VGND VGND VPWR VPWR _6362_/B sky130_fd_sc_hd__buf_8
Xfanout435 fanout456/X VGND VGND VPWR VPWR fanout435/X sky130_fd_sc_hd__buf_8
Xfanout424 _6454_/A VGND VGND VPWR VPWR fanout424/X sky130_fd_sc_hd__buf_8
X_7077_ _7124_/CLK _7077_/D fanout436/X VGND VGND VPWR VPWR _7077_/Q sky130_fd_sc_hd__dfstp_4
X_4289_ _6409_/A0 _4289_/A1 _4291_/S VGND VGND VPWR VPWR _6740_/D sky130_fd_sc_hd__mux2_1
X_3309_ _3309_/A hold52/X _3293_/B VGND VGND VPWR VPWR _3309_/X sky130_fd_sc_hd__or3b_4
X_6028_ _6037_/C _6033_/C _6035_/C VGND VGND VPWR VPWR _6028_/X sky130_fd_sc_hd__and3_4
XFILLER_100_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_340 hold78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_351 hold209/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_362 hold335/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_395 _6025_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_384 _5658_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_373 _5192_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3660_ _6750_/Q _4298_/A _4184_/A _6651_/Q _3659_/X VGND VGND VPWR VPWR _3663_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_186_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3591_ _6657_/Q _4190_/A _6406_/A _7224_/Q _3565_/X VGND VGND VPWR VPWR _3593_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_142_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5330_ _5600_/A0 hold449/X _5332_/S VGND VGND VPWR VPWR _5330_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5261_ _5261_/A _5576_/B VGND VGND VPWR VPWR _5269_/S sky130_fd_sc_hd__and2_4
X_4212_ _4212_/A0 hold459/X _4218_/S VGND VGND VPWR VPWR _4212_/X sky130_fd_sc_hd__mux2_1
X_7000_ _7152_/CLK _7000_/D fanout452/X VGND VGND VPWR VPWR _7000_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_142_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5192_ _5234_/C _5192_/A1 _5193_/S VGND VGND VPWR VPWR _5192_/X sky130_fd_sc_hd__mux2_1
X_4143_ _5289_/A0 _4143_/A1 _4147_/S VGND VGND VPWR VPWR _4143_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4074_ _6555_/Q _3794_/X _4081_/S VGND VGND VPWR VPWR _6555_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4976_ _4976_/A _4976_/B _4976_/C _4638_/X VGND VGND VPWR VPWR _4977_/D sky130_fd_sc_hd__or4b_1
X_6715_ _6715_/CLK _6715_/D fanout439/X VGND VGND VPWR VPWR _6715_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_137_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3927_ _6665_/Q _6668_/Q _3196_/Y VGND VGND VPWR VPWR _3928_/B sky130_fd_sc_hd__o21ai_1
XFILLER_192_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6646_ _7103_/CLK _6646_/D fanout436/X VGND VGND VPWR VPWR _6646_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_20_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3858_ _3864_/B VGND VGND VPWR VPWR _3858_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6577_ _6840_/CLK _6577_/D fanout424/X VGND VGND VPWR VPWR _6577_/Q sky130_fd_sc_hd__dfrtp_2
X_3789_ input93/X _3280_/Y _3308_/Y _4274_/A _6728_/Q VGND VGND VPWR VPWR _3789_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_192_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5528_ _5582_/A0 hold667/X hold55/X VGND VGND VPWR VPWR _5528_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5459_ _5459_/A _5576_/B VGND VGND VPWR VPWR _5467_/S sky130_fd_sc_hd__nand2_8
XFILLER_182_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7129_ _7129_/CLK _7129_/D fanout429/X VGND VGND VPWR VPWR _7129_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_87_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4830_ _4672_/B _4737_/Y _4829_/X _4758_/B VGND VGND VPWR VPWR _4834_/C sky130_fd_sc_hd__o31a_1
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_170 _6021_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_181 _6030_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_192 debug_mode VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4761_ _5062_/A _4832_/A VGND VGND VPWR VPWR _5073_/B sky130_fd_sc_hd__nor2_1
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4692_ _4711_/A _4758_/A _4758_/B VGND VGND VPWR VPWR _5035_/A sky130_fd_sc_hd__and3_2
XFILLER_119_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6500_ _6759_/CLK _6500_/D fanout419/X VGND VGND VPWR VPWR _6500_/Q sky130_fd_sc_hd__dfstp_4
X_3712_ _7110_/Q hold85/A _5200_/A _6806_/Q _3711_/X VGND VGND VPWR VPWR _3717_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6431_ _6446_/A _6446_/B VGND VGND VPWR VPWR _6431_/X sky130_fd_sc_hd__and2_1
X_3643_ input26/X _3283_/Y _4190_/A _6656_/Q VGND VGND VPWR VPWR _3643_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6362_ _6704_/D _6362_/B VGND VGND VPWR VPWR _6370_/S sky130_fd_sc_hd__and2_4
X_3574_ _7152_/Q _5594_/A _5558_/A _7120_/Q VGND VGND VPWR VPWR _3574_/X sky130_fd_sc_hd__a22o_1
X_5313_ _5601_/A0 hold659/X _5314_/S VGND VGND VPWR VPWR _5313_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6293_ _6626_/Q _6028_/X _6034_/Y _6725_/Q _6292_/X VGND VGND VPWR VPWR _6293_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_114_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5244_ _5254_/A0 hold936/X _5244_/S VGND VGND VPWR VPWR _5244_/X sky130_fd_sc_hd__mux2_1
X_5175_ _5175_/A _5175_/B _5175_/C _5175_/D VGND VGND VPWR VPWR _5175_/X sky130_fd_sc_hd__or4_1
Xhold29 hold29/A VGND VGND VPWR VPWR hold29/X sky130_fd_sc_hd__bufbuf_16
XFILLER_68_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold18 hold18/A VGND VGND VPWR VPWR hold18/X sky130_fd_sc_hd__bufbuf_16
X_4126_ hold531/X _5587_/A0 _4129_/S VGND VGND VPWR VPWR _4126_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4057_ _5254_/A0 hold893/X _4060_/S VGND VGND VPWR VPWR _4057_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4959_ _4959_/A _4959_/B VGND VGND VPWR VPWR _4959_/X sky130_fd_sc_hd__and2_4
XFILLER_177_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6629_ _6629_/CLK _6629_/D fanout456/X VGND VGND VPWR VPWR _6629_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_137_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3290_ hold83/X _3343_/A VGND VGND VPWR VPWR hold84/A sky130_fd_sc_hd__or2_4
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6980_ _7122_/CLK _6980_/D fanout443/X VGND VGND VPWR VPWR _6980_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_38_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5931_ _6542_/Q _5703_/X _5930_/X _5698_/B VGND VGND VPWR VPWR _5931_/X sky130_fd_sc_hd__a22o_4
XFILLER_53_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5862_ _7068_/Q _5669_/X _5692_/X _7076_/Q VGND VGND VPWR VPWR _5862_/X sky130_fd_sc_hd__a22o_1
X_4813_ _4395_/D _4470_/B _4656_/X _4494_/Y VGND VGND VPWR VPWR _4814_/C sky130_fd_sc_hd__a31o_1
X_5793_ _7001_/Q _5667_/X _5792_/X VGND VGND VPWR VPWR _5796_/C sky130_fd_sc_hd__a21o_1
X_4744_ _4672_/A _4566_/A _4745_/B _4742_/X _4743_/X VGND VGND VPWR VPWR _4753_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_178_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4675_ _4719_/B _4758_/B _4696_/B VGND VGND VPWR VPWR _4748_/B sky130_fd_sc_hd__and3_4
XFILLER_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3626_ _6919_/Q _5333_/A _4061_/A _6547_/Q _3615_/X VGND VGND VPWR VPWR _3629_/B
+ sky130_fd_sc_hd__a221o_1
X_6414_ _6446_/A _6446_/B VGND VGND VPWR VPWR _6414_/X sky130_fd_sc_hd__and2_1
XFILLER_115_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6345_ _6554_/Q _6020_/A _6021_/D _6633_/Q _6344_/X VGND VGND VPWR VPWR _6345_/X
+ sky130_fd_sc_hd__a221o_2
X_3557_ _7048_/Q _5477_/A _4172_/A _6642_/Q VGND VGND VPWR VPWR _3557_/X sky130_fd_sc_hd__a22o_1
XFILLER_163_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6276_ _6541_/Q _6023_/C _6025_/B _6564_/Q _6275_/X VGND VGND VPWR VPWR _6281_/B
+ sky130_fd_sc_hd__a221o_2
Xinput108 wb_adr_i[18] VGND VGND VPWR VPWR _4349_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_130_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3488_ _3488_/A _3488_/B _3488_/C _3488_/D VGND VGND VPWR VPWR _3548_/B sky130_fd_sc_hd__or4_2
X_5227_ _5227_/A _5576_/B VGND VGND VPWR VPWR _5233_/S sky130_fd_sc_hd__nand2_8
Xinput119 wb_adr_i[28] VGND VGND VPWR VPWR _3893_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_130_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5158_ _5158_/A _5158_/B VGND VGND VPWR VPWR _5158_/Y sky130_fd_sc_hd__nor2_2
XFILLER_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5089_ _4871_/A _4749_/C _4953_/A VGND VGND VPWR VPWR _5118_/D sky130_fd_sc_hd__a21oi_1
X_4109_ _6586_/Q _3452_/X _4111_/S VGND VGND VPWR VPWR _6586_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_70 _5558_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_81 _3488_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_92 _3606_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4460_ _4694_/A _4989_/A VGND VGND VPWR VPWR _5003_/A sky130_fd_sc_hd__or2_4
Xhold307 _7075_/Q VGND VGND VPWR VPWR hold307/X sky130_fd_sc_hd__bufbuf_16
Xhold318 _4243_/X VGND VGND VPWR VPWR _6691_/D sky130_fd_sc_hd__bufbuf_16
X_4391_ _4513_/A _4405_/B VGND VGND VPWR VPWR _4988_/A sky130_fd_sc_hd__or2_4
Xhold329 _3473_/B VGND VGND VPWR VPWR _3528_/B sky130_fd_sc_hd__bufbuf_16
X_3411_ _6995_/Q _3299_/Y _3978_/A _6494_/Q _3388_/X VGND VGND VPWR VPWR _3414_/C
+ sky130_fd_sc_hd__a221o_1
X_6130_ _6864_/Q _6025_/D _6029_/X _7048_/Q _6129_/X VGND VGND VPWR VPWR _6131_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3342_ hold327/X hold82/X VGND VGND VPWR VPWR _3342_/Y sky130_fd_sc_hd__nand2b_4
XFILLER_140_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3273_ hold90/X hold19/X VGND VGND VPWR VPWR hold91/A sky130_fd_sc_hd__or2_4
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _5663_/Y _6059_/X _6060_/X _6358_/B1 _7189_/Q VGND VGND VPWR VPWR _7189_/D
+ sky130_fd_sc_hd__a32o_1
X_5012_ _5012_/A _5105_/B _5011_/X VGND VGND VPWR VPWR _5016_/A sky130_fd_sc_hd__or3b_1
Xhold1029 _6885_/Q VGND VGND VPWR VPWR _5298_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1018 _4278_/X VGND VGND VPWR VPWR _6731_/D sky130_fd_sc_hd__bufbuf_16
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1007 _4059_/X VGND VGND VPWR VPWR _6543_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6963_ _7122_/CLK _6963_/D fanout443/X VGND VGND VPWR VPWR _6963_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6894_ _7153_/CLK _6894_/D _6421_/A VGND VGND VPWR VPWR _6894_/Q sky130_fd_sc_hd__dfstp_4
X_5914_ _6786_/Q _5690_/X _5693_/X _6655_/Q _5913_/X VGND VGND VPWR VPWR _5915_/D
+ sky130_fd_sc_hd__a221o_1
X_5845_ _7011_/Q _5678_/X _5682_/X _7019_/Q VGND VGND VPWR VPWR _5845_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5776_ _6976_/Q _5676_/X _5702_/X _6888_/Q _5775_/X VGND VGND VPWR VPWR _5777_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4727_ _4663_/A _4729_/C _4725_/A VGND VGND VPWR VPWR _4727_/Y sky130_fd_sc_hd__a21oi_1
X_4658_ _4470_/B _4656_/X _4653_/Y _4957_/A _5135_/A VGND VGND VPWR VPWR _4708_/C
+ sky130_fd_sc_hd__a2111o_1
XFILLER_190_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput90 spimemio_flash_io2_oeb VGND VGND VPWR VPWR input90/X sky130_fd_sc_hd__clkbuf_4
Xhold830 _4116_/X VGND VGND VPWR VPWR _6592_/D sky130_fd_sc_hd__bufbuf_16
X_3609_ _5234_/A _4241_/B VGND VGND VPWR VPWR _5238_/A sky130_fd_sc_hd__nor2_8
Xhold863 _7153_/Q VGND VGND VPWR VPWR hold863/X sky130_fd_sc_hd__bufbuf_16
X_4589_ _4593_/A _4693_/B VGND VGND VPWR VPWR _4590_/B sky130_fd_sc_hd__nand2_1
Xhold852 _5302_/X VGND VGND VPWR VPWR _6889_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_122_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold841 _6721_/Q VGND VGND VPWR VPWR hold841/X sky130_fd_sc_hd__bufbuf_16
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold874 _6675_/Q VGND VGND VPWR VPWR hold874/X sky130_fd_sc_hd__bufbuf_16
Xhold885 hold885/A VGND VGND VPWR VPWR hold885/X sky130_fd_sc_hd__bufbuf_16
XFILLER_115_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6328_ _6637_/Q _5653_/X _6022_/B _6612_/Q VGND VGND VPWR VPWR _6328_/X sky130_fd_sc_hd__a22o_1
Xhold896 _4168_/X VGND VGND VPWR VPWR _6635_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_131_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6259_ _5663_/A _7196_/Q _6358_/B1 VGND VGND VPWR VPWR _6259_/X sky130_fd_sc_hd__a21o_2
XFILLER_91_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3960_ _3960_/A VGND VGND VPWR VPWR _3960_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3891_ _4345_/A _4345_/B VGND VGND VPWR VPWR _4722_/B sky130_fd_sc_hd__or2_4
XFILLER_188_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5630_ _5633_/B VGND VGND VPWR VPWR _5630_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5561_ _5561_/A0 hold825/X _5566_/S VGND VGND VPWR VPWR _5561_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5492_ _5600_/A0 hold456/X _5494_/S VGND VGND VPWR VPWR _5492_/X sky130_fd_sc_hd__mux2_1
X_4512_ _4513_/A _4513_/B VGND VGND VPWR VPWR _4624_/B sky130_fd_sc_hd__nor2_8
XFILLER_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold104 _3253_/X VGND VGND VPWR VPWR hold104/X sky130_fd_sc_hd__bufbuf_16
Xhold115 _3292_/X VGND VGND VPWR VPWR hold27/A sky130_fd_sc_hd__bufbuf_16
Xhold126 _3341_/Y VGND VGND VPWR VPWR _5531_/A sky130_fd_sc_hd__bufbuf_16
Xhold159 _7212_/Q VGND VGND VPWR VPWR hold159/X sky130_fd_sc_hd__bufbuf_16
X_4443_ _4958_/B _4444_/B VGND VGND VPWR VPWR _4443_/X sky130_fd_sc_hd__and2_4
XFILLER_144_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold137 _5229_/X VGND VGND VPWR VPWR _6827_/D sky130_fd_sc_hd__bufbuf_16
Xhold148 _3359_/Y VGND VGND VPWR VPWR _5441_/A sky130_fd_sc_hd__bufbuf_16
X_4374_ _4507_/A _4992_/A VGND VGND VPWR VPWR _4400_/A sky130_fd_sc_hd__nand2_4
X_7162_ _3949_/A1 _7162_/D fanout443/X VGND VGND VPWR VPWR _7162_/Q sky130_fd_sc_hd__dfstp_4
X_6113_ _7064_/Q _5996_/X _6021_/C _6880_/Q VGND VGND VPWR VPWR _6131_/A sky130_fd_sc_hd__a22o_1
XFILLER_113_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3325_ _3473_/A hold20/X VGND VGND VPWR VPWR _5324_/A sky130_fd_sc_hd__nor2_8
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7093_ _7101_/CLK _7093_/D fanout430/X VGND VGND VPWR VPWR _7093_/Q sky130_fd_sc_hd__dfstp_4
X_6044_ _6917_/Q _6022_/D _6032_/X _7053_/Q VGND VGND VPWR VPWR _6044_/X sky130_fd_sc_hd__a22o_1
X_3256_ hold50/X _3845_/A hold223/X VGND VGND VPWR VPWR _3256_/Y sky130_fd_sc_hd__a21oi_4
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6946_ _7106_/CLK _6946_/D fanout438/X VGND VGND VPWR VPWR _6946_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6877_ _7150_/CLK _6877_/D fanout449/X VGND VGND VPWR VPWR _6877_/Q sky130_fd_sc_hd__dfstp_4
X_5828_ _6858_/Q _5722_/B _5826_/X _5827_/X _6308_/S VGND VGND VPWR VPWR _5828_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_10_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5759_ _6903_/Q _5689_/X _5707_/X _7023_/Q VGND VGND VPWR VPWR _5759_/X sky130_fd_sc_hd__a22o_1
XFILLER_108_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold660 _5313_/X VGND VGND VPWR VPWR _6899_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_78_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold671 _5519_/X VGND VGND VPWR VPWR _7082_/D sky130_fd_sc_hd__bufbuf_16
Xhold682 _4138_/X VGND VGND VPWR VPWR _6610_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_131_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold693 _7067_/Q VGND VGND VPWR VPWR hold693/X sky130_fd_sc_hd__bufbuf_16
XFILLER_134_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput209 _3234_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[6] sky130_fd_sc_hd__buf_8
XFILLER_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4090_ _6569_/Q _3727_/X _4096_/S VGND VGND VPWR VPWR _6569_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6800_ _6804_/CLK _6800_/D _6439_/A VGND VGND VPWR VPWR _6800_/Q sky130_fd_sc_hd__dfrtp_2
X_4992_ _4992_/A _4992_/B VGND VGND VPWR VPWR _4992_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6731_ _6804_/CLK _6731_/D _6439_/A VGND VGND VPWR VPWR _6731_/Q sky130_fd_sc_hd__dfrtp_2
X_3943_ _6475_/Q _3202_/Y _6473_/Q VGND VGND VPWR VPWR _3943_/Y sky130_fd_sc_hd__a21oi_2
X_3874_ _3875_/B hold64/A _3874_/S VGND VGND VPWR VPWR _6460_/D sky130_fd_sc_hd__mux2_1
XFILLER_149_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6662_ _6845_/CLK _6662_/D fanout417/X VGND VGND VPWR VPWR _6662_/Q sky130_fd_sc_hd__dfrtp_2
X_5613_ _3920_/Y _5610_/Y _5612_/Y _5605_/Y _7158_/Q VGND VGND VPWR VPWR _7158_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_31_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6593_ _6713_/CLK _6593_/D fanout426/X VGND VGND VPWR VPWR _6593_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_129_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5544_ hold136/X hold234/X hold22/X VGND VGND VPWR VPWR _7104_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5475_ _5583_/A0 hold643/X _5476_/S VGND VGND VPWR VPWR _5475_/X sky130_fd_sc_hd__mux2_1
X_7214_ _3949_/A1 _7214_/D fanout458/X VGND VGND VPWR VPWR _7214_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_160_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4426_ _4426_/A _4776_/A VGND VGND VPWR VPWR _4428_/C sky130_fd_sc_hd__nor2_4
XFILLER_132_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7145_ _7150_/CLK _7145_/D fanout446/X VGND VGND VPWR VPWR _7145_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout403 hold885/X VGND VGND VPWR VPWR _5289_/A0 sky130_fd_sc_hd__buf_8
Xfanout414 _6446_/A VGND VGND VPWR VPWR _6439_/A sky130_fd_sc_hd__buf_8
Xfanout447 fanout449/X VGND VGND VPWR VPWR fanout447/X sky130_fd_sc_hd__buf_8
X_4357_ _4372_/B _4372_/C VGND VGND VPWR VPWR _4484_/B sky130_fd_sc_hd__nand2_2
XFILLER_113_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout425 fanout426/X VGND VGND VPWR VPWR _6454_/A sky130_fd_sc_hd__buf_8
Xfanout436 fanout437/X VGND VGND VPWR VPWR fanout436/X sky130_fd_sc_hd__buf_8
XFILLER_101_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7076_ _7124_/CLK _7076_/D fanout438/X VGND VGND VPWR VPWR _7076_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout458 input164/X VGND VGND VPWR VPWR fanout458/X sky130_fd_sc_hd__buf_8
X_3308_ hold20/A VGND VGND VPWR VPWR _3308_/Y sky130_fd_sc_hd__inv_2
X_4288_ _6408_/A0 hold413/X _4291_/S VGND VGND VPWR VPWR _4288_/X sky130_fd_sc_hd__mux2_1
X_6027_ _6037_/C _6027_/B _6027_/C _6027_/D VGND VGND VPWR VPWR _6060_/B sky130_fd_sc_hd__or4_4
XFILLER_86_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3239_ _6856_/Q VGND VGND VPWR VPWR _3239_/Y sky130_fd_sc_hd__inv_2
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6929_ _7150_/CLK _6929_/D fanout449/X VGND VGND VPWR VPWR _6929_/Q sky130_fd_sc_hd__dfrtp_2
Xclkbuf_leaf_31_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7152_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_168_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_46_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7090_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_108_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold490 _4252_/X VGND VGND VPWR VPWR _6709_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_1_0_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_77_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1190 _5201_/X VGND VGND VPWR VPWR _6805_/D sky130_fd_sc_hd__bufbuf_16
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_341 hold78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_330 _6407_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_352 hold185/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_363 _6841_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_385 _5678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_374 _3996_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_396 _6025_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3590_ _6808_/Q _5200_/A _3551_/Y input95/X _3559_/X VGND VGND VPWR VPWR _3593_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_186_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5260_ _5584_/A0 hold429/X _5260_/S VGND VGND VPWR VPWR _5260_/X sky130_fd_sc_hd__mux2_1
X_4211_ hold458/X _5581_/A0 _4217_/S VGND VGND VPWR VPWR _4211_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5191_ _5191_/A _6406_/B VGND VGND VPWR VPWR _5193_/S sky130_fd_sc_hd__nand2_1
XFILLER_141_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4142_ _4142_/A _5558_/B VGND VGND VPWR VPWR _4147_/S sky130_fd_sc_hd__nand2_8
X_4073_ _6702_/Q _6362_/B VGND VGND VPWR VPWR _4081_/S sky130_fd_sc_hd__and2_4
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4975_ _5075_/A _5075_/C _4975_/C VGND VGND VPWR VPWR _4976_/B sky130_fd_sc_hd__or3_1
X_6714_ _6717_/CLK _6714_/D fanout426/X VGND VGND VPWR VPWR _6714_/Q sky130_fd_sc_hd__dfrtp_2
X_3926_ _3196_/Y _3898_/Y _3843_/B _6667_/Q VGND VGND VPWR VPWR _6666_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_165_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6645_ _7105_/CLK _6645_/D fanout427/X VGND VGND VPWR VPWR _6645_/Q sky130_fd_sc_hd__dfrtp_2
X_3857_ _3841_/B _6664_/Q _3857_/C _3857_/D VGND VGND VPWR VPWR _3864_/B sky130_fd_sc_hd__and4b_4
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3788_ _7053_/Q _5486_/A _4184_/A _6649_/Q _3787_/X VGND VGND VPWR VPWR _3792_/B
+ sky130_fd_sc_hd__a221o_4
X_6576_ _6717_/CLK _6576_/D fanout426/X VGND VGND VPWR VPWR _6576_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5527_ hold185/X hold250/X hold55/X VGND VGND VPWR VPWR _5527_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5458_ _5584_/A0 hold472/X _5458_/S VGND VGND VPWR VPWR _5458_/X sky130_fd_sc_hd__mux2_1
X_5389_ _5596_/A0 hold333/X _5395_/S VGND VGND VPWR VPWR _5389_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4409_ _4513_/B _4410_/D VGND VGND VPWR VPWR _4409_/Y sky130_fd_sc_hd__nor2_4
XFILLER_87_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7128_ _7130_/CLK _7128_/D fanout454/X VGND VGND VPWR VPWR _7128_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7059_ _7154_/CLK _7059_/D fanout451/X VGND VGND VPWR VPWR _7059_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_160 _5861_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_171 _6021_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_193 debug_oeb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_182 _6311_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4760_ _4947_/B _4832_/A VGND VGND VPWR VPWR _5047_/B sky130_fd_sc_hd__nor2_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4691_ _4746_/B _4707_/B _5050_/A VGND VGND VPWR VPWR _4756_/B sky130_fd_sc_hd__or3b_4
X_3711_ input53/X _4025_/A _4217_/S input44/X VGND VGND VPWR VPWR _3711_/X sky130_fd_sc_hd__a22o_4
XFILLER_147_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6430_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6430_/X sky130_fd_sc_hd__and2_1
X_3642_ _7055_/Q _5486_/A _5227_/A _6828_/Q _3641_/X VGND VGND VPWR VPWR _3645_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6361_ _7202_/Q _3896_/Y _6360_/Y _3916_/B _6704_/D VGND VGND VPWR VPWR _7202_/D
+ sky130_fd_sc_hd__a32o_1
X_5312_ _5600_/A0 hold552/X _5314_/S VGND VGND VPWR VPWR _5312_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3573_ _6960_/Q _5378_/A _3552_/Y _6823_/Q _3572_/X VGND VGND VPWR VPWR _3578_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_114_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6292_ _7223_/Q _6009_/X _6020_/D _6710_/Q VGND VGND VPWR VPWR _6292_/X sky130_fd_sc_hd__a22o_2
XFILLER_142_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5243_ _5234_/C _5243_/A1 _5244_/S VGND VGND VPWR VPWR _5243_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5174_ _5174_/A _5174_/B _5174_/C _5174_/D VGND VGND VPWR VPWR _5175_/D sky130_fd_sc_hd__or4_2
Xhold19 hold19/A VGND VGND VPWR VPWR hold19/X sky130_fd_sc_hd__bufbuf_16
X_4125_ _4125_/A0 _5289_/A0 _4129_/S VGND VGND VPWR VPWR _4125_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4056_ _5289_/A0 _4056_/A1 _4060_/S VGND VGND VPWR VPWR _4056_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4958_ _4958_/A _4958_/B VGND VGND VPWR VPWR _4959_/B sky130_fd_sc_hd__nor2_4
XFILLER_184_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4889_ _5005_/C _4832_/A _4575_/Y VGND VGND VPWR VPWR _5073_/C sky130_fd_sc_hd__o21ai_2
X_3909_ _5663_/A _3921_/B VGND VGND VPWR VPWR _3909_/Y sky130_fd_sc_hd__nand2_1
X_6628_ _6725_/CLK _6628_/D fanout440/X VGND VGND VPWR VPWR _6628_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_137_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6559_ _7209_/CLK _6559_/D VGND VGND VPWR VPWR _6559_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_193_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5930_ _6626_/Q _5963_/B VGND VGND VPWR VPWR _5930_/X sky130_fd_sc_hd__or2_1
XFILLER_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5861_ _5861_/A _5861_/B _5861_/C _5861_/D VGND VGND VPWR VPWR _5861_/X sky130_fd_sc_hd__or4_2
X_4812_ _4812_/A _5005_/A _4812_/C VGND VGND VPWR VPWR _4812_/X sky130_fd_sc_hd__or3_4
XFILLER_178_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5792_ _6905_/Q _5689_/X _5705_/X _6945_/Q VGND VGND VPWR VPWR _5792_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4743_ _4488_/X _4724_/A _4724_/B _4819_/B VGND VGND VPWR VPWR _4743_/X sky130_fd_sc_hd__a211o_1
XFILLER_166_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4674_ _4745_/A _4832_/A VGND VGND VPWR VPWR _5047_/A sky130_fd_sc_hd__nor2_4
X_6413_ _6446_/A _6446_/B VGND VGND VPWR VPWR _6413_/X sky130_fd_sc_hd__and2_1
XFILLER_147_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3625_ _6951_/Q _5369_/A _4262_/A _6720_/Q _3610_/X VGND VGND VPWR VPWR _3629_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3556_ _7056_/Q _5486_/A _5513_/A _7080_/Q VGND VGND VPWR VPWR _3556_/X sky130_fd_sc_hd__a22o_4
X_6344_ _6767_/Q _6027_/B _6021_/B _6722_/Q VGND VGND VPWR VPWR _6344_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6275_ _6620_/Q _6022_/C _6032_/X _6650_/Q VGND VGND VPWR VPWR _6275_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput109 wb_adr_i[19] VGND VGND VPWR VPWR _4349_/C sky130_fd_sc_hd__clkbuf_4
X_3487_ _7113_/Q hold85/A _5369_/A _6953_/Q _3486_/X VGND VGND VPWR VPWR _3488_/D
+ sky130_fd_sc_hd__a221o_4
XFILLER_130_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5226_ _5226_/A1 _3735_/Y _5576_/B _5225_/X VGND VGND VPWR VPWR _5226_/X sky130_fd_sc_hd__o211a_1
XFILLER_69_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5157_ _5157_/A _5157_/B _5157_/C VGND VGND VPWR VPWR _5158_/B sky130_fd_sc_hd__or3_4
XFILLER_130_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5088_ _4507_/A _5087_/X _4985_/Y VGND VGND VPWR VPWR _5140_/C sky130_fd_sc_hd__a21bo_1
X_4108_ _6585_/Q _4108_/A1 _4111_/S VGND VGND VPWR VPWR _6585_/D sky130_fd_sc_hd__mux2_1
X_4039_ _5581_/A0 hold267/X _4042_/S VGND VGND VPWR VPWR _4039_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_60 _5423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_82 _3504_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_93 _3645_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_71 _3404_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold308 _5511_/X VGND VGND VPWR VPWR _7075_/D sky130_fd_sc_hd__bufbuf_16
Xhold319 _6521_/Q VGND VGND VPWR VPWR hold319/X sky130_fd_sc_hd__bufbuf_16
XFILLER_183_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4390_ _4513_/A _4405_/B VGND VGND VPWR VPWR _4622_/B sky130_fd_sc_hd__nor2_8
X_3410_ _6931_/Q _5342_/A _5387_/A _6971_/Q _3409_/X VGND VGND VPWR VPWR _3414_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_171_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3341_ _3501_/A _5225_/B VGND VGND VPWR VPWR _3341_/Y sky130_fd_sc_hd__nor2_8
XFILLER_98_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3272_ hold18/X hold82/X VGND VGND VPWR VPWR hold19/A sky130_fd_sc_hd__or2_4
X_6060_ _6853_/Q _6060_/B VGND VGND VPWR VPWR _6060_/X sky130_fd_sc_hd__or2_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5011_ _5005_/C _4832_/B _5144_/B _5010_/X VGND VGND VPWR VPWR _5011_/X sky130_fd_sc_hd__o211a_1
Xhold1008 _6750_/Q VGND VGND VPWR VPWR _4301_/A1 sky130_fd_sc_hd__bufbuf_16
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1019 _6642_/Q VGND VGND VPWR VPWR _4176_/A0 sky130_fd_sc_hd__bufbuf_16
XFILLER_93_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6962_ _6971_/CLK _6962_/D fanout451/X VGND VGND VPWR VPWR _6962_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_179_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6893_ _7141_/CLK _6893_/D fanout448/X VGND VGND VPWR VPWR _6893_/Q sky130_fd_sc_hd__dfstp_4
X_5913_ _6749_/Q _5682_/X _5703_/X _6541_/Q VGND VGND VPWR VPWR _5913_/X sky130_fd_sc_hd__a22o_1
X_5844_ _7035_/Q _5688_/X _5690_/X _7099_/Q _5843_/X VGND VGND VPWR VPWR _5849_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5775_ _7064_/Q _5669_/X _5698_/B _6984_/Q _5697_/X VGND VGND VPWR VPWR _5775_/X
+ sky130_fd_sc_hd__a221o_1
X_4726_ _4740_/B _4832_/A VGND VGND VPWR VPWR _4729_/C sky130_fd_sc_hd__nor2_1
XFILLER_175_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4657_ _4758_/B _4657_/B VGND VGND VPWR VPWR _4754_/B sky130_fd_sc_hd__nand2_8
XFILLER_147_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold820 _5554_/X VGND VGND VPWR VPWR _7113_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_174_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput91 spimemio_flash_io3_do VGND VGND VPWR VPWR input91/X sky130_fd_sc_hd__clkbuf_4
XFILLER_116_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput80 spi_sck VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__clkbuf_4
X_3608_ _3607_/X _6793_/Q _3928_/A VGND VGND VPWR VPWR _6793_/D sky130_fd_sc_hd__mux2_1
X_4588_ _4663_/A _4740_/B VGND VGND VPWR VPWR _4588_/X sky130_fd_sc_hd__or2_4
Xhold853 _7057_/Q VGND VGND VPWR VPWR hold853/X sky130_fd_sc_hd__bufbuf_16
Xhold864 _5599_/X VGND VGND VPWR VPWR _7153_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_162_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6327_ _6543_/Q _6023_/C _6025_/B _6566_/Q _6310_/X VGND VGND VPWR VPWR _6330_/C
+ sky130_fd_sc_hd__a221o_1
Xhold842 _4266_/X VGND VGND VPWR VPWR _6721_/D sky130_fd_sc_hd__bufbuf_16
Xhold831 _6757_/Q VGND VGND VPWR VPWR hold831/X sky130_fd_sc_hd__bufbuf_16
Xhold875 _4216_/X VGND VGND VPWR VPWR _6675_/D sky130_fd_sc_hd__bufbuf_16
Xhold886 _5379_/X VGND VGND VPWR VPWR _6957_/D sky130_fd_sc_hd__bufbuf_16
X_3539_ _3540_/A _3732_/B VGND VGND VPWR VPWR _4250_/A sky130_fd_sc_hd__nor2_8
Xhold897 _6655_/Q VGND VGND VPWR VPWR hold897/X sky130_fd_sc_hd__bufbuf_16
XFILLER_130_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6258_ _6530_/Q _6060_/B _6248_/X _6257_/X _6308_/S VGND VGND VPWR VPWR _6258_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_103_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5209_ hold372/X _5578_/A0 _5215_/S VGND VGND VPWR VPWR _6812_/D sky130_fd_sc_hd__mux2_1
X_6189_ _7083_/Q _6311_/B _6036_/Y _7019_/Q _6186_/X VGND VGND VPWR VPWR _6194_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_29_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3890_ _4368_/A _4722_/A VGND VGND VPWR VPWR _4529_/A sky130_fd_sc_hd__nand2_4
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5560_ hold67/X _5560_/A1 _5566_/S VGND VGND VPWR VPWR hold37/A sky130_fd_sc_hd__mux2_1
X_5491_ _5599_/A0 hold853/X _5494_/S VGND VGND VPWR VPWR _5491_/X sky130_fd_sc_hd__mux2_1
X_4511_ _4956_/A _4538_/A VGND VGND VPWR VPWR _4953_/A sky130_fd_sc_hd__nand2_4
XFILLER_157_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4442_ _4529_/C _4442_/B VGND VGND VPWR VPWR _4444_/B sky130_fd_sc_hd__nand2b_4
XFILLER_156_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold105 hold145/X VGND VGND VPWR VPWR _3293_/B sky130_fd_sc_hd__bufbuf_16
Xhold116 hold27/X VGND VGND VPWR VPWR _3668_/A sky130_fd_sc_hd__bufbuf_16
Xhold127 _5534_/X VGND VGND VPWR VPWR _7095_/D sky130_fd_sc_hd__bufbuf_16
Xhold138 _7010_/Q VGND VGND VPWR VPWR hold138/X sky130_fd_sc_hd__bufbuf_16
Xhold149 _5441_/Y VGND VGND VPWR VPWR _5449_/S sky130_fd_sc_hd__bufbuf_16
XFILLER_172_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4373_ _4655_/A _4478_/C VGND VGND VPWR VPWR _4992_/A sky130_fd_sc_hd__nor2_4
XFILLER_144_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7161_ _7193_/CLK _7161_/D fanout435/X VGND VGND VPWR VPWR _7161_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_112_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6112_ _7136_/Q _6020_/B _6011_/X _7096_/Q VGND VGND VPWR VPWR _6112_/X sky130_fd_sc_hd__a22o_1
X_3324_ hold84/X _3473_/A VGND VGND VPWR VPWR _5333_/A sky130_fd_sc_hd__nor2_8
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7092_ _7101_/CLK _7092_/D fanout430/X VGND VGND VPWR VPWR _7092_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_112_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6043_ _6997_/Q _5987_/Y _6036_/Y _7013_/Q _6042_/X VGND VGND VPWR VPWR _6059_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _3845_/A _3255_/B VGND VGND VPWR VPWR _3255_/X sky130_fd_sc_hd__and2b_2
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6945_ _7134_/CLK _6945_/D fanout429/X VGND VGND VPWR VPWR _6945_/Q sky130_fd_sc_hd__dfrtp_2
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
X_6876_ _7122_/CLK _6876_/D fanout443/X VGND VGND VPWR VPWR _6876_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5827_ _5827_/A _5827_/B _5827_/C VGND VGND VPWR VPWR _5827_/X sky130_fd_sc_hd__or3_2
XFILLER_50_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5758_ _6999_/Q _5667_/X _5683_/X _7039_/Q _5757_/X VGND VGND VPWR VPWR _5763_/B
+ sky130_fd_sc_hd__a221o_4
XFILLER_182_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4709_ _4436_/B _5165_/A _4702_/A _4704_/X _4708_/X VGND VGND VPWR VPWR _4713_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_147_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5689_ _5864_/B _5704_/B _5707_/C VGND VGND VPWR VPWR _5689_/X sky130_fd_sc_hd__and3_4
XFILLER_135_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold650 _5267_/X VGND VGND VPWR VPWR _6858_/D sky130_fd_sc_hd__bufbuf_16
Xhold661 _7138_/Q VGND VGND VPWR VPWR hold661/X sky130_fd_sc_hd__bufbuf_16
XFILLER_78_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold672 _6830_/Q VGND VGND VPWR VPWR hold672/X sky130_fd_sc_hd__bufbuf_16
Xhold694 _5502_/X VGND VGND VPWR VPWR _7067_/D sky130_fd_sc_hd__bufbuf_16
Xhold683 _7039_/Q VGND VGND VPWR VPWR hold683/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4991_ _4818_/A _4672_/A _4566_/A _4648_/B VGND VGND VPWR VPWR _4991_/X sky130_fd_sc_hd__a211o_2
XFILLER_63_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6730_ _6804_/CLK _6730_/D _6439_/A VGND VGND VPWR VPWR _6730_/Q sky130_fd_sc_hd__dfstp_4
X_3942_ _6475_/Q _3942_/B VGND VGND VPWR VPWR _3942_/X sky130_fd_sc_hd__or2_1
X_3873_ hold64/A hold38/A _3874_/S VGND VGND VPWR VPWR _6461_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6661_ _6845_/CLK _6661_/D fanout417/X VGND VGND VPWR VPWR _6661_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_177_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6592_ _6713_/CLK _6592_/D fanout426/X VGND VGND VPWR VPWR _6592_/Q sky130_fd_sc_hd__dfrtp_2
X_5612_ _5612_/A _5612_/B VGND VGND VPWR VPWR _5612_/Y sky130_fd_sc_hd__nor2_1
XFILLER_192_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5543_ _5561_/A0 hold859/X hold22/X VGND VGND VPWR VPWR _5543_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5474_ _5582_/A0 hold577/X _5476_/S VGND VGND VPWR VPWR _5474_/X sky130_fd_sc_hd__mux2_1
X_7213_ _3949_/A1 _7213_/D fanout458/X VGND VGND VPWR VPWR _7213_/Q sky130_fd_sc_hd__dfrtp_1
X_4425_ _4422_/Y _4423_/X _4424_/Y _4414_/B VGND VGND VPWR VPWR _4776_/A sky130_fd_sc_hd__a211o_4
XFILLER_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7144_ _7152_/CLK _7144_/D fanout454/X VGND VGND VPWR VPWR _7144_/Q sky130_fd_sc_hd__dfrtp_2
X_4356_ _4722_/A _4529_/B _4486_/B VGND VGND VPWR VPWR _4372_/C sky130_fd_sc_hd__nand3b_4
Xfanout404 _5963_/B VGND VGND VPWR VPWR _5864_/B sky130_fd_sc_hd__buf_8
Xfanout448 fanout449/X VGND VGND VPWR VPWR fanout448/X sky130_fd_sc_hd__buf_8
XFILLER_113_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3307_ hold19/X _3343_/A VGND VGND VPWR VPWR hold20/A sky130_fd_sc_hd__or2_4
Xfanout415 fanout423/X VGND VGND VPWR VPWR _6446_/A sky130_fd_sc_hd__buf_8
Xfanout426 fanout427/X VGND VGND VPWR VPWR fanout426/X sky130_fd_sc_hd__buf_8
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout437 fanout456/X VGND VGND VPWR VPWR fanout437/X sky130_fd_sc_hd__buf_8
Xfanout459 _5007_/A1 VGND VGND VPWR VPWR _4707_/B sky130_fd_sc_hd__buf_8
X_7075_ _7075_/CLK _7075_/D fanout438/X VGND VGND VPWR VPWR _7075_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_59_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4287_ _6407_/A0 _4287_/A1 _4291_/S VGND VGND VPWR VPWR _4287_/X sky130_fd_sc_hd__mux2_1
X_6026_ _6037_/C _6027_/B _6027_/C _6027_/D VGND VGND VPWR VPWR _6232_/A sky130_fd_sc_hd__nor4_4
XFILLER_73_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3238_ _6864_/Q VGND VGND VPWR VPWR _3238_/Y sky130_fd_sc_hd__inv_2
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6928_ _7130_/CLK _6928_/D fanout453/X VGND VGND VPWR VPWR _6928_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_154_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6859_ _7131_/CLK _6859_/D fanout432/X VGND VGND VPWR VPWR _6859_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_183_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold480 _7124_/Q VGND VGND VPWR VPWR hold480/X sky130_fd_sc_hd__bufbuf_16
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold491 _6840_/Q VGND VGND VPWR VPWR hold491/X sky130_fd_sc_hd__bufbuf_16
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1191 _6542_/Q VGND VGND VPWR VPWR _4058_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1180 _4083_/X VGND VGND VPWR VPWR _6563_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_73_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_331 _5595_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_342 hold80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_320 _3944_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_353 hold309/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_364 _6841_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_375 _5276_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_386 _5684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_397 _6028_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_3_0_mgmt_gpio_in[4] clkbuf_2_3_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _3938_/A1
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_9_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4210_ hold916/X _4209_/X _4218_/S VGND VGND VPWR VPWR _4210_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5190_ _6411_/A0 hold733/X _5190_/S VGND VGND VPWR VPWR _5190_/X sky130_fd_sc_hd__mux2_1
X_4141_ _5599_/A0 hold794/X _4141_/S VGND VGND VPWR VPWR _4141_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4072_ _5599_/A0 hold878/X _4072_/S VGND VGND VPWR VPWR _4072_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4974_ _4974_/A _5145_/B _5073_/D _4974_/D VGND VGND VPWR VPWR _4975_/C sky130_fd_sc_hd__or4_1
X_6713_ _6713_/CLK _6713_/D fanout426/X VGND VGND VPWR VPWR _6713_/Q sky130_fd_sc_hd__dfrtp_2
X_3925_ _6667_/Q _3898_/A _3924_/X VGND VGND VPWR VPWR _6667_/D sky130_fd_sc_hd__a21bo_1
XFILLER_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6644_ _7103_/CLK _6644_/D fanout427/X VGND VGND VPWR VPWR _6644_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3856_ _3875_/B _6470_/Q _3856_/S VGND VGND VPWR VPWR _6470_/D sky130_fd_sc_hd__mux2_1
X_3787_ _6853_/Q _3315_/Y _5238_/A _6836_/Q VGND VGND VPWR VPWR _3787_/X sky130_fd_sc_hd__a22o_2
X_6575_ _7220_/CLK _6575_/D VGND VGND VPWR VPWR _6575_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_118_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5526_ hold136/X hold290/X hold55/X VGND VGND VPWR VPWR _7088_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5457_ _5583_/A0 hold729/X _5458_/S VGND VGND VPWR VPWR _5457_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4408_ _4408_/A _4408_/B VGND VGND VPWR VPWR _4410_/D sky130_fd_sc_hd__nand2_4
XFILLER_105_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5388_ _5595_/A0 _5388_/A1 _5395_/S VGND VGND VPWR VPWR _6965_/D sky130_fd_sc_hd__mux2_1
X_7127_ _7127_/CLK _7127_/D fanout449/X VGND VGND VPWR VPWR _7127_/Q sky130_fd_sc_hd__dfrtp_2
X_4339_ _4696_/A _4413_/C VGND VGND VPWR VPWR _4340_/B sky130_fd_sc_hd__nand2_8
XFILLER_132_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7058_ _7154_/CLK _7058_/D fanout454/X VGND VGND VPWR VPWR _7058_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_101_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6009_ _6037_/B _6037_/C _6032_/C VGND VGND VPWR VPWR _6009_/X sky130_fd_sc_hd__and3_4
XFILLER_131_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_150 _5704_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_161 _5861_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_172 _6023_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_194 debug_out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_183 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3710_ _6635_/Q _4166_/A _3701_/X _3709_/X VGND VGND VPWR VPWR _3726_/B sky130_fd_sc_hd__a211o_1
XFILLER_186_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4690_ _4690_/A _4746_/A _5062_/B VGND VGND VPWR VPWR _4757_/B sky130_fd_sc_hd__or3_4
XFILLER_41_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3641_ _6765_/Q _4316_/A _4304_/A _6755_/Q VGND VGND VPWR VPWR _3641_/X sky130_fd_sc_hd__a22o_1
X_3572_ _6607_/Q _4130_/A _4148_/A _6622_/Q VGND VGND VPWR VPWR _3572_/X sky130_fd_sc_hd__a22o_4
X_6360_ _6360_/A _6704_/Q VGND VGND VPWR VPWR _6360_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5311_ _5599_/A0 hold827/X _5314_/S VGND VGND VPWR VPWR _5311_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6291_ _6755_/Q _6023_/D _6030_/Y _6770_/Q _6290_/X VGND VGND VPWR VPWR _6291_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_102_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5242_ _5242_/A _6406_/B VGND VGND VPWR VPWR _5244_/S sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_30_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7141_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_130_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5173_ _5120_/C _5171_/X _5172_/Y VGND VGND VPWR VPWR _5184_/A sky130_fd_sc_hd__o21a_1
X_4124_ _4124_/A _5558_/B VGND VGND VPWR VPWR _4129_/S sky130_fd_sc_hd__and2_4
XFILLER_96_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput1 debug_mode VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__buf_4
XFILLER_56_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4055_ _4055_/A _5558_/B VGND VGND VPWR VPWR _4060_/S sky130_fd_sc_hd__nand2_8
XFILLER_83_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_45_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7088_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_64_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4957_ _4957_/A _5099_/C _4976_/C VGND VGND VPWR VPWR _5128_/D sky130_fd_sc_hd__or3_1
XFILLER_52_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4888_ _4956_/C _4758_/B _4652_/B _5078_/B VGND VGND VPWR VPWR _4909_/B sky130_fd_sc_hd__a31o_1
X_3908_ _6308_/S _3920_/B VGND VGND VPWR VPWR _5665_/A sky130_fd_sc_hd__nor2_4
XFILLER_20_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6627_ _6951_/CLK _6627_/D fanout440/X VGND VGND VPWR VPWR _6627_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_137_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3839_ _3191_/Y _3875_/B _3845_/A VGND VGND VPWR VPWR _3839_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6558_ _7209_/CLK _6558_/D VGND VGND VPWR VPWR _6558_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_146_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5509_ hold185/X hold248/X hold93/X VGND VGND VPWR VPWR _5509_/X sky130_fd_sc_hd__mux2_1
X_6489_ _6759_/CLK _6489_/D fanout421/X VGND VGND VPWR VPWR _6489_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_105_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5860_ _7004_/Q _5667_/X _5702_/X _6892_/Q _5859_/X VGND VGND VPWR VPWR _5861_/D
+ sky130_fd_sc_hd__a221o_4
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4811_ _4736_/B _4758_/B _4695_/X _5105_/A _4810_/Y VGND VGND VPWR VPWR _4817_/A
+ sky130_fd_sc_hd__a311o_1
X_5791_ _7033_/Q _5688_/X _5702_/X _6889_/Q _5790_/X VGND VGND VPWR VPWR _5796_/B
+ sky130_fd_sc_hd__a221o_4
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4742_ _4740_/A _4740_/B _4832_/B _4740_/X _4881_/B VGND VGND VPWR VPWR _4742_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_159_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4673_ _4697_/A _4832_/A VGND VGND VPWR VPWR _4920_/C sky130_fd_sc_hd__nor2_1
XFILLER_119_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3624_ _6631_/Q _4160_/A _3613_/X _3622_/X _3623_/X VGND VGND VPWR VPWR _3636_/B
+ sky130_fd_sc_hd__a2111o_2
X_6412_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6412_/X sky130_fd_sc_hd__and2_1
XFILLER_174_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3555_ _3202_/A _4023_/S _4292_/A _6746_/Q VGND VGND VPWR VPWR _3555_/X sky130_fd_sc_hd__a22o_1
X_6343_ _6343_/A _6343_/B _6343_/C _6343_/D VGND VGND VPWR VPWR _6356_/B sky130_fd_sc_hd__or4_1
X_6274_ _6577_/Q _6021_/A _6025_/A _6605_/Q _6273_/X VGND VGND VPWR VPWR _6281_/A
+ sky130_fd_sc_hd__a221o_1
X_3486_ _6549_/Q _4061_/A _4043_/A _6534_/Q VGND VGND VPWR VPWR _3486_/X sky130_fd_sc_hd__a22o_4
XFILLER_103_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5225_ _5225_/A _5225_/B _5234_/C VGND VGND VPWR VPWR _5225_/X sky130_fd_sc_hd__or3_1
XFILLER_130_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5156_ _6376_/A _5156_/B _5156_/C VGND VGND VPWR VPWR _5157_/C sky130_fd_sc_hd__or3_1
XFILLER_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5087_ _5087_/A _5087_/B _5087_/C _5087_/D VGND VGND VPWR VPWR _5087_/X sky130_fd_sc_hd__or4_4
XFILLER_111_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4107_ _6584_/Q _3606_/X _4111_/S VGND VGND VPWR VPWR _6584_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4038_ _5571_/A0 hold715/X _4042_/S VGND VGND VPWR VPWR _4038_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5989_ _7170_/Q _7171_/Q VGND VGND VPWR VPWR _6014_/A sky130_fd_sc_hd__or2_4
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_50 _5333_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_61 _5423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_83 _3522_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 _3415_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_94 _3664_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput190 _3217_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[23] sky130_fd_sc_hd__buf_8
XFILLER_153_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold309 _6515_/Q VGND VGND VPWR VPWR hold309/X sky130_fd_sc_hd__bufbuf_16
XFILLER_109_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A VGND VGND VPWR VPWR _7220_/CLK sky130_fd_sc_hd__clkbuf_8
X_3340_ _6908_/Q _5315_/A _5459_/A _7036_/Q VGND VGND VPWR VPWR _3340_/X sky130_fd_sc_hd__a22o_1
XFILLER_152_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _4697_/A _4832_/B _4812_/C _4505_/X VGND VGND VPWR VPWR _5010_/X sky130_fd_sc_hd__o22a_1
XFILLER_98_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ hold81/X hold357/X _3991_/S VGND VGND VPWR VPWR _3271_/X sky130_fd_sc_hd__mux2_8
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1009 _6636_/Q VGND VGND VPWR VPWR _4169_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_78_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6961_ _7133_/CLK _6961_/D fanout443/X VGND VGND VPWR VPWR _6961_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_93_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6892_ _7156_/CLK _6892_/D fanout444/X VGND VGND VPWR VPWR _6892_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_81_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5912_ _6577_/Q _5689_/X _5901_/X _5911_/X VGND VGND VPWR VPWR _5915_/C sky130_fd_sc_hd__a211o_1
XFILLER_34_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5843_ _7059_/Q _5706_/X _5842_/X _5698_/B VGND VGND VPWR VPWR _5843_/X sky130_fd_sc_hd__a22o_2
XFILLER_34_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5774_ _6880_/Q _5674_/X _5688_/X _7032_/Q _5773_/X VGND VGND VPWR VPWR _5777_/C
+ sky130_fd_sc_hd__a221o_1
X_4725_ _4725_/A VGND VGND VPWR VPWR _4725_/Y sky130_fd_sc_hd__inv_2
X_4656_ _4758_/B _4657_/B VGND VGND VPWR VPWR _4656_/X sky130_fd_sc_hd__and2_4
XFILLER_147_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4587_ _4663_/A _4740_/B VGND VGND VPWR VPWR _4956_/C sky130_fd_sc_hd__nor2_8
Xinput70 mgmt_gpio_in[7] VGND VGND VPWR VPWR _3972_/B sky130_fd_sc_hd__buf_8
Xinput81 spi_sdo VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__clkbuf_4
Xhold821 _6663_/Q VGND VGND VPWR VPWR hold821/X sky130_fd_sc_hd__bufbuf_16
Xhold810 _6456_/Q VGND VGND VPWR VPWR hold97/A sky130_fd_sc_hd__bufbuf_16
X_3607_ _3606_/X _6792_/Q _3857_/C VGND VGND VPWR VPWR _3607_/X sky130_fd_sc_hd__mux2_1
Xhold843 _6881_/Q VGND VGND VPWR VPWR hold843/X sky130_fd_sc_hd__bufbuf_16
Xhold854 _5491_/X VGND VGND VPWR VPWR _7057_/D sky130_fd_sc_hd__bufbuf_16
Xinput92 spimemio_flash_io3_oeb VGND VGND VPWR VPWR input92/X sky130_fd_sc_hd__clkbuf_4
XFILLER_131_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3538_ _6865_/Q hold28/A _5387_/A _6969_/Q _3537_/X VGND VGND VPWR VPWR _3546_/B
+ sky130_fd_sc_hd__a221o_2
X_6326_ _6579_/Q _6021_/A _6025_/A _6607_/Q _6325_/X VGND VGND VPWR VPWR _6331_/C
+ sky130_fd_sc_hd__a221o_1
Xhold832 _4309_/X VGND VGND VPWR VPWR _6757_/D sky130_fd_sc_hd__bufbuf_16
Xhold876 _6508_/Q VGND VGND VPWR VPWR hold876/X sky130_fd_sc_hd__bufbuf_16
Xhold887 _6671_/Q VGND VGND VPWR VPWR hold887/X sky130_fd_sc_hd__bufbuf_16
XFILLER_107_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold898 _4192_/X VGND VGND VPWR VPWR _6655_/D sky130_fd_sc_hd__bufbuf_16
Xhold865 _6736_/Q VGND VGND VPWR VPWR hold865/X sky130_fd_sc_hd__bufbuf_16
X_6257_ _6356_/A _6257_/B _6257_/C _6257_/D VGND VGND VPWR VPWR _6257_/X sky130_fd_sc_hd__or4_2
XFILLER_67_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3469_ _6752_/Q _4298_/A _4184_/A _6653_/Q VGND VGND VPWR VPWR _3469_/X sky130_fd_sc_hd__a22o_1
XFILLER_190_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5208_ _5208_/A0 _6407_/A0 _5215_/S VGND VGND VPWR VPWR _5208_/X sky130_fd_sc_hd__mux2_1
X_6188_ _7027_/Q _6010_/Y _6031_/X _7091_/Q _6187_/X VGND VGND VPWR VPWR _6194_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_184_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5139_ _4400_/A _4410_/D _4997_/B _5138_/Y VGND VGND VPWR VPWR _5139_/X sky130_fd_sc_hd__o31a_1
XFILLER_111_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5490_ hold71/X _5490_/A1 _5494_/S VGND VGND VPWR VPWR _5490_/X sky130_fd_sc_hd__mux2_1
X_4510_ _4534_/B _4510_/B VGND VGND VPWR VPWR _4538_/A sky130_fd_sc_hd__and2_4
XFILLER_129_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4441_ _4654_/A _4696_/A _4446_/B _4958_/A VGND VGND VPWR VPWR _4442_/B sky130_fd_sc_hd__a31o_2
XFILLER_171_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold106 _3278_/X VGND VGND VPWR VPWR _3314_/B sky130_fd_sc_hd__bufbuf_16
Xhold117 _3299_/Y VGND VGND VPWR VPWR _5414_/A sky130_fd_sc_hd__bufbuf_16
Xhold128 hold204/X VGND VGND VPWR VPWR hold205/A sky130_fd_sc_hd__bufbuf_16
XFILLER_172_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold139 _5438_/X VGND VGND VPWR VPWR _7010_/D sky130_fd_sc_hd__bufbuf_16
X_7160_ _7196_/CLK _7160_/D fanout433/X VGND VGND VPWR VPWR _7160_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_171_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4372_ _4533_/A _4372_/B _4372_/C _4484_/C VGND VGND VPWR VPWR _4410_/C sky130_fd_sc_hd__nand4b_4
X_6111_ _7080_/Q _6311_/B VGND VGND VPWR VPWR _6111_/X sky130_fd_sc_hd__and2_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3323_ input10/X _3320_/Y _4025_/A input60/X _3318_/X VGND VGND VPWR VPWR _3331_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7091_ _7131_/CLK _7091_/D fanout432/X VGND VGND VPWR VPWR _7091_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_112_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6042_ _7101_/Q _5653_/X _6028_/X _6981_/Q VGND VGND VPWR VPWR _6042_/X sky130_fd_sc_hd__a22o_1
XFILLER_98_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3254_ hold104/X hold144/X _3991_/S VGND VGND VPWR VPWR _3254_/X sky130_fd_sc_hd__mux2_8
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6944_ _7138_/CLK _6944_/D fanout438/X VGND VGND VPWR VPWR _6944_/Q sky130_fd_sc_hd__dfrtp_2
X_6875_ _6971_/CLK _6875_/D fanout450/X VGND VGND VPWR VPWR _6875_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_139_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5826_ _5826_/A _5826_/B _5826_/C _5826_/D VGND VGND VPWR VPWR _5826_/X sky130_fd_sc_hd__or4_2
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5757_ _6887_/Q _5702_/X _5756_/X _5698_/B VGND VGND VPWR VPWR _5757_/X sky130_fd_sc_hd__a22o_4
XFILLER_22_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4708_ _4708_/A _4708_/B _4708_/C _4708_/D VGND VGND VPWR VPWR _4708_/X sky130_fd_sc_hd__or4_1
XFILLER_108_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5688_ _7165_/Q _5704_/B _5707_/C VGND VGND VPWR VPWR _5688_/X sky130_fd_sc_hd__and3_4
X_4639_ _4871_/A _4965_/A _4574_/Y _4637_/X _4638_/X VGND VGND VPWR VPWR _4639_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_135_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold662 _5582_/X VGND VGND VPWR VPWR _7138_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_1_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold651 _7131_/Q VGND VGND VPWR VPWR hold651/X sky130_fd_sc_hd__bufbuf_16
Xhold640 _5547_/X VGND VGND VPWR VPWR _7107_/D sky130_fd_sc_hd__bufbuf_16
Xhold695 _6950_/Q VGND VGND VPWR VPWR hold695/X sky130_fd_sc_hd__bufbuf_16
XFILLER_143_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold673 _5232_/X VGND VGND VPWR VPWR _6830_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold684 _5471_/X VGND VGND VPWR VPWR _7039_/D sky130_fd_sc_hd__bufbuf_16
X_6309_ _7199_/Q _6308_/X _6309_/S VGND VGND VPWR VPWR _7199_/D sky130_fd_sc_hd__mux2_1
XFILLER_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4990_ _4990_/A _4997_/B VGND VGND VPWR VPWR _5114_/C sky130_fd_sc_hd__nor2_1
XFILLER_90_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3941_ _6682_/Q _6797_/Q _6455_/B VGND VGND VPWR VPWR _3942_/B sky130_fd_sc_hd__mux2_1
X_3872_ hold38/A _6462_/Q _3874_/S VGND VGND VPWR VPWR _6462_/D sky130_fd_sc_hd__mux2_1
XFILLER_149_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6660_ _6845_/CLK _6660_/D fanout417/X VGND VGND VPWR VPWR _6660_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6591_ _6649_/CLK _6591_/D fanout439/X VGND VGND VPWR VPWR _6591_/Q sky130_fd_sc_hd__dfstp_2
X_5611_ _5611_/A _6680_/Q VGND VGND VPWR VPWR _5612_/B sky130_fd_sc_hd__nor2_1
XFILLER_145_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5542_ hold67/X _7102_/Q hold22/X VGND VGND VPWR VPWR hold68/A sky130_fd_sc_hd__mux2_1
XFILLER_8_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5473_ hold185/X _5473_/A1 _5476_/S VGND VGND VPWR VPWR _5473_/X sky130_fd_sc_hd__mux2_1
X_7212_ _3949_/A1 _7212_/D fanout458/X VGND VGND VPWR VPWR _7212_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_172_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4424_ _4711_/A _4422_/B _4958_/A VGND VGND VPWR VPWR _4424_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_145_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7143_ _7150_/CLK _7143_/D fanout449/X VGND VGND VPWR VPWR _7143_/Q sky130_fd_sc_hd__dfrtp_2
X_4355_ _4529_/B _4486_/B _4722_/A VGND VGND VPWR VPWR _4372_/B sky130_fd_sc_hd__a21bo_4
XFILLER_132_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout405 _3197_/Y VGND VGND VPWR VPWR _6308_/S sky130_fd_sc_hd__buf_8
XFILLER_99_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7074_ _7075_/CLK _7074_/D fanout438/X VGND VGND VPWR VPWR _7074_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout438 fanout456/X VGND VGND VPWR VPWR fanout438/X sky130_fd_sc_hd__buf_8
Xfanout416 fanout423/X VGND VGND VPWR VPWR _6455_/A sky130_fd_sc_hd__buf_8
X_3306_ _3668_/A _3457_/A VGND VGND VPWR VPWR _5342_/A sky130_fd_sc_hd__nor2_8
Xfanout427 fanout456/X VGND VGND VPWR VPWR fanout427/X sky130_fd_sc_hd__buf_8
Xfanout449 fanout455/X VGND VGND VPWR VPWR fanout449/X sky130_fd_sc_hd__buf_8
XFILLER_113_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4286_ _4286_/A _6406_/B VGND VGND VPWR VPWR _4291_/S sky130_fd_sc_hd__nand2_4
X_6025_ _6025_/A _6025_/B _6025_/C _6025_/D VGND VGND VPWR VPWR _6027_/D sky130_fd_sc_hd__or4_4
XFILLER_100_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3237_ _6872_/Q VGND VGND VPWR VPWR _3237_/Y sky130_fd_sc_hd__inv_2
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6927_ _7150_/CLK _6927_/D fanout446/X VGND VGND VPWR VPWR _6927_/Q sky130_fd_sc_hd__dfrtp_2
X_6858_ _7090_/CLK _6858_/D fanout438/X VGND VGND VPWR VPWR _6858_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_80_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5809_ _7180_/Q _6309_/S _5808_/X VGND VGND VPWR VPWR _7180_/D sky130_fd_sc_hd__o21a_1
XFILLER_50_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6789_ _7225_/CLK _6789_/D fanout422/X VGND VGND VPWR VPWR _6789_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_135_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold481 _5566_/X VGND VGND VPWR VPWR _7124_/D sky130_fd_sc_hd__bufbuf_16
Xhold470 _6492_/Q VGND VGND VPWR VPWR hold470/X sky130_fd_sc_hd__bufbuf_16
XFILLER_145_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold492 _5247_/X VGND VGND VPWR VPWR _6840_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_131_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1170 _4265_/X VGND VGND VPWR VPWR _6720_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_310 input120/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1181 _6951_/Q VGND VGND VPWR VPWR _5372_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_73_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1192 _6748_/Q VGND VGND VPWR VPWR _4299_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_45_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_332 _5289_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_321 _3940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_343 hold80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_354 hold309/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_365 hold617/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_376 _7184_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_398 _6030_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_387 _5685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4140_ hold71/X hold242/X _4141_/S VGND VGND VPWR VPWR _4140_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4071_ hold71/X hold305/X _4072_/S VGND VGND VPWR VPWR _4071_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4973_ _5174_/D _5071_/D _4973_/C _4973_/D VGND VGND VPWR VPWR _4974_/D sky130_fd_sc_hd__or4_1
XFILLER_36_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6712_ _6717_/CLK _6712_/D fanout426/X VGND VGND VPWR VPWR _6712_/Q sky130_fd_sc_hd__dfrtp_2
X_3924_ _6457_/Q _6459_/Q _3924_/C VGND VGND VPWR VPWR _3924_/X sky130_fd_sc_hd__or3_1
XFILLER_189_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6643_ _6786_/CLK _6643_/D fanout417/X VGND VGND VPWR VPWR _6643_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_32_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3855_ _3857_/D _6487_/Q _6664_/Q VGND VGND VPWR VPWR _3856_/S sky130_fd_sc_hd__or3b_1
X_6574_ _7209_/CLK _6574_/D VGND VGND VPWR VPWR _6574_/Q sky130_fd_sc_hd__dfxtp_2
X_3786_ _6811_/Q _5207_/A _5191_/A _6798_/Q _3744_/X VGND VGND VPWR VPWR _3792_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_117_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5525_ hold43/X _5525_/A1 hold55/X VGND VGND VPWR VPWR hold56/A sky130_fd_sc_hd__mux2_1
XFILLER_133_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5456_ _5582_/A0 hold691/X _5458_/S VGND VGND VPWR VPWR _5456_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4407_ _4408_/A _4408_/B VGND VGND VPWR VPWR _4499_/C sky130_fd_sc_hd__and2_4
XFILLER_105_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5387_ _5387_/A _5594_/B VGND VGND VPWR VPWR _5395_/S sky130_fd_sc_hd__nand2_8
XFILLER_160_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4338_ _4564_/A _4566_/A VGND VGND VPWR VPWR _4501_/A sky130_fd_sc_hd__or2_4
XFILLER_115_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7126_ _7129_/CLK _7126_/D fanout428/X VGND VGND VPWR VPWR _7126_/Q sky130_fd_sc_hd__dfstp_4
X_7057_ _7153_/CLK _7057_/D fanout442/X VGND VGND VPWR VPWR _7057_/Q sky130_fd_sc_hd__dfrtp_2
X_4269_ _4269_/A0 _5289_/A0 _4273_/S VGND VGND VPWR VPWR _4269_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6008_ _6037_/A _6037_/B _6018_/A VGND VGND VPWR VPWR _6020_/C sky130_fd_sc_hd__and3_4
XFILLER_101_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_140 _5694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_151 _5704_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_173 _6025_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_184 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_162 _5916_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_195 _6972_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3640_ input5/X _3320_/Y _3344_/Y _6498_/Q _3639_/X VGND VGND VPWR VPWR _3645_/B
+ sky130_fd_sc_hd__a221o_4
XFILLER_174_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3571_ input46/X _4217_/S hold61/A _7136_/Q _3570_/X VGND VGND VPWR VPWR _3578_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_155_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5310_ _5571_/A0 hold583/X _5314_/S VGND VGND VPWR VPWR _6896_/D sky130_fd_sc_hd__mux2_1
X_6290_ _6730_/Q _5987_/Y _6022_/D _6596_/Q VGND VGND VPWR VPWR _6290_/X sky130_fd_sc_hd__a22o_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5241_ _5595_/A0 _5241_/A1 _5241_/S VGND VGND VPWR VPWR _5241_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5172_ _5172_/A _5172_/B VGND VGND VPWR VPWR _5172_/Y sky130_fd_sc_hd__nor2_1
XFILLER_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4123_ _4123_/A0 _5545_/A0 _4123_/S VGND VGND VPWR VPWR _4123_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput2 debug_oeb VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_4
XFILLER_68_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4054_ _4054_/A0 _5545_/A0 _4054_/S VGND VGND VPWR VPWR _6539_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_opt_1_0_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR clkbuf_opt_1_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4956_ _4956_/A _4956_/B _4956_/C VGND VGND VPWR VPWR _4976_/C sky130_fd_sc_hd__and3_2
XFILLER_51_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4887_ _4980_/A _4887_/B VGND VGND VPWR VPWR _4978_/B sky130_fd_sc_hd__or2_1
X_3907_ _3920_/B _5612_/A _7159_/Q _7160_/Q VGND VGND VPWR VPWR _3921_/B sky130_fd_sc_hd__and4b_4
X_6626_ _6725_/CLK _6626_/D fanout440/X VGND VGND VPWR VPWR _6626_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_137_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3838_ hold80/A _3837_/Y _3836_/X VGND VGND VPWR VPWR _6478_/D sky130_fd_sc_hd__a21o_1
XFILLER_165_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6557_ _7209_/CLK _6557_/D VGND VGND VPWR VPWR _6557_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_192_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3769_ _6545_/Q _4061_/A _3764_/X _3768_/X _3476_/Y VGND VGND VPWR VPWR _3794_/C
+ sky130_fd_sc_hd__a2111o_1
X_5508_ hold136/X hold239/X hold93/X VGND VGND VPWR VPWR _7072_/D sky130_fd_sc_hd__mux2_1
XFILLER_193_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6488_ _6759_/CLK _6488_/D fanout421/X VGND VGND VPWR VPWR _6488_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_161_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5439_ _5583_/A0 hold696/X _5440_/S VGND VGND VPWR VPWR _5439_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7109_ _7141_/CLK _7109_/D fanout447/X VGND VGND VPWR VPWR _7109_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_113_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4810_ _4745_/B _4660_/X _4809_/X VGND VGND VPWR VPWR _4810_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5790_ _6969_/Q _5691_/X _5701_/X _6953_/Q VGND VGND VPWR VPWR _5790_/X sky130_fd_sc_hd__a22o_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4741_ _4956_/C _4748_/B VGND VGND VPWR VPWR _4881_/B sky130_fd_sc_hd__nand2_4
XFILLER_159_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4672_ _4672_/A _4672_/B _4758_/B VGND VGND VPWR VPWR _5024_/A sky130_fd_sc_hd__and3_1
X_3623_ _6621_/Q _4148_/A _4268_/A _6725_/Q _3619_/X VGND VGND VPWR VPWR _3623_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6411_ _6411_/A0 hold750/X _6411_/S VGND VGND VPWR VPWR _6411_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3554_ _6944_/Q _5360_/A _5369_/A _6952_/Q VGND VGND VPWR VPWR _3554_/X sky130_fd_sc_hd__a22o_1
X_6342_ _6628_/Q _6028_/X _6034_/Y _6727_/Q _6341_/X VGND VGND VPWR VPWR _6343_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_170_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6273_ _6615_/Q _6022_/A _6025_/C _6600_/Q VGND VGND VPWR VPWR _6273_/X sky130_fd_sc_hd__a22o_2
X_3485_ _5234_/A _5252_/B VGND VGND VPWR VPWR _4043_/A sky130_fd_sc_hd__nor2_8
XFILLER_103_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5224_ _5234_/C _5224_/A1 _5224_/S VGND VGND VPWR VPWR _5224_/X sky130_fd_sc_hd__mux2_1
X_5155_ _5155_/A _5155_/B _5178_/C VGND VGND VPWR VPWR _5155_/X sky130_fd_sc_hd__or3_2
XFILLER_69_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5086_ _5086_/A _5086_/B VGND VGND VPWR VPWR _5121_/D sky130_fd_sc_hd__or2_1
XFILLER_84_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4106_ _6583_/Q _3665_/X _4111_/S VGND VGND VPWR VPWR _6583_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4037_ _5597_/A0 hold525/X _4042_/S VGND VGND VPWR VPWR _4037_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5988_ _7170_/Q _7171_/Q VGND VGND VPWR VPWR _6018_/A sky130_fd_sc_hd__nor2_8
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4939_ _4622_/B _4772_/A _4849_/A _4938_/Y VGND VGND VPWR VPWR _4940_/D sky130_fd_sc_hd__a211o_2
XANTENNA_40 _5963_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6609_ _6725_/CLK _6609_/D fanout440/X VGND VGND VPWR VPWR _6609_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_138_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_84 _3522_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 _3415_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 _3331_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 _3378_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_95 _3671_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput191 _3216_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[24] sky130_fd_sc_hd__buf_8
Xoutput180 _3226_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[14] sky130_fd_sc_hd__buf_8
XFILLER_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_44_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7124_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_140_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3270_ hold80/X _3875_/B _3845_/A VGND VGND VPWR VPWR hold81/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_59_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7134_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6960_ _6971_/CLK _6960_/D fanout443/X VGND VGND VPWR VPWR _6960_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5911_ _6590_/Q _5680_/X _5700_/X _6536_/Q _5897_/X VGND VGND VPWR VPWR _5911_/X
+ sky130_fd_sc_hd__a221o_1
X_6891_ _6987_/CLK _6891_/D fanout450/X VGND VGND VPWR VPWR _6891_/Q sky130_fd_sc_hd__dfrtp_2
X_5842_ _6987_/Q _5864_/B VGND VGND VPWR VPWR _5842_/X sky130_fd_sc_hd__or2_1
XFILLER_62_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5773_ _7104_/Q _5675_/X _5684_/X _6992_/Q VGND VGND VPWR VPWR _5773_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4724_ _4724_/A _4724_/B _4812_/C VGND VGND VPWR VPWR _4725_/A sky130_fd_sc_hd__nor3_4
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4655_ _4655_/A _5050_/A _4696_/B VGND VGND VPWR VPWR _4657_/B sky130_fd_sc_hd__and3_4
XFILLER_135_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput60 mgmt_gpio_in[31] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__buf_6
X_4586_ _4868_/A _4586_/B VGND VGND VPWR VPWR _4881_/A sky130_fd_sc_hd__nand2_4
Xinput71 mgmt_gpio_in[8] VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__clkbuf_4
Xinput82 spi_sdoenb VGND VGND VPWR VPWR input82/X sky130_fd_sc_hd__clkbuf_4
Xhold800 _6771_/Q VGND VGND VPWR VPWR hold800/X sky130_fd_sc_hd__bufbuf_16
Xhold811 hold97/X VGND VGND VPWR VPWR hold45/A sky130_fd_sc_hd__bufbuf_16
X_3606_ _3606_/A _3606_/B _3606_/C _3606_/D VGND VGND VPWR VPWR _3606_/X sky130_fd_sc_hd__or4_4
XFILLER_190_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold833 _7121_/Q VGND VGND VPWR VPWR hold833/X sky130_fd_sc_hd__bufbuf_16
Xhold844 _5293_/X VGND VGND VPWR VPWR _6881_/D sky130_fd_sc_hd__bufbuf_16
Xhold855 _6873_/Q VGND VGND VPWR VPWR hold855/X sky130_fd_sc_hd__bufbuf_16
X_3537_ _6929_/Q _5342_/A _5396_/A _6977_/Q VGND VGND VPWR VPWR _3537_/X sky130_fd_sc_hd__a22o_1
X_6325_ _6617_/Q _6022_/A _6025_/C _6602_/Q VGND VGND VPWR VPWR _6325_/X sky130_fd_sc_hd__a22o_1
Xinput93 trap VGND VGND VPWR VPWR input93/X sky130_fd_sc_hd__buf_8
Xhold822 _4201_/X VGND VGND VPWR VPWR _6663_/D sky130_fd_sc_hd__bufbuf_16
Xhold888 _4208_/X VGND VGND VPWR VPWR _6671_/D sky130_fd_sc_hd__bufbuf_16
Xhold877 _4014_/X VGND VGND VPWR VPWR _6508_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold866 _4284_/X VGND VGND VPWR VPWR _6736_/D sky130_fd_sc_hd__bufbuf_16
X_6256_ _7221_/Q _6009_/X _6253_/X _6255_/X VGND VGND VPWR VPWR _6257_/D sky130_fd_sc_hd__a211o_1
XFILLER_107_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3468_ _3514_/A _3733_/B VGND VGND VPWR VPWR _4184_/A sky130_fd_sc_hd__nor2_8
Xhold899 _6531_/Q VGND VGND VPWR VPWR hold899/X sky130_fd_sc_hd__bufbuf_16
XFILLER_191_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5207_ _5207_/A _5576_/B VGND VGND VPWR VPWR _5215_/S sky130_fd_sc_hd__and2_4
X_3399_ _7099_/Q _3341_/Y _5513_/A _7083_/Q _3391_/X VGND VGND VPWR VPWR _3399_/X
+ sky130_fd_sc_hd__a221o_1
X_6187_ _7139_/Q _6020_/B _6011_/X _7099_/Q VGND VGND VPWR VPWR _6187_/X sky130_fd_sc_hd__a22o_1
X_5138_ _4868_/A _4634_/B _4581_/B VGND VGND VPWR VPWR _5138_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_84_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5069_ _5069_/A _5069_/B _5069_/C _5069_/D VGND VGND VPWR VPWR _5076_/B sky130_fd_sc_hd__or4_1
XFILLER_57_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4440_ _4654_/A _4440_/B VGND VGND VPWR VPWR _4958_/B sky130_fd_sc_hd__xor2_4
XFILLER_172_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold107 _3551_/A VGND VGND VPWR VPWR _5234_/A sky130_fd_sc_hd__bufbuf_16
Xhold129 hold206/X VGND VGND VPWR VPWR hold207/A sky130_fd_sc_hd__bufbuf_16
Xhold118 _5420_/X VGND VGND VPWR VPWR _6994_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_171_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4371_ _4533_/A _4372_/B _4372_/C _4484_/C VGND VGND VPWR VPWR _4507_/A sky130_fd_sc_hd__and4b_4
XFILLER_125_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6110_ _7191_/Q _6109_/X _6309_/S VGND VGND VPWR VPWR _7191_/D sky130_fd_sc_hd__mux2_1
X_7090_ _7090_/CLK _7090_/D fanout438/X VGND VGND VPWR VPWR _7090_/Q sky130_fd_sc_hd__dfrtp_2
X_3322_ _5252_/A _5225_/B VGND VGND VPWR VPWR _4025_/A sky130_fd_sc_hd__nor2_8
XFILLER_3_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6041_ _7109_/Q _6027_/B _6039_/X _6040_/X VGND VGND VPWR VPWR _6059_/A sky130_fd_sc_hd__a211o_1
XFILLER_98_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _6482_/Q _3249_/B _3845_/A VGND VGND VPWR VPWR _3253_/X sky130_fd_sc_hd__mux2_2
XFILLER_112_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6943_ _7134_/CLK hold44/X fanout429/X VGND VGND VPWR VPWR _6943_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_179_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6874_ _6874_/CLK _6874_/D fanout443/X VGND VGND VPWR VPWR _6874_/Q sky130_fd_sc_hd__dfrtp_2
X_5825_ _6978_/Q _5676_/X _5702_/X _6890_/Q _5824_/X VGND VGND VPWR VPWR _5826_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_167_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5756_ _6983_/Q _5963_/B VGND VGND VPWR VPWR _5756_/X sky130_fd_sc_hd__or2_1
XFILLER_148_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4707_ _4707_/A _4707_/B _4773_/A _4930_/C VGND VGND VPWR VPWR _5031_/B sky130_fd_sc_hd__or4bb_4
X_5687_ _7165_/Q _5702_/B _5706_/B VGND VGND VPWR VPWR _5687_/X sky130_fd_sc_hd__and3_4
X_4638_ _4819_/B _4819_/D _4947_/B VGND VGND VPWR VPWR _4638_/X sky130_fd_sc_hd__or3_4
XFILLER_163_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold630 _6968_/Q VGND VGND VPWR VPWR hold630/X sky130_fd_sc_hd__bufbuf_16
XFILLER_118_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold663 _6920_/Q VGND VGND VPWR VPWR hold663/X sky130_fd_sc_hd__bufbuf_16
XFILLER_162_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold641 hold641/A VGND VGND VPWR VPWR hold641/X sky130_fd_sc_hd__bufbuf_16
XFILLER_104_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4569_ _4749_/C _4990_/A VGND VGND VPWR VPWR _5071_/A sky130_fd_sc_hd__nor2_4
XFILLER_78_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold652 _5574_/X VGND VGND VPWR VPWR _7131_/D sky130_fd_sc_hd__bufbuf_16
Xmax_cap360 _3506_/A VGND VGND VPWR VPWR _3514_/A sky130_fd_sc_hd__buf_8
X_6308_ _7198_/Q _6307_/X _6308_/S VGND VGND VPWR VPWR _6308_/X sky130_fd_sc_hd__mux2_1
Xhold685 _7019_/Q VGND VGND VPWR VPWR hold685/X sky130_fd_sc_hd__bufbuf_16
Xhold696 _7011_/Q VGND VGND VPWR VPWR hold696/X sky130_fd_sc_hd__bufbuf_16
Xhold674 _6537_/Q VGND VGND VPWR VPWR hold674/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6239_ _6659_/Q _5996_/X _6023_/B _6713_/Q VGND VGND VPWR VPWR _6239_/X sky130_fd_sc_hd__a22o_1
XFILLER_77_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3940_ _6687_/Q input77/X _3969_/B VGND VGND VPWR VPWR _3940_/X sky130_fd_sc_hd__mux2_8
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3871_ _6462_/Q _6463_/Q _3874_/S VGND VGND VPWR VPWR _6463_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6590_ _6713_/CLK _6590_/D fanout426/X VGND VGND VPWR VPWR _6590_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5610_ _7157_/Q _7158_/Q VGND VGND VPWR VPWR _5610_/Y sky130_fd_sc_hd__nand2_1
XFILLER_129_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5541_ _5541_/A0 _5541_/A1 hold22/X VGND VGND VPWR VPWR _7101_/D sky130_fd_sc_hd__mux2_1
XFILLER_157_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7211_ _3949_/A1 _7211_/D fanout458/X VGND VGND VPWR VPWR _7211_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_144_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5472_ hold136/X _7040_/Q _5476_/S VGND VGND VPWR VPWR _5472_/X sky130_fd_sc_hd__mux2_1
X_4423_ _4696_/A _4711_/A _4654_/A VGND VGND VPWR VPWR _4423_/X sky130_fd_sc_hd__a21o_1
XFILLER_144_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7142_ _7151_/CLK _7142_/D fanout446/X VGND VGND VPWR VPWR _7142_/Q sky130_fd_sc_hd__dfstp_4
X_4354_ _4696_/A _4413_/C _4436_/B VGND VGND VPWR VPWR _4486_/B sky130_fd_sc_hd__and3_4
XFILLER_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout439 fanout456/X VGND VGND VPWR VPWR fanout439/X sky130_fd_sc_hd__buf_8
X_3305_ _3673_/B _3540_/A VGND VGND VPWR VPWR _5378_/A sky130_fd_sc_hd__nor2_8
X_7073_ _7136_/CLK _7073_/D fanout436/X VGND VGND VPWR VPWR _7073_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout406 _3979_/S VGND VGND VPWR VPWR _3991_/S sky130_fd_sc_hd__buf_8
Xfanout428 fanout429/X VGND VGND VPWR VPWR fanout428/X sky130_fd_sc_hd__buf_8
Xfanout417 fanout423/X VGND VGND VPWR VPWR fanout417/X sky130_fd_sc_hd__buf_8
X_6024_ _6024_/A _6024_/B _6024_/C _6024_/D VGND VGND VPWR VPWR _6027_/C sky130_fd_sc_hd__or4_4
XFILLER_98_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4285_ _5545_/A0 hold925/X _4285_/S VGND VGND VPWR VPWR _4285_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3236_ _6888_/Q VGND VGND VPWR VPWR _3236_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6926_ _7151_/CLK _6926_/D fanout446/X VGND VGND VPWR VPWR _6926_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_81_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6857_ _7097_/CLK _6857_/D fanout437/X VGND VGND VPWR VPWR _6857_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_167_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6788_ _7225_/CLK _6788_/D fanout422/X VGND VGND VPWR VPWR _6788_/Q sky130_fd_sc_hd__dfrtp_2
X_5808_ _5663_/A _7179_/Q _6358_/B1 _5807_/X VGND VGND VPWR VPWR _5808_/X sky130_fd_sc_hd__a211o_1
X_5739_ _7006_/Q _5678_/X _5692_/X _7070_/Q VGND VGND VPWR VPWR _5739_/X sky130_fd_sc_hd__a22o_1
XFILLER_108_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold460 _4212_/X VGND VGND VPWR VPWR _6673_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold471 _3988_/X VGND VGND VPWR VPWR _6492_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold493 _6980_/Q VGND VGND VPWR VPWR hold493/X sky130_fd_sc_hd__bufbuf_16
Xhold482 _6996_/Q VGND VGND VPWR VPWR hold482/X sky130_fd_sc_hd__bufbuf_16
XFILLER_49_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1160 _6871_/Q VGND VGND VPWR VPWR _5282_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_161_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1182 _5372_/X VGND VGND VPWR VPWR _6951_/D sky130_fd_sc_hd__bufbuf_16
XANTENNA_300 input56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1193 _4299_/X VGND VGND VPWR VPWR _6748_/D sky130_fd_sc_hd__bufbuf_16
Xhold1171 _6811_/Q VGND VGND VPWR VPWR _5208_/A0 sky130_fd_sc_hd__bufbuf_16
XANTENNA_311 input169/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_322 _6356_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_333 _5611_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_355 hold309/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_377 _5963_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_366 hold641/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_344 _3249_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_388 _5688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_399 _6034_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4070_ _5588_/A0 _4070_/A1 _4072_/S VGND VGND VPWR VPWR _6552_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4972_ _4536_/X _4959_/A _5129_/B _4971_/X _4903_/A VGND VGND VPWR VPWR _4973_/D
+ sky130_fd_sc_hd__a2111o_4
XFILLER_64_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6711_ _6717_/CLK _6711_/D fanout426/X VGND VGND VPWR VPWR _6711_/Q sky130_fd_sc_hd__dfrtp_2
X_3923_ _6459_/Q _6664_/Q _3843_/B _6668_/Q VGND VGND VPWR VPWR _6668_/D sky130_fd_sc_hd__a31o_1
XFILLER_149_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3854_ _6486_/Q _6485_/Q VGND VGND VPWR VPWR _3857_/D sky130_fd_sc_hd__nand2b_1
X_6642_ _6845_/CLK _6642_/D fanout417/X VGND VGND VPWR VPWR _6642_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_177_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6573_ _7209_/CLK _6573_/D VGND VGND VPWR VPWR _6573_/Q sky130_fd_sc_hd__dfxtp_2
X_3785_ _3785_/A _3785_/B _3785_/C _3785_/D VGND VGND VPWR VPWR _3793_/C sky130_fd_sc_hd__or4_1
XFILLER_118_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR clkbuf_2_3_0_mgmt_gpio_in[4]/A
+ sky130_fd_sc_hd__clkbuf_8
X_5524_ _5578_/A0 hold339/X hold55/X VGND VGND VPWR VPWR _7086_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5455_ hold185/X hold297/X _5458_/S VGND VGND VPWR VPWR _5455_/X sky130_fd_sc_hd__mux2_1
X_4406_ _4707_/B _4478_/C _4410_/C VGND VGND VPWR VPWR _4513_/B sky130_fd_sc_hd__or3_4
XFILLER_133_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7125_ _7127_/CLK _7125_/D fanout448/X VGND VGND VPWR VPWR _7125_/Q sky130_fd_sc_hd__dfstp_4
X_5386_ hold14/X _5386_/A1 _5386_/S VGND VGND VPWR VPWR _5386_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4337_ _4818_/A _4469_/A _4395_/D VGND VGND VPWR VPWR _4413_/C sky130_fd_sc_hd__and3_4
XFILLER_141_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7056_ _7152_/CLK _7056_/D fanout448/X VGND VGND VPWR VPWR _7056_/Q sky130_fd_sc_hd__dfrtp_2
X_4268_ _4268_/A _5486_/B VGND VGND VPWR VPWR _4273_/S sky130_fd_sc_hd__and2_4
XFILLER_115_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3219_ _7024_/Q VGND VGND VPWR VPWR _3219_/Y sky130_fd_sc_hd__inv_2
X_6007_ _6032_/A _6018_/A _6032_/C VGND VGND VPWR VPWR _6025_/C sky130_fd_sc_hd__and3_4
X_4199_ _6409_/A0 _4199_/A1 _4201_/S VGND VGND VPWR VPWR _6661_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6909_ _7054_/CLK _6909_/D fanout445/X VGND VGND VPWR VPWR _6909_/Q sky130_fd_sc_hd__dfstp_4
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold290 _7088_/Q VGND VGND VPWR VPWR hold290/X sky130_fd_sc_hd__bufbuf_16
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_141 _5694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_152 _5705_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_130 _5566_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_163 _5987_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_174 _6011_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_185 _6084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_196 _6989_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3570_ _6736_/Q _4280_/A _4268_/A _6726_/Q VGND VGND VPWR VPWR _3570_/X sky130_fd_sc_hd__a22o_4
XFILLER_161_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5240_ _5596_/A0 hold425/X _5241_/S VGND VGND VPWR VPWR _5240_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5171_ _5171_/A _5171_/B _5171_/C _5170_/X VGND VGND VPWR VPWR _5171_/X sky130_fd_sc_hd__or4b_1
XFILLER_69_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4122_ hold761/X _4326_/A0 _4123_/S VGND VGND VPWR VPWR _4122_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4053_ hold989/X _6410_/A0 _4054_/S VGND VGND VPWR VPWR _6538_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput3 debug_out VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_4
XFILLER_64_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4955_ _4443_/X _4537_/X _4956_/C _5136_/B _5075_/C VGND VGND VPWR VPWR _5128_/C
+ sky130_fd_sc_hd__a311o_1
XFILLER_101_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3906_ _7157_/Q _7158_/Q VGND VGND VPWR VPWR _5612_/A sky130_fd_sc_hd__nor2_1
XFILLER_51_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4886_ _5005_/C _4886_/B VGND VGND VPWR VPWR _4886_/Y sky130_fd_sc_hd__nor2_1
XFILLER_177_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6625_ _6725_/CLK _6625_/D fanout440/X VGND VGND VPWR VPWR _6625_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_137_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3837_ hold16/A _3825_/B _3840_/S VGND VGND VPWR VPWR _3837_/Y sky130_fd_sc_hd__a21oi_1
X_6556_ _7209_/CLK _6556_/D VGND VGND VPWR VPWR _6556_/Q sky130_fd_sc_hd__dfxtp_4
X_3768_ _6748_/Q _4298_/A _5242_/A _6837_/Q _3767_/X VGND VGND VPWR VPWR _3768_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_152_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5507_ hold43/X _5507_/A1 hold93/X VGND VGND VPWR VPWR hold94/A sky130_fd_sc_hd__mux2_1
XFILLER_145_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6487_ _3957_/A1 _6487_/D _6442_/X VGND VGND VPWR VPWR _6487_/Q sky130_fd_sc_hd__dfrtp_2
X_3699_ _3699_/A _3699_/B _3699_/C _3699_/D VGND VGND VPWR VPWR _3727_/C sky130_fd_sc_hd__or4_2
XFILLER_160_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput340 _6583_/Q VGND VGND VPWR VPWR wb_dat_o[2] sky130_fd_sc_hd__buf_8
X_5438_ hold78/X hold138/X _5440_/S VGND VGND VPWR VPWR _5438_/X sky130_fd_sc_hd__mux2_1
X_5369_ _5369_/A _5594_/B VGND VGND VPWR VPWR _5377_/S sky130_fd_sc_hd__nand2_8
XFILLER_126_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7108_ _7136_/CLK hold23/X fanout436/X VGND VGND VPWR VPWR _7108_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_75_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7039_ _7134_/CLK _7039_/D fanout429/X VGND VGND VPWR VPWR _7039_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_90_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4740_ _4740_/A _4740_/B _4832_/C VGND VGND VPWR VPWR _4740_/X sky130_fd_sc_hd__or3_4
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4671_ _4671_/A _4745_/B VGND VGND VPWR VPWR _5099_/A sky130_fd_sc_hd__nor2_2
XFILLER_186_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3622_ _6591_/Q _4112_/A _4250_/A _6710_/Q _3614_/X VGND VGND VPWR VPWR _3622_/X
+ sky130_fd_sc_hd__a221o_1
X_6410_ _6410_/A0 hold977/X _6411_/S VGND VGND VPWR VPWR _6410_/X sky130_fd_sc_hd__mux2_1
X_6341_ _7225_/Q _6009_/X _6020_/D _6712_/Q VGND VGND VPWR VPWR _6341_/X sky130_fd_sc_hd__a22o_1
X_3553_ _7104_/Q hold21/A _4316_/A _6766_/Q VGND VGND VPWR VPWR _3553_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3484_ _3543_/A _5234_/B VGND VGND VPWR VPWR _4061_/A sky130_fd_sc_hd__nor2_8
X_6272_ _6744_/Q _6023_/A _6033_/X _6739_/Q _6271_/X VGND VGND VPWR VPWR _6282_/B
+ sky130_fd_sc_hd__a221o_2
X_5223_ _5223_/A _6406_/B VGND VGND VPWR VPWR _5224_/S sky130_fd_sc_hd__nand2_1
X_5154_ _5154_/A _5154_/B VGND VGND VPWR VPWR _5178_/C sky130_fd_sc_hd__or2_1
XFILLER_111_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4105_ _6582_/Q _3727_/X _4111_/S VGND VGND VPWR VPWR _6582_/D sky130_fd_sc_hd__mux2_1
X_5085_ _4986_/A _4844_/B _4935_/D VGND VGND VPWR VPWR _5086_/B sky130_fd_sc_hd__o21ai_1
X_4036_ _5596_/A0 hold321/X _4042_/S VGND VGND VPWR VPWR _4036_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5987_ _6036_/A _6004_/A VGND VGND VPWR VPWR _5987_/Y sky130_fd_sc_hd__nor2_8
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4938_ _4745_/A _4697_/A _4757_/B VGND VGND VPWR VPWR _4938_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_178_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_30 _7003_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4869_ _4737_/Y _5087_/D _4949_/C VGND VGND VPWR VPWR _4870_/A sky130_fd_sc_hd__o21ai_2
XFILLER_138_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_41 hold58/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_63 _5288_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_74 _3415_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6608_ _6777_/CLK _6608_/D _6454_/A VGND VGND VPWR VPWR _6608_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_52 _3331_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_85 _3522_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_96 _3687_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6539_ _6777_/CLK _6539_/D fanout424/X VGND VGND VPWR VPWR _6539_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_4_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput192 _3215_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[25] sky130_fd_sc_hd__buf_8
Xoutput181 _3225_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[15] sky130_fd_sc_hd__buf_8
XFILLER_101_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5910_ _5910_/A _5910_/B _5910_/C _5910_/D VGND VGND VPWR VPWR _5915_/B sky130_fd_sc_hd__or4_2
XFILLER_19_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6890_ _7154_/CLK _6890_/D fanout451/X VGND VGND VPWR VPWR _6890_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5841_ _7067_/Q _5669_/X _5703_/X _6875_/Q _5840_/X VGND VGND VPWR VPWR _5849_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_62_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5772_ _6960_/Q _5673_/X _5681_/X _6920_/Q _5771_/X VGND VGND VPWR VPWR _5777_/B
+ sky130_fd_sc_hd__a221o_1
X_4723_ _4947_/B _4898_/B _4886_/B VGND VGND VPWR VPWR _4723_/X sky130_fd_sc_hd__a21o_1
XFILLER_175_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4654_ _4654_/A _4654_/B VGND VGND VPWR VPWR _4696_/B sky130_fd_sc_hd__nor2_8
Xinput50 mgmt_gpio_in[22] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__buf_6
XFILLER_174_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput61 mgmt_gpio_in[32] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__clkbuf_4
XFILLER_128_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4585_ _4634_/B _4586_/B VGND VGND VPWR VPWR _5123_/C sky130_fd_sc_hd__nand2_4
Xinput72 mgmt_gpio_in[9] VGND VGND VPWR VPWR input72/X sky130_fd_sc_hd__buf_4
Xhold812 _3977_/Y VGND VGND VPWR VPWR hold812/X sky130_fd_sc_hd__bufbuf_16
Xhold801 _4326_/X VGND VGND VPWR VPWR _6771_/D sky130_fd_sc_hd__bufbuf_16
X_3605_ _3605_/A _3605_/B _3605_/C _3605_/D VGND VGND VPWR VPWR _3606_/D sky130_fd_sc_hd__or4_1
Xhold834 _5563_/X VGND VGND VPWR VPWR _7121_/D sky130_fd_sc_hd__bufbuf_16
Xhold845 _6937_/Q VGND VGND VPWR VPWR hold845/X sky130_fd_sc_hd__bufbuf_16
Xinput83 spimemio_flash_clk VGND VGND VPWR VPWR input83/X sky130_fd_sc_hd__buf_6
X_6324_ _6746_/Q _6023_/A _6033_/X _6741_/Q _6323_/X VGND VGND VPWR VPWR _6331_/B
+ sky130_fd_sc_hd__a221o_2
X_3536_ _7049_/Q _5477_/A _4262_/A _6722_/Q _3535_/X VGND VGND VPWR VPWR _3546_/A
+ sky130_fd_sc_hd__a221o_1
Xhold823 _6804_/Q VGND VGND VPWR VPWR hold823/X sky130_fd_sc_hd__bufbuf_16
Xinput94 uart_enabled VGND VGND VPWR VPWR _3969_/B sky130_fd_sc_hd__clkbuf_4
Xhold878 _6554_/Q VGND VGND VPWR VPWR hold878/X sky130_fd_sc_hd__bufbuf_16
Xhold856 _5284_/X VGND VGND VPWR VPWR _6873_/D sky130_fd_sc_hd__bufbuf_16
Xhold889 _6512_/Q VGND VGND VPWR VPWR hold889/X sky130_fd_sc_hd__bufbuf_16
X_6255_ _6550_/Q _6020_/A _6034_/Y _6723_/Q _6254_/X VGND VGND VPWR VPWR _6255_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_131_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold867 _6715_/Q VGND VGND VPWR VPWR hold867/X sky130_fd_sc_hd__bufbuf_16
XFILLER_170_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3467_ _3506_/A _3528_/B VGND VGND VPWR VPWR _4298_/A sky130_fd_sc_hd__nor2_8
X_5206_ _5582_/A0 hold605/X _5206_/S VGND VGND VPWR VPWR _5206_/X sky130_fd_sc_hd__mux2_1
X_3398_ _3398_/A _3398_/B _3398_/C _3398_/D VGND VGND VPWR VPWR _3415_/A sky130_fd_sc_hd__or4_2
X_6186_ _7043_/Q _6335_/B VGND VGND VPWR VPWR _6186_/X sky130_fd_sc_hd__and2_1
XFILLER_130_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5137_ _5137_/A _5137_/B _5137_/C VGND VGND VPWR VPWR _5172_/B sky130_fd_sc_hd__or3_1
X_5068_ _5069_/B _5068_/B _5067_/X VGND VGND VPWR VPWR _5132_/C sky130_fd_sc_hd__or3b_1
X_4019_ hold411/X _5600_/A0 _4023_/S VGND VGND VPWR VPWR _4019_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold108 _3315_/Y VGND VGND VPWR VPWR _5261_/A sky130_fd_sc_hd__bufbuf_16
X_4370_ _4484_/C VGND VGND VPWR VPWR _4370_/Y sky130_fd_sc_hd__inv_2
XFILLER_156_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold119 _7106_/Q VGND VGND VPWR VPWR hold119/X sky130_fd_sc_hd__bufbuf_16
XFILLER_125_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3321_ _3419_/A hold83/X VGND VGND VPWR VPWR _3551_/B sky130_fd_sc_hd__or2_4
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6893_/Q _6025_/B _6025_/D _6861_/Q _6038_/X VGND VGND VPWR VPWR _6040_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ hold59/X VGND VGND VPWR VPWR _3314_/A sky130_fd_sc_hd__inv_2
XFILLER_66_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6942_ _7132_/CLK _6942_/D fanout428/X VGND VGND VPWR VPWR _6942_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6873_ _7153_/CLK _6873_/D _6421_/A VGND VGND VPWR VPWR _6873_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5824_ _7066_/Q _5669_/X _5698_/B _6986_/Q _5697_/X VGND VGND VPWR VPWR _5824_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5755_ _6879_/Q _5674_/X _5681_/X _6919_/Q _5754_/X VGND VGND VPWR VPWR _5763_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_147_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4706_ _5165_/A _4453_/Y _4695_/X _5166_/A VGND VGND VPWR VPWR _4706_/X sky130_fd_sc_hd__a31o_1
X_5686_ _6989_/Q _5684_/X _5685_/X _7085_/Q VGND VGND VPWR VPWR _5686_/X sky130_fd_sc_hd__a22o_1
XFILLER_190_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4637_ _4636_/A _4844_/A _4591_/X _4635_/X VGND VGND VPWR VPWR _4637_/X sky130_fd_sc_hd__o211a_1
XFILLER_135_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold620 _6865_/Q VGND VGND VPWR VPWR hold620/X sky130_fd_sc_hd__bufbuf_16
XFILLER_135_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold631 _5391_/X VGND VGND VPWR VPWR _6968_/D sky130_fd_sc_hd__bufbuf_16
Xhold642 _4245_/X VGND VGND VPWR VPWR _6693_/D sky130_fd_sc_hd__bufbuf_16
Xmax_cap350 _6306_/A VGND VGND VPWR VPWR _6356_/A sky130_fd_sc_hd__buf_6
X_4568_ _4868_/A _4624_/B VGND VGND VPWR VPWR _4623_/A sky130_fd_sc_hd__nand2_4
XFILLER_104_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold653 _7035_/Q VGND VGND VPWR VPWR hold653/X sky130_fd_sc_hd__bufbuf_16
Xhold664 _5337_/X VGND VGND VPWR VPWR _6920_/D sky130_fd_sc_hd__bufbuf_16
X_3519_ _7121_/Q _5558_/A _4124_/A _6603_/Q VGND VGND VPWR VPWR _3519_/X sky130_fd_sc_hd__a22o_2
X_4499_ _4553_/B _4507_/A _4499_/C VGND VGND VPWR VPWR _4586_/B sky130_fd_sc_hd__and3b_4
XFILLER_104_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6307_ _6288_/X _6294_/X _6306_/X _6060_/B _6532_/Q VGND VGND VPWR VPWR _6307_/X
+ sky130_fd_sc_hd__o32a_4
Xhold686 _5448_/X VGND VGND VPWR VPWR _7019_/D sky130_fd_sc_hd__bufbuf_16
Xhold697 _5439_/X VGND VGND VPWR VPWR _7011_/D sky130_fd_sc_hd__bufbuf_16
Xhold675 _4052_/X VGND VGND VPWR VPWR _6537_/D sky130_fd_sc_hd__bufbuf_16
X_6238_ _6563_/Q _6025_/B _6020_/C _6589_/Q _6237_/X VGND VGND VPWR VPWR _6248_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6169_ _6986_/Q _6028_/X _6034_/Y _6994_/Q _6168_/X VGND VGND VPWR VPWR _6170_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_43_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7097_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_58_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7129_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3870_ _6463_/Q hold73/A _3874_/S VGND VGND VPWR VPWR _6464_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5540_ hold21/X _5576_/B VGND VGND VPWR VPWR hold22/A sky130_fd_sc_hd__nand2_8
XFILLER_172_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5471_ _5561_/A0 hold683/X _5476_/S VGND VGND VPWR VPWR _5471_/X sky130_fd_sc_hd__mux2_1
X_4422_ _4711_/A _4422_/B VGND VGND VPWR VPWR _4422_/Y sky130_fd_sc_hd__nand2_2
XFILLER_117_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7210_ _7220_/CLK _7210_/D VGND VGND VPWR VPWR _7210_/Q sky130_fd_sc_hd__dfxtp_4
X_7141_ _7141_/CLK _7141_/D fanout448/X VGND VGND VPWR VPWR _7141_/Q sky130_fd_sc_hd__dfstp_4
X_4353_ _4654_/A _4958_/A VGND VGND VPWR VPWR _4436_/B sky130_fd_sc_hd__and2_4
XFILLER_113_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7072_ _7136_/CLK _7072_/D fanout436/X VGND VGND VPWR VPWR _7072_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout429 fanout431/X VGND VGND VPWR VPWR fanout429/X sky130_fd_sc_hd__buf_8
X_3304_ _3314_/A _3304_/B VGND VGND VPWR VPWR _3457_/A sky130_fd_sc_hd__or2_4
Xfanout407 _5611_/A VGND VGND VPWR VPWR _5663_/A sky130_fd_sc_hd__buf_8
Xfanout418 fanout423/X VGND VGND VPWR VPWR fanout418/X sky130_fd_sc_hd__buf_8
X_4284_ _4326_/A0 hold865/X _4285_/S VGND VGND VPWR VPWR _4284_/X sky130_fd_sc_hd__mux2_1
X_6023_ _6023_/A _6023_/B _6023_/C _6023_/D VGND VGND VPWR VPWR _6024_/D sky130_fd_sc_hd__or4_1
XFILLER_98_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3235_ _6896_/Q VGND VGND VPWR VPWR _3235_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6925_ _7127_/CLK _6925_/D fanout448/X VGND VGND VPWR VPWR _6925_/Q sky130_fd_sc_hd__dfstp_4
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6856_ _7140_/CLK _6856_/D fanout428/X VGND VGND VPWR VPWR _6856_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_167_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5807_ _6857_/Q _5722_/B _5796_/X _5806_/X _6308_/S VGND VGND VPWR VPWR _5807_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6787_ _7225_/CLK _6787_/D fanout422/X VGND VGND VPWR VPWR _6787_/Q sky130_fd_sc_hd__dfstp_4
X_3999_ _3999_/A0 _6410_/A0 _4003_/S VGND VGND VPWR VPWR _6499_/D sky130_fd_sc_hd__mux2_1
XFILLER_167_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5738_ _7094_/Q _5690_/X _5693_/X _7078_/Q _5737_/X VGND VGND VPWR VPWR _5741_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_129_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5669_ _7165_/Q _5704_/B _5706_/B VGND VGND VPWR VPWR _5669_/X sky130_fd_sc_hd__and3_4
XFILLER_136_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold461 _7142_/Q VGND VGND VPWR VPWR hold461/X sky130_fd_sc_hd__bufbuf_16
Xhold450 _5330_/X VGND VGND VPWR VPWR _6914_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_150_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold472 _7028_/Q VGND VGND VPWR VPWR hold472/X sky130_fd_sc_hd__bufbuf_16
Xhold494 _5404_/X VGND VGND VPWR VPWR _6980_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_77_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold483 _5422_/X VGND VGND VPWR VPWR _6996_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_145_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1150 _6718_/Q VGND VGND VPWR VPWR _4263_/A0 sky130_fd_sc_hd__bufbuf_16
XFILLER_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1161 _5282_/X VGND VGND VPWR VPWR _6871_/D sky130_fd_sc_hd__bufbuf_16
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1183 _6833_/Q VGND VGND VPWR VPWR _5237_/A1 sky130_fd_sc_hd__bufbuf_16
XANTENNA_301 input56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1194 _6738_/Q VGND VGND VPWR VPWR _4287_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1172 _5208_/X VGND VGND VPWR VPWR _6811_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_312 input169/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_334 _7137_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_323 _5584_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_356 hold309/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_367 hold752/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_345 hold209/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_389 _5688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_378 _3249_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_96_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4971_ _5130_/A _4971_/B _4970_/X VGND VGND VPWR VPWR _4971_/X sky130_fd_sc_hd__or3b_2
XFILLER_91_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6710_ _6717_/CLK _6710_/D fanout426/X VGND VGND VPWR VPWR _6710_/Q sky130_fd_sc_hd__dfstp_4
X_3922_ _6679_/Q _5606_/B VGND VGND VPWR VPWR _6678_/D sky130_fd_sc_hd__or2_1
XFILLER_32_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3853_ _3875_/B _6471_/Q _3853_/S VGND VGND VPWR VPWR _6471_/D sky130_fd_sc_hd__mux2_1
X_6641_ _7225_/CLK _6641_/D fanout417/X VGND VGND VPWR VPWR _6641_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_32_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6572_ _7209_/CLK _6572_/D VGND VGND VPWR VPWR _6572_/Q sky130_fd_sc_hd__dfxtp_2
X_3784_ input11/X _3368_/Y _4286_/A _6738_/Q _3783_/X VGND VGND VPWR VPWR _3785_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_157_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5523_ _5541_/A0 _5523_/A1 hold55/X VGND VGND VPWR VPWR _7085_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5454_ hold136/X hold228/X _5458_/S VGND VGND VPWR VPWR _5454_/X sky130_fd_sc_hd__mux2_1
X_4405_ _4553_/A _4405_/B VGND VGND VPWR VPWR _4636_/A sky130_fd_sc_hd__or2_4
X_5385_ hold209/X hold291/X _5386_/S VGND VGND VPWR VPWR _5385_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4336_ _4469_/A _4395_/D VGND VGND VPWR VPWR _4566_/A sky130_fd_sc_hd__nand2_8
XFILLER_99_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7124_ _7124_/CLK _7124_/D fanout437/X VGND VGND VPWR VPWR _7124_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_5_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7055_ _7150_/CLK _7055_/D fanout446/X VGND VGND VPWR VPWR _7055_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_140_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4267_ _4267_/A0 _5545_/A0 _4267_/S VGND VGND VPWR VPWR _6722_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3218_ _7032_/Q VGND VGND VPWR VPWR _3218_/Y sky130_fd_sc_hd__inv_2
X_6006_ _6035_/A _6018_/A _6035_/C VGND VGND VPWR VPWR _6022_/A sky130_fd_sc_hd__and3_4
XFILLER_74_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4198_ _5254_/A0 hold940/X _4201_/S VGND VGND VPWR VPWR _4198_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6908_ _6964_/CLK _6908_/D fanout445/X VGND VGND VPWR VPWR _6908_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6839_ _6840_/CLK _6839_/D _6454_/A VGND VGND VPWR VPWR _6839_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_183_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold280 _5410_/X VGND VGND VPWR VPWR _6985_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_151_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold291 _6963_/Q VGND VGND VPWR VPWR hold291/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_120 _4763_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 _5575_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_142 _5694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_164 _5987_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_153 _5706_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_175 _6011_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_186 _6144_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_197 _6997_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5170_ _4871_/A _4988_/A _4617_/A _4997_/B _4893_/A VGND VGND VPWR VPWR _5170_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_110_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4121_ hold712/X _5561_/A0 _4123_/S VGND VGND VPWR VPWR _6596_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4052_ hold674/X _5561_/A0 _4054_/S VGND VGND VPWR VPWR _4052_/X sky130_fd_sc_hd__mux2_1
Xinput4 mask_rev_in[0] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_4
XFILLER_52_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4954_ _4636_/A _4986_/C _5005_/C _4591_/B VGND VGND VPWR VPWR _5075_/C sky130_fd_sc_hd__o22ai_4
XFILLER_101_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3905_ _6019_/A _6030_/A VGND VGND VPWR VPWR _3905_/X sky130_fd_sc_hd__or2_4
X_4885_ _4986_/A _4997_/A _4740_/X _4395_/D VGND VGND VPWR VPWR _5123_/D sky130_fd_sc_hd__o22a_1
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6624_ _6725_/CLK _6624_/D fanout440/X VGND VGND VPWR VPWR _6624_/Q sky130_fd_sc_hd__dfrtp_2
X_3836_ _3191_/Y _3840_/S _3825_/B hold16/A VGND VGND VPWR VPWR _3836_/X sky130_fd_sc_hd__o211a_1
XFILLER_118_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6555_ _7208_/CLK _6555_/D VGND VGND VPWR VPWR _6555_/Q sky130_fd_sc_hd__dfxtp_2
X_3767_ _6504_/Q _4004_/A _3765_/X _3766_/X VGND VGND VPWR VPWR _3767_/X sky130_fd_sc_hd__a211o_2
XFILLER_118_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5506_ _5578_/A0 hold420/X hold93/X VGND VGND VPWR VPWR _7070_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6486_ _3957_/A1 _6486_/D _6441_/X VGND VGND VPWR VPWR _6486_/Q sky130_fd_sc_hd__dfrtp_2
X_3698_ _7094_/Q _3341_/Y _4304_/A _6754_/Q _3675_/X VGND VGND VPWR VPWR _3699_/D
+ sky130_fd_sc_hd__a221o_1
Xoutput341 _7209_/Q VGND VGND VPWR VPWR wb_dat_o[30] sky130_fd_sc_hd__buf_8
XFILLER_126_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput330 _6559_/Q VGND VGND VPWR VPWR wb_dat_o[20] sky130_fd_sc_hd__buf_8
X_5437_ hold185/X hold275/X _5440_/S VGND VGND VPWR VPWR _5437_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5368_ _5584_/A0 hold398/X _5368_/S VGND VGND VPWR VPWR _5368_/X sky130_fd_sc_hd__mux2_1
X_5299_ _5587_/A0 hold507/X _5305_/S VGND VGND VPWR VPWR _6886_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7107_ _7107_/CLK _7107_/D fanout435/X VGND VGND VPWR VPWR _7107_/Q sky130_fd_sc_hd__dfrtp_2
X_4319_ _4319_/A0 _6409_/A0 _4321_/S VGND VGND VPWR VPWR _6765_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7038_ _7129_/CLK _7038_/D fanout428/X VGND VGND VPWR VPWR _7038_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4670_ _4832_/B _4660_/X _4664_/X _4669_/X VGND VGND VPWR VPWR _4670_/X sky130_fd_sc_hd__o211a_1
XFILLER_119_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3621_ _6911_/Q _5324_/A _4217_/S input45/X _3620_/X VGND VGND VPWR VPWR _3636_/A
+ sky130_fd_sc_hd__a221o_4
XFILLER_119_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6340_ _6732_/Q _5987_/Y _6022_/D _6598_/Q _6339_/X VGND VGND VPWR VPWR _6343_/C
+ sky130_fd_sc_hd__a221o_1
X_3552_ hold84/X _3552_/B VGND VGND VPWR VPWR _3552_/Y sky130_fd_sc_hd__nor2_8
X_3483_ _7089_/Q hold54/A _4118_/A _6598_/Q _3482_/X VGND VGND VPWR VPWR _3488_/C
+ sky130_fd_sc_hd__a221o_1
X_6271_ _6764_/Q _6027_/B _6021_/B _6719_/Q _6270_/X VGND VGND VPWR VPWR _6271_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5222_ _5222_/A0 hold136/X _5222_/S VGND VGND VPWR VPWR _5222_/X sky130_fd_sc_hd__mux2_1
X_5153_ _4737_/Y _5152_/X _4758_/B VGND VGND VPWR VPWR _5154_/B sky130_fd_sc_hd__o21a_1
XFILLER_111_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4104_ _6581_/Q _3794_/X _4111_/S VGND VGND VPWR VPWR _6581_/D sky130_fd_sc_hd__mux2_1
X_5084_ _5084_/A _5084_/B VGND VGND VPWR VPWR _5119_/B sky130_fd_sc_hd__or2_1
XFILLER_111_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4035_ hold885/X _4035_/A1 _4042_/S VGND VGND VPWR VPWR _4035_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5986_ _6012_/A _6033_/C VGND VGND VPWR VPWR _6004_/A sky130_fd_sc_hd__nand2_8
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4937_ _5033_/A _5033_/B _5033_/C _5035_/C VGND VGND VPWR VPWR _4940_/C sky130_fd_sc_hd__or4_1
XANTENNA_31 _5494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4868_ _4868_/A _4949_/B _4956_/B VGND VGND VPWR VPWR _5087_/D sky130_fd_sc_hd__and3_2
XANTENNA_20 _5196_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_64 _5288_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6607_ _6722_/CLK _6607_/D _6454_/A VGND VGND VPWR VPWR _6607_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_75 _3415_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_42 _5477_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3819_ _6482_/Q _6481_/Q _3828_/S hold50/A VGND VGND VPWR VPWR _3820_/C sky130_fd_sc_hd__a31o_1
XANTENNA_53 _3978_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4799_ _4799_/A _4799_/B _5180_/A _4799_/D VGND VGND VPWR VPWR _4800_/D sky130_fd_sc_hd__or4_1
XANTENNA_97 _3693_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_86 _3562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6538_ _6786_/CLK _6538_/D fanout417/X VGND VGND VPWR VPWR _6538_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_173_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6469_ _3957_/A1 _6469_/D _6424_/X VGND VGND VPWR VPWR _6469_/Q sky130_fd_sc_hd__dfrtp_2
Xoutput193 _3214_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[26] sky130_fd_sc_hd__buf_8
Xoutput182 _3224_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[16] sky130_fd_sc_hd__buf_8
XFILLER_133_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput171 _3971_/X VGND VGND VPWR VPWR debug_in sky130_fd_sc_hd__buf_8
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5840_ _6883_/Q _5674_/X _5692_/X _7075_/Q VGND VGND VPWR VPWR _5840_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5771_ _6968_/Q _5691_/X _5701_/X _6952_/Q VGND VGND VPWR VPWR _5771_/X sky130_fd_sc_hd__a22o_1
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4722_ _4722_/A _4722_/B _4368_/A VGND VGND VPWR VPWR _4812_/C sky130_fd_sc_hd__or3b_4
XFILLER_159_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput40 mgmt_gpio_in[13] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__clkbuf_4
X_4653_ _5164_/B _4832_/A VGND VGND VPWR VPWR _4653_/Y sky130_fd_sc_hd__nor2_4
X_4584_ _4584_/A _4740_/B VGND VGND VPWR VPWR _5005_/C sky130_fd_sc_hd__or2_4
Xinput51 mgmt_gpio_in[23] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__clkbuf_4
Xhold802 _6511_/Q VGND VGND VPWR VPWR hold802/X sky130_fd_sc_hd__bufbuf_16
Xinput62 mgmt_gpio_in[33] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__buf_4
Xinput73 pad_flash_io0_di VGND VGND VPWR VPWR _3964_/B sky130_fd_sc_hd__clkbuf_4
X_3604_ _7096_/Q _3341_/Y _4322_/A _6771_/Q _3603_/X VGND VGND VPWR VPWR _3605_/D
+ sky130_fd_sc_hd__a221o_1
Xinput95 usr1_vcc_pwrgood VGND VGND VPWR VPWR input95/X sky130_fd_sc_hd__buf_6
Xhold846 _5356_/X VGND VGND VPWR VPWR _6937_/D sky130_fd_sc_hd__bufbuf_16
Xinput84 spimemio_flash_csb VGND VGND VPWR VPWR input84/X sky130_fd_sc_hd__buf_6
XFILLER_155_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold813 _5252_/D VGND VGND VPWR VPWR _4241_/D sky130_fd_sc_hd__bufbuf_16
Xhold835 _6746_/Q VGND VGND VPWR VPWR hold835/X sky130_fd_sc_hd__bufbuf_16
X_6323_ _6766_/Q _6027_/B _6021_/B _6721_/Q _6322_/X VGND VGND VPWR VPWR _6323_/X
+ sky130_fd_sc_hd__a221o_1
Xhold824 _5199_/X VGND VGND VPWR VPWR _6804_/D sky130_fd_sc_hd__bufbuf_16
X_3535_ input30/X _3283_/Y _5567_/A _7129_/Q VGND VGND VPWR VPWR _3535_/X sky130_fd_sc_hd__a22o_4
Xhold879 _4072_/X VGND VGND VPWR VPWR _6554_/D sky130_fd_sc_hd__bufbuf_16
X_6254_ _6718_/Q _6021_/B _6028_/X _6624_/Q VGND VGND VPWR VPWR _6254_/X sky130_fd_sc_hd__a22o_1
Xhold868 _7137_/Q VGND VGND VPWR VPWR hold868/X sky130_fd_sc_hd__bufbuf_16
XFILLER_115_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3466_ _6961_/Q _5378_/A hold61/A _7137_/Q _3465_/X VGND VGND VPWR VPWR _3472_/C
+ sky130_fd_sc_hd__a221o_4
XFILLER_107_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold857 _7033_/Q VGND VGND VPWR VPWR hold857/X sky130_fd_sc_hd__bufbuf_16
XFILLER_170_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5205_ _6411_/A0 hold787/X _5206_/S VGND VGND VPWR VPWR _6809_/D sky130_fd_sc_hd__mux2_1
XFILLER_97_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3397_ input9/X _3320_/Y _5459_/A _7035_/Q _3392_/X VGND VGND VPWR VPWR _3398_/D
+ sky130_fd_sc_hd__a221o_4
X_6185_ _7194_/Q _5665_/Y _6183_/X _6184_/X VGND VGND VPWR VPWR _7194_/D sky130_fd_sc_hd__o22a_1
X_5136_ _5136_/A _5136_/B _5136_/C _5136_/D VGND VGND VPWR VPWR _5137_/C sky130_fd_sc_hd__or4_1
XFILLER_111_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5067_ _4469_/A _4819_/A _4603_/B _4740_/B VGND VGND VPWR VPWR _5067_/X sky130_fd_sc_hd__a211o_1
XFILLER_123_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4018_ hold770/X _4017_/X _4024_/S VGND VGND VPWR VPWR _4018_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5969_ _6777_/Q _5683_/X _5704_/X _6608_/Q _5968_/X VGND VGND VPWR VPWR _5976_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_52_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold109 _5269_/X VGND VGND VPWR VPWR _6860_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_171_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3320_ _5225_/A _3375_/B VGND VGND VPWR VPWR _3320_/Y sky130_fd_sc_hd__nor2_8
XFILLER_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ hold58/X hold173/X _3991_/S VGND VGND VPWR VPWR _3251_/X sky130_fd_sc_hd__mux2_8
XFILLER_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6941_ _7132_/CLK _6941_/D fanout428/X VGND VGND VPWR VPWR _6941_/Q sky130_fd_sc_hd__dfstp_4
X_6872_ _6874_/CLK _6872_/D fanout443/X VGND VGND VPWR VPWR _6872_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5823_ _7106_/Q _5675_/X _5684_/X _6994_/Q _5822_/X VGND VGND VPWR VPWR _5826_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5754_ _6959_/Q _5673_/X _5691_/X _6967_/Q VGND VGND VPWR VPWR _5754_/X sky130_fd_sc_hd__a22o_1
XFILLER_175_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4705_ _5023_/B _4724_/B VGND VGND VPWR VPWR _5166_/A sky130_fd_sc_hd__nor2_2
X_5685_ _7165_/Q _5707_/B _5701_/C VGND VGND VPWR VPWR _5685_/X sky130_fd_sc_hd__and3_4
XFILLER_163_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4636_ _4636_/A _4989_/A VGND VGND VPWR VPWR _5136_/B sky130_fd_sc_hd__nor2_4
XFILLER_118_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold621 _5275_/X VGND VGND VPWR VPWR _6865_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_162_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold610 _4270_/X VGND VGND VPWR VPWR _6724_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_190_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4567_ _4694_/A _4947_/B _6707_/Q VGND VGND VPWR VPWR _4567_/X sky130_fd_sc_hd__o21a_2
X_6306_ _6306_/A _6306_/B _6306_/C VGND VGND VPWR VPWR _6306_/X sky130_fd_sc_hd__or3_4
Xhold643 _7043_/Q VGND VGND VPWR VPWR hold643/X sky130_fd_sc_hd__bufbuf_16
Xhold654 _5466_/X VGND VGND VPWR VPWR _7035_/D sky130_fd_sc_hd__bufbuf_16
Xhold632 _7018_/Q VGND VGND VPWR VPWR hold632/X sky130_fd_sc_hd__bufbuf_16
X_4498_ _4986_/A _4745_/B VGND VGND VPWR VPWR _5119_/A sky130_fd_sc_hd__nor2_4
XFILLER_143_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3518_ _3543_/A _3733_/B VGND VGND VPWR VPWR _4124_/A sky130_fd_sc_hd__nor2_8
Xhold665 _7015_/Q VGND VGND VPWR VPWR hold665/X sky130_fd_sc_hd__bufbuf_16
Xhold687 _6847_/Q VGND VGND VPWR VPWR hold687/X sky130_fd_sc_hd__bufbuf_16
Xhold676 _6991_/Q VGND VGND VPWR VPWR hold676/X sky130_fd_sc_hd__bufbuf_16
X_6237_ _6728_/Q _5987_/Y _6022_/B _6609_/Q VGND VGND VPWR VPWR _6237_/X sky130_fd_sc_hd__a22o_1
X_3449_ input49/X _4217_/S hold61/A _7138_/Q _3448_/X VGND VGND VPWR VPWR _3450_/D
+ sky130_fd_sc_hd__a221o_4
XFILLER_77_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold698 _7123_/Q VGND VGND VPWR VPWR hold698/X sky130_fd_sc_hd__bufbuf_16
XFILLER_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6168_ _7074_/Q _6009_/X _6020_/D _6970_/Q VGND VGND VPWR VPWR _6168_/X sky130_fd_sc_hd__a22o_1
XFILLER_76_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5119_ _5119_/A _5119_/B _5119_/C VGND VGND VPWR VPWR _5135_/C sky130_fd_sc_hd__or3_1
XFILLER_94_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6099_ _7127_/Q _6023_/A _6033_/X _7007_/Q _6098_/X VGND VGND VPWR VPWR _6107_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A VGND VGND VPWR VPWR _7193_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5470_ _5578_/A0 hold346/X _5476_/S VGND VGND VPWR VPWR _7038_/D sky130_fd_sc_hd__mux2_1
X_4421_ _4728_/A _4671_/A VGND VGND VPWR VPWR _4702_/A sky130_fd_sc_hd__nor2_2
XFILLER_117_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4352_ _4352_/A _4352_/B _4352_/C VGND VGND VPWR VPWR _4529_/B sky130_fd_sc_hd__and3_4
X_7140_ _7140_/CLK _7140_/D fanout428/X VGND VGND VPWR VPWR _7140_/Q sky130_fd_sc_hd__dfrtp_2
X_4283_ _5588_/A0 hold947/X _4285_/S VGND VGND VPWR VPWR _6735_/D sky130_fd_sc_hd__mux2_1
XFILLER_152_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7071_ _7136_/CLK hold94/X fanout436/X VGND VGND VPWR VPWR _7071_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout419 fanout421/X VGND VGND VPWR VPWR fanout419/X sky130_fd_sc_hd__buf_8
Xfanout408 _6678_/Q VGND VGND VPWR VPWR _5611_/A sky130_fd_sc_hd__buf_8
X_3303_ _7028_/Q _5450_/A _3302_/Y input28/X _3300_/X VGND VGND VPWR VPWR _3331_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_140_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6022_ _6022_/A _6022_/B _6022_/C _6022_/D VGND VGND VPWR VPWR _6024_/C sky130_fd_sc_hd__or4_1
XFILLER_98_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3234_ _6904_/Q VGND VGND VPWR VPWR _3234_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6924_ _7152_/CLK _6924_/D fanout452/X VGND VGND VPWR VPWR _6924_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6855_ _7097_/CLK _6855_/D fanout437/X VGND VGND VPWR VPWR _6855_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5806_ _5806_/A _5806_/B _5806_/C _5806_/D VGND VGND VPWR VPWR _5806_/X sky130_fd_sc_hd__or4_2
X_6786_ _6786_/CLK _6786_/D fanout422/X VGND VGND VPWR VPWR _6786_/Q sky130_fd_sc_hd__dfrtp_2
X_3998_ _3998_/A0 _6409_/A0 _4003_/S VGND VGND VPWR VPWR _6498_/D sky130_fd_sc_hd__mux2_1
XFILLER_148_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5737_ _7014_/Q _5682_/X _5703_/X _6870_/Q VGND VGND VPWR VPWR _5737_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5668_ _7163_/Q _7164_/Q VGND VGND VPWR VPWR _5706_/B sky130_fd_sc_hd__and2b_4
XFILLER_135_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5599_ _5599_/A0 hold863/X _5602_/S VGND VGND VPWR VPWR _5599_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4619_ _4619_/A _4619_/B _4619_/C _4619_/D VGND VGND VPWR VPWR _4619_/X sky130_fd_sc_hd__and4_1
XFILLER_190_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold451 _7146_/Q VGND VGND VPWR VPWR hold451/X sky130_fd_sc_hd__bufbuf_16
Xhold462 _7065_/Q VGND VGND VPWR VPWR hold462/X sky130_fd_sc_hd__bufbuf_16
Xhold440 _5575_/X VGND VGND VPWR VPWR _7132_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_145_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold484 _7068_/Q VGND VGND VPWR VPWR hold484/X sky130_fd_sc_hd__bufbuf_16
XFILLER_104_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold495 _6577_/Q VGND VGND VPWR VPWR hold495/X sky130_fd_sc_hd__bufbuf_16
Xhold473 _5458_/X VGND VGND VPWR VPWR _7028_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_77_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1151 _4263_/X VGND VGND VPWR VPWR _6718_/D sky130_fd_sc_hd__bufbuf_16
Xhold1140 _6604_/Q VGND VGND VPWR VPWR _4131_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_85_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1162 _6745_/Q VGND VGND VPWR VPWR _4295_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1184 _5237_/X VGND VGND VPWR VPWR _6833_/D sky130_fd_sc_hd__bufbuf_16
Xhold1173 _6629_/Q VGND VGND VPWR VPWR _4161_/A1 sky130_fd_sc_hd__bufbuf_16
XANTENNA_313 input169/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_324 _5601_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_302 input50/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1195 _4287_/X VGND VGND VPWR VPWR _6738_/D sky130_fd_sc_hd__bufbuf_16
XANTENNA_357 hold335/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_368 _6671_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_346 hold209/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_335 hold7/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_379 _3253_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4970_ _5147_/A _4970_/B _4959_/A VGND VGND VPWR VPWR _4970_/X sky130_fd_sc_hd__or3b_2
XFILLER_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3921_ _6308_/S _3921_/B VGND VGND VPWR VPWR _5606_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3852_ _6487_/Q _6486_/Q _6485_/Q _6664_/Q VGND VGND VPWR VPWR _3853_/S sky130_fd_sc_hd__or4b_1
X_6640_ _6786_/CLK _6640_/D fanout417/X VGND VGND VPWR VPWR _6640_/Q sky130_fd_sc_hd__dfrtp_2
X_6571_ _7209_/CLK _6571_/D VGND VGND VPWR VPWR _6571_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_20_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5522_ hold54/X _5576_/B VGND VGND VPWR VPWR hold55/A sky130_fd_sc_hd__nand2_8
X_3783_ _6989_/Q _3299_/Y _3341_/Y _7093_/Q VGND VGND VPWR VPWR _3783_/X sky130_fd_sc_hd__a22o_2
XFILLER_118_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5453_ hold43/A _5453_/A1 _5458_/S VGND VGND VPWR VPWR hold34/A sky130_fd_sc_hd__mux2_1
X_5384_ _5600_/A0 hold579/X _5386_/S VGND VGND VPWR VPWR _5384_/X sky130_fd_sc_hd__mux2_1
X_4404_ _4553_/A _4405_/B VGND VGND VPWR VPWR _4845_/A sky130_fd_sc_hd__nor2_2
Xclkbuf_leaf_42_csclk _7137_/CLK VGND VGND VPWR VPWR _7122_/CLK sky130_fd_sc_hd__clkbuf_8
X_4335_ _4707_/B _5050_/A VGND VGND VPWR VPWR _4728_/A sky130_fd_sc_hd__nand2_8
XFILLER_125_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7123_ _7123_/CLK _7123_/D fanout434/X VGND VGND VPWR VPWR _7123_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_115_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7054_ _7054_/CLK _7054_/D fanout445/X VGND VGND VPWR VPWR _7054_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_140_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4266_ hold841/X _4326_/A0 _4267_/S VGND VGND VPWR VPWR _4266_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3217_ _7040_/Q VGND VGND VPWR VPWR _3217_/Y sky130_fd_sc_hd__inv_2
X_6005_ _6014_/A _6010_/B VGND VGND VPWR VPWR _6025_/B sky130_fd_sc_hd__nor2_8
XFILLER_55_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_57_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7132_/CLK sky130_fd_sc_hd__clkbuf_8
X_4197_ _5234_/C _4197_/A1 _4201_/S VGND VGND VPWR VPWR _4197_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6907_ _6976_/CLK _6907_/D fanout450/X VGND VGND VPWR VPWR _6907_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6838_ _6845_/CLK _6838_/D fanout417/X VGND VGND VPWR VPWR _6838_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6769_ _7222_/CLK _6769_/D fanout422/X VGND VGND VPWR VPWR _6769_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold270 _5536_/X VGND VGND VPWR VPWR _7097_/D sky130_fd_sc_hd__bufbuf_16
Xhold281 _6513_/Q VGND VGND VPWR VPWR hold281/X sky130_fd_sc_hd__bufbuf_16
Xhold292 _5385_/X VGND VGND VPWR VPWR _6963_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_132 _5593_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_121 _4906_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_143 _5702_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_110 _3830_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 _6020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_154 _5734_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_176 _6011_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_198 _7000_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_187 _6146_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4120_ hold513/X _6408_/A0 _4123_/S VGND VGND VPWR VPWR _4120_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4051_ hold891/X _5254_/A0 _4054_/S VGND VGND VPWR VPWR _4051_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput5 mask_rev_in[10] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_4
XFILLER_37_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4953_ _4953_/A _5062_/A VGND VGND VPWR VPWR _5068_/B sky130_fd_sc_hd__nor2_1
XFILLER_51_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3904_ _6012_/A _6037_/A VGND VGND VPWR VPWR _6030_/A sky130_fd_sc_hd__nand2_8
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4884_ _4898_/B _4756_/B _4623_/A VGND VGND VPWR VPWR _4907_/A sky130_fd_sc_hd__o21ai_4
X_6623_ _6715_/CLK _6623_/D fanout439/X VGND VGND VPWR VPWR _6623_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_60_670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3835_ _3834_/X hold24/A _3840_/S VGND VGND VPWR VPWR _6479_/D sky130_fd_sc_hd__mux2_1
X_6554_ _6745_/CLK _6554_/D _6421_/A VGND VGND VPWR VPWR _6554_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_118_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3766_ _7005_/Q _5432_/A _4322_/A _6768_/Q VGND VGND VPWR VPWR _3766_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5505_ _5541_/A0 _5505_/A1 hold93/X VGND VGND VPWR VPWR _7069_/D sky130_fd_sc_hd__mux2_1
X_6485_ _6668_/CLK _6485_/D _6440_/X VGND VGND VPWR VPWR _6485_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_161_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3697_ _6655_/Q _4190_/A _6406_/A _7222_/Q _3674_/X VGND VGND VPWR VPWR _3699_/C
+ sky130_fd_sc_hd__a221o_2
X_5436_ hold136/X hold258/X _5440_/S VGND VGND VPWR VPWR _5436_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput342 _7210_/Q VGND VGND VPWR VPWR wb_dat_o[31] sky130_fd_sc_hd__buf_8
XFILLER_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput331 _6560_/Q VGND VGND VPWR VPWR wb_dat_o[21] sky130_fd_sc_hd__buf_8
XFILLER_105_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput320 _6571_/Q VGND VGND VPWR VPWR wb_dat_o[11] sky130_fd_sc_hd__buf_8
XFILLER_120_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5367_ _5583_/A0 hold622/X _5368_/S VGND VGND VPWR VPWR _5367_/X sky130_fd_sc_hd__mux2_1
X_5298_ _5595_/A0 _5298_/A1 _5305_/S VGND VGND VPWR VPWR _6885_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7106_ _7106_/CLK _7106_/D fanout438/X VGND VGND VPWR VPWR _7106_/Q sky130_fd_sc_hd__dfrtp_2
X_4318_ hold914/X _5254_/A0 _4321_/S VGND VGND VPWR VPWR _4318_/X sky130_fd_sc_hd__mux2_1
X_4249_ hold3/X _4249_/A1 _4249_/S VGND VGND VPWR VPWR hold4/A sky130_fd_sc_hd__mux2_1
XFILLER_75_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7037_ _7132_/CLK _7037_/D fanout428/X VGND VGND VPWR VPWR _7037_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_142_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3620_ _7143_/Q _5585_/A _4280_/A _6735_/Q VGND VGND VPWR VPWR _3620_/X sky130_fd_sc_hd__a22o_1
XFILLER_128_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3551_ _3551_/A _3551_/B VGND VGND VPWR VPWR _3551_/Y sky130_fd_sc_hd__nor2_4
XFILLER_155_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3482_ _7057_/Q _5486_/A _4082_/A _6567_/Q VGND VGND VPWR VPWR _3482_/X sky130_fd_sc_hd__a22o_1
X_6270_ _6551_/Q _6020_/A _6021_/D _6630_/Q VGND VGND VPWR VPWR _6270_/X sky130_fd_sc_hd__a22o_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5221_ hold680/X _5561_/A0 _5222_/S VGND VGND VPWR VPWR _6822_/D sky130_fd_sc_hd__mux2_1
X_5152_ _5062_/C _5050_/C _5041_/X _4668_/B VGND VGND VPWR VPWR _5152_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_111_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4103_ _6701_/Q _6362_/B VGND VGND VPWR VPWR _4111_/S sky130_fd_sc_hd__and2_4
X_5083_ _5137_/A _5171_/B _5115_/A _5117_/A VGND VGND VPWR VPWR _5083_/X sky130_fd_sc_hd__or4_2
XFILLER_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4034_ hold20/X _4241_/A _6421_/B _5252_/D VGND VGND VPWR VPWR _4042_/S sky130_fd_sc_hd__or4_4
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5985_ _7169_/Q _7168_/Q VGND VGND VPWR VPWR _6033_/C sky130_fd_sc_hd__nor2_8
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4936_ _4936_/A _4936_/B _4936_/C VGND VGND VPWR VPWR _5035_/C sky130_fd_sc_hd__or3_2
XFILLER_52_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_10 _4028_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_32 _5499_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4867_ _4818_/A _4740_/A _4452_/Y _4866_/X VGND VGND VPWR VPWR _4867_/X sky130_fd_sc_hd__a31o_1
XFILLER_138_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_21 _6802_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6606_ _6649_/CLK _6606_/D fanout439/X VGND VGND VPWR VPWR _6606_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA_65 _5288_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_54 _3978_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 _5477_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3818_ _6484_/Q _3840_/S _3817_/Y VGND VGND VPWR VPWR _6484_/D sky130_fd_sc_hd__a21o_1
XFILLER_119_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4798_ _4798_/A _5022_/B _4798_/C _4798_/D VGND VGND VPWR VPWR _4799_/D sky130_fd_sc_hd__or4_1
XANTENNA_87 _3587_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 _3415_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_98 _3711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6537_ _6840_/CLK _6537_/D fanout424/X VGND VGND VPWR VPWR _6537_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_180_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3749_ _6965_/Q _5387_/A _4154_/A _6624_/Q _3748_/X VGND VGND VPWR VPWR _3754_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6468_ _6668_/CLK _6468_/D _6423_/X VGND VGND VPWR VPWR _6468_/Q sky130_fd_sc_hd__dfrtp_2
X_6399_ _6705_/Q _6399_/A2 _6399_/B1 _4238_/B _6398_/X VGND VGND VPWR VPWR _6399_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5419_ hold185/X hold230/X _5422_/S VGND VGND VPWR VPWR _5419_/X sky130_fd_sc_hd__mux2_1
Xoutput194 _3213_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[27] sky130_fd_sc_hd__buf_8
Xoutput183 _3223_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[17] sky130_fd_sc_hd__buf_8
Xoutput172 _6825_/Q VGND VGND VPWR VPWR irq[0] sky130_fd_sc_hd__buf_8
XFILLER_153_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5770_ _7040_/Q _5683_/X _5704_/X _6936_/Q _5769_/X VGND VGND VPWR VPWR _5777_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4721_ _4818_/C _4724_/B _4238_/B VGND VGND VPWR VPWR _5003_/B sky130_fd_sc_hd__o21a_4
XFILLER_159_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4652_ _4758_/B _4652_/B VGND VGND VPWR VPWR _4832_/A sky130_fd_sc_hd__nand2_8
X_3603_ _3877_/C _4234_/S _4262_/A _6721_/Q _3602_/X VGND VGND VPWR VPWR _3603_/X
+ sky130_fd_sc_hd__a221o_4
Xinput30 mask_rev_in[4] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__clkbuf_4
Xinput52 mgmt_gpio_in[24] VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__clkbuf_4
Xinput63 mgmt_gpio_in[34] VGND VGND VPWR VPWR _3970_/A sky130_fd_sc_hd__buf_8
X_4583_ _4584_/A _4740_/B VGND VGND VPWR VPWR _4736_/B sky130_fd_sc_hd__nor2_8
Xhold803 _4020_/X VGND VGND VPWR VPWR _6511_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_162_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput41 mgmt_gpio_in[14] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__clkbuf_4
XFILLER_116_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput96 usr1_vdd_pwrgood VGND VGND VPWR VPWR input96/X sky130_fd_sc_hd__buf_6
Xhold814 _4246_/X VGND VGND VPWR VPWR _6694_/D sky130_fd_sc_hd__bufbuf_16
Xinput85 spimemio_flash_io0_do VGND VGND VPWR VPWR input85/X sky130_fd_sc_hd__buf_6
XFILLER_143_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6322_ _6553_/Q _6020_/A _6021_/D _6632_/Q VGND VGND VPWR VPWR _6322_/X sky130_fd_sc_hd__a22o_1
Xhold836 _4296_/X VGND VGND VPWR VPWR _6746_/D sky130_fd_sc_hd__bufbuf_16
Xhold825 _7119_/Q VGND VGND VPWR VPWR hold825/X sky130_fd_sc_hd__bufbuf_16
Xinput74 pad_flash_io1_di VGND VGND VPWR VPWR _3965_/B sky130_fd_sc_hd__clkbuf_4
X_3534_ _3534_/A _5252_/A VGND VGND VPWR VPWR _4262_/A sky130_fd_sc_hd__nor2_8
Xhold869 _5581_/X VGND VGND VPWR VPWR _7137_/D sky130_fd_sc_hd__bufbuf_16
X_6253_ _6629_/Q _6021_/D _6030_/Y _6768_/Q VGND VGND VPWR VPWR _6253_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3465_ _6897_/Q _5306_/A _4190_/A _6658_/Q VGND VGND VPWR VPWR _3465_/X sky130_fd_sc_hd__a22o_1
Xhold858 _5464_/X VGND VGND VPWR VPWR _7033_/D sky130_fd_sc_hd__bufbuf_16
Xhold847 _6688_/Q VGND VGND VPWR VPWR hold847/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5204_ _6410_/A0 hold980/X _5206_/S VGND VGND VPWR VPWR _5204_/X sky130_fd_sc_hd__mux2_1
X_3396_ _6939_/Q _5351_/A _5369_/A _6955_/Q _3387_/X VGND VGND VPWR VPWR _3398_/C
+ sky130_fd_sc_hd__a221o_4
XFILLER_130_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6184_ _5663_/A _7193_/Q _5664_/X VGND VGND VPWR VPWR _6184_/X sky130_fd_sc_hd__a21o_1
X_5135_ _5135_/A _5135_/B _5135_/C _5135_/D VGND VGND VPWR VPWR _5172_/A sky130_fd_sc_hd__or4_2
XFILLER_97_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5066_ _5066_/A _5124_/B VGND VGND VPWR VPWR _5074_/A sky130_fd_sc_hd__nand2_2
XFILLER_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4017_ hold267/X _5581_/A0 _4023_/S VGND VGND VPWR VPWR _4017_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5968_ _6732_/Q _5667_/X _5687_/X _6643_/Q VGND VGND VPWR VPWR _5968_/X sky130_fd_sc_hd__a22o_1
X_4919_ _4395_/D _4469_/Y _4656_/X _4796_/B _4412_/Y VGND VGND VPWR VPWR _5095_/B
+ sky130_fd_sc_hd__a311o_2
XFILLER_32_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5899_ _6625_/Q _5963_/B VGND VGND VPWR VPWR _5899_/X sky130_fd_sc_hd__or2_1
XFILLER_21_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ hold111/X _3845_/A _3249_/Y VGND VGND VPWR VPWR hold58/A sky130_fd_sc_hd__a21bo_2
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6940_ _6975_/CLK _6940_/D fanout443/X VGND VGND VPWR VPWR _6940_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_81_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6871_ _7153_/CLK _6871_/D fanout444/X VGND VGND VPWR VPWR _6871_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_179_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5822_ _6882_/Q _5674_/X _5688_/X _7034_/Q VGND VGND VPWR VPWR _5822_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5753_ _5753_/A _5753_/B _5753_/C _5753_/D VGND VGND VPWR VPWR _5753_/X sky130_fd_sc_hd__or4_4
XFILLER_34_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4704_ _4772_/A _4711_/C _4772_/C VGND VGND VPWR VPWR _4704_/X sky130_fd_sc_hd__and3_4
XFILLER_148_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5684_ _7165_/Q _5703_/B _5707_/B VGND VGND VPWR VPWR _5684_/X sky130_fd_sc_hd__and3_4
XFILLER_147_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4635_ _4996_/A _4844_/A _4631_/X _4633_/X _5144_/A VGND VGND VPWR VPWR _4635_/X
+ sky130_fd_sc_hd__o2111a_1
X_4566_ _4566_/A _4740_/B VGND VGND VPWR VPWR _4947_/B sky130_fd_sc_hd__or2_4
Xhold600 _5295_/X VGND VGND VPWR VPWR _6883_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold611 _6719_/Q VGND VGND VPWR VPWR hold611/X sky130_fd_sc_hd__bufbuf_16
XFILLER_150_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6305_ _6305_/A _6305_/B _6305_/C _6305_/D VGND VGND VPWR VPWR _6306_/C sky130_fd_sc_hd__or4_1
X_3517_ _7009_/Q _5432_/A _3317_/Y _7065_/Q _3516_/X VGND VGND VPWR VPWR _3522_/C
+ sky130_fd_sc_hd__a221o_1
Xhold644 _5475_/X VGND VGND VPWR VPWR _7043_/D sky130_fd_sc_hd__bufbuf_16
Xhold633 _5447_/X VGND VGND VPWR VPWR _7018_/D sky130_fd_sc_hd__bufbuf_16
Xhold622 _6947_/Q VGND VGND VPWR VPWR hold622/X sky130_fd_sc_hd__bufbuf_16
XFILLER_171_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4497_ _5164_/B _4745_/B VGND VGND VPWR VPWR _5013_/A sky130_fd_sc_hd__nor2_4
XFILLER_143_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold655 _7050_/Q VGND VGND VPWR VPWR hold655/X sky130_fd_sc_hd__bufbuf_16
Xhold666 _5444_/X VGND VGND VPWR VPWR _7015_/D sky130_fd_sc_hd__bufbuf_16
Xhold688 _5255_/X VGND VGND VPWR VPWR _6847_/D sky130_fd_sc_hd__bufbuf_16
Xhold677 _5417_/X VGND VGND VPWR VPWR _6991_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_134_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6236_ _6743_/Q _6023_/A _6020_/D _6708_/Q VGND VGND VPWR VPWR _6248_/A sky130_fd_sc_hd__a22o_1
X_3448_ _7050_/Q _5477_/A _5297_/A _6890_/Q VGND VGND VPWR VPWR _3448_/X sky130_fd_sc_hd__a22o_1
Xhold699 _5565_/X VGND VGND VPWR VPWR _7123_/D sky130_fd_sc_hd__bufbuf_16
X_6167_ _7122_/Q _6023_/D _6030_/Y _7034_/Q _6166_/X VGND VGND VPWR VPWR _6170_/C
+ sky130_fd_sc_hd__a221o_1
X_3379_ _3379_/A _3379_/B _3379_/C VGND VGND VPWR VPWR _3379_/X sky130_fd_sc_hd__or3_4
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _5118_/A _5118_/B _5118_/C _5118_/D VGND VGND VPWR VPWR _5119_/C sky130_fd_sc_hd__or4_1
XFILLER_97_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6098_ _6887_/Q _6020_/A _6021_/D _7143_/Q _6097_/X VGND VGND VPWR VPWR _6098_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_84_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5049_ _4956_/C _4668_/B _5041_/X _4657_/B VGND VGND VPWR VPWR _5049_/X sky130_fd_sc_hd__a22o_1
XFILLER_150_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4420_ _4654_/A _4707_/B _5050_/A VGND VGND VPWR VPWR _4422_/B sky130_fd_sc_hd__and3_2
XFILLER_8_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4351_ _4351_/A _4351_/B _4351_/C _4351_/D VGND VGND VPWR VPWR _4352_/C sky130_fd_sc_hd__and4_1
XFILLER_153_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7070_ _7136_/CLK _7070_/D fanout436/X VGND VGND VPWR VPWR _7070_/Q sky130_fd_sc_hd__dfstp_2
X_3302_ hold91/A _5225_/A VGND VGND VPWR VPWR _3302_/Y sky130_fd_sc_hd__nor2_8
Xfanout409 _6667_/Q VGND VGND VPWR VPWR _3845_/A sky130_fd_sc_hd__buf_8
X_4282_ _6408_/A0 hold566/X _4285_/S VGND VGND VPWR VPWR _4282_/X sky130_fd_sc_hd__mux2_1
X_6021_ _6021_/A _6021_/B _6021_/C _6021_/D VGND VGND VPWR VPWR _6024_/B sky130_fd_sc_hd__or4_1
X_3233_ _6912_/Q VGND VGND VPWR VPWR _3233_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_101_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_1_csclk clkbuf_1_1_1_csclk/A VGND VGND VPWR VPWR clkbuf_2_3_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_79_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6923_ _7154_/CLK _6923_/D fanout452/X VGND VGND VPWR VPWR _6923_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_82_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6854_ _7101_/CLK _6854_/D fanout430/X VGND VGND VPWR VPWR _6854_/Q sky130_fd_sc_hd__dfstp_2
X_5805_ _6977_/Q _5676_/X _5685_/X _7089_/Q _5804_/X VGND VGND VPWR VPWR _5806_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3997_ hold909/X _5254_/A0 _4003_/S VGND VGND VPWR VPWR _6497_/D sky130_fd_sc_hd__mux2_1
X_6785_ _7225_/CLK _6785_/D fanout422/X VGND VGND VPWR VPWR _6785_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5736_ _6902_/Q _5689_/X _5725_/X _5735_/X VGND VGND VPWR VPWR _5741_/A sky130_fd_sc_hd__a211o_4
XFILLER_13_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5667_ _7165_/Q _5703_/B _5704_/B VGND VGND VPWR VPWR _5667_/X sky130_fd_sc_hd__and3_4
XFILLER_190_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4618_ _4844_/A _4749_/C _4617_/A VGND VGND VPWR VPWR _4619_/D sky130_fd_sc_hd__a21o_1
XFILLER_190_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5598_ hold71/X hold140/X _5602_/S VGND VGND VPWR VPWR _5598_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold452 _5591_/X VGND VGND VPWR VPWR _7146_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_163_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold463 _5500_/X VGND VGND VPWR VPWR _7065_/D sky130_fd_sc_hd__bufbuf_16
X_4549_ _4987_/B _4624_/B _5114_/A _4548_/X VGND VGND VPWR VPWR _4549_/X sky130_fd_sc_hd__a211o_1
XFILLER_104_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold430 _5260_/X VGND VGND VPWR VPWR _6852_/D sky130_fd_sc_hd__bufbuf_16
Xhold441 _7022_/Q VGND VGND VPWR VPWR hold441/X sky130_fd_sc_hd__bufbuf_16
XFILLER_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold485 _5503_/X VGND VGND VPWR VPWR _7068_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_104_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold496 _4099_/X VGND VGND VPWR VPWR _6577_/D sky130_fd_sc_hd__bufbuf_16
Xhold474 _7012_/Q VGND VGND VPWR VPWR hold474/X sky130_fd_sc_hd__bufbuf_16
XFILLER_104_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6219_ _6219_/A _6219_/B _6219_/C _6219_/D VGND VGND VPWR VPWR _6219_/X sky130_fd_sc_hd__or4_1
X_7199_ _7201_/CLK _7199_/D _6446_/A VGND VGND VPWR VPWR _7199_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1130 _4125_/X VGND VGND VPWR VPWR _6599_/D sky130_fd_sc_hd__bufbuf_16
Xhold1141 _4131_/X VGND VGND VPWR VPWR _6604_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_100_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1152 _6919_/Q VGND VGND VPWR VPWR _5336_/A0 sky130_fd_sc_hd__bufbuf_16
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1174 _4161_/X VGND VGND VPWR VPWR _6629_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_85_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1163 _6708_/Q VGND VGND VPWR VPWR _4251_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_58_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1185 _6785_/Q VGND VGND VPWR VPWR _5186_/A1 sky130_fd_sc_hd__bufbuf_16
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_303 input49/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_314 input169/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1196 _6800_/Q VGND VGND VPWR VPWR _5195_/A1 sky130_fd_sc_hd__bufbuf_16
XANTENNA_325 _5582_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_358 hold335/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_336 hold14/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_347 hold209/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_369 _6672_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3920_ _5663_/A _3920_/B VGND VGND VPWR VPWR _3920_/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3851_ _3797_/X _3898_/A _3850_/Y _6664_/Q VGND VGND VPWR VPWR _6472_/D sky130_fd_sc_hd__a211oi_1
X_6570_ _7209_/CLK _6570_/D VGND VGND VPWR VPWR _6570_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3782_ _7061_/Q _3317_/Y hold21/A _7101_/Q _3781_/X VGND VGND VPWR VPWR _3785_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_164_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5521_ _5584_/A0 hold400/X _5521_/S VGND VGND VPWR VPWR _5521_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5452_ _5578_/A0 hold441/X _5458_/S VGND VGND VPWR VPWR _7022_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5383_ _5581_/A0 hold433/X _5386_/S VGND VGND VPWR VPWR _5383_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4403_ _4671_/A _4617_/A VGND VGND VPWR VPWR _4847_/A sky130_fd_sc_hd__nor2_2
X_4334_ _4707_/B _5050_/A VGND VGND VPWR VPWR _4696_/A sky130_fd_sc_hd__and2_4
XFILLER_141_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7122_ _7122_/CLK _7122_/D fanout443/X VGND VGND VPWR VPWR _7122_/Q sky130_fd_sc_hd__dfrtp_2
X_7053_ _7111_/CLK _7053_/D fanout445/X VGND VGND VPWR VPWR _7053_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_141_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4265_ _4265_/A0 _5588_/A0 _4267_/S VGND VGND VPWR VPWR _4265_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6004_ _6004_/A _6014_/A VGND VGND VPWR VPWR _6023_/C sky130_fd_sc_hd__nor2_8
X_3216_ _7048_/Q VGND VGND VPWR VPWR _3216_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4196_ _4196_/A _6406_/B VGND VGND VPWR VPWR _4201_/S sky130_fd_sc_hd__nand2_4
XFILLER_82_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6906_ _6971_/CLK _6906_/D fanout451/X VGND VGND VPWR VPWR _6906_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_70_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6837_ _6845_/CLK _6837_/D fanout417/X VGND VGND VPWR VPWR _6837_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6768_ _7222_/CLK _6768_/D fanout422/X VGND VGND VPWR VPWR _6768_/Q sky130_fd_sc_hd__dfrtp_2
X_5719_ _6917_/Q _5681_/X _5682_/X _7013_/Q _5677_/X VGND VGND VPWR VPWR _5720_/D
+ sky130_fd_sc_hd__a221o_1
X_6699_ _7220_/CLK _6699_/D _6362_/B VGND VGND VPWR VPWR _6704_/D sky130_fd_sc_hd__dfrtp_2
XFILLER_40_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold260 _6979_/Q VGND VGND VPWR VPWR hold260/X sky130_fd_sc_hd__bufbuf_16
Xhold271 _7049_/Q VGND VGND VPWR VPWR hold271/X sky130_fd_sc_hd__bufbuf_16
Xhold282 _4024_/X VGND VGND VPWR VPWR _6513_/D sky130_fd_sc_hd__bufbuf_16
Xhold293 _6849_/Q VGND VGND VPWR VPWR hold293/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_100 _3785_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_133 _5658_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_111 _3831_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_122 _5251_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_144 _5703_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_166 _6020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_155 _5734_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_177 _6020_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_199 _6729_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_188 _6196_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4050_ _4050_/A0 _6407_/A0 _4054_/S VGND VGND VPWR VPWR _4050_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput6 mask_rev_in[11] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4952_ _4949_/A _4956_/A _4736_/B _4983_/B VGND VGND VPWR VPWR _5142_/B sky130_fd_sc_hd__a31o_2
X_4883_ _4883_/A _4922_/A VGND VGND VPWR VPWR _4983_/B sky130_fd_sc_hd__or2_2
X_3903_ _7169_/Q _7168_/Q VGND VGND VPWR VPWR _6037_/A sky130_fd_sc_hd__and2b_4
XFILLER_189_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6622_ _6713_/CLK _6622_/D fanout426/X VGND VGND VPWR VPWR _6622_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_60_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3834_ hold16/A _3845_/A _3827_/Y _3833_/X VGND VGND VPWR VPWR _3834_/X sky130_fd_sc_hd__a22o_1
X_6553_ _6745_/CLK _6553_/D fanout440/X VGND VGND VPWR VPWR _6553_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_118_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3765_ input4/X _3283_/Y _3359_/Y _7013_/Q VGND VGND VPWR VPWR _3765_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5504_ hold92/X hold47/X VGND VGND VPWR VPWR hold93/A sky130_fd_sc_hd__nand2_8
X_6484_ _6668_/CLK _6484_/D _6439_/X VGND VGND VPWR VPWR _6484_/Q sky130_fd_sc_hd__dfrtp_4
X_3696_ input21/X _3302_/Y _3359_/Y _7014_/Q _3695_/X VGND VGND VPWR VPWR _3699_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_145_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput310 _3952_/X VGND VGND VPWR VPWR serial_load sky130_fd_sc_hd__buf_8
X_5435_ _5561_/A0 hold717/X _5440_/S VGND VGND VPWR VPWR _5435_/X sky130_fd_sc_hd__mux2_1
Xoutput332 _6561_/Q VGND VGND VPWR VPWR wb_dat_o[22] sky130_fd_sc_hd__buf_8
Xoutput321 _6572_/Q VGND VGND VPWR VPWR wb_dat_o[12] sky130_fd_sc_hd__buf_8
Xoutput343 _6584_/Q VGND VGND VPWR VPWR wb_dat_o[3] sky130_fd_sc_hd__buf_8
XFILLER_10_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5366_ _5582_/A0 hold710/X _5368_/S VGND VGND VPWR VPWR _5366_/X sky130_fd_sc_hd__mux2_1
X_5297_ _5297_/A _5594_/B VGND VGND VPWR VPWR _5305_/S sky130_fd_sc_hd__nand2_8
XFILLER_99_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4317_ _4317_/A0 _5234_/C _4321_/S VGND VGND VPWR VPWR _4317_/X sky130_fd_sc_hd__mux2_1
X_7105_ _7105_/CLK _7105_/D fanout436/X VGND VGND VPWR VPWR _7105_/Q sky130_fd_sc_hd__dfrtp_2
X_4248_ _5601_/A0 hold521/X _4249_/S VGND VGND VPWR VPWR _4248_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7036_ _7132_/CLK _7036_/D fanout428/X VGND VGND VPWR VPWR _7036_/Q sky130_fd_sc_hd__dfrtp_2
X_4179_ _4179_/A0 _6407_/A0 _4183_/S VGND VGND VPWR VPWR _4179_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_56_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7140_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_128_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3550_ _3549_/X _6794_/Q _3928_/A VGND VGND VPWR VPWR _6794_/D sky130_fd_sc_hd__mux2_1
XFILLER_155_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3481_ _3534_/A _3543_/A VGND VGND VPWR VPWR _4082_/A sky130_fd_sc_hd__nor2_8
X_5220_ hold353/X _5578_/A0 _5222_/S VGND VGND VPWR VPWR _5220_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5151_ _5151_/A _5151_/B _5150_/X VGND VGND VPWR VPWR _5155_/B sky130_fd_sc_hd__or3b_1
XFILLER_69_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5082_ _4581_/B _4987_/X _4950_/A _4411_/Y _4846_/X VGND VGND VPWR VPWR _5117_/A
+ sky130_fd_sc_hd__a2111o_2
XFILLER_111_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4102_ _5545_/A0 _4102_/A1 _4102_/S VGND VGND VPWR VPWR _4102_/X sky130_fd_sc_hd__mux2_1
X_4033_ _5602_/A0 hold319/X _4033_/S VGND VGND VPWR VPWR _4033_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5984_ _7188_/Q _6309_/S _5982_/X _5983_/X VGND VGND VPWR VPWR _7188_/D sky130_fd_sc_hd__o22a_1
Xclkbuf_3_7_0_csclk clkbuf_3_7_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_7_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
X_4935_ _4802_/A _5102_/D _4935_/C _4935_/D VGND VGND VPWR VPWR _4941_/C sky130_fd_sc_hd__nand4b_1
XANTENNA_11 _4030_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4866_ _5013_/A _4922_/A _5086_/A _4866_/D VGND VGND VPWR VPWR _4866_/X sky130_fd_sc_hd__or4_1
XANTENNA_22 _5203_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_33 _7112_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4797_ _5116_/A _4797_/B _4797_/C _4797_/D VGND VGND VPWR VPWR _4798_/D sky130_fd_sc_hd__or4_1
X_6605_ _6777_/CLK _6605_/D _6454_/A VGND VGND VPWR VPWR _6605_/Q sky130_fd_sc_hd__dfrtp_2
X_3817_ _3840_/S _3817_/B VGND VGND VPWR VPWR _3817_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_66 _4234_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_55 _3978_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_44 _5477_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_77 _5245_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3748_ _6609_/Q _4136_/A _3511_/Y _6614_/Q VGND VGND VPWR VPWR _3748_/X sky130_fd_sc_hd__a22o_1
XANTENNA_99 _3725_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6536_ _6786_/CLK _6536_/D fanout417/X VGND VGND VPWR VPWR _6536_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_88 _3606_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3679_ _7118_/Q _5558_/A _4160_/A _6630_/Q VGND VGND VPWR VPWR _3679_/X sky130_fd_sc_hd__a22o_1
X_6467_ _6668_/CLK _6467_/D _6422_/X VGND VGND VPWR VPWR _6467_/Q sky130_fd_sc_hd__dfrtp_2
X_6398_ _6707_/Q _6398_/A2 _6398_/B1 _6706_/Q VGND VGND VPWR VPWR _6398_/X sky130_fd_sc_hd__a22o_1
X_5418_ hold136/X hold220/X _5422_/S VGND VGND VPWR VPWR _6992_/D sky130_fd_sc_hd__mux2_1
Xoutput195 _3212_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[28] sky130_fd_sc_hd__buf_8
Xoutput184 _3222_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[18] sky130_fd_sc_hd__buf_8
X_5349_ _5601_/A0 hold545/X _5350_/S VGND VGND VPWR VPWR _5349_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput173 _3972_/X VGND VGND VPWR VPWR irq[1] sky130_fd_sc_hd__buf_8
XFILLER_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7019_ _7104_/CLK _7019_/D fanout434/X VGND VGND VPWR VPWR _7019_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_55_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _4706_/X _4713_/X _4917_/B VGND VGND VPWR VPWR _4720_/X sky130_fd_sc_hd__o21a_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4651_ _4728_/A _4651_/B VGND VGND VPWR VPWR _4652_/B sky130_fd_sc_hd__nor2_8
XFILLER_159_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3602_ _7144_/Q _5585_/A _4118_/A _6597_/Q VGND VGND VPWR VPWR _3602_/X sky130_fd_sc_hd__a22o_1
Xinput31 mask_rev_in[5] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__clkbuf_4
XFILLER_30_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput20 mask_rev_in[24] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__clkbuf_4
Xinput53 mgmt_gpio_in[25] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__clkbuf_4
Xinput64 mgmt_gpio_in[35] VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__buf_4
Xinput42 mgmt_gpio_in[15] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__clkbuf_4
X_4582_ _4988_/A _4749_/C VGND VGND VPWR VPWR _5174_/A sky130_fd_sc_hd__nor2_1
Xinput97 usr2_vcc_pwrgood VGND VGND VPWR VPWR input97/X sky130_fd_sc_hd__buf_6
Xhold837 _6921_/Q VGND VGND VPWR VPWR hold837/X sky130_fd_sc_hd__bufbuf_16
Xinput86 spimemio_flash_io0_oeb VGND VGND VPWR VPWR _3959_/B sky130_fd_sc_hd__buf_8
Xhold815 _6628_/Q VGND VGND VPWR VPWR hold815/X sky130_fd_sc_hd__bufbuf_16
XFILLER_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold826 _5561_/X VGND VGND VPWR VPWR _7119_/D sky130_fd_sc_hd__bufbuf_16
X_3533_ _3533_/A _3533_/B _3533_/C VGND VGND VPWR VPWR _3547_/C sky130_fd_sc_hd__or3_1
Xinput75 porb VGND VGND VPWR VPWR input75/X sky130_fd_sc_hd__clkbuf_4
Xhold804 _6652_/Q VGND VGND VPWR VPWR hold804/X sky130_fd_sc_hd__bufbuf_16
X_6321_ _6321_/A _6321_/B _6321_/C _6321_/D VGND VGND VPWR VPWR _6321_/X sky130_fd_sc_hd__or4_1
X_6252_ _6758_/Q _6010_/Y _6023_/D _6753_/Q _6251_/X VGND VGND VPWR VPWR _6257_/C
+ sky130_fd_sc_hd__a221o_1
Xhold859 _7103_/Q VGND VGND VPWR VPWR hold859/X sky130_fd_sc_hd__bufbuf_16
X_3464_ hold53/X _3528_/B VGND VGND VPWR VPWR _4190_/A sky130_fd_sc_hd__nor2_8
Xhold848 _4235_/X VGND VGND VPWR VPWR _6688_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_170_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6183_ _6858_/Q _6060_/B _6170_/X _6182_/X _3197_/Y VGND VGND VPWR VPWR _6183_/X
+ sky130_fd_sc_hd__o221a_4
X_5203_ _6409_/A0 _5203_/A1 _5206_/S VGND VGND VPWR VPWR _5203_/X sky130_fd_sc_hd__mux2_1
X_5134_ _5077_/Y _5120_/X _5133_/Y _5112_/X VGND VGND VPWR VPWR _6782_/D sky130_fd_sc_hd__a211o_4
X_3395_ _6867_/Q hold28/A _3334_/Y _7043_/Q _3394_/X VGND VGND VPWR VPWR _3398_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_123_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5065_ _5065_/A _5130_/B VGND VGND VPWR VPWR _5124_/B sky130_fd_sc_hd__nor2_4
X_4016_ hold943/X _4015_/X _4024_/S VGND VGND VPWR VPWR _4016_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5967_ _6567_/Q _5694_/X _5706_/X _6653_/Q VGND VGND VPWR VPWR _5967_/X sky130_fd_sc_hd__a22o_1
XFILLER_25_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4918_ _5069_/B _5132_/A VGND VGND VPWR VPWR _5102_/D sky130_fd_sc_hd__nor2_4
XFILLER_21_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5898_ _6610_/Q _5705_/X _5707_/X _6759_/Q VGND VGND VPWR VPWR _5898_/X sky130_fd_sc_hd__a22o_1
X_4849_ _4849_/A _5071_/A VGND VGND VPWR VPWR _5081_/B sky130_fd_sc_hd__or2_1
XFILLER_180_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6519_ _7130_/CLK _6519_/D fanout452/X VGND VGND VPWR VPWR _6519_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_106_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7172__460 VGND VGND VPWR VPWR _7172_/D _7172__460/LO sky130_fd_sc_hd__conb_1
XFILLER_188_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6870_ _7121_/CLK _6870_/D _6421_/A VGND VGND VPWR VPWR _6870_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_81_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5821_ _6962_/Q _5673_/X _5681_/X _6922_/Q _5820_/X VGND VGND VPWR VPWR _5826_/B
+ sky130_fd_sc_hd__a221o_4
XFILLER_62_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5752_ _6863_/Q _5700_/X _5705_/X _6943_/Q _5751_/X VGND VGND VPWR VPWR _5753_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_188_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4703_ _4773_/A _4930_/C _4773_/B VGND VGND VPWR VPWR _4772_/C sky130_fd_sc_hd__and3b_2
XFILLER_187_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5683_ _7165_/Q _5705_/B _5707_/C VGND VGND VPWR VPWR _5683_/X sky130_fd_sc_hd__and3_4
X_4634_ _4845_/A _4634_/B VGND VGND VPWR VPWR _5144_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold601 _7128_/Q VGND VGND VPWR VPWR hold601/X sky130_fd_sc_hd__bufbuf_16
X_4565_ _4566_/A _4740_/B VGND VGND VPWR VPWR _4565_/Y sky130_fd_sc_hd__nor2_4
Xhold612 _4264_/X VGND VGND VPWR VPWR _6719_/D sky130_fd_sc_hd__bufbuf_16
Xhold645 _7115_/Q VGND VGND VPWR VPWR hold645/X sky130_fd_sc_hd__bufbuf_16
X_6304_ _6715_/Q _6023_/B _6021_/C _6547_/Q _6303_/X VGND VGND VPWR VPWR _6305_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold623 _5367_/X VGND VGND VPWR VPWR _6947_/D sky130_fd_sc_hd__bufbuf_16
X_3516_ _6772_/Q _4322_/A _5194_/A _6804_/Q VGND VGND VPWR VPWR _3516_/X sky130_fd_sc_hd__a22o_2
Xhold634 _7098_/Q VGND VGND VPWR VPWR hold634/X sky130_fd_sc_hd__bufbuf_16
X_4496_ _4819_/B _4724_/A VGND VGND VPWR VPWR _4745_/B sky130_fd_sc_hd__or2_4
XFILLER_116_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold667 _7090_/Q VGND VGND VPWR VPWR hold667/X sky130_fd_sc_hd__bufbuf_16
Xhold656 _5483_/X VGND VGND VPWR VPWR _7050_/D sky130_fd_sc_hd__bufbuf_16
Xhold678 _6578_/Q VGND VGND VPWR VPWR hold678/X sky130_fd_sc_hd__bufbuf_16
XFILLER_104_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold689 _6651_/Q VGND VGND VPWR VPWR hold689/X sky130_fd_sc_hd__bufbuf_16
X_3447_ _7018_/Q _3359_/Y _5396_/A _6978_/Q _3446_/X VGND VGND VPWR VPWR _3450_/C
+ sky130_fd_sc_hd__a221o_1
X_6235_ _7196_/Q _5665_/Y _6233_/X _6234_/X VGND VGND VPWR VPWR _7196_/D sky130_fd_sc_hd__o22a_1
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6166_ _7002_/Q _5987_/Y _6022_/D _6922_/Q VGND VGND VPWR VPWR _6166_/X sky130_fd_sc_hd__a22o_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3378_ _3378_/A _3378_/B _3378_/C _3378_/D VGND VGND VPWR VPWR _3379_/C sky130_fd_sc_hd__or4_2
X_6097_ _7111_/Q _6027_/B _6021_/B _7151_/Q VGND VGND VPWR VPWR _6097_/X sky130_fd_sc_hd__a22o_1
X_5117_ _5117_/A _5117_/B VGND VGND VPWR VPWR _5120_/C sky130_fd_sc_hd__or2_2
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5048_ _5048_/A _5151_/B VGND VGND VPWR VPWR _5056_/A sky130_fd_sc_hd__or2_1
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6999_ _7134_/CLK hold49/X fanout429/X VGND VGND VPWR VPWR _6999_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_159_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4350_ _4350_/A _4350_/B _4350_/C _4350_/D VGND VGND VPWR VPWR _4352_/B sky130_fd_sc_hd__and4_1
X_3301_ _3506_/A _3673_/B VGND VGND VPWR VPWR _5450_/A sky130_fd_sc_hd__nor2_8
X_4281_ _5289_/A0 hold905/X _4285_/S VGND VGND VPWR VPWR _4281_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6020_ _6020_/A _6020_/B _6020_/C _6020_/D VGND VGND VPWR VPWR _6024_/A sky130_fd_sc_hd__or4_1
X_3232_ _6920_/Q VGND VGND VPWR VPWR _3232_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6922_ _7130_/CLK _6922_/D fanout452/X VGND VGND VPWR VPWR _6922_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_82_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6853_ _7140_/CLK _6853_/D fanout430/X VGND VGND VPWR VPWR _6853_/Q sky130_fd_sc_hd__dfstp_4
X_5804_ _7065_/Q _5669_/X _5687_/X _7049_/Q VGND VGND VPWR VPWR _5804_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6784_ _7208_/CLK _6784_/D fanout458/X VGND VGND VPWR VPWR _6784_/Q sky130_fd_sc_hd__dfrtp_2
X_3996_ _3996_/A0 _5234_/C _4003_/S VGND VGND VPWR VPWR _6496_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5735_ _6910_/Q _5680_/X _5700_/X _6862_/Q _5726_/X VGND VGND VPWR VPWR _5735_/X
+ sky130_fd_sc_hd__a221o_1
X_5666_ _7161_/Q _7162_/Q VGND VGND VPWR VPWR _5704_/B sky130_fd_sc_hd__and2b_4
XFILLER_129_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4617_ _4617_/A _4989_/A VGND VGND VPWR VPWR _4617_/Y sky130_fd_sc_hd__nor2_2
X_5597_ _5597_/A0 hold533/X _5602_/S VGND VGND VPWR VPWR _5597_/X sky130_fd_sc_hd__mux2_1
Xhold420 _7070_/Q VGND VGND VPWR VPWR hold420/X sky130_fd_sc_hd__bufbuf_16
Xhold431 _7063_/Q VGND VGND VPWR VPWR hold431/X sky130_fd_sc_hd__bufbuf_16
Xhold442 _6938_/Q VGND VGND VPWR VPWR hold442/X sky130_fd_sc_hd__bufbuf_16
XFILLER_145_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4548_ _5081_/A _4849_/A _4548_/C _4548_/D VGND VGND VPWR VPWR _4548_/X sky130_fd_sc_hd__or4_1
XFILLER_104_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold453 _6759_/Q VGND VGND VPWR VPWR hold453/X sky130_fd_sc_hd__bufbuf_16
Xhold464 _7154_/Q VGND VGND VPWR VPWR hold464/X sky130_fd_sc_hd__bufbuf_16
X_4479_ _4775_/A _4636_/A VGND VGND VPWR VPWR _4766_/A sky130_fd_sc_hd__nor2_2
XFILLER_104_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold486 _7076_/Q VGND VGND VPWR VPWR hold486/X sky130_fd_sc_hd__bufbuf_16
Xhold475 _5440_/X VGND VGND VPWR VPWR _7012_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6218_ _6988_/Q _6028_/X _6034_/Y _6996_/Q _6217_/X VGND VGND VPWR VPWR _6219_/D
+ sky130_fd_sc_hd__a221o_2
Xhold497 _6754_/Q VGND VGND VPWR VPWR hold497/X sky130_fd_sc_hd__bufbuf_16
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7198_ _7201_/CLK _7198_/D _6446_/A VGND VGND VPWR VPWR _7198_/Q sky130_fd_sc_hd__dfrtp_1
Xhold1131 _7143_/Q VGND VGND VPWR VPWR _5588_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1120 _4293_/X VGND VGND VPWR VPWR _6743_/D sky130_fd_sc_hd__bufbuf_16
X_6149_ _6905_/Q _6021_/A _6025_/A _6937_/Q _6148_/X VGND VGND VPWR VPWR _6156_/A
+ sky130_fd_sc_hd__a221o_2
Xhold1142 _6649_/Q VGND VGND VPWR VPWR _4185_/A0 sky130_fd_sc_hd__bufbuf_16
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1153 _5336_/X VGND VGND VPWR VPWR _6919_/D sky130_fd_sc_hd__bufbuf_16
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1164 _4251_/X VGND VGND VPWR VPWR _6708_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_58_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1175 _6728_/Q VGND VGND VPWR VPWR _4275_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_45_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_304 input46/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_315 input169/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1197 _5195_/X VGND VGND VPWR VPWR _6800_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_26_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1186 _5186_/X VGND VGND VPWR VPWR _6785_/D sky130_fd_sc_hd__bufbuf_16
XANTENNA_359 hold335/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_348 hold209/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_337 hold43/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_326 _5545_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3850_ _6470_/Q _3797_/X _6472_/Q VGND VGND VPWR VPWR _3850_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_177_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3781_ input20/X _3302_/Y _3320_/Y input34/X VGND VGND VPWR VPWR _3781_/X sky130_fd_sc_hd__a22o_2
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5520_ _5583_/A0 hold713/X _5521_/S VGND VGND VPWR VPWR _5520_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5451_ _5541_/A0 _5451_/A1 _5458_/S VGND VGND VPWR VPWR _7021_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5382_ hold71/X hold295/X _5386_/S VGND VGND VPWR VPWR _5382_/X sky130_fd_sc_hd__mux2_1
X_4402_ _4553_/B _4410_/C _4513_/A VGND VGND VPWR VPWR _4995_/A sky130_fd_sc_hd__or3_4
X_7121_ _7121_/CLK _7121_/D fanout442/X VGND VGND VPWR VPWR _7121_/Q sky130_fd_sc_hd__dfrtp_2
X_4333_ _5545_/A0 _4333_/A1 _4333_/S VGND VGND VPWR VPWR _4333_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4264_ hold611/X _6408_/A0 _4267_/S VGND VGND VPWR VPWR _4264_/X sky130_fd_sc_hd__mux2_1
X_7052_ _7124_/CLK _7052_/D fanout436/X VGND VGND VPWR VPWR _7052_/Q sky130_fd_sc_hd__dfrtp_2
X_3215_ _7056_/Q VGND VGND VPWR VPWR _3215_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6003_ _6037_/B _6033_/C _6018_/A VGND VGND VPWR VPWR _6021_/C sky130_fd_sc_hd__and3_4
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4195_ _6411_/A0 hold731/X _4195_/S VGND VGND VPWR VPWR _4195_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6905_ _6959_/CLK _6905_/D fanout442/X VGND VGND VPWR VPWR _6905_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_82_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6836_ _6964_/CLK _6836_/D fanout444/X VGND VGND VPWR VPWR _6836_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6767_ _6840_/CLK _6767_/D fanout424/X VGND VGND VPWR VPWR _6767_/Q sky130_fd_sc_hd__dfrtp_2
X_3979_ _3875_/B hold883/X _3979_/S VGND VGND VPWR VPWR _3979_/X sky130_fd_sc_hd__mux2_8
XFILLER_148_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5718_ _7037_/Q _5683_/X _5699_/X _6925_/Q _5717_/X VGND VGND VPWR VPWR _5720_/C
+ sky130_fd_sc_hd__a221o_2
X_6698_ _7220_/CLK _6698_/D _6362_/B VGND VGND VPWR VPWR _6698_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_156_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5649_ _7170_/Q _5654_/A VGND VGND VPWR VPWR _5649_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold250 _7089_/Q VGND VGND VPWR VPWR hold250/X sky130_fd_sc_hd__bufbuf_16
Xhold261 _5403_/X VGND VGND VPWR VPWR _6979_/D sky130_fd_sc_hd__bufbuf_16
Xhold283 _6969_/Q VGND VGND VPWR VPWR hold283/X sky130_fd_sc_hd__bufbuf_16
XFILLER_104_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold272 _5482_/X VGND VGND VPWR VPWR _7049_/D sky130_fd_sc_hd__bufbuf_16
Xhold294 _5257_/X VGND VGND VPWR VPWR _6849_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_172_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 _5680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_112 _3857_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_123 _5251_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_101 _3792_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_167 _6020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_145 _5703_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 _5734_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_189 _6221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_178 _6060_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_1_1_1_csclk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_155_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput7 mask_rev_in[12] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4951_ _4949_/B _4536_/B _4959_/A _4903_/A VGND VGND VPWR VPWR _5148_/A sky130_fd_sc_hd__a31o_1
XFILLER_91_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4882_ _4736_/B _4758_/B _4657_/B _4581_/B _4987_/A VGND VGND VPWR VPWR _4903_/C
+ sky130_fd_sc_hd__a32o_2
X_3902_ _7166_/Q _7167_/Q VGND VGND VPWR VPWR _6012_/A sky130_fd_sc_hd__and2b_4
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6621_ _6649_/CLK _6621_/D fanout456/X VGND VGND VPWR VPWR _6621_/Q sky130_fd_sc_hd__dfstp_2
X_3833_ hold16/A hold80/A hold24/A VGND VGND VPWR VPWR _3833_/X sky130_fd_sc_hd__a21o_1
XFILLER_60_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6552_ _6725_/CLK _6552_/D fanout440/X VGND VGND VPWR VPWR _6552_/Q sky130_fd_sc_hd__dfstp_4
X_3764_ _3764_/A _3764_/B _3764_/C _3764_/D VGND VGND VPWR VPWR _3764_/X sky130_fd_sc_hd__or4_4
XFILLER_118_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5503_ _5602_/A0 hold484/X _5503_/S VGND VGND VPWR VPWR _5503_/X sky130_fd_sc_hd__mux2_1
X_3695_ _7070_/Q hold92/A _4292_/A _6744_/Q VGND VGND VPWR VPWR _3695_/X sky130_fd_sc_hd__a22o_2
X_6483_ _6668_/CLK _6483_/D _6438_/X VGND VGND VPWR VPWR hold50/A sky130_fd_sc_hd__dfrtp_2
XFILLER_160_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput300 _6489_/Q VGND VGND VPWR VPWR pll_trim[9] sky130_fd_sc_hd__buf_8
X_5434_ _5578_/A0 hold448/X _5440_/S VGND VGND VPWR VPWR _7006_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput333 _6562_/Q VGND VGND VPWR VPWR wb_dat_o[23] sky130_fd_sc_hd__buf_8
XFILLER_126_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput322 _6573_/Q VGND VGND VPWR VPWR wb_dat_o[13] sky130_fd_sc_hd__buf_8
Xoutput344 _6585_/Q VGND VGND VPWR VPWR wb_dat_o[4] sky130_fd_sc_hd__buf_8
Xoutput311 _3951_/X VGND VGND VPWR VPWR serial_resetn sky130_fd_sc_hd__buf_8
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_3_0_csclk clkbuf_3_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_3_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
X_5365_ hold185/X hold237/X _5368_/S VGND VGND VPWR VPWR _5365_/X sky130_fd_sc_hd__mux2_1
X_7104_ _7104_/CLK _7104_/D fanout434/X VGND VGND VPWR VPWR _7104_/Q sky130_fd_sc_hd__dfrtp_2
X_5296_ _5602_/A0 hold377/X _5296_/S VGND VGND VPWR VPWR _5296_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4316_ _4316_/A _6406_/B VGND VGND VPWR VPWR _4321_/S sky130_fd_sc_hd__and2_4
X_4247_ hold7/X _4247_/A1 _4249_/S VGND VGND VPWR VPWR hold8/A sky130_fd_sc_hd__mux2_1
X_7035_ _7035_/CLK _7035_/D fanout432/X VGND VGND VPWR VPWR _7035_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_19_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4178_ _4178_/A hold47/X VGND VGND VPWR VPWR _4183_/S sky130_fd_sc_hd__and2_4
XFILLER_67_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6819_ _7134_/CLK _6819_/D fanout429/X VGND VGND VPWR VPWR _6819_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_51_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3480_ _3543_/A _5252_/B VGND VGND VPWR VPWR _4118_/A sky130_fd_sc_hd__nor2_8
XFILLER_170_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5150_ _4947_/B _4832_/B _5050_/C _4832_/A _4835_/X VGND VGND VPWR VPWR _5150_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_111_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5081_ _5081_/A _5081_/B _5081_/C _4623_/A VGND VGND VPWR VPWR _5115_/A sky130_fd_sc_hd__or4b_2
X_4101_ _4326_/A0 hold780/X _4102_/S VGND VGND VPWR VPWR _4101_/X sky130_fd_sc_hd__mux2_1
X_4032_ _5601_/A0 hold537/X _4033_/S VGND VGND VPWR VPWR _4032_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5983_ _5611_/A _7187_/Q _6358_/B1 VGND VGND VPWR VPWR _5983_/X sky130_fd_sc_hd__a21o_1
XFILLER_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4934_ _4398_/Y _5023_/B _5062_/C _4933_/Y VGND VGND VPWR VPWR _4935_/C sky130_fd_sc_hd__o22a_1
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_12 _4033_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4865_ _5118_/B _4865_/B _4865_/C VGND VGND VPWR VPWR _4866_/D sky130_fd_sc_hd__or3_1
XANTENNA_23 _6822_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 _5571_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6604_ _6649_/CLK _6604_/D fanout439/X VGND VGND VPWR VPWR _6604_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_56 _5585_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4796_ _5140_/B _4796_/B _4796_/C _4796_/D VGND VGND VPWR VPWR _4797_/D sky130_fd_sc_hd__or4_1
XANTENNA_45 _5486_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3816_ _3255_/X _3256_/Y _3820_/B VGND VGND VPWR VPWR _3817_/B sky130_fd_sc_hd__mux2_1
XANTENNA_78 _5245_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3747_ _6861_/Q hold28/A _5306_/A _6893_/Q _3746_/X VGND VGND VPWR VPWR _3754_/A
+ sky130_fd_sc_hd__a221o_2
XANTENNA_67 _5396_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_89 _3606_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6535_ _6777_/CLK _6535_/D fanout424/X VGND VGND VPWR VPWR _6535_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6466_ _3938_/A1 _6466_/D _6421_/X VGND VGND VPWR VPWR hold9/A sky130_fd_sc_hd__dfrtp_2
XFILLER_173_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3678_ _6831_/Q _5227_/A _4298_/A _6749_/Q VGND VGND VPWR VPWR _3678_/X sky130_fd_sc_hd__a22o_1
X_6397_ _6396_/X _7217_/Q _6400_/S VGND VGND VPWR VPWR _7217_/D sky130_fd_sc_hd__mux2_1
X_5417_ _5561_/A0 hold676/X _5422_/S VGND VGND VPWR VPWR _5417_/X sky130_fd_sc_hd__mux2_1
Xoutput185 _3221_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[19] sky130_fd_sc_hd__buf_8
X_5348_ _5600_/A0 hold374/X _5350_/S VGND VGND VPWR VPWR _5348_/X sky130_fd_sc_hd__mux2_1
Xoutput174 _3973_/X VGND VGND VPWR VPWR irq[2] sky130_fd_sc_hd__buf_8
Xoutput196 _3211_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[29] sky130_fd_sc_hd__buf_8
XFILLER_87_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5279_ _5279_/A _5558_/B VGND VGND VPWR VPWR _5287_/S sky130_fd_sc_hd__nand2_8
XFILLER_87_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7018_ _7104_/CLK _7018_/D fanout434/X VGND VGND VPWR VPWR _7018_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_47_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout390 _5300_/A0 VGND VGND VPWR VPWR _5588_/A0 sky130_fd_sc_hd__buf_8
XFILLER_19_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4650_ _4722_/B _4650_/B VGND VGND VPWR VPWR _5062_/B sky130_fd_sc_hd__or2_4
XFILLER_175_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3601_ _7024_/Q _5450_/A _4328_/A _6776_/Q _3561_/X VGND VGND VPWR VPWR _3605_/C
+ sky130_fd_sc_hd__a221o_1
Xinput10 mask_rev_in[15] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__clkbuf_4
Xinput21 mask_rev_in[25] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__clkbuf_4
XFILLER_190_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput54 mgmt_gpio_in[26] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__clkbuf_4
X_4581_ _4987_/A _4581_/B VGND VGND VPWR VPWR _4612_/B sky130_fd_sc_hd__nand2_1
Xinput43 mgmt_gpio_in[16] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__clkbuf_4
X_6320_ _6627_/Q _6028_/X _6034_/Y _6726_/Q _6319_/X VGND VGND VPWR VPWR _6321_/D
+ sky130_fd_sc_hd__a221o_2
Xinput32 mask_rev_in[6] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__clkbuf_4
Xinput98 usr2_vdd_pwrgood VGND VGND VPWR VPWR input98/X sky130_fd_sc_hd__buf_6
Xhold827 _6897_/Q VGND VGND VPWR VPWR hold827/X sky130_fd_sc_hd__bufbuf_16
Xinput87 spimemio_flash_io1_do VGND VGND VPWR VPWR _7227_/A sky130_fd_sc_hd__buf_8
Xhold816 _4159_/X VGND VGND VPWR VPWR _6628_/D sky130_fd_sc_hd__bufbuf_16
Xinput65 mgmt_gpio_in[36] VGND VGND VPWR VPWR _7228_/A sky130_fd_sc_hd__buf_4
XFILLER_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3532_ _7097_/Q _3341_/Y _4097_/A _6580_/Q _3530_/X VGND VGND VPWR VPWR _3533_/C
+ sky130_fd_sc_hd__a221o_1
Xhold805 _4188_/X VGND VGND VPWR VPWR _6652_/D sky130_fd_sc_hd__bufbuf_16
Xinput76 qspi_enabled VGND VGND VPWR VPWR _3932_/S sky130_fd_sc_hd__buf_8
Xhold838 _5338_/X VGND VGND VPWR VPWR _6921_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_170_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold849 _6953_/Q VGND VGND VPWR VPWR hold849/X sky130_fd_sc_hd__bufbuf_16
X_6251_ _6619_/Q _6022_/C _6033_/X _6738_/Q VGND VGND VPWR VPWR _6251_/X sky130_fd_sc_hd__a22o_1
XFILLER_89_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3463_ _6905_/Q _5315_/A _4256_/A _6717_/Q _3461_/X VGND VGND VPWR VPWR _3472_/B
+ sky130_fd_sc_hd__a221o_1
X_6182_ _6306_/A _6182_/B _6182_/C VGND VGND VPWR VPWR _6182_/X sky130_fd_sc_hd__or3_4
XFILLER_88_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5202_ _5254_/A0 hold919/X _5206_/S VGND VGND VPWR VPWR _6806_/D sky130_fd_sc_hd__mux2_1
X_5133_ _5133_/A _5133_/B VGND VGND VPWR VPWR _5133_/Y sky130_fd_sc_hd__nor2_2
X_3394_ _7059_/Q _5486_/A _5423_/A _7003_/Q VGND VGND VPWR VPWR _3394_/X sky130_fd_sc_hd__a22o_1
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5064_ _4949_/C _4748_/A _4657_/B _4903_/C _4846_/B VGND VGND VPWR VPWR _5130_/B
+ sky130_fd_sc_hd__a311o_4
XFILLER_123_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4015_ hold715/X _5571_/A0 _4023_/S VGND VGND VPWR VPWR _4015_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5966_ _6613_/Q _5705_/X _5707_/X _6762_/Q VGND VGND VPWR VPWR _5981_/B sky130_fd_sc_hd__a22o_1
XFILLER_12_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4917_ _4917_/A _4917_/B _5003_/C VGND VGND VPWR VPWR _5102_/C sky130_fd_sc_hd__and3_2
X_5897_ _6645_/Q _5685_/X _5699_/X _6600_/Q VGND VGND VPWR VPWR _5897_/X sky130_fd_sc_hd__a22o_1
XFILLER_40_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4848_ _4845_/A _4634_/B _4920_/A VGND VGND VPWR VPWR _5136_/C sky130_fd_sc_hd__a21o_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4779_ _4724_/B _4757_/B _5081_/A VGND VGND VPWR VPWR _4799_/A sky130_fd_sc_hd__o21bai_1
X_6518_ _7152_/CLK _6518_/D fanout452/X VGND VGND VPWR VPWR _6518_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_180_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6449_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6449_/X sky130_fd_sc_hd__and2_1
XFILLER_134_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_40_csclk _7137_/CLK VGND VGND VPWR VPWR _6874_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_0_0_csclk clkbuf_2_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_1_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_102_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_55_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7123_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_113_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5820_ _6970_/Q _5691_/X _5701_/X _6954_/Q VGND VGND VPWR VPWR _5820_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5751_ _7031_/Q _5688_/X _5693_/X _7079_/Q VGND VGND VPWR VPWR _5751_/X sky130_fd_sc_hd__a22o_2
XFILLER_62_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4702_ _4702_/A _4702_/B VGND VGND VPWR VPWR _4773_/B sky130_fd_sc_hd__or2_1
XFILLER_147_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5682_ _7165_/Q _5702_/B _5707_/C VGND VGND VPWR VPWR _5682_/X sky130_fd_sc_hd__and3_4
XFILLER_175_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4633_ _4986_/A _4996_/A VGND VGND VPWR VPWR _4633_/X sky130_fd_sc_hd__or2_2
X_4564_ _4564_/A _4672_/A VGND VGND VPWR VPWR _4740_/B sky130_fd_sc_hd__nand2_8
Xhold602 _5571_/X VGND VGND VPWR VPWR _7128_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_128_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold624 _6939_/Q VGND VGND VPWR VPWR hold624/X sky130_fd_sc_hd__bufbuf_16
X_6303_ _6661_/Q _5996_/X _6020_/C _6591_/Q VGND VGND VPWR VPWR _6303_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold613 _6493_/Q VGND VGND VPWR VPWR hold613/X sky130_fd_sc_hd__bufbuf_16
X_3515_ _5234_/A _3515_/B VGND VGND VPWR VPWR _5194_/A sky130_fd_sc_hd__nor2_8
Xhold635 _5537_/X VGND VGND VPWR VPWR _7098_/D sky130_fd_sc_hd__bufbuf_16
X_4495_ _4651_/B _4707_/B _5050_/A VGND VGND VPWR VPWR _4724_/A sky130_fd_sc_hd__or3b_4
Xhold657 _6551_/Q VGND VGND VPWR VPWR hold657/X sky130_fd_sc_hd__bufbuf_16
Xhold646 _5556_/X VGND VGND VPWR VPWR _7115_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_131_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold668 _5528_/X VGND VGND VPWR VPWR _7090_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_89_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold679 _6817_/Q VGND VGND VPWR VPWR hold679/X sky130_fd_sc_hd__bufbuf_16
X_6234_ _5663_/A _7195_/Q _5664_/X VGND VGND VPWR VPWR _6234_/X sky130_fd_sc_hd__a21o_1
XFILLER_103_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3446_ _6930_/Q _5342_/A _5200_/A _6810_/Q VGND VGND VPWR VPWR _3446_/X sky130_fd_sc_hd__a22o_1
XFILLER_112_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3377_ _3377_/A _3377_/B _3377_/C _3377_/D VGND VGND VPWR VPWR _3378_/D sky130_fd_sc_hd__or4_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _7018_/Q _6036_/Y _6335_/B _7042_/Q _6162_/X VGND VGND VPWR VPWR _6170_/B
+ sky130_fd_sc_hd__a221o_4
X_5116_ _5116_/A _5116_/B _5116_/C _4881_/A VGND VGND VPWR VPWR _5117_/B sky130_fd_sc_hd__or4b_1
X_6096_ _7079_/Q _6311_/B _6091_/X _6093_/X _6095_/X VGND VGND VPWR VPWR _6096_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_85_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5047_ _5047_/A _5047_/B _5047_/C _5047_/D VGND VGND VPWR VPWR _5151_/B sky130_fd_sc_hd__or4_1
XFILLER_85_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6998_ _7134_/CLK _6998_/D fanout429/X VGND VGND VPWR VPWR _6998_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_41_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5949_ _6548_/Q _5674_/X _5688_/X _6771_/Q VGND VGND VPWR VPWR _5949_/X sky130_fd_sc_hd__a22o_1
XFILLER_41_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3300_ _7060_/Q _5486_/A _3299_/Y _6996_/Q VGND VGND VPWR VPWR _3300_/X sky130_fd_sc_hd__a22o_1
X_4280_ _4280_/A _5486_/B VGND VGND VPWR VPWR _4285_/S sky130_fd_sc_hd__nand2_8
XFILLER_140_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3231_ _6928_/Q VGND VGND VPWR VPWR _3231_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_634 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6921_ _7121_/CLK _6921_/D fanout442/X VGND VGND VPWR VPWR _6921_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6852_ _7107_/CLK _6852_/D fanout434/X VGND VGND VPWR VPWR _6852_/Q sky130_fd_sc_hd__dfrtp_1
X_5803_ _7105_/Q _5675_/X _5683_/X _7041_/Q _5802_/X VGND VGND VPWR VPWR _5806_/C
+ sky130_fd_sc_hd__a221o_1
X_6783_ _7208_/CLK _6783_/D fanout458/X VGND VGND VPWR VPWR _6783_/Q sky130_fd_sc_hd__dfrtp_2
X_3995_ _3995_/A _6406_/B VGND VGND VPWR VPWR _4003_/S sky130_fd_sc_hd__and2_4
X_5734_ _5734_/A _5734_/B _5734_/C _5734_/D VGND VGND VPWR VPWR _5734_/X sky130_fd_sc_hd__or4_2
XFILLER_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5665_ _5665_/A _5665_/B VGND VGND VPWR VPWR _5665_/Y sky130_fd_sc_hd__nor2_8
XFILLER_148_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4616_ _4986_/A _4997_/A _5123_/C _4881_/A VGND VGND VPWR VPWR _4619_/C sky130_fd_sc_hd__o211a_1
Xhold410 _5411_/X VGND VGND VPWR VPWR _6986_/D sky130_fd_sc_hd__bufbuf_16
X_5596_ _5596_/A0 hold383/X _5602_/S VGND VGND VPWR VPWR _7150_/D sky130_fd_sc_hd__mux2_1
XFILLER_163_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold432 _5498_/X VGND VGND VPWR VPWR _7063_/D sky130_fd_sc_hd__bufbuf_16
Xhold443 _5357_/X VGND VGND VPWR VPWR _6938_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_145_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4547_ _4986_/B _4988_/A VGND VGND VPWR VPWR _4548_/D sky130_fd_sc_hd__nor2_1
Xhold454 _4312_/X VGND VGND VPWR VPWR _6759_/D sky130_fd_sc_hd__bufbuf_16
Xhold421 _7020_/Q VGND VGND VPWR VPWR hold421/X sky130_fd_sc_hd__bufbuf_16
XFILLER_171_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold465 _5600_/X VGND VGND VPWR VPWR _7154_/D sky130_fd_sc_hd__bufbuf_16
Xhold476 _6970_/Q VGND VGND VPWR VPWR hold476/X sky130_fd_sc_hd__bufbuf_16
X_4478_ _4707_/B _4478_/B _4478_/C VGND VGND VPWR VPWR _4844_/B sky130_fd_sc_hd__or3_4
XFILLER_104_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold487 _5512_/X VGND VGND VPWR VPWR _7076_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_104_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6217_ _7076_/Q _6009_/X _6020_/D _6972_/Q VGND VGND VPWR VPWR _6217_/X sky130_fd_sc_hd__a22o_1
XFILLER_58_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7197_ _7197_/CLK _7197_/D fanout421/X VGND VGND VPWR VPWR _7197_/Q sky130_fd_sc_hd__dfrtp_2
X_3429_ _7042_/Q _3334_/Y _5423_/A _7002_/Q _3428_/X VGND VGND VPWR VPWR _3450_/B
+ sky130_fd_sc_hd__a221o_1
Xhold498 _4306_/X VGND VGND VPWR VPWR _6754_/D sky130_fd_sc_hd__bufbuf_16
X_6148_ _6953_/Q _6022_/A _6025_/C _6929_/Q VGND VGND VPWR VPWR _6148_/X sky130_fd_sc_hd__a22o_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1132 _5588_/X VGND VGND VPWR VPWR _7143_/D sky130_fd_sc_hd__bufbuf_16
Xhold1121 _6550_/Q VGND VGND VPWR VPWR _4068_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1110 _4137_/X VGND VGND VPWR VPWR _6609_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_58_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1143 _4185_/X VGND VGND VPWR VPWR _6649_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_100_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6079_ _6862_/Q _6025_/D _6029_/X _7046_/Q _6078_/X VGND VGND VPWR VPWR _6082_/C
+ sky130_fd_sc_hd__a221o_4
XFILLER_72_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1176 _4275_/X VGND VGND VPWR VPWR _6728_/D sky130_fd_sc_hd__bufbuf_16
Xhold1154 _6634_/Q VGND VGND VPWR VPWR _4167_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1165 _6654_/Q VGND VGND VPWR VPWR _4191_/A1 sky130_fd_sc_hd__bufbuf_16
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1187 _6959_/Q VGND VGND VPWR VPWR _5381_/A1 sky130_fd_sc_hd__bufbuf_16
XANTENNA_305 input43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_316 input169/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1198 _6832_/Q VGND VGND VPWR VPWR _5235_/A1 sky130_fd_sc_hd__bufbuf_16
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_338 hold71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_349 hold209/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_327 _5581_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3780_ _6805_/Q _5200_/A _4166_/A _6634_/Q _3779_/X VGND VGND VPWR VPWR _3785_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_185_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5450_ _5450_/A hold47/X VGND VGND VPWR VPWR _5458_/S sky130_fd_sc_hd__nand2_8
XFILLER_172_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4401_ _4553_/B _4410_/C _4513_/A VGND VGND VPWR VPWR _4575_/B sky130_fd_sc_hd__nor3_4
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5381_ _5588_/A0 _5381_/A1 _5386_/S VGND VGND VPWR VPWR _5381_/X sky130_fd_sc_hd__mux2_1
X_7120_ _7130_/CLK _7120_/D fanout454/X VGND VGND VPWR VPWR _7120_/Q sky130_fd_sc_hd__dfrtp_2
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A VGND VGND VPWR VPWR _7196_/CLK sky130_fd_sc_hd__clkbuf_8
X_4332_ _6410_/A0 _4332_/A1 _4333_/S VGND VGND VPWR VPWR _4332_/X sky130_fd_sc_hd__mux2_1
X_4263_ _4263_/A0 _5289_/A0 _4267_/S VGND VGND VPWR VPWR _4263_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7051_ _7123_/CLK _7051_/D fanout434/X VGND VGND VPWR VPWR _7051_/Q sky130_fd_sc_hd__dfrtp_2
X_3214_ _7064_/Q VGND VGND VPWR VPWR _3214_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6002_ _6019_/A _6010_/B VGND VGND VPWR VPWR _6021_/B sky130_fd_sc_hd__nor2_8
X_4194_ _6410_/A0 hold972/X _4195_/S VGND VGND VPWR VPWR _4194_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6904_ _6976_/CLK _6904_/D fanout450/X VGND VGND VPWR VPWR _6904_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6835_ _6964_/CLK _6835_/D fanout444/X VGND VGND VPWR VPWR _6835_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3978_ _3978_/A hold47/X VGND VGND VPWR VPWR _3994_/S sky130_fd_sc_hd__and2_4
X_6766_ _6851_/CLK _6766_/D fanout418/X VGND VGND VPWR VPWR _6766_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5717_ _6909_/Q _5680_/X _5703_/X _6869_/Q VGND VGND VPWR VPWR _5717_/X sky130_fd_sc_hd__a22o_1
X_6697_ _7127_/CLK hold4/X fanout448/X VGND VGND VPWR VPWR _6697_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5648_ _7170_/Q _5648_/B _6035_/A VGND VGND VPWR VPWR _5654_/B sky130_fd_sc_hd__and3_1
XFILLER_156_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5579_ hold43/X _5579_/A1 hold62/X VGND VGND VPWR VPWR hold63/A sky130_fd_sc_hd__mux2_1
XFILLER_116_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold251 _5527_/X VGND VGND VPWR VPWR _7089_/D sky130_fd_sc_hd__bufbuf_16
Xhold240 _7032_/Q VGND VGND VPWR VPWR hold240/X sky130_fd_sc_hd__bufbuf_16
Xhold262 _6944_/Q VGND VGND VPWR VPWR hold262/X sky130_fd_sc_hd__bufbuf_16
Xhold273 _6674_/Q VGND VGND VPWR VPWR hold273/X sky130_fd_sc_hd__bufbuf_16
XFILLER_172_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold284 _5392_/X VGND VGND VPWR VPWR _6969_/D sky130_fd_sc_hd__bufbuf_16
Xhold295 _6960_/Q VGND VGND VPWR VPWR hold295/X sky130_fd_sc_hd__bufbuf_16
XFILLER_132_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_124 _5251_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 _3879_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_102 _3801_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_135 _5681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_146 _5703_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_157 _5741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 _6025_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_179 _6030_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 mask_rev_in[13] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4950_ _4950_/A _4950_/B _4950_/C VGND VGND VPWR VPWR _5129_/B sky130_fd_sc_hd__or3_4
XFILLER_64_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4881_ _4881_/A _4881_/B VGND VGND VPWR VPWR _4905_/B sky130_fd_sc_hd__nand2_1
X_3901_ _7170_/Q _7171_/Q VGND VGND VPWR VPWR _6019_/A sky130_fd_sc_hd__nand2b_4
X_6620_ _6649_/CLK _6620_/D fanout439/X VGND VGND VPWR VPWR _6620_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_32_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3832_ _3831_/X _6480_/Q _3840_/S VGND VGND VPWR VPWR _6480_/D sky130_fd_sc_hd__mux2_1
X_6551_ _6843_/CLK _6551_/D _6421_/A VGND VGND VPWR VPWR _6551_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3763_ _6885_/Q _5297_/A hold61/A _7133_/Q _3738_/X VGND VGND VPWR VPWR _3764_/D
+ sky130_fd_sc_hd__a221o_1
X_5502_ _5583_/A0 hold693/X _5503_/S VGND VGND VPWR VPWR _5502_/X sky130_fd_sc_hd__mux2_1
X_6482_ _6668_/CLK _6482_/D _6437_/X VGND VGND VPWR VPWR _6482_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_9_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3694_ _6812_/Q _5207_/A hold61/A _7134_/Q _3678_/X VGND VGND VPWR VPWR _3699_/A
+ sky130_fd_sc_hd__a221o_1
Xoutput301 _6820_/Q VGND VGND VPWR VPWR pwr_ctrl_out[0] sky130_fd_sc_hd__buf_8
X_5433_ _5541_/A0 _5433_/A1 _5440_/S VGND VGND VPWR VPWR _7005_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput334 _7203_/Q VGND VGND VPWR VPWR wb_dat_o[24] sky130_fd_sc_hd__buf_8
XFILLER_105_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput323 _6574_/Q VGND VGND VPWR VPWR wb_dat_o[14] sky130_fd_sc_hd__buf_8
X_5364_ hold136/X hold262/X _5368_/S VGND VGND VPWR VPWR _5364_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput312 _3970_/X VGND VGND VPWR VPWR spi_sdi sky130_fd_sc_hd__buf_8
XFILLER_126_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput345 _6586_/Q VGND VGND VPWR VPWR wb_dat_o[5] sky130_fd_sc_hd__buf_8
X_7103_ _7103_/CLK _7103_/D fanout436/X VGND VGND VPWR VPWR _7103_/Q sky130_fd_sc_hd__dfrtp_2
X_4315_ hold763/X _6411_/A0 _4315_/S VGND VGND VPWR VPWR _4315_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5295_ _5601_/A0 hold599/X _5296_/S VGND VGND VPWR VPWR _5295_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4246_ _5599_/A0 hold458/X _4249_/S VGND VGND VPWR VPWR _4246_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7034_ _7131_/CLK _7034_/D fanout432/X VGND VGND VPWR VPWR _7034_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_67_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4177_ hold744/X _6411_/A0 _4177_/S VGND VGND VPWR VPWR _4177_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6818_ _7132_/CLK _6818_/D fanout428/X VGND VGND VPWR VPWR _6818_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_51_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6749_ _6810_/CLK _6749_/D fanout419/X VGND VGND VPWR VPWR _6749_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5080_ _4586_/B _4987_/X _4850_/X _4617_/Y _4798_/A VGND VGND VPWR VPWR _5171_/B
+ sky130_fd_sc_hd__a2111o_1
X_4100_ _5561_/A0 hold678/X _4102_/S VGND VGND VPWR VPWR _6578_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4031_ _5600_/A0 hold384/X _4033_/S VGND VGND VPWR VPWR _4031_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5982_ _6534_/Q _5722_/B _5976_/X _5981_/X _6308_/S VGND VGND VPWR VPWR _5982_/X
+ sky130_fd_sc_hd__o221a_4
X_4933_ _5165_/A _4933_/B VGND VGND VPWR VPWR _4933_/Y sky130_fd_sc_hd__nand2_1
XFILLER_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_13 _4041_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4864_ _4648_/B _5164_/B _4638_/X VGND VGND VPWR VPWR _4865_/C sky130_fd_sc_hd__o21ai_1
XANTENNA_24 _5248_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6603_ _6725_/CLK _6603_/D fanout440/X VGND VGND VPWR VPWR _6603_/Q sky130_fd_sc_hd__dfrtp_2
X_4795_ _4772_/A _5165_/A _4428_/C _4794_/X VGND VGND VPWR VPWR _4796_/D sky130_fd_sc_hd__a31o_1
XANTENNA_46 _5486_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_57 _5585_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_35 _3191_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3815_ hold50/A _6482_/Q _6481_/Q _3828_/S VGND VGND VPWR VPWR _3820_/B sky130_fd_sc_hd__nand4_2
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_79 _5245_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3746_ _6941_/Q _5360_/A _4268_/A _6723_/Q VGND VGND VPWR VPWR _3746_/X sky130_fd_sc_hd__a22o_1
XANTENNA_68 _5396_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6534_ _6777_/CLK _6534_/D fanout424/X VGND VGND VPWR VPWR _6534_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_180_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6465_ _3938_/A1 _6465_/D _6420_/X VGND VGND VPWR VPWR _6465_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_137_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3677_ _6489_/Q _3978_/A _4322_/A _6769_/Q _3676_/X VGND VGND VPWR VPWR _3717_/A
+ sky130_fd_sc_hd__a221o_1
X_5416_ _5578_/A0 hold397/X _5422_/S VGND VGND VPWR VPWR _6990_/D sky130_fd_sc_hd__mux2_1
X_6396_ _6707_/Q _6396_/A2 _6396_/B1 _4238_/B _6395_/X VGND VGND VPWR VPWR _6396_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5347_ _5581_/A0 hold301/X _5350_/S VGND VGND VPWR VPWR _5347_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput175 _3947_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[0] sky130_fd_sc_hd__buf_8
Xoutput186 _3946_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[1] sky130_fd_sc_hd__buf_8
XFILLER_102_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5278_ hold14/X _5278_/A1 hold29/X VGND VGND VPWR VPWR hold30/A sky130_fd_sc_hd__mux2_1
Xoutput197 _3237_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[2] sky130_fd_sc_hd__buf_8
X_7017_ _7135_/CLK _7017_/D fanout429/X VGND VGND VPWR VPWR _7017_/Q sky130_fd_sc_hd__dfrtp_2
X_4229_ hold548/X _4228_/X _4235_/S VGND VGND VPWR VPWR _4229_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout391 _5597_/A0 VGND VGND VPWR VPWR _5300_/A0 sky130_fd_sc_hd__buf_8
XFILLER_120_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout380 hold183/X VGND VGND VPWR VPWR hold184/A sky130_fd_sc_hd__buf_8
XFILLER_62_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4580_ _4581_/B _4634_/B _4536_/X _4987_/A VGND VGND VPWR VPWR _4612_/A sky130_fd_sc_hd__a22oi_4
XFILLER_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3600_ _6756_/Q _4304_/A _4049_/A _6538_/Q _3560_/X VGND VGND VPWR VPWR _3605_/B
+ sky130_fd_sc_hd__a221o_1
Xinput11 mask_rev_in[16] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__clkbuf_4
XFILLER_52_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput22 mask_rev_in[26] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__clkbuf_4
Xinput44 mgmt_gpio_in[17] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__clkbuf_4
Xinput55 mgmt_gpio_in[27] VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__buf_4
XFILLER_162_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3531_ _3543_/A _3732_/B VGND VGND VPWR VPWR _4097_/A sky130_fd_sc_hd__nor2_8
Xinput33 mask_rev_in[7] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__clkbuf_4
Xhold828 _5311_/X VGND VGND VPWR VPWR _6897_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_183_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput66 mgmt_gpio_in[37] VGND VGND VPWR VPWR _7229_/A sky130_fd_sc_hd__buf_8
Xinput88 spimemio_flash_io1_oeb VGND VGND VPWR VPWR _3961_/B sky130_fd_sc_hd__buf_8
Xhold806 _6603_/Q VGND VGND VPWR VPWR hold806/X sky130_fd_sc_hd__bufbuf_16
Xhold817 _6622_/Q VGND VGND VPWR VPWR hold817/X sky130_fd_sc_hd__bufbuf_16
Xinput77 ser_tx VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__clkbuf_4
Xinput99 wb_adr_i[0] VGND VGND VPWR VPWR _4672_/A sky130_fd_sc_hd__buf_8
Xhold839 _7145_/Q VGND VGND VPWR VPWR hold839/X sky130_fd_sc_hd__bufbuf_16
X_3462_ _3540_/A _4241_/B VGND VGND VPWR VPWR _4256_/A sky130_fd_sc_hd__nor2_8
XFILLER_115_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6250_ _6594_/Q _6022_/D _6036_/Y _6748_/Q _6249_/X VGND VGND VPWR VPWR _6257_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6181_ _6181_/A _6181_/B _6181_/C _6181_/D VGND VGND VPWR VPWR _6182_/C sky130_fd_sc_hd__or4_1
X_3393_ _6963_/Q _5378_/A hold61/A _7139_/Q _3390_/X VGND VGND VPWR VPWR _3398_/A
+ sky130_fd_sc_hd__a221o_1
X_5201_ _5234_/C _5201_/A1 _5206_/S VGND VGND VPWR VPWR _5201_/X sky130_fd_sc_hd__mux2_1
X_5132_ _5132_/A _5133_/A _5132_/C VGND VGND VPWR VPWR _5143_/B sky130_fd_sc_hd__or3_1
XFILLER_69_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5063_ _4505_/X _5062_/B _4963_/Y _5062_/X _4612_/C VGND VGND VPWR VPWR _5066_/A
+ sky130_fd_sc_hd__o2111a_2
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4014_ hold876/X _4013_/X _4024_/S VGND VGND VPWR VPWR _4014_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5965_ _6742_/Q _5678_/X _5692_/X _7225_/Q VGND VGND VPWR VPWR _5981_/A sky130_fd_sc_hd__a22o_1
X_4916_ _6779_/Q _4239_/X _4807_/X _4915_/X VGND VGND VPWR VPWR _6779_/D sky130_fd_sc_hd__o22a_1
X_5896_ _7184_/Q _6309_/S _5895_/X VGND VGND VPWR VPWR _7184_/D sky130_fd_sc_hd__o21a_1
XFILLER_40_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4847_ _4847_/A _5174_/A VGND VGND VPWR VPWR _5171_/A sky130_fd_sc_hd__or2_1
XFILLER_119_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4778_ _5165_/A _4778_/B VGND VGND VPWR VPWR _5033_/C sky130_fd_sc_hd__and2_1
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6517_ _7152_/CLK _6517_/D fanout452/X VGND VGND VPWR VPWR _6517_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_107_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3729_ _3728_/X _6791_/Q _3928_/A VGND VGND VPWR VPWR _6791_/D sky130_fd_sc_hd__mux2_1
XFILLER_164_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6448_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6448_/X sky130_fd_sc_hd__and2_1
X_6379_ _6378_/X _7211_/Q _6400_/S VGND VGND VPWR VPWR _7211_/D sky130_fd_sc_hd__mux2_1
XFILLER_164_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5750_ _6895_/Q _5694_/X _5749_/X VGND VGND VPWR VPWR _5753_/C sky130_fd_sc_hd__a21o_1
XFILLER_97_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4701_ _5050_/A _4711_/A _4707_/B VGND VGND VPWR VPWR _4702_/B sky130_fd_sc_hd__a21oi_1
X_5681_ _5864_/B _5702_/B _5706_/B VGND VGND VPWR VPWR _5681_/X sky130_fd_sc_hd__and3_4
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4632_ _4996_/A _4989_/A VGND VGND VPWR VPWR _5078_/B sky130_fd_sc_hd__nor2_2
XFILLER_190_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold603 _7155_/Q VGND VGND VPWR VPWR hold603/X sky130_fd_sc_hd__bufbuf_16
XFILLER_162_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4563_ _4763_/B _4980_/A _4559_/X _4980_/B _4367_/X VGND VGND VPWR VPWR _4563_/X
+ sky130_fd_sc_hd__o41a_4
X_4494_ _4501_/A _4648_/B VGND VGND VPWR VPWR _4494_/Y sky130_fd_sc_hd__nor2_2
Xhold625 _5358_/X VGND VGND VPWR VPWR _6939_/D sky130_fd_sc_hd__bufbuf_16
Xhold636 _6880_/Q VGND VGND VPWR VPWR hold636/X sky130_fd_sc_hd__bufbuf_16
X_6302_ _6537_/Q _6025_/D _6029_/X _6641_/Q _6301_/X VGND VGND VPWR VPWR _6305_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_116_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold614 _6816_/Q VGND VGND VPWR VPWR hold614/X sky130_fd_sc_hd__bufbuf_16
X_3514_ _3514_/A _3732_/B VGND VGND VPWR VPWR _4322_/A sky130_fd_sc_hd__nor2_8
Xhold658 _4069_/X VGND VGND VPWR VPWR _6551_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_171_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3445_ _7010_/Q _5432_/A _5324_/A _6914_/Q _3444_/X VGND VGND VPWR VPWR _3451_/C
+ sky130_fd_sc_hd__a221o_1
Xhold647 _7091_/Q VGND VGND VPWR VPWR hold647/X sky130_fd_sc_hd__bufbuf_16
Xhold669 _6775_/Q VGND VGND VPWR VPWR hold669/X sky130_fd_sc_hd__bufbuf_16
X_6233_ _6860_/Q _6060_/B _6219_/X _6232_/X _3197_/Y VGND VGND VPWR VPWR _6233_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_170_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6164_ _7026_/Q _6010_/Y _6031_/X _7090_/Q _6163_/X VGND VGND VPWR VPWR _6170_/A
+ sky130_fd_sc_hd__a221o_1
X_3376_ _6876_/Q _5279_/A _5369_/A _6956_/Q _3373_/X VGND VGND VPWR VPWR _3377_/D
+ sky130_fd_sc_hd__a221o_4
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5115_ _5115_/A _5115_/B VGND VGND VPWR VPWR _5137_/B sky130_fd_sc_hd__or2_2
XFILLER_85_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6095_ _6983_/Q _6028_/X _6034_/Y _6991_/Q _6094_/X VGND VGND VPWR VPWR _6095_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5046_ _5046_/A _5108_/A _5154_/A VGND VGND VPWR VPWR _5057_/A sky130_fd_sc_hd__or3_1
XFILLER_85_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6997_ _7129_/CLK _6997_/D fanout428/X VGND VGND VPWR VPWR _6997_/Q sky130_fd_sc_hd__dfstp_4
X_5948_ _6622_/Q _5673_/X _5681_/X _6597_/Q _5947_/X VGND VGND VPWR VPWR _5953_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5879_ _6634_/Q _5675_/X _5683_/X _6773_/Q VGND VGND VPWR VPWR _5879_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3230_ _6936_/Q VGND VGND VPWR VPWR _3230_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6920_ _7154_/CLK _6920_/D fanout452/X VGND VGND VPWR VPWR _6920_/Q sky130_fd_sc_hd__dfrtp_2
X_6851_ _6851_/CLK _6851_/D fanout417/X VGND VGND VPWR VPWR _6851_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5802_ _6913_/Q _5680_/X _5700_/X _6865_/Q VGND VGND VPWR VPWR _5802_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6782_ _7208_/CLK _6782_/D fanout458/X VGND VGND VPWR VPWR _6782_/Q sky130_fd_sc_hd__dfrtp_2
X_3994_ hold408/X _5584_/A0 _3994_/S VGND VGND VPWR VPWR _6495_/D sky130_fd_sc_hd__mux2_1
XFILLER_188_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5733_ _6974_/Q _5676_/X _5702_/X _6886_/Q _5732_/X VGND VGND VPWR VPWR _5734_/D
+ sky130_fd_sc_hd__a221o_4
XFILLER_176_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5664_ _5665_/A _5665_/B VGND VGND VPWR VPWR _5664_/X sky130_fd_sc_hd__or2_4
X_5595_ _5595_/A0 _5595_/A1 _5602_/S VGND VGND VPWR VPWR _7149_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4615_ _4846_/B _4615_/B _4615_/C VGND VGND VPWR VPWR _4619_/B sky130_fd_sc_hd__and3b_1
XFILLER_108_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_54_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7104_/CLK sky130_fd_sc_hd__clkbuf_8
Xhold411 _6527_/Q VGND VGND VPWR VPWR hold411/X sky130_fd_sc_hd__bufbuf_16
X_4546_ _4850_/A _5022_/A _4546_/C _4546_/D VGND VGND VPWR VPWR _4548_/C sky130_fd_sc_hd__or4_1
Xhold400 _7084_/Q VGND VGND VPWR VPWR hold400/X sky130_fd_sc_hd__bufbuf_16
Xhold444 _6905_/Q VGND VGND VPWR VPWR hold444/X sky130_fd_sc_hd__bufbuf_16
Xhold433 _6961_/Q VGND VGND VPWR VPWR hold433/X sky130_fd_sc_hd__bufbuf_16
Xhold422 _5449_/X VGND VGND VPWR VPWR _7020_/D sky130_fd_sc_hd__bufbuf_16
Xhold477 _5393_/X VGND VGND VPWR VPWR _6970_/D sky130_fd_sc_hd__bufbuf_16
X_4477_ _4603_/B _4749_/C VGND VGND VPWR VPWR _4883_/A sky130_fd_sc_hd__nor2_1
XFILLER_143_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold466 _6815_/Q VGND VGND VPWR VPWR hold466/X sky130_fd_sc_hd__bufbuf_16
Xhold455 _7046_/Q VGND VGND VPWR VPWR hold455/X sky130_fd_sc_hd__bufbuf_16
Xhold499 _6956_/Q VGND VGND VPWR VPWR hold499/X sky130_fd_sc_hd__bufbuf_16
Xclkbuf_leaf_69_csclk _6722_/CLK VGND VGND VPWR VPWR _6744_/CLK sky130_fd_sc_hd__clkbuf_8
X_3428_ input31/X _3283_/Y _3978_/A _6493_/Q VGND VGND VPWR VPWR _3428_/X sky130_fd_sc_hd__a22o_2
Xhold488 _6503_/Q VGND VGND VPWR VPWR hold488/X sky130_fd_sc_hd__bufbuf_16
X_7196_ _7196_/CLK _7196_/D fanout435/X VGND VGND VPWR VPWR _7196_/Q sky130_fd_sc_hd__dfrtp_1
X_6216_ _7124_/Q _6023_/D _6030_/Y _7036_/Q _6215_/X VGND VGND VPWR VPWR _6219_/C
+ sky130_fd_sc_hd__a221o_1
Xhold1100 _4056_/X VGND VGND VPWR VPWR _6540_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_131_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6147_ _7129_/Q _6023_/A _6033_/X _7009_/Q _6146_/X VGND VGND VPWR VPWR _6157_/B
+ sky130_fd_sc_hd__a221o_1
X_3359_ _3506_/A _3375_/B VGND VGND VPWR VPWR _3359_/Y sky130_fd_sc_hd__nor2_8
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1122 _4068_/X VGND VGND VPWR VPWR _6550_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_97_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1111 _7077_/Q VGND VGND VPWR VPWR _5514_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_58_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1133 _6825_/Q VGND VGND VPWR VPWR _5226_/A1 sky130_fd_sc_hd__bufbuf_16
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1144 _6619_/Q VGND VGND VPWR VPWR _4149_/A0 sky130_fd_sc_hd__bufbuf_16
X_6078_ _7102_/Q _5653_/X _6022_/B _6942_/Q VGND VGND VPWR VPWR _6078_/X sky130_fd_sc_hd__a22o_2
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1155 _4167_/X VGND VGND VPWR VPWR _6634_/D sky130_fd_sc_hd__bufbuf_16
Xhold1166 _4191_/X VGND VGND VPWR VPWR _6654_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_45_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5029_ _4414_/B _4711_/C _4704_/X _4802_/A _4932_/B VGND VGND VPWR VPWR _5101_/A
+ sky130_fd_sc_hd__a2111o_1
Xhold1188 _5381_/X VGND VGND VPWR VPWR _6959_/D sky130_fd_sc_hd__bufbuf_16
XANTENNA_306 _3971_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1199 _5235_/X VGND VGND VPWR VPWR _6832_/D sky130_fd_sc_hd__bufbuf_16
Xhold1177 _6659_/Q VGND VGND VPWR VPWR _4197_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_317 _3932_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_339 hold71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_328 _6409_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4400_ _4400_/A _4513_/A VGND VGND VPWR VPWR _4617_/A sky130_fd_sc_hd__or2_4
XFILLER_160_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5380_ _5596_/A0 hold382/X _5386_/S VGND VGND VPWR VPWR _6958_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4331_ _5561_/A0 hold669/X _4333_/S VGND VGND VPWR VPWR _6775_/D sky130_fd_sc_hd__mux2_1
X_4262_ _4262_/A _5558_/B VGND VGND VPWR VPWR _4267_/S sky130_fd_sc_hd__and2_4
XFILLER_113_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7050_ _7090_/CLK _7050_/D fanout438/X VGND VGND VPWR VPWR _7050_/Q sky130_fd_sc_hd__dfrtp_2
X_3213_ _7072_/Q VGND VGND VPWR VPWR _3213_/Y sky130_fd_sc_hd__inv_2
X_6001_ _6037_/A _6032_/A VGND VGND VPWR VPWR _6010_/B sky130_fd_sc_hd__nand2_8
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4193_ _6409_/A0 _4193_/A1 _4195_/S VGND VGND VPWR VPWR _6656_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6903_ _7153_/CLK _6903_/D fanout444/X VGND VGND VPWR VPWR _6903_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6834_ _6964_/CLK _6834_/D fanout444/X VGND VGND VPWR VPWR _6834_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3977_ hold98/X _3975_/B hold155/X VGND VGND VPWR VPWR _3977_/Y sky130_fd_sc_hd__o21ai_4
X_6765_ _6851_/CLK _6765_/D fanout418/X VGND VGND VPWR VPWR _6765_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_50_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5716_ _6861_/Q _5700_/X _5706_/X _7053_/Q _5686_/X VGND VGND VPWR VPWR _5720_/B
+ sky130_fd_sc_hd__a221o_1
X_6696_ _7127_/CLK _6696_/D fanout448/X VGND VGND VPWR VPWR _6696_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5647_ _7169_/Q _5635_/B _5645_/Y _5646_/X VGND VGND VPWR VPWR _7169_/D sky130_fd_sc_hd__a31o_1
XFILLER_163_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5578_ _5578_/A0 hold362/X hold62/X VGND VGND VPWR VPWR _7134_/D sky130_fd_sc_hd__mux2_1
Xhold252 _6518_/Q VGND VGND VPWR VPWR hold252/X sky130_fd_sc_hd__bufbuf_16
X_4529_ _4529_/A _4529_/B _4529_/C VGND VGND VPWR VPWR _4533_/B sky130_fd_sc_hd__and3_4
XFILLER_144_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold241 _5463_/X VGND VGND VPWR VPWR _7032_/D sky130_fd_sc_hd__bufbuf_16
Xhold230 _6993_/Q VGND VGND VPWR VPWR hold230/X sky130_fd_sc_hd__bufbuf_16
Xhold274 _4214_/X VGND VGND VPWR VPWR _6674_/D sky130_fd_sc_hd__bufbuf_16
Xhold296 _5382_/X VGND VGND VPWR VPWR _6960_/D sky130_fd_sc_hd__bufbuf_16
Xhold285 _6781_/Q VGND VGND VPWR VPWR hold88/A sky130_fd_sc_hd__bufbuf_16
XFILLER_104_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold263 _5364_/X VGND VGND VPWR VPWR _6944_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_172_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7179_ _7196_/CLK _7179_/D fanout432/X VGND VGND VPWR VPWR _7179_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_114 _3994_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_103 _3801_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_125 _5251_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_136 _5682_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_158 _5764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_147 _5703_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_169 _6021_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 mask_rev_in[14] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_4
XFILLER_45_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4880_ _4875_/A _4588_/X _4593_/Y VGND VGND VPWR VPWR _4962_/A sky130_fd_sc_hd__o21ai_1
X_3900_ _6707_/Q _3883_/X _6702_/Q VGND VGND VPWR VPWR _6707_/D sky130_fd_sc_hd__a21o_1
XFILLER_177_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3831_ hold24/A _3845_/A _3824_/B _3830_/X VGND VGND VPWR VPWR _3831_/X sky130_fd_sc_hd__a22o_1
X_6550_ _6745_/CLK _6550_/D _6421_/A VGND VGND VPWR VPWR _6550_/Q sky130_fd_sc_hd__dfrtp_2
X_3762_ _6917_/Q _5333_/A _4292_/A _6743_/Q _3737_/X VGND VGND VPWR VPWR _3764_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_32_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5501_ _5600_/A0 hold402/X _5503_/S VGND VGND VPWR VPWR _5501_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3693_ _3693_/A _3693_/B _3693_/C _3693_/D VGND VGND VPWR VPWR _3727_/B sky130_fd_sc_hd__or4_2
XFILLER_9_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6481_ _6668_/CLK _6481_/D _6436_/X VGND VGND VPWR VPWR _6481_/Q sky130_fd_sc_hd__dfrtp_2
X_5432_ _5432_/A _5576_/B VGND VGND VPWR VPWR _5440_/S sky130_fd_sc_hd__nand2_8
Xoutput313 _3964_/X VGND VGND VPWR VPWR spimemio_flash_io0_di sky130_fd_sc_hd__buf_8
XFILLER_161_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput335 _7204_/Q VGND VGND VPWR VPWR wb_dat_o[25] sky130_fd_sc_hd__buf_8
Xoutput324 _6575_/Q VGND VGND VPWR VPWR wb_dat_o[15] sky130_fd_sc_hd__buf_8
XFILLER_99_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5363_ hold43/X _5363_/A1 _5368_/S VGND VGND VPWR VPWR hold44/A sky130_fd_sc_hd__mux2_1
Xoutput302 _6821_/Q VGND VGND VPWR VPWR pwr_ctrl_out[1] sky130_fd_sc_hd__buf_8
Xoutput346 _6587_/Q VGND VGND VPWR VPWR wb_dat_o[6] sky130_fd_sc_hd__buf_8
X_7102_ _7118_/CLK hold68/X fanout436/X VGND VGND VPWR VPWR _7102_/Q sky130_fd_sc_hd__dfstp_2
X_4314_ hold798/X _4326_/A0 _4315_/S VGND VGND VPWR VPWR _4314_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5294_ _5600_/A0 hold393/X _5296_/S VGND VGND VPWR VPWR _5294_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4245_ _5571_/A0 hold641/X _4249_/S VGND VGND VPWR VPWR _4245_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7033_ _7118_/CLK _7033_/D fanout436/X VGND VGND VPWR VPWR _7033_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4176_ _4176_/A0 _6410_/A0 _4177_/S VGND VGND VPWR VPWR _4176_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6817_ _7132_/CLK _6817_/D fanout432/X VGND VGND VPWR VPWR _6817_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6748_ _6810_/CLK _6748_/D fanout419/X VGND VGND VPWR VPWR _6748_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6679_ _7196_/CLK _6679_/D fanout433/X VGND VGND VPWR VPWR _6679_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_3_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4030_ _5581_/A0 hold252/X _4033_/S VGND VGND VPWR VPWR _4030_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5981_ _5981_/A _5981_/B _5981_/C _5981_/D VGND VGND VPWR VPWR _5981_/X sky130_fd_sc_hd__or4_1
X_4932_ _4932_/A _4932_/B _4932_/C VGND VGND VPWR VPWR _4940_/B sky130_fd_sc_hd__or3_2
XFILLER_45_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_14 _4218_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6602_ _6725_/CLK _6602_/D fanout440/X VGND VGND VPWR VPWR _6602_/Q sky130_fd_sc_hd__dfrtp_2
X_4863_ _5118_/A _4863_/B _4863_/C _5084_/A VGND VGND VPWR VPWR _4865_/B sky130_fd_sc_hd__or4_1
XANTENNA_25 _6888_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4794_ _5165_/A _4793_/Y _4791_/X _5035_/B VGND VGND VPWR VPWR _4794_/X sky130_fd_sc_hd__a211o_1
XANTENNA_47 _5342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_36 _5659_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3814_ _6480_/Q _3830_/B VGND VGND VPWR VPWR _3828_/S sky130_fd_sc_hd__and2_2
XANTENNA_69 _5558_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 _5423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3745_ _7085_/Q hold54/A _5459_/A _7029_/Q VGND VGND VPWR VPWR _3745_/X sky130_fd_sc_hd__a22o_2
X_6533_ _6777_/CLK _6533_/D fanout424/X VGND VGND VPWR VPWR _6533_/Q sky130_fd_sc_hd__dfstp_4
X_6464_ _3938_/A1 _6464_/D _6419_/X VGND VGND VPWR VPWR hold73/A sky130_fd_sc_hd__dfrtp_2
XFILLER_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5415_ _5541_/A0 _5415_/A1 _5422_/S VGND VGND VPWR VPWR _6989_/D sky130_fd_sc_hd__mux2_1
X_3676_ input35/X _3320_/Y _4049_/A _6536_/Q VGND VGND VPWR VPWR _3676_/X sky130_fd_sc_hd__a22o_1
X_6395_ _6705_/Q _6395_/A2 _6395_/B1 _6706_/Q VGND VGND VPWR VPWR _6395_/X sky130_fd_sc_hd__a22o_1
X_5346_ _5571_/A0 hold591/X _5350_/S VGND VGND VPWR VPWR _5346_/X sky130_fd_sc_hd__mux2_1
Xoutput176 _3230_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[10] sky130_fd_sc_hd__buf_8
XFILLER_102_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput187 _3220_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[20] sky130_fd_sc_hd__buf_8
Xoutput198 _3210_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[30] sky130_fd_sc_hd__buf_8
XFILLER_153_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5277_ hold209/X hold256/X hold29/X VGND VGND VPWR VPWR _5277_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7016_ _7140_/CLK _7016_/D fanout430/X VGND VGND VPWR VPWR _7016_/Q sky130_fd_sc_hd__dfrtp_2
X_4228_ hold293/X hold185/A _4234_/S VGND VGND VPWR VPWR _4228_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4159_ hold815/X _5599_/A0 _4159_/S VGND VGND VPWR VPWR _4159_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout381 _5581_/A0 VGND VGND VPWR VPWR _5599_/A0 sky130_fd_sc_hd__buf_8
Xfanout370 hold14/X VGND VGND VPWR VPWR _5602_/A0 sky130_fd_sc_hd__buf_8
Xfanout392 hold43/A VGND VGND VPWR VPWR _5597_/A0 sky130_fd_sc_hd__buf_8
XFILLER_143_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_1_0_mgmt_gpio_in[4] clkbuf_2_1_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _6668_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_93_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput12 mask_rev_in[17] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput45 mgmt_gpio_in[18] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__clkbuf_4
XFILLER_168_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3530_ _6633_/Q _4160_/A _4112_/A _6593_/Q VGND VGND VPWR VPWR _3530_/X sky130_fd_sc_hd__a22o_1
Xinput34 mask_rev_in[8] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__clkbuf_4
Xinput23 mask_rev_in[27] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__clkbuf_4
Xinput56 mgmt_gpio_in[28] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__buf_6
Xinput89 spimemio_flash_io2_do VGND VGND VPWR VPWR input89/X sky130_fd_sc_hd__clkbuf_4
Xhold807 _4129_/X VGND VGND VPWR VPWR _6603_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_143_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold818 _4152_/X VGND VGND VPWR VPWR _6622_/D sky130_fd_sc_hd__bufbuf_16
Xinput78 spi_csb VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__clkbuf_4
Xinput67 mgmt_gpio_in[3] VGND VGND VPWR VPWR _3877_/C sky130_fd_sc_hd__buf_8
XFILLER_116_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold829 _6592_/Q VGND VGND VPWR VPWR hold829/X sky130_fd_sc_hd__bufbuf_16
X_3461_ _6767_/Q _4316_/A _4328_/A _6777_/Q VGND VGND VPWR VPWR _3461_/X sky130_fd_sc_hd__a22o_2
XFILLER_170_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6180_ _7066_/Q _5996_/X _6020_/C _6914_/Q _6161_/X VGND VGND VPWR VPWR _6181_/D
+ sky130_fd_sc_hd__a221o_1
X_5200_ _5200_/A _6406_/B VGND VGND VPWR VPWR _5206_/S sky130_fd_sc_hd__nand2_8
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3392_ _7091_/Q hold54/A _3359_/Y _7019_/Q VGND VGND VPWR VPWR _3392_/X sky130_fd_sc_hd__a22o_1
X_5131_ _5131_/A _5146_/A _5143_/A VGND VGND VPWR VPWR _5133_/B sky130_fd_sc_hd__nor3_2
XFILLER_123_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5062_ _5062_/A _5062_/B _5062_/C VGND VGND VPWR VPWR _5062_/X sky130_fd_sc_hd__or3_1
X_4013_ hold525/X _5597_/A0 _4023_/S VGND VGND VPWR VPWR _4013_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5964_ _6648_/Q _5685_/X _5699_/X _6603_/Q VGND VGND VPWR VPWR _5964_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4915_ _4367_/X _4867_/X _4914_/X VGND VGND VPWR VPWR _4915_/X sky130_fd_sc_hd__a21o_2
XFILLER_33_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5895_ _5611_/A _7183_/Q _6358_/B1 _5894_/X VGND VGND VPWR VPWR _5895_/X sky130_fd_sc_hd__a211o_1
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4846_ _5033_/A _4846_/B VGND VGND VPWR VPWR _4846_/X sky130_fd_sc_hd__or2_1
XFILLER_32_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6516_ _7152_/CLK _6516_/D fanout447/X VGND VGND VPWR VPWR _6516_/Q sky130_fd_sc_hd__dfrtp_2
X_4777_ _4772_/A _5165_/B _4698_/Y VGND VGND VPWR VPWR _4778_/B sky130_fd_sc_hd__a21o_1
XFILLER_119_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3728_ _3727_/X _6790_/Q _3857_/C VGND VGND VPWR VPWR _3728_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6447_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6447_/X sky130_fd_sc_hd__and2_1
X_3659_ _6775_/Q _4328_/A _4172_/A _6641_/Q VGND VGND VPWR VPWR _3659_/X sky130_fd_sc_hd__a22o_1
X_6378_ _6707_/Q _6378_/A2 _6378_/B1 _4238_/B _6377_/X VGND VGND VPWR VPWR _6378_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_164_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5329_ _5599_/A0 hold735/X _5332_/S VGND VGND VPWR VPWR _5329_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4700_ _4422_/Y _4423_/X _4424_/Y _4414_/B VGND VGND VPWR VPWR _4930_/C sky130_fd_sc_hd__o2bb2a_2
X_5680_ _5864_/B _5705_/B _5707_/C VGND VGND VPWR VPWR _5680_/X sky130_fd_sc_hd__and3_4
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4631_ _4995_/A _4844_/A _4575_/Y _4627_/X _4630_/Y VGND VGND VPWR VPWR _4631_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_30_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4562_ _4819_/B _4562_/B VGND VGND VPWR VPWR _4980_/B sky130_fd_sc_hd__nor2_8
XFILLER_128_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold604 _5601_/X VGND VGND VPWR VPWR _7155_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_155_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4493_ _4648_/B _5164_/B VGND VGND VPWR VPWR _4840_/A sky130_fd_sc_hd__nor2_2
XFILLER_143_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6301_ _6636_/Q _5653_/X _6022_/B _6611_/Q VGND VGND VPWR VPWR _6301_/X sky130_fd_sc_hd__a22o_1
X_3513_ input56/X _4025_/A _4049_/A _6539_/Q _3512_/X VGND VGND VPWR VPWR _3522_/B
+ sky130_fd_sc_hd__a221o_1
Xhold615 _7034_/Q VGND VGND VPWR VPWR hold615/X sky130_fd_sc_hd__bufbuf_16
Xhold626 _6494_/Q VGND VGND VPWR VPWR hold626/X sky130_fd_sc_hd__bufbuf_16
Xhold659 _6899_/Q VGND VGND VPWR VPWR hold659/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold637 _6620_/Q VGND VGND VPWR VPWR hold637/X sky130_fd_sc_hd__bufbuf_16
XFILLER_116_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6232_ _6232_/A _6232_/B _6232_/C VGND VGND VPWR VPWR _6232_/X sky130_fd_sc_hd__or3_1
X_3444_ input25/X _3302_/Y _3320_/Y input8/X VGND VGND VPWR VPWR _3444_/X sky130_fd_sc_hd__a22o_4
Xhold648 _5529_/X VGND VGND VPWR VPWR _7091_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_170_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3375_ _3540_/A _3375_/B VGND VGND VPWR VPWR _5369_/A sky130_fd_sc_hd__nor2_8
X_6163_ _7138_/Q _6020_/B _6011_/X _7098_/Q VGND VGND VPWR VPWR _6163_/X sky130_fd_sc_hd__a22o_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5114_ _5114_/A _5114_/B _5114_/C _5114_/D VGND VGND VPWR VPWR _5115_/B sky130_fd_sc_hd__or4_1
X_6094_ _7071_/Q _6009_/X _6020_/D _6967_/Q VGND VGND VPWR VPWR _6094_/X sky130_fd_sc_hd__a22o_1
XFILLER_57_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _4758_/B _5042_/Y _5016_/C _5035_/A VGND VGND VPWR VPWR _5154_/A sky130_fd_sc_hd__a211o_1
XFILLER_111_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6996_ _7123_/CLK _6996_/D fanout434/X VGND VGND VPWR VPWR _6996_/Q sky130_fd_sc_hd__dfrtp_2
X_5947_ _6711_/Q _5691_/X _5701_/X _6617_/Q VGND VGND VPWR VPWR _5947_/X sky130_fd_sc_hd__a22o_1
XFILLER_43_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5878_ _6659_/Q _5669_/X _5678_/X _6738_/Q _5877_/X VGND VGND VPWR VPWR _5883_/B
+ sky130_fd_sc_hd__a221o_1
X_4829_ _4736_/B _4657_/B _4697_/Y _4828_/Y VGND VGND VPWR VPWR _4829_/X sky130_fd_sc_hd__a211o_1
XFILLER_166_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1 hold9/X VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__bufbuf_16
XFILLER_94_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6850_ _7138_/CLK _6850_/D fanout438/X VGND VGND VPWR VPWR _6850_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6781_ _3949_/A1 _6781_/D fanout458/X VGND VGND VPWR VPWR _6781_/Q sky130_fd_sc_hd__dfrtp_2
X_5801_ _7017_/Q _5682_/X _5706_/X _7057_/Q _5800_/X VGND VGND VPWR VPWR _5806_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3993_ hold10/X _7218_/Q _6689_/Q VGND VGND VPWR VPWR hold11/A sky130_fd_sc_hd__mux2_8
X_5732_ _7062_/Q _5669_/X _5698_/B _6982_/Q _5697_/X VGND VGND VPWR VPWR _5732_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5663_ _5663_/A _5663_/B VGND VGND VPWR VPWR _5663_/Y sky130_fd_sc_hd__nor2_2
X_5594_ _5594_/A _5594_/B VGND VGND VPWR VPWR _5602_/S sky130_fd_sc_hd__nand2_8
X_4614_ _4997_/A _4844_/A VGND VGND VPWR VPWR _4615_/C sky130_fd_sc_hd__or2_1
XFILLER_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4545_ _4500_/A _4622_/B _4772_/A _4399_/Y _4847_/A VGND VGND VPWR VPWR _4546_/D
+ sky130_fd_sc_hd__a221o_1
Xhold401 _5521_/X VGND VGND VPWR VPWR _7084_/D sky130_fd_sc_hd__bufbuf_16
Xhold412 _4040_/X VGND VGND VPWR VPWR _6527_/D sky130_fd_sc_hd__bufbuf_16
Xhold445 _5320_/X VGND VGND VPWR VPWR _6905_/D sky130_fd_sc_hd__bufbuf_16
Xhold434 _5383_/X VGND VGND VPWR VPWR _6961_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_116_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold423 _7044_/Q VGND VGND VPWR VPWR hold423/X sky130_fd_sc_hd__bufbuf_16
Xhold456 _7058_/Q VGND VGND VPWR VPWR hold456/X sky130_fd_sc_hd__bufbuf_16
X_4476_ _4558_/B _4584_/A VGND VGND VPWR VPWR _4749_/C sky130_fd_sc_hd__or2_4
XFILLER_131_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold478 _6977_/Q VGND VGND VPWR VPWR hold478/X sky130_fd_sc_hd__bufbuf_16
XFILLER_89_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold467 _5212_/X VGND VGND VPWR VPWR _6815_/D sky130_fd_sc_hd__bufbuf_16
X_6215_ _7004_/Q _5987_/Y _6022_/D _6924_/Q VGND VGND VPWR VPWR _6215_/X sky130_fd_sc_hd__a22o_4
XFILLER_143_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold489 _6709_/Q VGND VGND VPWR VPWR hold489/X sky130_fd_sc_hd__bufbuf_16
X_7195_ _7196_/CLK _7195_/D fanout435/X VGND VGND VPWR VPWR _7195_/Q sky130_fd_sc_hd__dfrtp_4
X_3427_ _6816_/Q _5207_/A _5459_/A _7034_/Q _3426_/X VGND VGND VPWR VPWR _3450_/A
+ sky130_fd_sc_hd__a221o_1
X_6146_ _6889_/Q _6020_/A _6021_/D _7145_/Q _6145_/X VGND VGND VPWR VPWR _6146_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_112_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3358_ _5252_/A _3515_/B VGND VGND VPWR VPWR _5567_/A sky130_fd_sc_hd__nor2_8
Xhold1123 _6927_/Q VGND VGND VPWR VPWR _5345_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_97_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1112 _7029_/Q VGND VGND VPWR VPWR _5460_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1101 _6648_/Q VGND VGND VPWR VPWR _4183_/A0 sky130_fd_sc_hd__bufbuf_16
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1156 _6903_/Q VGND VGND VPWR VPWR _5318_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1167 _6614_/Q VGND VGND VPWR VPWR _4143_/A1 sky130_fd_sc_hd__bufbuf_16
X_6077_ _6870_/Q _6023_/C _6025_/B _6894_/Q _6076_/X VGND VGND VPWR VPWR _6082_/B
+ sky130_fd_sc_hd__a221o_1
Xhold1145 _4149_/X VGND VGND VPWR VPWR _6619_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_100_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1134 _5226_/X VGND VGND VPWR VPWR _6825_/D sky130_fd_sc_hd__bufbuf_16
X_3289_ hold26/X _3421_/B VGND VGND VPWR VPWR _3343_/A sky130_fd_sc_hd__nand2_2
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5028_ _5180_/C _5028_/B _5098_/B _5163_/B VGND VGND VPWR VPWR _5036_/A sky130_fd_sc_hd__or4_1
Xhold1189 _6805_/Q VGND VGND VPWR VPWR _5201_/A1 sky130_fd_sc_hd__bufbuf_16
XANTENNA_307 input22/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1178 _4197_/X VGND VGND VPWR VPWR _6659_/D sky130_fd_sc_hd__bufbuf_16
XANTENNA_318 _3931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_329 _6408_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6979_ _7138_/CLK _6979_/D fanout438/X VGND VGND VPWR VPWR _6979_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_110_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold990 _6741_/Q VGND VGND VPWR VPWR hold990/X sky130_fd_sc_hd__bufbuf_16
XFILLER_1_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4330_ _5254_/A0 hold928/X _4333_/S VGND VGND VPWR VPWR _4330_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4261_ _4261_/A0 _5545_/A0 _4261_/S VGND VGND VPWR VPWR _4261_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3212_ _7080_/Q VGND VGND VPWR VPWR _3212_/Y sky130_fd_sc_hd__inv_2
X_6000_ _6037_/B _6035_/A _6018_/A VGND VGND VPWR VPWR _6023_/B sky130_fd_sc_hd__and3_4
XFILLER_79_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4192_ _5254_/A0 hold897/X _4195_/S VGND VGND VPWR VPWR _4192_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6902_ _6959_/CLK _6902_/D fanout444/X VGND VGND VPWR VPWR _6902_/Q sky130_fd_sc_hd__dfstp_4
X_6833_ _6833_/CLK _6833_/D fanout456/X VGND VGND VPWR VPWR _6833_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3976_ hold98/X _3991_/S hold155/X VGND VGND VPWR VPWR hold99/A sky130_fd_sc_hd__o21a_4
XFILLER_23_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6764_ _6851_/CLK _6764_/D fanout418/X VGND VGND VPWR VPWR _6764_/Q sky130_fd_sc_hd__dfrtp_2
X_6695_ _7127_/CLK hold8/X fanout446/X VGND VGND VPWR VPWR _6695_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5715_ _6965_/Q _5691_/X _5704_/X _6933_/Q _5714_/X VGND VGND VPWR VPWR _5720_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_50_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5646_ _6679_/Q _6037_/A _6037_/B VGND VGND VPWR VPWR _5646_/X sky130_fd_sc_hd__and3_1
XFILLER_191_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5577_ hold885/X hold923/X hold62/X VGND VGND VPWR VPWR _7133_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold220 _6992_/Q VGND VGND VPWR VPWR hold220/X sky130_fd_sc_hd__bufbuf_16
X_4528_ _4444_/B _4958_/B VGND VGND VPWR VPWR _4949_/B sky130_fd_sc_hd__and2b_4
Xhold242 _6612_/Q VGND VGND VPWR VPWR hold242/X sky130_fd_sc_hd__bufbuf_16
Xhold253 _4030_/X VGND VGND VPWR VPWR _6518_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_144_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold231 _5419_/X VGND VGND VPWR VPWR _6993_/D sky130_fd_sc_hd__bufbuf_16
X_4459_ _4694_/A _4989_/A VGND VGND VPWR VPWR _4763_/B sky130_fd_sc_hd__nor2_1
Xhold264 _6874_/Q VGND VGND VPWR VPWR hold264/X sky130_fd_sc_hd__bufbuf_16
Xhold275 _7009_/Q VGND VGND VPWR VPWR hold275/X sky130_fd_sc_hd__bufbuf_16
Xhold286 hold88/X VGND VGND VPWR VPWR hold286/X sky130_fd_sc_hd__bufbuf_16
XFILLER_104_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold297 _7025_/Q VGND VGND VPWR VPWR hold297/X sky130_fd_sc_hd__bufbuf_16
X_7178_ _7197_/CLK _7178_/D fanout431/X VGND VGND VPWR VPWR _7178_/Q sky130_fd_sc_hd__dfrtp_4
X_6129_ _7104_/Q _5653_/X _6022_/B _6944_/Q VGND VGND VPWR VPWR _6129_/X sky130_fd_sc_hd__a22o_1
XFILLER_105_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_115 _4033_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_104 _3801_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 _5404_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_148 _5703_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_137 _5682_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_159 _5807_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_53_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7131_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_68_csclk _6722_/CLK VGND VGND VPWR VPWR _7105_/CLK sky130_fd_sc_hd__clkbuf_8
X_3830_ _6480_/Q _3830_/B VGND VGND VPWR VPWR _3830_/X sky130_fd_sc_hd__or2_1
X_3761_ _6909_/Q _5324_/A _4160_/A _6629_/Q _3736_/X VGND VGND VPWR VPWR _3764_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_185_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5500_ _5581_/A0 hold462/X _5503_/S VGND VGND VPWR VPWR _5500_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6480_ _6668_/CLK _6480_/D _6435_/X VGND VGND VPWR VPWR _6480_/Q sky130_fd_sc_hd__dfrtp_2
X_3692_ _6640_/Q _4172_/A _3551_/Y input96/X _3669_/X VGND VGND VPWR VPWR _3693_/D
+ sky130_fd_sc_hd__a221o_1
X_5431_ _5602_/A0 hold380/X hold48/X VGND VGND VPWR VPWR _5431_/X sky130_fd_sc_hd__mux2_1
Xoutput314 _3965_/X VGND VGND VPWR VPWR spimemio_flash_io1_di sky130_fd_sc_hd__buf_8
XFILLER_145_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput325 _6555_/Q VGND VGND VPWR VPWR wb_dat_o[16] sky130_fd_sc_hd__buf_8
Xoutput303 _6822_/Q VGND VGND VPWR VPWR pwr_ctrl_out[2] sky130_fd_sc_hd__buf_8
X_5362_ _5578_/A0 hold379/X _5368_/S VGND VGND VPWR VPWR _6942_/D sky130_fd_sc_hd__mux2_1
Xoutput336 _7205_/Q VGND VGND VPWR VPWR wb_dat_o[26] sky130_fd_sc_hd__buf_8
Xoutput347 _6588_/Q VGND VGND VPWR VPWR wb_dat_o[7] sky130_fd_sc_hd__buf_8
X_4313_ _4313_/A0 _6409_/A0 _4315_/S VGND VGND VPWR VPWR _6760_/D sky130_fd_sc_hd__mux2_1
X_7101_ _7101_/CLK _7101_/D fanout430/X VGND VGND VPWR VPWR _7101_/Q sky130_fd_sc_hd__dfstp_4
X_5293_ _5599_/A0 hold843/X _5296_/S VGND VGND VPWR VPWR _5293_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7032_ _7136_/CLK _7032_/D fanout436/X VGND VGND VPWR VPWR _7032_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_141_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4244_ _5597_/A0 hold554/X _4249_/S VGND VGND VPWR VPWR _4244_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4175_ hold992/X _6409_/A0 _4177_/S VGND VGND VPWR VPWR _6641_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6816_ _7132_/CLK _6816_/D fanout432/X VGND VGND VPWR VPWR _6816_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6747_ _6747_/CLK _6747_/D fanout456/X VGND VGND VPWR VPWR _6747_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3959_ _6474_/Q _3959_/B VGND VGND VPWR VPWR _3960_/A sky130_fd_sc_hd__nand2b_4
XFILLER_176_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6678_ _7196_/CLK _6678_/D fanout433/X VGND VGND VPWR VPWR _6678_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5629_ _7163_/Q _5629_/B VGND VGND VPWR VPWR _5633_/B sky130_fd_sc_hd__or2_2
XFILLER_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5980_ _6789_/Q _5690_/X _5693_/X _6658_/Q _5979_/X VGND VGND VPWR VPWR _5981_/D
+ sky130_fd_sc_hd__a221o_1
X_4931_ _4735_/B _4494_/Y _4957_/A _4930_/X VGND VGND VPWR VPWR _4932_/C sky130_fd_sc_hd__a211o_1
XFILLER_80_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4862_ _4735_/B _4486_/B _4554_/A _4554_/X VGND VGND VPWR VPWR _5084_/A sky130_fd_sc_hd__a31o_1
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6601_ _6725_/CLK _6601_/D fanout440/X VGND VGND VPWR VPWR _6601_/Q sky130_fd_sc_hd__dfstp_4
X_3813_ hold24/A hold16/A hold80/A VGND VGND VPWR VPWR _3830_/B sky130_fd_sc_hd__and3_1
XANTENNA_26 _5304_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_15 _4245_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4793_ _4793_/A VGND VGND VPWR VPWR _4793_/Y sky130_fd_sc_hd__inv_2
XANTENNA_37 _5963_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 _3331_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_59 _5423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3744_ _6488_/Q _3978_/A _3730_/X _5223_/A VGND VGND VPWR VPWR _3744_/X sky130_fd_sc_hd__a22o_1
X_6532_ _6786_/CLK _6532_/D fanout422/X VGND VGND VPWR VPWR _6532_/Q sky130_fd_sc_hd__dfrtp_2
X_6463_ _3938_/A1 _6463_/D _6418_/X VGND VGND VPWR VPWR _6463_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_146_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3675_ _7126_/Q _5567_/A _4234_/S input47/X VGND VGND VPWR VPWR _3675_/X sky130_fd_sc_hd__a22o_1
X_5414_ _5414_/A _5576_/B VGND VGND VPWR VPWR _5422_/S sky130_fd_sc_hd__nand2_8
X_6394_ _6393_/X _7216_/Q _6400_/S VGND VGND VPWR VPWR _7216_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5345_ _5588_/A0 _5345_/A1 _5350_/S VGND VGND VPWR VPWR _5345_/X sky130_fd_sc_hd__mux2_1
Xoutput177 _3229_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[11] sky130_fd_sc_hd__buf_8
Xoutput199 _3209_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[31] sky130_fd_sc_hd__buf_8
Xoutput188 _3219_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[21] sky130_fd_sc_hd__buf_8
X_5276_ hold78/X _5276_/A1 hold29/X VGND VGND VPWR VPWR hold79/A sky130_fd_sc_hd__mux2_1
XFILLER_102_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7015_ _7135_/CLK _7015_/D fanout431/X VGND VGND VPWR VPWR _7015_/Q sky130_fd_sc_hd__dfrtp_2
X_4227_ hold446/X _4226_/X _4235_/S VGND VGND VPWR VPWR _4227_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4158_ hold312/X hold71/X _4159_/S VGND VGND VPWR VPWR _4158_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4089_ _6568_/Q _3794_/X _4096_/S VGND VGND VPWR VPWR _6568_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout371 hold12/X VGND VGND VPWR VPWR hold13/A sky130_fd_sc_hd__buf_8
Xfanout382 hold183/X VGND VGND VPWR VPWR _5581_/A0 sky130_fd_sc_hd__buf_8
Xfanout393 hold41/X VGND VGND VPWR VPWR hold42/A sky130_fd_sc_hd__buf_8
XFILLER_120_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput13 mask_rev_in[18] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput46 mgmt_gpio_in[19] VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__buf_6
Xinput35 mask_rev_in[9] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__clkbuf_4
Xinput24 mask_rev_in[28] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__clkbuf_4
Xinput57 mgmt_gpio_in[29] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__clkbuf_4
Xhold819 _7113_/Q VGND VGND VPWR VPWR hold819/X sky130_fd_sc_hd__bufbuf_16
Xhold808 _6617_/Q VGND VGND VPWR VPWR hold808/X sky130_fd_sc_hd__bufbuf_16
Xinput68 mgmt_gpio_in[5] VGND VGND VPWR VPWR _3969_/A sky130_fd_sc_hd__buf_8
XFILLER_10_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput79 spi_enabled VGND VGND VPWR VPWR _3970_/B sky130_fd_sc_hd__buf_6
XFILLER_143_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3460_ _3514_/A _4241_/B VGND VGND VPWR VPWR _4328_/A sky130_fd_sc_hd__nor2_8
XFILLER_124_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3391_ _7027_/Q _5450_/A hold21/A _7107_/Q VGND VGND VPWR VPWR _3391_/X sky130_fd_sc_hd__a22o_1
X_5130_ _5130_/A _5130_/B _5130_/C _4970_/X VGND VGND VPWR VPWR _5175_/B sky130_fd_sc_hd__or4b_4
XFILLER_111_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5061_ _5132_/A _5133_/A VGND VGND VPWR VPWR _5061_/Y sky130_fd_sc_hd__nor2_1
XFILLER_123_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4012_ hold719/X _4011_/X _4024_/S VGND VGND VPWR VPWR _4012_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5963_ _6628_/Q _5963_/B VGND VGND VPWR VPWR _5963_/X sky130_fd_sc_hd__or2_1
XFILLER_53_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4914_ _5003_/B _4838_/X _4913_/X _4567_/X _6376_/A VGND VGND VPWR VPWR _4914_/X
+ sky130_fd_sc_hd__a221o_1
Xclkbuf_opt_4_0_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR clkbuf_opt_4_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
X_5894_ _6530_/Q _5722_/B _5883_/X _5893_/X _6308_/S VGND VGND VPWR VPWR _5894_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_80_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4845_ _4845_/A _4845_/B VGND VGND VPWR VPWR _4863_/B sky130_fd_sc_hd__and2_2
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4776_ _4776_/A _4776_/B VGND VGND VPWR VPWR _5165_/B sky130_fd_sc_hd__nor2_2
XFILLER_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6515_ _7141_/CLK _6515_/D fanout447/X VGND VGND VPWR VPWR _6515_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_165_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3727_ _3727_/A _3727_/B _3727_/C _3727_/D VGND VGND VPWR VPWR _3727_/X sky130_fd_sc_hd__or4_4
XFILLER_173_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3658_ _7111_/Q hold85/A _3315_/Y _6855_/Q _3657_/X VGND VGND VPWR VPWR _3664_/C
+ sky130_fd_sc_hd__a221o_4
X_6446_ _6446_/A _6446_/B VGND VGND VPWR VPWR _6446_/X sky130_fd_sc_hd__and2_1
X_6377_ _6705_/Q _6377_/A2 _6377_/B1 _6706_/Q VGND VGND VPWR VPWR _6377_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3589_ input23/X _3302_/Y _5459_/A _7032_/Q _3553_/X VGND VGND VPWR VPWR _3593_/A
+ sky130_fd_sc_hd__a221o_1
X_5328_ _5571_/A0 hold573/X _5332_/S VGND VGND VPWR VPWR _5328_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5259_ hold209/X hold246/X _5260_/S VGND VGND VPWR VPWR _5259_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4630_ _5079_/B VGND VGND VPWR VPWR _4630_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4561_ _4562_/B VGND VGND VPWR VPWR _4561_/Y sky130_fd_sc_hd__inv_2
X_6300_ _6542_/Q _6023_/C _6025_/B _6565_/Q _6299_/X VGND VGND VPWR VPWR _6305_/B
+ sky130_fd_sc_hd__a221o_1
X_4492_ _4566_/A _4663_/B VGND VGND VPWR VPWR _4687_/A sky130_fd_sc_hd__or2_4
Xhold627 _6894_/Q VGND VGND VPWR VPWR hold627/X sky130_fd_sc_hd__bufbuf_16
X_3512_ _7081_/Q _5513_/A _3511_/Y _6618_/Q VGND VGND VPWR VPWR _3512_/X sky130_fd_sc_hd__a22o_1
Xhold605 _6810_/Q VGND VGND VPWR VPWR hold605/X sky130_fd_sc_hd__bufbuf_16
Xhold616 _5465_/X VGND VGND VPWR VPWR _7034_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_170_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold638 _4150_/X VGND VGND VPWR VPWR _6620_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_116_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6231_ _6231_/A _6231_/B _6231_/C _6231_/D VGND VGND VPWR VPWR _6232_/C sky130_fd_sc_hd__or4_4
Xhold649 _6858_/Q VGND VGND VPWR VPWR hold649/X sky130_fd_sc_hd__bufbuf_16
X_3443_ _6906_/Q _5315_/A _5513_/A _7082_/Q _3430_/X VGND VGND VPWR VPWR _3451_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _7082_/Q _6311_/B VGND VGND VPWR VPWR _6162_/X sky130_fd_sc_hd__and2_1
X_5113_ _4871_/A _4989_/A _4995_/A VGND VGND VPWR VPWR _5114_/D sky130_fd_sc_hd__a21oi_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _3473_/A _3515_/B VGND VGND VPWR VPWR _5279_/A sky130_fd_sc_hd__nor2_8
XFILLER_112_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6093_ _7119_/Q _6023_/D _6030_/Y _7031_/Q _6092_/X VGND VGND VPWR VPWR _6093_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _4745_/A _4756_/B _5050_/C _4757_/B _5043_/X VGND VGND VPWR VPWR _5108_/A
+ sky130_fd_sc_hd__o221ai_2
XFILLER_111_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6995_ _7106_/CLK _6995_/D fanout434/X VGND VGND VPWR VPWR _6995_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_53_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5946_ _6776_/Q _5683_/X _5704_/X _6607_/Q _5945_/X VGND VGND VPWR VPWR _5953_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5877_ _6748_/Q _5682_/X _5700_/X _6535_/Q VGND VGND VPWR VPWR _5877_/X sky130_fd_sc_hd__a22o_1
X_4828_ _4687_/A _4898_/B _5147_/B VGND VGND VPWR VPWR _4828_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_139_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4759_ _5062_/B _4739_/X _4753_/X _4733_/X VGND VGND VPWR VPWR _4759_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_175_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6429_ _6446_/A _6446_/B VGND VGND VPWR VPWR _6429_/X sky130_fd_sc_hd__and2_1
XFILLER_134_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2 hold2/A VGND VGND VPWR VPWR hold2/X sky130_fd_sc_hd__bufbuf_16
XFILLER_67_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5800_ _6937_/Q _5704_/X _5799_/X _5698_/B VGND VGND VPWR VPWR _5800_/X sky130_fd_sc_hd__a22o_2
XFILLER_90_662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6780_ _7208_/CLK _6780_/D fanout458/X VGND VGND VPWR VPWR _6780_/Q sky130_fd_sc_hd__dfrtp_2
X_3992_ hold626/X _5583_/A0 _3994_/S VGND VGND VPWR VPWR _6494_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5731_ _7102_/Q _5675_/X _5684_/X _6990_/Q _5730_/X VGND VGND VPWR VPWR _5734_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5662_ _6832_/Q _5626_/A _6680_/Q _3918_/X _5661_/X VGND VGND VPWR VPWR _7175_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_191_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5593_ _5602_/A0 hold349/X _5593_/S VGND VGND VPWR VPWR _5593_/X sky130_fd_sc_hd__mux2_1
X_4613_ _4997_/A _4989_/A VGND VGND VPWR VPWR _4950_/A sky130_fd_sc_hd__nor2_4
Xhold402 _7066_/Q VGND VGND VPWR VPWR hold402/X sky130_fd_sc_hd__bufbuf_16
XFILLER_163_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4544_ _4987_/B _4586_/B _4542_/X _4543_/X VGND VGND VPWR VPWR _4546_/C sky130_fd_sc_hd__a211o_1
XFILLER_116_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold413 _6739_/Q VGND VGND VPWR VPWR hold413/X sky130_fd_sc_hd__bufbuf_16
Xhold424 _5476_/X VGND VGND VPWR VPWR _7044_/D sky130_fd_sc_hd__bufbuf_16
Xhold435 _7092_/Q VGND VGND VPWR VPWR hold435/X sky130_fd_sc_hd__bufbuf_16
Xhold457 _5492_/X VGND VGND VPWR VPWR _7058_/D sky130_fd_sc_hd__bufbuf_16
X_4475_ _4558_/B _4584_/A VGND VGND VPWR VPWR _4634_/B sky130_fd_sc_hd__nor2_8
Xhold468 _6890_/Q VGND VGND VPWR VPWR hold468/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold446 _6684_/Q VGND VGND VPWR VPWR hold446/X sky130_fd_sc_hd__bufbuf_16
X_6214_ _7020_/Q _6036_/Y _6335_/B _7044_/Q _6211_/X VGND VGND VPWR VPWR _6219_/B
+ sky130_fd_sc_hd__a221o_1
X_3426_ _7058_/Q _5486_/A hold85/A _7114_/Q VGND VGND VPWR VPWR _3426_/X sky130_fd_sc_hd__a22o_4
Xhold479 _5401_/X VGND VGND VPWR VPWR _6977_/D sky130_fd_sc_hd__bufbuf_16
X_7194_ _7196_/CLK _7194_/D fanout435/X VGND VGND VPWR VPWR _7194_/Q sky130_fd_sc_hd__dfrtp_4
X_6145_ _7113_/Q _6027_/B _6021_/B _7153_/Q VGND VGND VPWR VPWR _6145_/X sky130_fd_sc_hd__a22o_1
XFILLER_112_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3357_ _7108_/Q hold21/A _5351_/A _6940_/Q _3354_/X VGND VGND VPWR VPWR _3377_/A
+ sky130_fd_sc_hd__a221o_2
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1113 _6877_/Q VGND VGND VPWR VPWR _5289_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1124 _5345_/X VGND VGND VPWR VPWR _6927_/D sky130_fd_sc_hd__bufbuf_16
X_6076_ _6958_/Q _6022_/C _6032_/X _7054_/Q VGND VGND VPWR VPWR _6076_/X sky130_fd_sc_hd__a22o_1
XFILLER_112_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1102 _4183_/X VGND VGND VPWR VPWR _6648_/D sky130_fd_sc_hd__bufbuf_16
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1146 _6935_/Q VGND VGND VPWR VPWR _5354_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1157 _5318_/X VGND VGND VPWR VPWR _6903_/D sky130_fd_sc_hd__bufbuf_16
Xhold1135 _6601_/Q VGND VGND VPWR VPWR _4127_/A0 sky130_fd_sc_hd__bufbuf_16
X_5027_ _4758_/C _4684_/Y _4941_/B _4653_/Y _4386_/Y VGND VGND VPWR VPWR _5163_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_85_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3288_ hold82/X hold18/X VGND VGND VPWR VPWR hold83/A sky130_fd_sc_hd__nand2b_4
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1168 _4143_/X VGND VGND VPWR VPWR _6614_/D sky130_fd_sc_hd__bufbuf_16
Xhold1179 _6563_/Q VGND VGND VPWR VPWR _4083_/A0 sky130_fd_sc_hd__bufbuf_16
XFILLER_73_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_308 input16/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_319 _3945_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6978_ _7122_/CLK _6978_/D fanout443/X VGND VGND VPWR VPWR _6978_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5929_ _6646_/Q _5685_/X _5706_/X _6651_/Q _5928_/X VGND VGND VPWR VPWR _5937_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_186_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold991 _4290_/X VGND VGND VPWR VPWR _6741_/D sky130_fd_sc_hd__bufbuf_16
Xhold980 _6808_/Q VGND VGND VPWR VPWR hold980/X sky130_fd_sc_hd__bufbuf_16
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4260_ hold742/X _4326_/A0 _4261_/S VGND VGND VPWR VPWR _4260_/X sky130_fd_sc_hd__mux2_1
X_3211_ _7088_/Q VGND VGND VPWR VPWR _3211_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4191_ _5234_/C _4191_/A1 _4195_/S VGND VGND VPWR VPWR _4191_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6901_ _6964_/CLK _6901_/D fanout445/X VGND VGND VPWR VPWR _6901_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_47_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6832_ _7104_/CLK _6832_/D fanout433/X VGND VGND VPWR VPWR _6832_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3975_ hold154/X _3975_/B VGND VGND VPWR VPWR _3975_/Y sky130_fd_sc_hd__nand2b_4
X_6763_ _6851_/CLK _6763_/D fanout417/X VGND VGND VPWR VPWR _6763_/Q sky130_fd_sc_hd__dfrtp_2
X_6694_ _7150_/CLK _6694_/D fanout446/X VGND VGND VPWR VPWR _6694_/Q sky130_fd_sc_hd__dfrtp_1
X_5714_ _6981_/Q _5698_/B _5705_/X _6941_/Q _5697_/X VGND VGND VPWR VPWR _5714_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5645_ _5648_/B _6035_/A VGND VGND VPWR VPWR _5645_/Y sky130_fd_sc_hd__nand2_1
XFILLER_176_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold210 _5592_/X VGND VGND VPWR VPWR _7147_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5576_ hold61/X _5576_/B VGND VGND VPWR VPWR hold62/A sky130_fd_sc_hd__nand2_8
XFILLER_191_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold243 _4140_/X VGND VGND VPWR VPWR _6612_/D sky130_fd_sc_hd__bufbuf_16
Xhold232 _6602_/Q VGND VGND VPWR VPWR hold232/X sky130_fd_sc_hd__bufbuf_16
X_4527_ _4986_/A _4648_/B VGND VGND VPWR VPWR _4805_/A sky130_fd_sc_hd__nor2_1
XFILLER_117_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold221 _7096_/Q VGND VGND VPWR VPWR hold221/X sky130_fd_sc_hd__bufbuf_16
Xhold254 _6676_/Q VGND VGND VPWR VPWR hold254/X sky130_fd_sc_hd__bufbuf_16
X_4458_ _4558_/B _4818_/B VGND VGND VPWR VPWR _4989_/A sky130_fd_sc_hd__or2_4
XFILLER_132_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold265 _5285_/X VGND VGND VPWR VPWR _6874_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_116_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold276 _5437_/X VGND VGND VPWR VPWR _7009_/D sky130_fd_sc_hd__bufbuf_16
Xhold287 _3386_/B VGND VGND VPWR VPWR _3515_/B sky130_fd_sc_hd__bufbuf_16
X_3409_ _6899_/Q _5306_/A _5227_/A _3385_/X VGND VGND VPWR VPWR _3409_/X sky130_fd_sc_hd__a22o_1
Xhold298 _5455_/X VGND VGND VPWR VPWR _7025_/D sky130_fd_sc_hd__bufbuf_16
X_7177_ _7197_/CLK _7177_/D fanout431/X VGND VGND VPWR VPWR _7177_/Q sky130_fd_sc_hd__dfrtp_4
X_4389_ _4507_/A _4851_/B VGND VGND VPWR VPWR _4405_/B sky130_fd_sc_hd__nand2_8
X_6128_ _6872_/Q _6023_/C _6025_/B _6896_/Q _6127_/X VGND VGND VPWR VPWR _6131_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _6059_/A _6059_/B _6059_/C _6059_/D VGND VGND VPWR VPWR _6059_/X sky130_fd_sc_hd__or4_4
XFILLER_105_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_116 _4033_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_105 _3802_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 _5503_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 _5691_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_149 _5703_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3760_ _7117_/Q _5558_/A _5245_/A input61/X _3741_/X VGND VGND VPWR VPWR _3764_/A
+ sky130_fd_sc_hd__a221o_4
XFILLER_192_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5430_ _5601_/A0 hold628/X hold48/X VGND VGND VPWR VPWR _7003_/D sky130_fd_sc_hd__mux2_1
X_3691_ _7062_/Q _3317_/Y _4130_/A _6605_/Q _3671_/X VGND VGND VPWR VPWR _3693_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput315 _7228_/X VGND VGND VPWR VPWR spimemio_flash_io2_di sky130_fd_sc_hd__buf_8
XFILLER_173_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput326 _6556_/Q VGND VGND VPWR VPWR wb_dat_o[17] sky130_fd_sc_hd__buf_8
X_5361_ _5541_/A0 _5361_/A1 _5368_/S VGND VGND VPWR VPWR _6941_/D sky130_fd_sc_hd__mux2_1
Xoutput304 _6823_/Q VGND VGND VPWR VPWR pwr_ctrl_out[3] sky130_fd_sc_hd__buf_8
Xoutput337 _7206_/Q VGND VGND VPWR VPWR wb_dat_o[27] sky130_fd_sc_hd__buf_8
X_5292_ _5571_/A0 hold636/X _5296_/S VGND VGND VPWR VPWR _6880_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput348 _6568_/Q VGND VGND VPWR VPWR wb_dat_o[8] sky130_fd_sc_hd__buf_8
X_4312_ hold453/X _6408_/A0 _4315_/S VGND VGND VPWR VPWR _4312_/X sky130_fd_sc_hd__mux2_1
X_7100_ _7101_/CLK _7100_/D fanout431/X VGND VGND VPWR VPWR _7100_/Q sky130_fd_sc_hd__dfrtp_2
X_4243_ _5596_/A0 hold317/X _4249_/S VGND VGND VPWR VPWR _4243_/X sky130_fd_sc_hd__mux2_1
X_7031_ _7118_/CLK _7031_/D fanout436/X VGND VGND VPWR VPWR _7031_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_113_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4174_ hold910/X _5254_/A0 _4177_/S VGND VGND VPWR VPWR _4174_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6815_ _6825_/CLK _6815_/D fanout429/X VGND VGND VPWR VPWR _6815_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_23_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6746_ _6746_/CLK _6746_/D fanout427/X VGND VGND VPWR VPWR _6746_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3958_ _6473_/Q _6446_/A VGND VGND VPWR VPWR _3958_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3889_ _4368_/A _4722_/A VGND VGND VPWR VPWR _4346_/S sky130_fd_sc_hd__and2_2
XFILLER_137_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6677_ _7196_/CLK _6677_/D fanout433/X VGND VGND VPWR VPWR _6677_/Q sky130_fd_sc_hd__dfstp_4
X_5628_ _5663_/B _5702_/B _5705_/B _7162_/Q _5621_/X VGND VGND VPWR VPWR _7162_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_164_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5559_ _5595_/A0 hold984/X _5566_/S VGND VGND VPWR VPWR _7117_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7229_ _7229_/A VGND VGND VPWR VPWR _7229_/X sky130_fd_sc_hd__buf_2
XFILLER_132_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A VGND VGND VPWR VPWR _7197_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4930_ _4426_/A _4707_/A _4930_/C _4930_/D VGND VGND VPWR VPWR _4930_/X sky130_fd_sc_hd__and4bb_1
XFILLER_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4861_ _4376_/Y _4845_/B _5136_/C _4859_/X _4860_/X VGND VGND VPWR VPWR _4863_/C
+ sky130_fd_sc_hd__a2111o_2
XFILLER_17_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6600_ _6725_/CLK _6600_/D fanout440/X VGND VGND VPWR VPWR _6600_/Q sky130_fd_sc_hd__dfrtp_2
X_3812_ _6664_/Q _3812_/B VGND VGND VPWR VPWR _3840_/S sky130_fd_sc_hd__nand2b_4
XFILLER_32_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4792_ _4775_/A _4776_/A _4776_/B _5147_/B _4745_/A VGND VGND VPWR VPWR _4793_/A
+ sky130_fd_sc_hd__o32a_1
XANTENNA_27 _6893_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 _5963_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_16 _6782_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_49 _3331_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3743_ _7037_/Q _3334_/Y _5216_/A _6819_/Q VGND VGND VPWR VPWR _3743_/X sky130_fd_sc_hd__a22o_1
X_6531_ _6786_/CLK _6531_/D fanout417/X VGND VGND VPWR VPWR _6531_/Q sky130_fd_sc_hd__dfrtp_2
X_6462_ _3938_/A1 _6462_/D _6417_/X VGND VGND VPWR VPWR _6462_/Q sky130_fd_sc_hd__dfrtp_2
X_3674_ _7150_/Q _5594_/A _5245_/A input62/X VGND VGND VPWR VPWR _3674_/X sky130_fd_sc_hd__a22o_4
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6393_ _6707_/Q _6393_/A2 _6393_/B1 _4238_/B _6392_/X VGND VGND VPWR VPWR _6393_/X
+ sky130_fd_sc_hd__a221o_1
X_5413_ hold370/X _5602_/A0 _5413_/S VGND VGND VPWR VPWR _5413_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5344_ _5596_/A0 hold311/X _5350_/S VGND VGND VPWR VPWR _6926_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5275_ _5599_/A0 hold620/X hold29/X VGND VGND VPWR VPWR _5275_/X sky130_fd_sc_hd__mux2_1
Xoutput189 _3218_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[22] sky130_fd_sc_hd__buf_8
XFILLER_141_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput178 _3228_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[12] sky130_fd_sc_hd__buf_8
XFILLER_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7014_ _7135_/CLK _7014_/D fanout430/X VGND VGND VPWR VPWR _7014_/Q sky130_fd_sc_hd__dfstp_2
X_4226_ _5256_/A1 hold136/X _4234_/S VGND VGND VPWR VPWR _4226_/X sky130_fd_sc_hd__mux2_1
X_4157_ _4157_/A0 _5588_/A0 _4159_/S VGND VGND VPWR VPWR _6626_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4088_ _6700_/Q _6362_/B VGND VGND VPWR VPWR _4096_/S sky130_fd_sc_hd__and2_4
XFILLER_56_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6729_ _6804_/CLK _6729_/D _6439_/A VGND VGND VPWR VPWR _6729_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_52_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7035_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_127_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_67_csclk _6722_/CLK VGND VGND VPWR VPWR _7103_/CLK sky130_fd_sc_hd__clkbuf_8
Xfanout361 _4588_/X VGND VGND VPWR VPWR _4898_/B sky130_fd_sc_hd__buf_8
XFILLER_120_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout383 _4326_/A0 VGND VGND VPWR VPWR _6410_/A0 sky130_fd_sc_hd__buf_8
Xfanout372 hold209/A VGND VGND VPWR VPWR _5583_/A0 sky130_fd_sc_hd__buf_8
XFILLER_143_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout394 _6408_/A0 VGND VGND VPWR VPWR _5254_/A0 sky130_fd_sc_hd__buf_8
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput36 mgmt_gpio_in[0] VGND VGND VPWR VPWR _3971_/A sky130_fd_sc_hd__buf_8
Xinput14 mask_rev_in[19] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__clkbuf_4
Xinput25 mask_rev_in[29] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__clkbuf_4
XFILLER_183_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold809 _4146_/X VGND VGND VPWR VPWR _6617_/D sky130_fd_sc_hd__bufbuf_16
Xinput69 mgmt_gpio_in[6] VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__clkbuf_4
Xinput58 mgmt_gpio_in[2] VGND VGND VPWR VPWR _3875_/B sky130_fd_sc_hd__buf_8
Xinput47 mgmt_gpio_in[1] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__clkbuf_4
XFILLER_182_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3390_ _6891_/Q _5297_/A _5405_/A _6987_/Q VGND VGND VPWR VPWR _3390_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5060_ _5060_/A _5060_/B VGND VGND VPWR VPWR _5133_/A sky130_fd_sc_hd__or2_4
XFILLER_111_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4011_ hold321/X _5596_/A0 _4023_/S VGND VGND VPWR VPWR _4011_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5962_ _7187_/Q _6309_/S _5961_/X VGND VGND VPWR VPWR _7187_/D sky130_fd_sc_hd__o21a_1
XFILLER_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4913_ _4978_/B _4913_/B _4913_/C _5069_/C VGND VGND VPWR VPWR _4913_/X sky130_fd_sc_hd__or4_1
XFILLER_178_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5893_ _5893_/A _5893_/B _5893_/C _5893_/D VGND VGND VPWR VPWR _5893_/X sky130_fd_sc_hd__or4_2
X_4844_ _4844_/A _4844_/B VGND VGND VPWR VPWR _5086_/A sky130_fd_sc_hd__nor2_1
XFILLER_60_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4775_ _4775_/A _4927_/B VGND VGND VPWR VPWR _5099_/B sky130_fd_sc_hd__nor2_1
XFILLER_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6514_ _7141_/CLK _6514_/D fanout447/X VGND VGND VPWR VPWR _6514_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_165_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3726_ _3726_/A _3726_/B _3726_/C _3726_/D VGND VGND VPWR VPWR _3727_/D sky130_fd_sc_hd__or4_1
XFILLER_174_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3657_ _7063_/Q _3317_/Y _3341_/Y _7095_/Q VGND VGND VPWR VPWR _3657_/X sky130_fd_sc_hd__a22o_1
X_6445_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6445_/X sky130_fd_sc_hd__and2_1
X_6376_ _6376_/A _6376_/B _6376_/C _6374_/X VGND VGND VPWR VPWR _6400_/S sky130_fd_sc_hd__or4b_4
XFILLER_164_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3588_ _3588_/A _3588_/B _3588_/C _3588_/D VGND VGND VPWR VPWR _3606_/A sky130_fd_sc_hd__or4_4
X_5327_ _5597_/A0 hold511/X _5332_/S VGND VGND VPWR VPWR _5327_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5258_ _5582_/A0 hold700/X _5260_/S VGND VGND VPWR VPWR _5258_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4209_ hold641/X _5571_/A0 _4217_/S VGND VGND VPWR VPWR _4209_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5189_ _6410_/A0 hold970/X _5190_/S VGND VGND VPWR VPWR _5189_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4560_ _4812_/A _4697_/A VGND VGND VPWR VPWR _4562_/B sky130_fd_sc_hd__or2_4
XFILLER_156_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold617 _6984_/Q VGND VGND VPWR VPWR hold617/X sky130_fd_sc_hd__bufbuf_16
X_4491_ _5004_/A _4659_/A VGND VGND VPWR VPWR _4648_/B sky130_fd_sc_hd__nand2_8
X_3511_ _3540_/A _3528_/B VGND VGND VPWR VPWR _3511_/Y sky130_fd_sc_hd__nor2_8
Xhold606 _5206_/X VGND VGND VPWR VPWR _6810_/D sky130_fd_sc_hd__bufbuf_16
Xhold628 _7003_/Q VGND VGND VPWR VPWR hold628/X sky130_fd_sc_hd__bufbuf_16
X_3442_ _7146_/Q _5585_/A _5369_/A _6954_/Q _3441_/X VGND VGND VPWR VPWR _3451_/A
+ sky130_fd_sc_hd__a221o_4
X_6230_ _6980_/Q _6023_/B _6021_/C _6884_/Q _6229_/X VGND VGND VPWR VPWR _6231_/D
+ sky130_fd_sc_hd__a221o_1
Xhold639 _7107_/Q VGND VGND VPWR VPWR hold639/X sky130_fd_sc_hd__bufbuf_16
X_6161_ _6978_/Q _6023_/B _6021_/C _6882_/Q VGND VGND VPWR VPWR _6161_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3373_ _7124_/Q _5558_/A _5405_/A _6988_/Q VGND VGND VPWR VPWR _3373_/X sky130_fd_sc_hd__a22o_1
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5112_ _6782_/Q _6376_/A _5038_/Y _5111_/X _5103_/X VGND VGND VPWR VPWR _5112_/X
+ sky130_fd_sc_hd__a221o_4
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _6999_/Q _5987_/Y _6022_/D _6919_/Q VGND VGND VPWR VPWR _6092_/X sky130_fd_sc_hd__a22o_1
XFILLER_85_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _4818_/A _4566_/A _4756_/B _4893_/B VGND VGND VPWR VPWR _5043_/X sky130_fd_sc_hd__o31a_2
XFILLER_78_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_wbbd_sck _7219_/Q VGND VGND VPWR VPWR clkbuf_0_wbbd_sck/X sky130_fd_sc_hd__clkbuf_8
XFILLER_80_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6994_ _7106_/CLK _6994_/D fanout438/X VGND VGND VPWR VPWR _6994_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_80_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5945_ _6731_/Q _5667_/X _5687_/X _6642_/Q VGND VGND VPWR VPWR _5945_/X sky130_fd_sc_hd__a22o_1
XFILLER_43_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5876_ _6785_/Q _5690_/X _5705_/X _6609_/Q _5875_/X VGND VGND VPWR VPWR _5883_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4827_ _4827_/A _5013_/B _5047_/C _4826_/X VGND VGND VPWR VPWR _4834_/B sky130_fd_sc_hd__or4b_1
XFILLER_178_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4758_ _4758_/A _4758_/B _4758_/C VGND VGND VPWR VPWR _5105_/A sky130_fd_sc_hd__and3_1
XFILLER_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3709_ _3709_/A _3709_/B _3709_/C _3709_/D VGND VGND VPWR VPWR _3709_/X sky130_fd_sc_hd__or4_4
X_4689_ _4717_/B VGND VGND VPWR VPWR _4689_/Y sky130_fd_sc_hd__inv_6
XFILLER_4_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6428_ _6455_/A _6446_/B VGND VGND VPWR VPWR _6428_/X sky130_fd_sc_hd__and2_1
XFILLER_162_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6359_ _7201_/Q _6309_/S _6357_/X _6358_/X VGND VGND VPWR VPWR _7201_/D sky130_fd_sc_hd__o22a_1
XFILLER_191_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3 hold3/A VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__bufbuf_16
XFILLER_121_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3991_ hold205/X _7217_/Q _3991_/S VGND VGND VPWR VPWR _3991_/X sky130_fd_sc_hd__mux2_8
XFILLER_90_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5730_ _6878_/Q _5674_/X _5688_/X _7030_/Q VGND VGND VPWR VPWR _5730_/X sky130_fd_sc_hd__a22o_1
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5661_ _6677_/Q _5659_/C _7175_/Q VGND VGND VPWR VPWR _5661_/X sky130_fd_sc_hd__a21o_1
X_4612_ _4612_/A _4612_/B _4612_/C _4612_/D VGND VGND VPWR VPWR _4615_/B sky130_fd_sc_hd__and4_4
X_5592_ hold209/X _5592_/A1 _5593_/S VGND VGND VPWR VPWR _5592_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4543_ _4772_/A _4409_/Y _4412_/Y _5116_/A VGND VGND VPWR VPWR _4543_/X sky130_fd_sc_hd__a211o_1
XFILLER_116_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold403 _5501_/X VGND VGND VPWR VPWR _7066_/D sky130_fd_sc_hd__bufbuf_16
Xhold425 _6835_/Q VGND VGND VPWR VPWR hold425/X sky130_fd_sc_hd__bufbuf_16
XFILLER_144_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold414 _4288_/X VGND VGND VPWR VPWR _6739_/D sky130_fd_sc_hd__bufbuf_16
Xhold436 _5530_/X VGND VGND VPWR VPWR _7092_/D sky130_fd_sc_hd__bufbuf_16
Xhold458 _6694_/Q VGND VGND VPWR VPWR hold458/X sky130_fd_sc_hd__bufbuf_16
Xhold469 _5303_/X VGND VGND VPWR VPWR _6890_/D sky130_fd_sc_hd__bufbuf_16
X_4474_ _4949_/A _4956_/A VGND VGND VPWR VPWR _4603_/B sky130_fd_sc_hd__nand2_8
XFILLER_144_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold447 _4227_/X VGND VGND VPWR VPWR _6684_/D sky130_fd_sc_hd__bufbuf_16
X_6213_ _7028_/Q _6010_/Y _6031_/X _7092_/Q _6212_/X VGND VGND VPWR VPWR _6219_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3425_ _6938_/Q _5351_/A _5279_/A _6874_/Q VGND VGND VPWR VPWR _3425_/X sky130_fd_sc_hd__a22o_1
X_7193_ _7193_/CLK _7193_/D fanout435/X VGND VGND VPWR VPWR _7193_/Q sky130_fd_sc_hd__dfrtp_4
X_6144_ _6144_/A _6144_/B _6144_/C _6144_/D VGND VGND VPWR VPWR _6144_/X sky130_fd_sc_hd__or4_2
XFILLER_98_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3356_ _3457_/A _3515_/B VGND VGND VPWR VPWR _5351_/A sky130_fd_sc_hd__nor2_8
XFILLER_161_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6075_ _6902_/Q _6021_/A _6025_/A _6934_/Q _6074_/X VGND VGND VPWR VPWR _6082_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_100_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1103 _6646_/Q VGND VGND VPWR VPWR _4181_/A0 sky130_fd_sc_hd__bufbuf_16
XFILLER_58_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1114 _6773_/Q VGND VGND VPWR VPWR _4329_/A1 sky130_fd_sc_hd__bufbuf_16
X_3287_ input33/X _3283_/Y hold54/A _7092_/Q VGND VGND VPWR VPWR _3287_/X sky130_fd_sc_hd__a22o_1
Xhold1136 _6895_/Q VGND VGND VPWR VPWR _5309_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1147 _5354_/X VGND VGND VPWR VPWR _6935_/D sky130_fd_sc_hd__bufbuf_16
X_5026_ _5164_/A _4990_/A _4926_/X _5025_/X VGND VGND VPWR VPWR _5098_/B sky130_fd_sc_hd__o211ai_4
XFILLER_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1125 _6576_/Q VGND VGND VPWR VPWR _4098_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1158 _7221_/Q VGND VGND VPWR VPWR _6407_/A1 sky130_fd_sc_hd__bufbuf_16
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1169 _6720_/Q VGND VGND VPWR VPWR _4265_/A0 sky130_fd_sc_hd__bufbuf_16
XFILLER_38_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_309 input116/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6977_ _7133_/CLK _6977_/D fanout443/X VGND VGND VPWR VPWR _6977_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5928_ _6636_/Q _5675_/X _5683_/X _6775_/Q VGND VGND VPWR VPWR _5928_/X sky130_fd_sc_hd__a22o_1
XFILLER_41_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5859_ _6916_/Q _5680_/X _5689_/X _6908_/Q VGND VGND VPWR VPWR _5859_/X sky130_fd_sc_hd__a22o_1
XFILLER_182_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold981 _5204_/X VGND VGND VPWR VPWR _6808_/D sky130_fd_sc_hd__bufbuf_16
Xhold970 _6788_/Q VGND VGND VPWR VPWR hold970/X sky130_fd_sc_hd__bufbuf_16
XFILLER_135_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold992 _6641_/Q VGND VGND VPWR VPWR hold992/X sky130_fd_sc_hd__bufbuf_16
XFILLER_103_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3210_ _7096_/Q VGND VGND VPWR VPWR _3210_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4190_ _4190_/A _6406_/B VGND VGND VPWR VPWR _4195_/S sky130_fd_sc_hd__nand2_4
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6900_ _7156_/CLK _6900_/D fanout444/X VGND VGND VPWR VPWR _6900_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_63_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6831_ _7035_/CLK _6831_/D fanout433/X VGND VGND VPWR VPWR _6831_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3974_ _6707_/Q _3974_/B VGND VGND VPWR VPWR _6699_/D sky130_fd_sc_hd__and2_1
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6762_ _7225_/CLK _6762_/D fanout420/X VGND VGND VPWR VPWR _6762_/Q sky130_fd_sc_hd__dfrtp_2
X_6693_ _6939_/CLK _6693_/D fanout453/X VGND VGND VPWR VPWR _6693_/Q sky130_fd_sc_hd__dfrtp_1
X_5713_ _6901_/Q _5689_/X _5710_/X _5712_/X VGND VGND VPWR VPWR _5713_/X sky130_fd_sc_hd__a211o_4
XFILLER_148_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5644_ _7169_/Q _7168_/Q VGND VGND VPWR VPWR _6035_/A sky130_fd_sc_hd__and2_4
XFILLER_191_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold200 _7215_/Q VGND VGND VPWR VPWR hold200/X sky130_fd_sc_hd__bufbuf_16
XFILLER_163_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold211 _6567_/Q VGND VGND VPWR VPWR hold211/X sky130_fd_sc_hd__bufbuf_16
X_5575_ _5584_/A0 hold439/X _5575_/S VGND VGND VPWR VPWR _5575_/X sky130_fd_sc_hd__mux2_1
X_4526_ _4749_/C _4965_/A VGND VGND VPWR VPWR _4557_/C sky130_fd_sc_hd__nor2_1
Xhold233 _4128_/X VGND VGND VPWR VPWR _6602_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_117_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold222 _6484_/Q VGND VGND VPWR VPWR _3255_/B sky130_fd_sc_hd__bufbuf_16
Xhold244 _7136_/Q VGND VGND VPWR VPWR hold244/X sky130_fd_sc_hd__bufbuf_16
Xhold255 _4218_/X VGND VGND VPWR VPWR _6676_/D sky130_fd_sc_hd__bufbuf_16
X_4457_ _4558_/B _4818_/B VGND VGND VPWR VPWR _4868_/A sky130_fd_sc_hd__nor2_8
XFILLER_171_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold277 _6857_/Q VGND VGND VPWR VPWR hold277/X sky130_fd_sc_hd__bufbuf_16
Xhold266 _7048_/Q VGND VGND VPWR VPWR hold266/X sky130_fd_sc_hd__bufbuf_16
XFILLER_172_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold299 _7081_/Q VGND VGND VPWR VPWR hold299/X sky130_fd_sc_hd__bufbuf_16
X_3408_ _6859_/Q _3315_/Y _4217_/S input50/X _3407_/X VGND VGND VPWR VPWR _3414_/A
+ sky130_fd_sc_hd__a221o_1
Xhold288 _3317_/Y VGND VGND VPWR VPWR _5495_/A sky130_fd_sc_hd__bufbuf_16
X_7176_ _7197_/CLK _7176_/D fanout431/X VGND VGND VPWR VPWR _7176_/Q sky130_fd_sc_hd__dfrtp_4
X_4388_ _4478_/C _4388_/B VGND VGND VPWR VPWR _4851_/B sky130_fd_sc_hd__and2_4
XFILLER_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6127_ _6960_/Q _6022_/C _6032_/X _7056_/Q VGND VGND VPWR VPWR _6127_/X sky130_fd_sc_hd__a22o_1
XFILLER_86_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _3514_/A _5225_/B VGND VGND VPWR VPWR _5459_/A sky130_fd_sc_hd__nor2_8
X_6058_ _6306_/A _6058_/B _6058_/C VGND VGND VPWR VPWR _6059_/D sky130_fd_sc_hd__or3_1
XFILLER_100_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5009_ _5004_/A _4469_/Y _4652_/B _4494_/Y VGND VGND VPWR VPWR _5105_/B sky130_fd_sc_hd__a31o_1
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_106 _3841_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_128 _5503_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_139 _5694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_117 _4209_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3690_ _6910_/Q _5324_/A _5297_/A _6886_/Q _3689_/X VGND VGND VPWR VPWR _3693_/B
+ sky130_fd_sc_hd__a221o_4
XFILLER_161_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput316 _7229_/X VGND VGND VPWR VPWR spimemio_flash_io3_di sky130_fd_sc_hd__buf_8
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput305 _3730_/X VGND VGND VPWR VPWR reset sky130_fd_sc_hd__buf_8
X_5360_ _5360_/A _5576_/B VGND VGND VPWR VPWR _5368_/S sky130_fd_sc_hd__nand2_8
X_5291_ _5588_/A0 _5291_/A1 _5296_/S VGND VGND VPWR VPWR _5291_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput338 _7207_/Q VGND VGND VPWR VPWR wb_dat_o[28] sky130_fd_sc_hd__buf_8
Xoutput327 _6557_/Q VGND VGND VPWR VPWR wb_dat_o[18] sky130_fd_sc_hd__buf_8
XFILLER_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput349 _6569_/Q VGND VGND VPWR VPWR wb_dat_o[9] sky130_fd_sc_hd__buf_8
X_4311_ _4311_/A0 _6407_/A0 _4315_/S VGND VGND VPWR VPWR _4311_/X sky130_fd_sc_hd__mux2_1
X_4242_ _5289_/A0 hold956/X _4249_/S VGND VGND VPWR VPWR _4242_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7030_ _7134_/CLK _7030_/D fanout429/X VGND VGND VPWR VPWR _7030_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_113_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4173_ _4173_/A0 _5234_/C _4177_/S VGND VGND VPWR VPWR _4173_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6814_ _6825_/CLK _6814_/D fanout421/X VGND VGND VPWR VPWR _6814_/Q sky130_fd_sc_hd__dfstp_2
X_6745_ _6745_/CLK _6745_/D fanout442/X VGND VGND VPWR VPWR _6745_/Q sky130_fd_sc_hd__dfstp_4
X_3957_ input83/X _3957_/A1 _6473_/Q VGND VGND VPWR VPWR _3957_/X sky130_fd_sc_hd__mux2_1
XFILLER_167_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6676_ _7127_/CLK _6676_/D fanout448/X VGND VGND VPWR VPWR _6676_/Q sky130_fd_sc_hd__dfrtp_2
X_3888_ _4350_/C _4350_/D _4349_/A _4349_/B VGND VGND VPWR VPWR _3895_/C sky130_fd_sc_hd__or4_2
XFILLER_136_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5627_ _6677_/Q _5663_/B VGND VGND VPWR VPWR _5635_/B sky130_fd_sc_hd__nand2_4
X_5558_ _5558_/A _5558_/B VGND VGND VPWR VPWR _5566_/S sky130_fd_sc_hd__nand2_8
XFILLER_132_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4509_ _4996_/A _4775_/A VGND VGND VPWR VPWR _4920_/B sky130_fd_sc_hd__nor2_1
XFILLER_117_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5489_ _5588_/A0 hold938/X _5494_/S VGND VGND VPWR VPWR _5489_/X sky130_fd_sc_hd__mux2_1
X_7228_ _7228_/A VGND VGND VPWR VPWR _7228_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_105_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7159_ _7196_/CLK _7159_/D fanout433/X VGND VGND VPWR VPWR _7159_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_100_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4860_ _4575_/B _4845_/B _5079_/B _5079_/A VGND VGND VPWR VPWR _4860_/X sky130_fd_sc_hd__a211o_1
XANTENNA_470 hold209/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3811_ _6666_/Q _3843_/B _3898_/B _3845_/A VGND VGND VPWR VPWR _3812_/B sky130_fd_sc_hd__a31o_4
XFILLER_33_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_28 _6896_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4791_ _4772_/A _5165_/A _4772_/C _4936_/A VGND VGND VPWR VPWR _4791_/X sky130_fd_sc_hd__a31o_1
XFILLER_119_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_17 _6782_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 _5963_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6530_ _6786_/CLK _6530_/D fanout417/X VGND VGND VPWR VPWR _6530_/Q sky130_fd_sc_hd__dfrtp_2
X_3742_ input52/X _4025_/A _5594_/A _7149_/Q VGND VGND VPWR VPWR _3742_/X sky130_fd_sc_hd__a22o_4
XFILLER_158_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6461_ _3938_/A1 _6461_/D _6416_/X VGND VGND VPWR VPWR hold38/A sky130_fd_sc_hd__dfrtp_2
XFILLER_146_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3673_ _5225_/A _3673_/B VGND VGND VPWR VPWR _5191_/A sky130_fd_sc_hd__nor2_4
X_6392_ _6705_/Q _6392_/A2 _6392_/B1 _6706_/Q VGND VGND VPWR VPWR _6392_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5412_ hold560/X _5601_/A0 _5413_/S VGND VGND VPWR VPWR _5412_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5343_ _5595_/A0 hold962/X _5350_/S VGND VGND VPWR VPWR _6925_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5274_ hold71/X hold171/X hold29/X VGND VGND VPWR VPWR _5274_/X sky130_fd_sc_hd__mux2_1
Xoutput179 _3227_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[13] sky130_fd_sc_hd__buf_8
XFILLER_68_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7013_ _7135_/CLK _7013_/D fanout428/X VGND VGND VPWR VPWR _7013_/Q sky130_fd_sc_hd__dfstp_4
X_4225_ hold921/X _4224_/X _4235_/S VGND VGND VPWR VPWR _4225_/X sky130_fd_sc_hd__mux2_1
X_4156_ hold535/X _5587_/A0 _4159_/S VGND VGND VPWR VPWR _4156_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4087_ hold211/X _5581_/A0 _4087_/S VGND VGND VPWR VPWR _4087_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4989_ _4989_/A _4989_/B VGND VGND VPWR VPWR _5121_/C sky130_fd_sc_hd__nor2_1
XFILLER_23_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6728_ _6804_/CLK _6728_/D _6439_/A VGND VGND VPWR VPWR _6728_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_176_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6659_ _6845_/CLK _6659_/D fanout417/X VGND VGND VPWR VPWR _6659_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout373 hold209/A VGND VGND VPWR VPWR _5601_/A0 sky130_fd_sc_hd__buf_8
XFILLER_120_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout384 hold136/X VGND VGND VPWR VPWR _4326_/A0 sky130_fd_sc_hd__buf_8
Xfanout362 hold47/X VGND VGND VPWR VPWR _6406_/B sky130_fd_sc_hd__buf_8
XFILLER_101_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout395 hold67/X VGND VGND VPWR VPWR _6408_/A0 sky130_fd_sc_hd__buf_8
XFILLER_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput37 mgmt_gpio_in[10] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput26 mask_rev_in[2] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__clkbuf_4
Xinput15 mask_rev_in[1] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__clkbuf_4
Xinput48 mgmt_gpio_in[20] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__clkbuf_4
XFILLER_143_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput59 mgmt_gpio_in[30] VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__buf_6
XFILLER_128_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4010_ hold948/X _4009_/X _4024_/S VGND VGND VPWR VPWR _4010_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5961_ _5611_/A _7186_/Q _6358_/B1 _5960_/X VGND VGND VPWR VPWR _5961_/X sky130_fd_sc_hd__a211o_1
XFILLER_52_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4912_ _5062_/A _4898_/B _4603_/B VGND VGND VPWR VPWR _5069_/C sky130_fd_sc_hd__a21oi_1
X_5892_ _6768_/Q _5688_/X _5692_/X _7221_/Q _5891_/X VGND VGND VPWR VPWR _5893_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4843_ _5023_/A _4986_/C VGND VGND VPWR VPWR _4845_/B sky130_fd_sc_hd__nand2_8
XFILLER_21_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4774_ _4774_/A _4776_/B _4774_/C _4930_/C VGND VGND VPWR VPWR _4927_/B sky130_fd_sc_hd__or4b_4
XFILLER_159_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6513_ _7156_/CLK _6513_/D fanout447/X VGND VGND VPWR VPWR _6513_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_165_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3725_ _3725_/A _3725_/B _3725_/C _3725_/D VGND VGND VPWR VPWR _3726_/D sky130_fd_sc_hd__or4_1
XFILLER_146_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6444_ _6446_/A _6446_/B VGND VGND VPWR VPWR _6444_/X sky130_fd_sc_hd__and2_1
XFILLER_173_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3656_ _7007_/Q _5432_/A _3359_/Y _7015_/Q _3655_/X VGND VGND VPWR VPWR _3664_/B
+ sky130_fd_sc_hd__a221o_1
X_6375_ _6402_/A2 _6372_/A _6707_/Q VGND VGND VPWR VPWR _6376_/B sky130_fd_sc_hd__a21boi_1
XFILLER_164_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3587_ _3587_/A _3587_/B _3587_/C _3587_/D VGND VGND VPWR VPWR _3588_/D sky130_fd_sc_hd__or4_1
X_5326_ _5596_/A0 hold315/X _5332_/S VGND VGND VPWR VPWR _5326_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5257_ hold185/X hold293/X _5260_/S VGND VGND VPWR VPWR _5257_/X sky130_fd_sc_hd__mux2_1
X_4208_ hold887/X _4207_/X _4218_/S VGND VGND VPWR VPWR _4208_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5188_ _6409_/A0 hold996/X _5190_/S VGND VGND VPWR VPWR _6787_/D sky130_fd_sc_hd__mux2_1
X_4139_ _5588_/A0 _4139_/A1 _4141_/S VGND VGND VPWR VPWR _6611_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3510_ _5234_/A _3733_/B VGND VGND VPWR VPWR _4049_/A sky130_fd_sc_hd__nor2_8
X_4490_ _4651_/B _4746_/A VGND VGND VPWR VPWR _4819_/D sky130_fd_sc_hd__or2_1
XFILLER_183_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold618 _5409_/X VGND VGND VPWR VPWR _6984_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_143_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold607 _6645_/Q VGND VGND VPWR VPWR hold607/X sky130_fd_sc_hd__bufbuf_16
XFILLER_7_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold629 _7000_/Q VGND VGND VPWR VPWR hold629/X sky130_fd_sc_hd__bufbuf_16
X_3441_ _6970_/Q _5387_/A _4234_/S _3969_/A VGND VGND VPWR VPWR _3441_/X sky130_fd_sc_hd__a22o_4
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap359 hold60/X VGND VGND VPWR VPWR _5252_/A sky130_fd_sc_hd__buf_8
X_3372_ hold84/X _3457_/A VGND VGND VPWR VPWR _5405_/A sky130_fd_sc_hd__nor2_8
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6160_ _7193_/Q _5665_/Y _6159_/X VGND VGND VPWR VPWR _7193_/D sky130_fd_sc_hd__o21a_1
X_5111_ _5157_/B _5155_/A _5178_/B _5156_/C VGND VGND VPWR VPWR _5111_/X sky130_fd_sc_hd__or4_4
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6091_ _7015_/Q _6036_/Y _6335_/B _7039_/Q VGND VGND VPWR VPWR _6091_/X sky130_fd_sc_hd__a22o_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _4745_/A _5062_/C _4734_/X VGND VGND VPWR VPWR _5042_/Y sky130_fd_sc_hd__o21ai_2
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6993_ _7135_/CLK _6993_/D fanout431/X VGND VGND VPWR VPWR _6993_/Q sky130_fd_sc_hd__dfrtp_2
Xclkbuf_leaf_51_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7107_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_53_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5944_ _6647_/Q _5685_/X _5699_/X _6602_/Q VGND VGND VPWR VPWR _5944_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5875_ _6713_/Q _5676_/X _5702_/X _6550_/Q VGND VGND VPWR VPWR _5875_/X sky130_fd_sc_hd__a22o_1
X_4826_ _4562_/B _5062_/B _4725_/Y _4823_/X _4825_/X VGND VGND VPWR VPWR _4826_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_178_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4757_ _5062_/A _4757_/B VGND VGND VPWR VPWR _5174_/B sky130_fd_sc_hd__nor2_1
X_4688_ _4728_/A _4690_/A _5062_/B VGND VGND VPWR VPWR _4717_/B sky130_fd_sc_hd__or3_4
XFILLER_147_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3708_ _6650_/Q _4184_/A _4055_/A _6541_/Q _3680_/X VGND VGND VPWR VPWR _3709_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_107_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3639_ input22/X _3302_/Y _4286_/A _6740_/Q VGND VGND VPWR VPWR _3639_/X sky130_fd_sc_hd__a22o_1
X_6427_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6427_/X sky130_fd_sc_hd__and2_1
X_6358_ _5611_/A _7200_/Q _6358_/B1 VGND VGND VPWR VPWR _6358_/X sky130_fd_sc_hd__a21o_1
X_5309_ _5588_/A0 _5309_/A1 _5314_/S VGND VGND VPWR VPWR _5309_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6289_ _6750_/Q _6036_/Y _6335_/B _6775_/Q VGND VGND VPWR VPWR _6289_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_19_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7153_/CLK sky130_fd_sc_hd__clkbuf_8
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold4 hold4/A VGND VGND VPWR VPWR hold4/X sky130_fd_sc_hd__bufbuf_16
XFILLER_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3990_ hold613/X _5582_/A0 _3994_/S VGND VGND VPWR VPWR _6493_/D sky130_fd_sc_hd__mux2_1
Xnet399_2 _3545_/A1 VGND VGND VPWR VPWR _3953_/B sky130_fd_sc_hd__inv_2
XFILLER_90_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5660_ _7158_/Q _5659_/X _5658_/S _7174_/Q VGND VGND VPWR VPWR _7174_/D sky130_fd_sc_hd__a2bb2o_1
X_4611_ _4875_/A _5005_/C _4610_/Y _4564_/A _4593_/Y VGND VGND VPWR VPWR _4612_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5591_ _5600_/A0 hold451/X _5593_/S VGND VGND VPWR VPWR _5591_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4542_ _5033_/A _4542_/B _4542_/C _4542_/D VGND VGND VPWR VPWR _4542_/X sky130_fd_sc_hd__or4_1
XFILLER_128_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4473_ _4525_/A _4572_/A VGND VGND VPWR VPWR _4956_/A sky130_fd_sc_hd__nor2_8
Xhold426 _5240_/X VGND VGND VPWR VPWR _6835_/D sky130_fd_sc_hd__bufbuf_16
Xhold404 _6922_/Q VGND VGND VPWR VPWR hold404/X sky130_fd_sc_hd__bufbuf_16
XFILLER_7_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold415 _7078_/Q VGND VGND VPWR VPWR hold415/X sky130_fd_sc_hd__bufbuf_16
Xhold459 _4211_/X VGND VGND VPWR VPWR hold459/X sky130_fd_sc_hd__bufbuf_16
Xhold437 _7127_/Q VGND VGND VPWR VPWR hold437/X sky130_fd_sc_hd__bufbuf_16
X_3424_ _6962_/Q _5378_/A _5306_/A _6898_/Q VGND VGND VPWR VPWR _3424_/X sky130_fd_sc_hd__a22o_1
Xhold448 _7006_/Q VGND VGND VPWR VPWR hold448/X sky130_fd_sc_hd__bufbuf_16
X_6212_ _7140_/Q _6020_/B _6011_/X _7100_/Q VGND VGND VPWR VPWR _6212_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7192_ _7196_/CLK _7192_/D fanout432/X VGND VGND VPWR VPWR _7192_/Q sky130_fd_sc_hd__dfrtp_4
X_6143_ _6985_/Q _6028_/X _6034_/Y _6993_/Q _6142_/X VGND VGND VPWR VPWR _6144_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3355_ _3501_/A hold20/X VGND VGND VPWR VPWR hold21/A sky130_fd_sc_hd__nor2_8
X_6074_ _6950_/Q _6022_/A _6025_/C _6926_/Q VGND VGND VPWR VPWR _6074_/X sky130_fd_sc_hd__a22o_1
XFILLER_97_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1104 _6747_/Q VGND VGND VPWR VPWR _4297_/A1 sky130_fd_sc_hd__bufbuf_16
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ hold53/X _3673_/B VGND VGND VPWR VPWR hold54/A sky130_fd_sc_hd__nor2_8
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1115 _4329_/X VGND VGND VPWR VPWR _6773_/D sky130_fd_sc_hd__bufbuf_16
Xhold1148 _6879_/Q VGND VGND VPWR VPWR _5291_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1137 _5309_/X VGND VGND VPWR VPWR _6895_/D sky130_fd_sc_hd__bufbuf_16
X_5025_ _5164_/B _4756_/B _4746_/X _4724_/B VGND VGND VPWR VPWR _5025_/X sky130_fd_sc_hd__o22a_2
Xhold1126 _4098_/X VGND VGND VPWR VPWR _6576_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_57_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1159 _6407_/X VGND VGND VPWR VPWR _7221_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_93_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6976_ _6976_/CLK _6976_/D fanout450/X VGND VGND VPWR VPWR _6976_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5927_ _5927_/A _5927_/B _5927_/C _5927_/D VGND VGND VPWR VPWR _5927_/X sky130_fd_sc_hd__or4_4
XFILLER_110_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5858_ _6868_/Q _5700_/X _5857_/X VGND VGND VPWR VPWR _5861_/C sky130_fd_sc_hd__a21o_1
XFILLER_22_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4809_ _4697_/A _5005_/C _4746_/X VGND VGND VPWR VPWR _4809_/X sky130_fd_sc_hd__a21o_1
X_5789_ _6881_/Q _5674_/X _5694_/X _6897_/Q _5788_/X VGND VGND VPWR VPWR _5796_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold982 _6514_/Q VGND VGND VPWR VPWR hold982/X sky130_fd_sc_hd__bufbuf_16
Xhold960 _6917_/Q VGND VGND VPWR VPWR hold960/X sky130_fd_sc_hd__bufbuf_16
Xhold971 _5189_/X VGND VGND VPWR VPWR _6788_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_115_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold993 _6751_/Q VGND VGND VPWR VPWR hold993/X sky130_fd_sc_hd__bufbuf_16
XFILLER_192_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6830_ _7035_/CLK _6830_/D fanout432/X VGND VGND VPWR VPWR _6830_/Q sky130_fd_sc_hd__dfrtp_2
X_6761_ _7222_/CLK _6761_/D fanout420/X VGND VGND VPWR VPWR _6761_/Q sky130_fd_sc_hd__dfrtp_2
X_5712_ _6877_/Q _5674_/X _5690_/X _7093_/Q _5711_/X VGND VGND VPWR VPWR _5712_/X
+ sky130_fd_sc_hd__a221o_2
X_3973_ _6838_/Q _3973_/B VGND VGND VPWR VPWR _3973_/X sky130_fd_sc_hd__and2_4
X_6692_ _6939_/CLK _6692_/D fanout453/X VGND VGND VPWR VPWR _6692_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5643_ _7168_/Q _5648_/B _5642_/Y VGND VGND VPWR VPWR _7168_/D sky130_fd_sc_hd__a21oi_1
XFILLER_117_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5574_ _5583_/A0 hold651/X _5575_/S VGND VGND VPWR VPWR _5574_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold201 _3987_/X VGND VGND VPWR VPWR hold201/X sky130_fd_sc_hd__bufbuf_16
X_4525_ _4525_/A _4572_/A _4538_/A VGND VGND VPWR VPWR _4965_/A sky130_fd_sc_hd__or3b_4
XFILLER_132_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold212 _4087_/X VGND VGND VPWR VPWR _6567_/D sky130_fd_sc_hd__bufbuf_16
Xhold223 _3255_/X VGND VGND VPWR VPWR hold223/X sky130_fd_sc_hd__bufbuf_16
Xhold234 _7104_/Q VGND VGND VPWR VPWR hold234/X sky130_fd_sc_hd__bufbuf_16
Xhold267 _6526_/Q VGND VGND VPWR VPWR hold267/X sky130_fd_sc_hd__bufbuf_16
X_4456_ _4469_/A _4558_/B VGND VGND VPWR VPWR _4844_/A sky130_fd_sc_hd__or2_4
XFILLER_131_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold256 _6867_/Q VGND VGND VPWR VPWR hold256/X sky130_fd_sc_hd__bufbuf_16
Xhold278 _5266_/X VGND VGND VPWR VPWR _6857_/D sky130_fd_sc_hd__bufbuf_16
Xhold245 _5580_/X VGND VGND VPWR VPWR _7136_/D sky130_fd_sc_hd__bufbuf_16
Xhold289 _5497_/X VGND VGND VPWR VPWR _7062_/D sky130_fd_sc_hd__bufbuf_16
X_4387_ _4958_/A _4408_/A VGND VGND VPWR VPWR _4513_/A sky130_fd_sc_hd__or2_4
X_3407_ _7075_/Q hold92/A _5333_/A _6923_/Q VGND VGND VPWR VPWR _3407_/X sky130_fd_sc_hd__a22o_1
X_7175_ _7193_/CLK _7175_/D fanout435/X VGND VGND VPWR VPWR _7175_/Q sky130_fd_sc_hd__dfrtp_2
X_6126_ _6904_/Q _6021_/A _6025_/A _6936_/Q _6125_/X VGND VGND VPWR VPWR _6132_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_86_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3338_ _3473_/A _5225_/B VGND VGND VPWR VPWR _5315_/A sky130_fd_sc_hd__nor2_8
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6057_ _6057_/A _6057_/B _6057_/C _6057_/D VGND VGND VPWR VPWR _6058_/C sky130_fd_sc_hd__or4_1
XFILLER_85_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3269_ hold17/X hold325/X _3991_/S VGND VGND VPWR VPWR _3269_/X sky130_fd_sc_hd__mux2_8
X_5008_ _5008_/A _5008_/B VGND VGND VPWR VPWR _5012_/A sky130_fd_sc_hd__nand2_1
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 _3830_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_129 _5503_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 _6376_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6959_ _6959_/CLK _6959_/D fanout444/X VGND VGND VPWR VPWR _6959_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_10_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold790 _6772_/Q VGND VGND VPWR VPWR hold790/X sky130_fd_sc_hd__bufbuf_16
XFILLER_150_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput317 _7202_/Q VGND VGND VPWR VPWR wb_ack_o sky130_fd_sc_hd__buf_8
Xoutput306 _3969_/X VGND VGND VPWR VPWR ser_rx sky130_fd_sc_hd__buf_8
X_5290_ _5587_/A0 hold587/X _5296_/S VGND VGND VPWR VPWR _5290_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput339 _7208_/Q VGND VGND VPWR VPWR wb_dat_o[29] sky130_fd_sc_hd__buf_8
Xoutput328 _6558_/Q VGND VGND VPWR VPWR wb_dat_o[19] sky130_fd_sc_hd__buf_8
XFILLER_113_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4310_ _4310_/A hold47/X VGND VGND VPWR VPWR _4315_/S sky130_fd_sc_hd__and2_4
X_4241_ _4241_/A _4241_/B _6421_/B _4241_/D VGND VGND VPWR VPWR _4249_/S sky130_fd_sc_hd__or4_4
XFILLER_114_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4172_ _4172_/A _6406_/B VGND VGND VPWR VPWR _4177_/S sky130_fd_sc_hd__and2_4
XFILLER_83_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6813_ _7134_/CLK _6813_/D fanout429/X VGND VGND VPWR VPWR _6813_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_51_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6744_ _6744_/CLK _6744_/D fanout427/X VGND VGND VPWR VPWR _6744_/Q sky130_fd_sc_hd__dfrtp_2
X_3956_ _6474_/Q _6446_/A VGND VGND VPWR VPWR _3956_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6675_ _7127_/CLK _6675_/D fanout447/X VGND VGND VPWR VPWR _6675_/Q sky130_fd_sc_hd__dfrtp_2
X_3887_ _4349_/C _4349_/D _3887_/C input116/X VGND VGND VPWR VPWR _3895_/B sky130_fd_sc_hd__or4b_4
X_5626_ _5626_/A _6679_/Q VGND VGND VPWR VPWR _5654_/A sky130_fd_sc_hd__nor2_4
XFILLER_136_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5557_ _5557_/A0 hold14/X hold86/A VGND VGND VPWR VPWR hold15/A sky130_fd_sc_hd__mux2_1
X_5488_ _5596_/A0 hold365/X _5494_/S VGND VGND VPWR VPWR _7054_/D sky130_fd_sc_hd__mux2_1
X_4508_ _4711_/A _4581_/B VGND VGND VPWR VPWR _5033_/A sky130_fd_sc_hd__and2_2
XFILLER_105_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4439_ _4774_/A _4593_/A VGND VGND VPWR VPWR _4525_/A sky130_fd_sc_hd__or2_4
XFILLER_132_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7227_ _7227_/A VGND VGND VPWR VPWR _7227_/X sky130_fd_sc_hd__buf_2
XFILLER_160_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7158_ _7196_/CLK _7158_/D fanout433/X VGND VGND VPWR VPWR _7158_/Q sky130_fd_sc_hd__dfrtp_2
X_7089_ _7097_/CLK _7089_/D fanout437/X VGND VGND VPWR VPWR _7089_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_58_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6109_ _7190_/Q _6108_/X _6308_/S VGND VGND VPWR VPWR _6109_/X sky130_fd_sc_hd__mux2_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_471 hold209/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_460 _6764_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4790_ _4758_/B _4758_/C _4668_/B _4411_/Y VGND VGND VPWR VPWR _4796_/C sky130_fd_sc_hd__a31o_1
XFILLER_82_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3810_ _6467_/Q _3810_/B VGND VGND VPWR VPWR _3898_/B sky130_fd_sc_hd__nand2_2
XFILLER_20_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_29 _5341_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3741_ _6901_/Q _5315_/A _5585_/A _7141_/Q VGND VGND VPWR VPWR _3741_/X sky130_fd_sc_hd__a22o_1
XANTENNA_18 _5192_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6460_ _3938_/A1 _6460_/D _6415_/X VGND VGND VPWR VPWR hold64/A sky130_fd_sc_hd__dfrtp_2
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3672_ hold20/X _5234_/A VGND VGND VPWR VPWR _5242_/A sky130_fd_sc_hd__nor2_8
X_6391_ _6390_/X _7215_/Q _6400_/S VGND VGND VPWR VPWR _7215_/D sky130_fd_sc_hd__mux2_1
X_5411_ hold409/X _5600_/A0 _5413_/S VGND VGND VPWR VPWR _5411_/X sky130_fd_sc_hd__mux2_1
X_5342_ _5342_/A _5594_/B VGND VGND VPWR VPWR _5350_/S sky130_fd_sc_hd__nand2_8
XFILLER_133_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5273_ _5588_/A0 _5273_/A1 hold29/X VGND VGND VPWR VPWR _5273_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7012_ _7136_/CLK _7012_/D fanout436/X VGND VGND VPWR VPWR _7012_/Q sky130_fd_sc_hd__dfrtp_2
X_4224_ hold687/X _5561_/A0 _4234_/S VGND VGND VPWR VPWR _4224_/X sky130_fd_sc_hd__mux2_1
X_4155_ _4155_/A0 _5289_/A0 _4159_/S VGND VGND VPWR VPWR _4155_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4086_ _4086_/A0 hold71/X _4087_/S VGND VGND VPWR VPWR hold72/A sky130_fd_sc_hd__mux2_1
XFILLER_55_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4988_ _4988_/A _4997_/B VGND VGND VPWR VPWR _5081_/C sky130_fd_sc_hd__nor2_2
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3939_ _6506_/Q _3877_/C _6476_/Q VGND VGND VPWR VPWR _3939_/X sky130_fd_sc_hd__mux2_2
X_6727_ _6746_/CLK _6727_/D fanout427/X VGND VGND VPWR VPWR _6727_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6658_ _7225_/CLK _6658_/D fanout422/X VGND VGND VPWR VPWR _6658_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_137_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5609_ _5617_/A _5609_/B _5609_/C VGND VGND VPWR VPWR _7157_/D sky130_fd_sc_hd__and3_1
XFILLER_164_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6589_ _6649_/CLK _6589_/D fanout439/X VGND VGND VPWR VPWR _6589_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout374 hold207/X VGND VGND VPWR VPWR hold208/A sky130_fd_sc_hd__buf_8
XFILLER_143_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout363 hold47/X VGND VGND VPWR VPWR _5576_/B sky130_fd_sc_hd__buf_8
Xfanout352 _5665_/Y VGND VGND VPWR VPWR _6309_/S sky130_fd_sc_hd__buf_8
Xfanout385 hold135/X VGND VGND VPWR VPWR hold136/A sky130_fd_sc_hd__buf_8
Xfanout396 hold67/X VGND VGND VPWR VPWR _5578_/A0 sky130_fd_sc_hd__buf_8
XFILLER_47_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput16 mask_rev_in[20] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__buf_4
Xinput27 mask_rev_in[30] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__clkbuf_4
Xinput49 mgmt_gpio_in[21] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__buf_6
XFILLER_182_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput38 mgmt_gpio_in[11] VGND VGND VPWR VPWR _3202_/A sky130_fd_sc_hd__buf_6
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5960_ _6533_/Q _5722_/B _5953_/X _5959_/X _6308_/S VGND VGND VPWR VPWR _5960_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_37_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4911_ _4983_/B _4911_/B _4976_/A _4911_/D VGND VGND VPWR VPWR _4913_/C sky130_fd_sc_hd__or4_1
X_5891_ _6545_/Q _5674_/X _5707_/X _6758_/Q VGND VGND VPWR VPWR _5891_/X sky130_fd_sc_hd__a22o_1
XANTENNA_290 wb_dat_i[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4842_ _4554_/A _5087_/A _4554_/B _4507_/A VGND VGND VPWR VPWR _4842_/X sky130_fd_sc_hd__a22o_2
XFILLER_60_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4773_ _4773_/A _4773_/B VGND VGND VPWR VPWR _4776_/B sky130_fd_sc_hd__or2_4
X_6512_ _6987_/CLK _6512_/D fanout450/X VGND VGND VPWR VPWR _6512_/Q sky130_fd_sc_hd__dfrtp_2
X_3724_ _6714_/Q _4256_/A _4118_/A _6595_/Q _3723_/X VGND VGND VPWR VPWR _3725_/D
+ sky130_fd_sc_hd__a221o_4
XFILLER_174_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6443_ _6455_/A _6446_/B VGND VGND VPWR VPWR _6443_/X sky130_fd_sc_hd__and2_1
X_3655_ _6991_/Q _3299_/Y _4310_/A _6760_/Q VGND VGND VPWR VPWR _3655_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6374_ _6372_/A _6374_/A2 _6703_/Q VGND VGND VPWR VPWR _6374_/X sky130_fd_sc_hd__a21bo_1
X_3586_ _6976_/Q _5396_/A _5245_/A input64/X _3585_/X VGND VGND VPWR VPWR _3587_/D
+ sky130_fd_sc_hd__a221o_4
XFILLER_115_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5325_ _5595_/A0 _5325_/A1 _5332_/S VGND VGND VPWR VPWR _6909_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5256_ hold136/X _5256_/A1 _5260_/S VGND VGND VPWR VPWR _5256_/X sky130_fd_sc_hd__mux2_1
X_4207_ hold554/X _5597_/A0 _4217_/S VGND VGND VPWR VPWR _4207_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5187_ _5254_/A0 hold901/X _5190_/S VGND VGND VPWR VPWR _5187_/X sky130_fd_sc_hd__mux2_1
X_4138_ _5587_/A0 hold681/X _4141_/S VGND VGND VPWR VPWR _4138_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4069_ _5587_/A0 hold657/X _4072_/S VGND VGND VPWR VPWR _4069_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold608 _4180_/X VGND VGND VPWR VPWR _6645_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_10_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3440_ _7098_/Q _3341_/Y _5360_/A _6946_/Q _3439_/X VGND VGND VPWR VPWR _3452_/C
+ sky130_fd_sc_hd__a221o_1
Xhold619 _6501_/Q VGND VGND VPWR VPWR hold619/X sky130_fd_sc_hd__bufbuf_16
XFILLER_112_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3371_ _3668_/A _5252_/A VGND VGND VPWR VPWR _5558_/A sky130_fd_sc_hd__nor2_8
X_5110_ _5004_/A _4469_/Y _4659_/A _5099_/A _5046_/A VGND VGND VPWR VPWR _5156_/C
+ sky130_fd_sc_hd__a311o_1
X_6090_ _7023_/Q _6010_/Y _6031_/X _7087_/Q _6088_/X VGND VGND VPWR VPWR _6090_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _4469_/A _4470_/B _4565_/Y VGND VGND VPWR VPWR _5041_/X sky130_fd_sc_hd__a21o_1
XFILLER_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_8
XFILLER_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6992_ _7107_/CLK _6992_/D fanout434/X VGND VGND VPWR VPWR _6992_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_53_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5943_ _6566_/Q _5694_/X _5706_/X _6652_/Q VGND VGND VPWR VPWR _5959_/A sky130_fd_sc_hd__a22o_2
XFILLER_80_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5874_ _7183_/Q _6309_/S _5872_/X _5873_/X VGND VGND VPWR VPWR _7183_/D sky130_fd_sc_hd__o22a_1
X_4825_ _4898_/B _4728_/X _4746_/X _5164_/B _4824_/X VGND VGND VPWR VPWR _4825_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_193_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4756_ _5062_/A _4756_/B VGND VGND VPWR VPWR _5071_/B sky130_fd_sc_hd__nor2_1
X_4687_ _4687_/A _4832_/C VGND VGND VPWR VPWR _5095_/A sky130_fd_sc_hd__nor2_4
XFILLER_147_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3707_ _6950_/Q _5369_/A _5185_/A _6786_/Q _3706_/X VGND VGND VPWR VPWR _3709_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_107_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3638_ _7031_/Q _5459_/A _5513_/A _7079_/Q _3637_/X VGND VGND VPWR VPWR _3645_/A
+ sky130_fd_sc_hd__a221o_2
X_6426_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6426_/X sky130_fd_sc_hd__and2_1
XFILLER_115_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3569_ _6928_/Q _5342_/A _3567_/X _3568_/X VGND VGND VPWR VPWR _3588_/B sky130_fd_sc_hd__a211o_1
X_6357_ _6534_/Q _6060_/B _6356_/X _6308_/S VGND VGND VPWR VPWR _6357_/X sky130_fd_sc_hd__o211a_4
X_5308_ _5587_/A0 hold627/X _5314_/S VGND VGND VPWR VPWR _6894_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6288_ _6760_/Q _6010_/Y _6031_/X _6646_/Q _6287_/X VGND VGND VPWR VPWR _6288_/X
+ sky130_fd_sc_hd__a221o_2
X_5239_ _5597_/A0 hold725/X _5241_/S VGND VGND VPWR VPWR _5239_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold5 hold5/A VGND VGND VPWR VPWR hold5/X sky130_fd_sc_hd__bufbuf_16
XFILLER_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4610_ _4536_/B _4537_/X _4735_/B _4740_/A _4949_/B VGND VGND VPWR VPWR _4610_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_175_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5590_ _5599_/A0 hold839/X _5593_/S VGND VGND VPWR VPWR _5590_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4541_ _5023_/A _4871_/A _4997_/A VGND VGND VPWR VPWR _4542_/D sky130_fd_sc_hd__a21oi_1
XFILLER_7_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold405 _5339_/X VGND VGND VPWR VPWR _6922_/D sky130_fd_sc_hd__bufbuf_16
X_4472_ _4707_/B _4534_/B VGND VGND VPWR VPWR _4949_/A sky130_fd_sc_hd__nor2_8
XFILLER_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold427 _7140_/Q VGND VGND VPWR VPWR hold427/X sky130_fd_sc_hd__bufbuf_16
Xhold416 _5515_/X VGND VGND VPWR VPWR _7078_/D sky130_fd_sc_hd__bufbuf_16
Xhold438 _5570_/X VGND VGND VPWR VPWR _7127_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_171_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold449 _6914_/Q VGND VGND VPWR VPWR hold449/X sky130_fd_sc_hd__bufbuf_16
XFILLER_143_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7191_ _7196_/CLK _7191_/D fanout432/X VGND VGND VPWR VPWR _7191_/Q sky130_fd_sc_hd__dfrtp_4
X_3423_ _7188_/Q _6829_/Q _6831_/Q VGND VGND VPWR VPWR _3423_/X sky130_fd_sc_hd__mux2_8
X_6211_ _7084_/Q _6311_/B VGND VGND VPWR VPWR _6211_/X sky130_fd_sc_hd__and2_1
XFILLER_112_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6142_ _7073_/Q _6009_/X _6020_/D _6969_/Q VGND VGND VPWR VPWR _6142_/X sky130_fd_sc_hd__a22o_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3354_ _6900_/Q _5306_/A _5288_/A _6884_/Q VGND VGND VPWR VPWR _3354_/X sky130_fd_sc_hd__a22o_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1105 _4297_/X VGND VGND VPWR VPWR _6747_/D sky130_fd_sc_hd__bufbuf_16
X_6073_ _7126_/Q _6023_/A _6033_/X _7006_/Q _6072_/X VGND VGND VPWR VPWR _6083_/B
+ sky130_fd_sc_hd__a221o_1
X_3285_ hold19/X _3419_/A VGND VGND VPWR VPWR _3673_/B sky130_fd_sc_hd__or2_4
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1149 _5291_/X VGND VGND VPWR VPWR _6879_/D sky130_fd_sc_hd__bufbuf_16
Xhold1116 _6611_/Q VGND VGND VPWR VPWR _4139_/A1 sky130_fd_sc_hd__bufbuf_16
X_5024_ _5024_/A _5035_/B _5024_/C _5035_/D VGND VGND VPWR VPWR _5028_/B sky130_fd_sc_hd__or4_2
Xhold1138 _6589_/Q VGND VGND VPWR VPWR _4113_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1127 _6545_/Q VGND VGND VPWR VPWR _4062_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_85_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6975_ _6975_/CLK _6975_/D fanout443/X VGND VGND VPWR VPWR _6975_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5926_ _6787_/Q _5690_/X _5699_/X _6601_/Q _5925_/X VGND VGND VPWR VPWR _5927_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_110_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5857_ _7108_/Q _5675_/X _5706_/X _7060_/Q VGND VGND VPWR VPWR _5857_/X sky130_fd_sc_hd__a22o_1
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4808_ _4808_/A _5069_/B VGND VGND VPWR VPWR _5037_/A sky130_fd_sc_hd__or2_2
X_5788_ _7009_/Q _5678_/X _5684_/X _6993_/Q VGND VGND VPWR VPWR _5788_/X sky130_fd_sc_hd__a22o_1
X_4739_ _4714_/B _5147_/C _4738_/Y _4734_/X _4505_/X VGND VGND VPWR VPWR _4739_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_147_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6409_ _6409_/A0 hold995/X _6411_/S VGND VGND VPWR VPWR _7223_/D sky130_fd_sc_hd__mux2_1
Xhold961 _7125_/Q VGND VGND VPWR VPWR hold961/X sky130_fd_sc_hd__bufbuf_16
Xhold950 _6621_/Q VGND VGND VPWR VPWR hold950/X sky130_fd_sc_hd__bufbuf_16
XFILLER_89_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold972 _6657_/Q VGND VGND VPWR VPWR hold972/X sky130_fd_sc_hd__bufbuf_16
Xhold983 _4026_/X VGND VGND VPWR VPWR _6514_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_103_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold994 _4302_/X VGND VGND VPWR VPWR _6751_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_50_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7139_/CLK sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_65_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7081_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_82_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6760_ _7222_/CLK _6760_/D fanout420/X VGND VGND VPWR VPWR _6760_/Q sky130_fd_sc_hd__dfstp_4
X_5711_ _7005_/Q _5678_/X _5702_/X _6885_/Q VGND VGND VPWR VPWR _5711_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3972_ _6837_/Q _3972_/B VGND VGND VPWR VPWR _3972_/X sky130_fd_sc_hd__and2_2
XFILLER_188_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6691_ _6939_/CLK _6691_/D fanout453/X VGND VGND VPWR VPWR _6691_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5642_ _7168_/Q _5635_/B _5648_/B VGND VGND VPWR VPWR _5642_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_176_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5573_ _5600_/A0 hold388/X _5575_/S VGND VGND VPWR VPWR _5573_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold202 hold202/A VGND VGND VPWR VPWR hold202/X sky130_fd_sc_hd__bufbuf_16
XFILLER_116_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4524_ _4988_/A _4671_/A VGND VGND VPWR VPWR _4849_/A sky130_fd_sc_hd__nor2_2
Xclkbuf_leaf_18_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7150_/CLK sky130_fd_sc_hd__clkbuf_8
Xhold235 _7080_/Q VGND VGND VPWR VPWR hold235/X sky130_fd_sc_hd__bufbuf_16
Xhold213 _6689_/Q VGND VGND VPWR VPWR _3979_/S sky130_fd_sc_hd__bufbuf_16
Xhold224 _3256_/Y VGND VGND VPWR VPWR hold51/A sky130_fd_sc_hd__bufbuf_16
X_4455_ _4694_/A _4745_/A VGND VGND VPWR VPWR _4808_/A sky130_fd_sc_hd__nor2_2
Xhold268 _4039_/X VGND VGND VPWR VPWR _6526_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_144_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold257 _5277_/X VGND VGND VPWR VPWR _6867_/D sky130_fd_sc_hd__bufbuf_16
Xhold246 _6851_/Q VGND VGND VPWR VPWR hold246/X sky130_fd_sc_hd__bufbuf_16
Xhold279 _6985_/Q VGND VGND VPWR VPWR hold279/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4386_ _4996_/A _5164_/A VGND VGND VPWR VPWR _4386_/Y sky130_fd_sc_hd__nor2_1
X_3406_ _6907_/Q _5315_/A _3726_/A _3403_/X _3405_/X VGND VGND VPWR VPWR _3415_/C
+ sky130_fd_sc_hd__a2111o_1
X_7174_ _7196_/CLK _7174_/D fanout433/X VGND VGND VPWR VPWR _7174_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6125_ _6952_/Q _6022_/A _6025_/C _6928_/Q VGND VGND VPWR VPWR _6125_/X sky130_fd_sc_hd__a22o_1
XFILLER_100_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3337_ _6818_/Q _5207_/A _3336_/X VGND VGND VPWR VPWR _3378_/A sky130_fd_sc_hd__a21o_2
XFILLER_100_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _6933_/Q _6025_/A _6023_/C _6869_/Q _6055_/X VGND VGND VPWR VPWR _6057_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_85_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3268_ hold16/X hold80/X _3845_/A VGND VGND VPWR VPWR hold17/A sky130_fd_sc_hd__mux2_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5007_ _5007_/A1 _4746_/B _5050_/C _4745_/A _4648_/B VGND VGND VPWR VPWR _5008_/B
+ sky130_fd_sc_hd__o32a_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3199_ _6680_/Q VGND VGND VPWR VPWR _5659_/C sky130_fd_sc_hd__inv_2
XFILLER_39_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_119 _4659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_108 _3820_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6958_ _7054_/CLK _6958_/D fanout445/X VGND VGND VPWR VPWR _6958_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6889_ _7153_/CLK _6889_/D fanout444/X VGND VGND VPWR VPWR _6889_/Q sky130_fd_sc_hd__dfrtp_2
X_5909_ _6714_/Q _5676_/X _5702_/X _6551_/Q _5908_/X VGND VGND VPWR VPWR _5910_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_139_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold780 _6579_/Q VGND VGND VPWR VPWR hold780/X sky130_fd_sc_hd__bufbuf_16
Xhold791 _4327_/X VGND VGND VPWR VPWR _6772_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_131_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput307 _3920_/B VGND VGND VPWR VPWR serial_clock sky130_fd_sc_hd__buf_8
XFILLER_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput329 _6582_/Q VGND VGND VPWR VPWR wb_dat_o[1] sky130_fd_sc_hd__buf_8
Xoutput318 _6581_/Q VGND VGND VPWR VPWR wb_dat_o[0] sky130_fd_sc_hd__buf_8
XFILLER_153_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4240_ _6360_/A _3991_/S _6704_/Q _4237_/X _4239_/X VGND VGND VPWR VPWR _6689_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4171_ _6411_/A0 hold754/X _4171_/S VGND VGND VPWR VPWR _4171_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6812_ _7134_/CLK _6812_/D fanout429/X VGND VGND VPWR VPWR _6812_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_168_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6743_ _6745_/CLK _6743_/D fanout442/X VGND VGND VPWR VPWR _6743_/Q sky130_fd_sc_hd__dfrtp_2
X_3955_ input84/X _3877_/C _6474_/Q VGND VGND VPWR VPWR _3955_/X sky130_fd_sc_hd__mux2_8
X_6674_ _7127_/CLK _6674_/D fanout446/X VGND VGND VPWR VPWR _6674_/Q sky130_fd_sc_hd__dfrtp_2
X_3886_ _4351_/A _4351_/B _3886_/C VGND VGND VPWR VPWR _3895_/A sky130_fd_sc_hd__or3_4
X_5625_ _7162_/Q _7161_/Q VGND VGND VPWR VPWR _5705_/B sky130_fd_sc_hd__and2_4
XFILLER_137_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5556_ hold645/X _5601_/A0 hold86/X VGND VGND VPWR VPWR _5556_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5487_ _5595_/A0 hold924/X _5494_/S VGND VGND VPWR VPWR _7053_/D sky130_fd_sc_hd__mux2_1
XFILLER_151_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4507_ _4507_/A _4711_/A _4659_/A VGND VGND VPWR VPWR _4920_/A sky130_fd_sc_hd__and3_4
X_4438_ _4722_/A _4438_/B VGND VGND VPWR VPWR _4593_/A sky130_fd_sc_hd__xor2_4
XFILLER_160_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4369_ _4529_/A _4650_/B VGND VGND VPWR VPWR _4484_/C sky130_fd_sc_hd__nand2_4
X_7157_ _7196_/CLK _7157_/D fanout433/X VGND VGND VPWR VPWR _7157_/Q sky130_fd_sc_hd__dfrtp_2
X_6108_ _6090_/X _6096_/X _6107_/X _6060_/B _6855_/Q VGND VGND VPWR VPWR _6108_/X
+ sky130_fd_sc_hd__o32a_4
X_7088_ _7088_/CLK _7088_/D fanout438/X VGND VGND VPWR VPWR _7088_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6039_ _6877_/Q _6021_/C _6022_/C _6957_/Q VGND VGND VPWR VPWR _6039_/X sky130_fd_sc_hd__a22o_1
XFILLER_74_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_450 _4287_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_461 _6485_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_472 _5260_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3740_ _6933_/Q _5351_/A _5279_/A _6869_/Q VGND VGND VPWR VPWR _3740_/X sky130_fd_sc_hd__a22o_1
XANTENNA_19 _6799_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3671_ _6739_/Q _4286_/A _5194_/A _6801_/Q VGND VGND VPWR VPWR _3671_/X sky130_fd_sc_hd__a22o_4
X_6390_ _6707_/Q _6390_/A2 _6390_/B1 _6706_/Q _6389_/X VGND VGND VPWR VPWR _6390_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_185_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5410_ hold279/X _5581_/A0 _5413_/S VGND VGND VPWR VPWR _5410_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5341_ hold337/X _5602_/A0 _5341_/S VGND VGND VPWR VPWR _5341_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5272_ _5587_/A0 hold392/X hold29/X VGND VGND VPWR VPWR _6862_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7011_ _7104_/CLK _7011_/D fanout434/X VGND VGND VPWR VPWR _7011_/Q sky130_fd_sc_hd__dfrtp_2
X_4223_ _4223_/A0 _4222_/X _4235_/S VGND VGND VPWR VPWR _4223_/X sky130_fd_sc_hd__mux2_1
X_4154_ _4154_/A _5558_/B VGND VGND VPWR VPWR _4159_/S sky130_fd_sc_hd__and2_4
XFILLER_56_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4085_ hold986/X _5300_/A0 _4087_/S VGND VGND VPWR VPWR _4085_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4987_ _4987_/A _4987_/B _4992_/B VGND VGND VPWR VPWR _4987_/X sky130_fd_sc_hd__or3_4
X_6726_ _6747_/CLK _6726_/D fanout427/X VGND VGND VPWR VPWR _6726_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_177_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3938_ _6507_/Q _3938_/A1 _6475_/Q VGND VGND VPWR VPWR _3938_/X sky130_fd_sc_hd__mux2_1
X_3869_ hold73/A _6465_/Q _3874_/S VGND VGND VPWR VPWR _6465_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6657_ _7225_/CLK _6657_/D fanout422/X VGND VGND VPWR VPWR _6657_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_176_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5608_ _7157_/Q _5615_/D VGND VGND VPWR VPWR _5609_/C sky130_fd_sc_hd__or2_1
X_6588_ _7201_/CLK _6588_/D VGND VGND VPWR VPWR _6588_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_191_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5539_ _5584_/A0 hold418/X _5539_/S VGND VGND VPWR VPWR _5539_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7209_ _7209_/CLK _7209_/D VGND VGND VPWR VPWR _7209_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_143_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout375 hold7/X VGND VGND VPWR VPWR _5582_/A0 sky130_fd_sc_hd__buf_8
Xfanout364 _5486_/B VGND VGND VPWR VPWR hold47/A sky130_fd_sc_hd__buf_8
Xfanout353 _5664_/X VGND VGND VPWR VPWR _6358_/B1 sky130_fd_sc_hd__buf_8
Xfanout386 hold71/X VGND VGND VPWR VPWR _5571_/A0 sky130_fd_sc_hd__buf_8
Xfanout397 hold67/X VGND VGND VPWR VPWR _5587_/A0 sky130_fd_sc_hd__buf_8
XFILLER_143_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput17 mask_rev_in[21] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__clkbuf_4
Xinput28 mask_rev_in[31] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__clkbuf_4
XFILLER_155_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput39 mgmt_gpio_in[12] VGND VGND VPWR VPWR _3973_/B sky130_fd_sc_hd__buf_8
XFILLER_182_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4910_ _5128_/A _5075_/B _4910_/C VGND VGND VPWR VPWR _4911_/D sky130_fd_sc_hd__or3_1
X_5890_ _6619_/Q _5673_/X _5693_/X _6654_/Q _5889_/X VGND VGND VPWR VPWR _5893_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_92_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4841_ _4412_/Y _5123_/C VGND VGND VPWR VPWR _5116_/B sky130_fd_sc_hd__nand2b_1
XFILLER_45_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_291 _4349_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_280 wb_dat_i[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4772_ _4772_/A _5165_/A _4772_/C VGND VGND VPWR VPWR _4936_/B sky130_fd_sc_hd__and3_1
X_6511_ _7141_/CLK _6511_/D fanout447/X VGND VGND VPWR VPWR _6511_/Q sky130_fd_sc_hd__dfrtp_2
X_3723_ _6577_/Q _4097_/A _5242_/A _6838_/Q VGND VGND VPWR VPWR _3723_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6442_ _6446_/A _6446_/B VGND VGND VPWR VPWR _6442_/X sky130_fd_sc_hd__and2_1
X_3654_ _3654_/A _3654_/B _3654_/C _3654_/D VGND VGND VPWR VPWR _3664_/A sky130_fd_sc_hd__or4_1
XFILLER_174_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6373_ _6706_/Q _6371_/Y _6372_/Y _6705_/Q VGND VGND VPWR VPWR _6376_/C sky130_fd_sc_hd__a22o_1
XFILLER_173_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3585_ _6553_/Q _4067_/A _4136_/A _6612_/Q VGND VGND VPWR VPWR _3585_/X sky130_fd_sc_hd__a22o_4
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A VGND VGND VPWR VPWR _7201_/CLK sky130_fd_sc_hd__clkbuf_8
X_5324_ _5324_/A _5594_/B VGND VGND VPWR VPWR _5332_/S sky130_fd_sc_hd__nand2_8
XFILLER_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5255_ _5561_/A0 hold687/X _5260_/S VGND VGND VPWR VPWR _5255_/X sky130_fd_sc_hd__mux2_1
X_4206_ hold727/X _4205_/X _4218_/S VGND VGND VPWR VPWR _4206_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5186_ _5234_/C _5186_/A1 _5190_/S VGND VGND VPWR VPWR _5186_/X sky130_fd_sc_hd__mux2_1
X_4137_ _5289_/A0 _4137_/A1 _4141_/S VGND VGND VPWR VPWR _4137_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4068_ _5289_/A0 _4068_/A1 _4072_/S VGND VGND VPWR VPWR _4068_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6709_ _6717_/CLK _6709_/D fanout426/X VGND VGND VPWR VPWR _6709_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_138_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold609 _6724_/Q VGND VGND VPWR VPWR hold609/X sky130_fd_sc_hd__bufbuf_16
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3370_ input19/X _3368_/Y _5396_/A _6980_/Q _3366_/X VGND VGND VPWR VPWR _3377_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _4565_/Y _4689_/Y _4817_/C _5039_/X VGND VGND VPWR VPWR _5048_/A sky130_fd_sc_hd__a211o_1
XFILLER_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6991_ _7135_/CLK _6991_/D fanout431/X VGND VGND VPWR VPWR _6991_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5942_ _6627_/Q _5963_/B VGND VGND VPWR VPWR _5942_/X sky130_fd_sc_hd__or2_1
X_5873_ _5663_/A _7182_/Q _6358_/B1 VGND VGND VPWR VPWR _5873_/X sky130_fd_sc_hd__a21o_1
X_4824_ _5164_/B _4756_/B _4746_/X _4898_/B VGND VGND VPWR VPWR _4824_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4755_ _4898_/B _4757_/B VGND VGND VPWR VPWR _4893_/B sky130_fd_sc_hd__or2_4
XFILLER_147_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3706_ _6870_/Q _5279_/A _4124_/A _6600_/Q VGND VGND VPWR VPWR _3706_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4686_ _4724_/B _4832_/C VGND VGND VPWR VPWR _5022_/B sky130_fd_sc_hd__nor2_1
XFILLER_119_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3637_ _7071_/Q hold92/A _4178_/A _6646_/Q VGND VGND VPWR VPWR _3637_/X sky130_fd_sc_hd__a22o_1
X_6425_ _6455_/A _6446_/B VGND VGND VPWR VPWR _6425_/X sky130_fd_sc_hd__and2_1
XFILLER_115_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3568_ _6602_/Q _4124_/A _4112_/A _6592_/Q _3555_/X VGND VGND VPWR VPWR _3568_/X
+ sky130_fd_sc_hd__a221o_4
X_6356_ _6356_/A _6356_/B _6356_/C _6356_/D VGND VGND VPWR VPWR _6356_/X sky130_fd_sc_hd__or4_2
X_5307_ _5595_/A0 hold965/X _5314_/S VGND VGND VPWR VPWR _6893_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6287_ _6735_/Q _6020_/B _6011_/X _6787_/Q VGND VGND VPWR VPWR _6287_/X sky130_fd_sc_hd__a22o_1
X_3499_ input7/X _3320_/Y _5200_/A _6809_/Q _3498_/X VGND VGND VPWR VPWR _3504_/C
+ sky130_fd_sc_hd__a221o_2
X_5238_ _5238_/A _5594_/B VGND VGND VPWR VPWR _5241_/S sky130_fd_sc_hd__nand2_2
XFILLER_29_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5169_ _5169_/A _5169_/B _5169_/C VGND VGND VPWR VPWR _6783_/D sky130_fd_sc_hd__or3_2
XFILLER_56_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__1132_ clkbuf_0__1132_/X VGND VGND VPWR VPWR _6367_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_193_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold6 hold6/A VGND VGND VPWR VPWR hold6/X sky130_fd_sc_hd__bufbuf_16
XFILLER_47_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4540_ _5140_/A _5140_/B _4520_/X VGND VGND VPWR VPWR _4542_/C sky130_fd_sc_hd__or3b_1
XFILLER_129_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4471_ _4818_/B _4663_/B VGND VGND VPWR VPWR _4697_/A sky130_fd_sc_hd__or2_4
XFILLER_183_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold406 _7036_/Q VGND VGND VPWR VPWR hold406/X sky130_fd_sc_hd__bufbuf_16
Xhold417 _6818_/Q VGND VGND VPWR VPWR hold417/X sky130_fd_sc_hd__bufbuf_16
XFILLER_144_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold439 _7132_/Q VGND VGND VPWR VPWR hold439/X sky130_fd_sc_hd__bufbuf_16
X_3422_ _5234_/A _3543_/B VGND VGND VPWR VPWR _5200_/A sky130_fd_sc_hd__nor2_8
X_7190_ _7197_/CLK _7190_/D fanout429/X VGND VGND VPWR VPWR _7190_/Q sky130_fd_sc_hd__dfrtp_1
Xhold428 _5584_/X VGND VGND VPWR VPWR _7140_/D sky130_fd_sc_hd__bufbuf_16
X_6210_ _7195_/Q _5665_/Y _6209_/X VGND VGND VPWR VPWR _7195_/D sky130_fd_sc_hd__o21a_1
X_6141_ _7121_/Q _6023_/D _6030_/Y _7033_/Q _6140_/X VGND VGND VPWR VPWR _6144_/C
+ sky130_fd_sc_hd__a221o_4
XFILLER_124_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ hold91/X _3473_/A VGND VGND VPWR VPWR _5288_/A sky130_fd_sc_hd__nor2_8
X_6072_ _6886_/Q _6020_/A _6021_/D _7142_/Q _6062_/X VGND VGND VPWR VPWR _6072_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_112_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_727 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1106 _7069_/Q VGND VGND VPWR VPWR _5505_/A1 sky130_fd_sc_hd__bufbuf_16
X_3284_ _3421_/A hold89/X VGND VGND VPWR VPWR _3284_/X sky130_fd_sc_hd__or2_4
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1117 _6626_/Q VGND VGND VPWR VPWR _4157_/A0 sky130_fd_sc_hd__bufbuf_16
X_5023_ _5023_/A _5023_/B VGND VGND VPWR VPWR _5035_/D sky130_fd_sc_hd__nor2_1
Xhold1139 _4113_/X VGND VGND VPWR VPWR _6589_/D sky130_fd_sc_hd__bufbuf_16
Xhold1128 _4062_/X VGND VGND VPWR VPWR _6545_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_85_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6974_ _7111_/CLK _6974_/D fanout444/X VGND VGND VPWR VPWR _6974_/Q sky130_fd_sc_hd__dfstp_4
X_5925_ _6537_/Q _5700_/X _5701_/X _6616_/Q VGND VGND VPWR VPWR _5925_/X sky130_fd_sc_hd__a22o_1
XFILLER_81_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5856_ _7100_/Q _5690_/X _5704_/X _6940_/Q _5855_/X VGND VGND VPWR VPWR _5861_/B
+ sky130_fd_sc_hd__a221o_1
X_4807_ _4980_/B _4980_/C _5132_/A _4806_/X _4917_/B VGND VGND VPWR VPWR _4807_/X
+ sky130_fd_sc_hd__o41a_4
XFILLER_139_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5787_ _7179_/Q _6309_/S _5785_/X _5786_/X VGND VGND VPWR VPWR _7179_/D sky130_fd_sc_hd__o22a_1
X_4738_ _4758_/A _4758_/C _4737_/Y VGND VGND VPWR VPWR _4738_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_119_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4669_ _4697_/A _5164_/B _4724_/B _4886_/B VGND VGND VPWR VPWR _4669_/X sky130_fd_sc_hd__a31o_1
XFILLER_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6408_ _6408_/A0 hold517/X _6411_/S VGND VGND VPWR VPWR _6408_/X sky130_fd_sc_hd__mux2_1
Xhold940 _6660_/Q VGND VGND VPWR VPWR hold940/X sky130_fd_sc_hd__bufbuf_16
Xhold962 _6925_/Q VGND VGND VPWR VPWR hold962/X sky130_fd_sc_hd__bufbuf_16
Xhold951 _4151_/X VGND VGND VPWR VPWR _6621_/D sky130_fd_sc_hd__bufbuf_16
Xhold973 _4194_/X VGND VGND VPWR VPWR _6657_/D sky130_fd_sc_hd__bufbuf_16
Xhold984 _7117_/Q VGND VGND VPWR VPWR hold984/X sky130_fd_sc_hd__bufbuf_16
Xhold995 _7223_/Q VGND VGND VPWR VPWR hold995/X sky130_fd_sc_hd__bufbuf_16
X_6339_ _6757_/Q _6023_/D _6030_/Y _6772_/Q VGND VGND VPWR VPWR _6339_/X sky130_fd_sc_hd__a22o_1
XFILLER_135_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3971_ _3971_/A input1/X VGND VGND VPWR VPWR _3971_/X sky130_fd_sc_hd__and2_2
X_5710_ _6957_/Q _5673_/X _5695_/X VGND VGND VPWR VPWR _5710_/X sky130_fd_sc_hd__a21o_1
XFILLER_62_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6690_ _6939_/CLK _6690_/D fanout453/X VGND VGND VPWR VPWR _6690_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5641_ _5663_/B _6012_/A _6032_/A _5621_/X _7167_/Q VGND VGND VPWR VPWR _7167_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_191_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5572_ hold185/X hold218/X _5575_/S VGND VGND VPWR VPWR _5572_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4523_ _4671_/A _4990_/A VGND VGND VPWR VPWR _5114_/A sky130_fd_sc_hd__nor2_4
Xclkbuf_1_0_1_csclk clkbuf_1_0_1_csclk/A VGND VGND VPWR VPWR clkbuf_2_1_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_116_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold203 _4153_/X VGND VGND VPWR VPWR _6623_/D sky130_fd_sc_hd__bufbuf_16
Xhold214 _3991_/S VGND VGND VPWR VPWR _3975_/B sky130_fd_sc_hd__bufbuf_16
Xhold225 _3277_/Y VGND VGND VPWR VPWR _3278_/B sky130_fd_sc_hd__bufbuf_16
X_4454_ _4584_/A _4663_/B VGND VGND VPWR VPWR _4745_/A sky130_fd_sc_hd__or2_4
Xhold236 _5517_/X VGND VGND VPWR VPWR _7080_/D sky130_fd_sc_hd__bufbuf_16
Xhold269 _7097_/Q VGND VGND VPWR VPWR hold269/X sky130_fd_sc_hd__bufbuf_16
Xhold247 _5259_/X VGND VGND VPWR VPWR _6851_/D sky130_fd_sc_hd__bufbuf_16
Xhold258 _7008_/Q VGND VGND VPWR VPWR hold258/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4385_ _5023_/A _4871_/A VGND VGND VPWR VPWR _5164_/A sky130_fd_sc_hd__and2_4
X_7173_ _7196_/CLK _7173_/D fanout433/X VGND VGND VPWR VPWR _7173_/Q sky130_fd_sc_hd__dfrtp_2
X_3405_ _7011_/Q _5432_/A _3344_/Y _6502_/Q _3404_/X VGND VGND VPWR VPWR _3405_/X
+ sky130_fd_sc_hd__a221o_1
X_6124_ _7128_/Q _6023_/A _6033_/X _7008_/Q _6123_/X VGND VGND VPWR VPWR _6132_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3336_ _7044_/Q _3334_/Y _3978_/A _6495_/Q VGND VGND VPWR VPWR _3336_/X sky130_fd_sc_hd__a22o_1
X_6055_ _6909_/Q _6020_/C _6030_/Y _7029_/Q VGND VGND VPWR VPWR _6055_/X sky130_fd_sc_hd__a22o_1
XFILLER_100_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _4832_/A _4728_/X _5050_/C VGND VGND VPWR VPWR _5008_/A sky130_fd_sc_hd__a21o_1
XFILLER_100_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3267_ hold26/X hold89/X VGND VGND VPWR VPWR hold90/A sky130_fd_sc_hd__nand2_2
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3198_ _6677_/Q VGND VGND VPWR VPWR _5626_/A sky130_fd_sc_hd__inv_2
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_109 _3820_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6957_ _7122_/CLK _6957_/D fanout443/X VGND VGND VPWR VPWR _6957_/Q sky130_fd_sc_hd__dfstp_2
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6888_ _6987_/CLK _6888_/D fanout450/X VGND VGND VPWR VPWR _6888_/Q sky130_fd_sc_hd__dfrtp_2
X_5908_ _6660_/Q _5669_/X _5698_/B _5899_/X VGND VGND VPWR VPWR _5908_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5839_ _5839_/A _5839_/B _5839_/C _5839_/D VGND VGND VPWR VPWR _5839_/X sky130_fd_sc_hd__or4_2
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold770 _6510_/Q VGND VGND VPWR VPWR hold770/X sky130_fd_sc_hd__bufbuf_16
Xhold781 _4101_/X VGND VGND VPWR VPWR _6579_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_1_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold792 _6533_/Q VGND VGND VPWR VPWR hold792/X sky130_fd_sc_hd__bufbuf_16
XFILLER_162_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput308 _3423_/X VGND VGND VPWR VPWR serial_data_1 sky130_fd_sc_hd__buf_8
XFILLER_113_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput319 _6570_/Q VGND VGND VPWR VPWR wb_dat_o[10] sky130_fd_sc_hd__buf_8
XFILLER_5_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4170_ _6410_/A0 hold966/X _4171_/S VGND VGND VPWR VPWR _4170_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6811_ _6825_/CLK _6811_/D fanout421/X VGND VGND VPWR VPWR _6811_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_51_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6742_ _6759_/CLK _6742_/D fanout419/X VGND VGND VPWR VPWR _6742_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3954_ _3991_/S _3954_/A2 _6455_/B _3953_/Y VGND VGND VPWR VPWR _3954_/X sky130_fd_sc_hd__a22o_2
XFILLER_51_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6673_ _7127_/CLK _6673_/D fanout446/X VGND VGND VPWR VPWR _6673_/Q sky130_fd_sc_hd__dfrtp_2
X_3885_ _4351_/C _4351_/D _4350_/A _4350_/B VGND VGND VPWR VPWR _3886_/C sky130_fd_sc_hd__or4_1
XFILLER_176_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5624_ _6679_/Q _5702_/B VGND VGND VPWR VPWR _5629_/B sky130_fd_sc_hd__nand2_1
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5555_ _5555_/A0 hold78/X hold86/X VGND VGND VPWR VPWR hold87/A sky130_fd_sc_hd__mux2_1
XFILLER_129_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4506_ _4986_/A _4749_/C _4687_/A _4812_/A VGND VGND VPWR VPWR _4506_/X sky130_fd_sc_hd__a31o_1
X_5486_ _5486_/A _5486_/B VGND VGND VPWR VPWR _5494_/S sky130_fd_sc_hd__nand2_8
X_4437_ _4529_/B _4529_/C VGND VGND VPWR VPWR _4438_/B sky130_fd_sc_hd__nand2_4
XFILLER_104_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7225_ _7225_/CLK _7225_/D fanout422/X VGND VGND VPWR VPWR _7225_/Q sky130_fd_sc_hd__dfrtp_2
X_7156_ _7156_/CLK _7156_/D fanout447/X VGND VGND VPWR VPWR _7156_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_132_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4368_ _4368_/A _4722_/A VGND VGND VPWR VPWR _4650_/B sky130_fd_sc_hd__or2_4
X_6107_ _6306_/A _6107_/B _6107_/C VGND VGND VPWR VPWR _6107_/X sky130_fd_sc_hd__or3_4
XFILLER_113_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3319_ hold90/X hold83/X VGND VGND VPWR VPWR _3375_/B sky130_fd_sc_hd__or2_4
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4299_ _5234_/C _4299_/A1 _4303_/S VGND VGND VPWR VPWR _4299_/X sky130_fd_sc_hd__mux2_1
X_7087_ _7135_/CLK hold56/X fanout428/X VGND VGND VPWR VPWR _7087_/Q sky130_fd_sc_hd__dfrtp_2
X_6038_ _7093_/Q _6011_/X _6031_/X _7085_/Q VGND VGND VPWR VPWR _6038_/X sky130_fd_sc_hd__a22o_1
XFILLER_100_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_64_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7118_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_41_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_440 hold273/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_17_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7121_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_451 _6501_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_462 _6487_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_473 hold431/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3670_ _6862_/Q hold28/A _5387_/A _6966_/Q VGND VGND VPWR VPWR _3670_/X sky130_fd_sc_hd__a22o_1
XFILLER_9_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5340_ hold589/X _5601_/A0 _5341_/S VGND VGND VPWR VPWR _5340_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5271_ _5595_/A0 hold985/X hold29/X VGND VGND VPWR VPWR _6861_/D sky130_fd_sc_hd__mux2_1
XFILLER_181_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7010_ _7088_/CLK _7010_/D fanout438/X VGND VGND VPWR VPWR _7010_/Q sky130_fd_sc_hd__dfrtp_2
X_4222_ hold912/X _5254_/A0 _4234_/S VGND VGND VPWR VPWR _4222_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4153_ _4153_/A0 _5581_/A0 _4153_/S VGND VGND VPWR VPWR _4153_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4084_ hold344/X _5587_/A0 _4087_/S VGND VGND VPWR VPWR _4084_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4986_ _4986_/A _4986_/B _4986_/C VGND VGND VPWR VPWR _4997_/B sky130_fd_sc_hd__and3_4
X_6725_ _6725_/CLK _6725_/D fanout440/X VGND VGND VPWR VPWR _6725_/Q sky130_fd_sc_hd__dfstp_4
X_3937_ _6508_/Q _3875_/B _6476_/Q VGND VGND VPWR VPWR _3937_/X sky130_fd_sc_hd__mux2_2
XFILLER_51_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3868_ _6465_/Q hold9/A _3874_/S VGND VGND VPWR VPWR _6466_/D sky130_fd_sc_hd__mux2_1
X_6656_ _7225_/CLK _6656_/D fanout422/X VGND VGND VPWR VPWR _6656_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_191_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6587_ _7220_/CLK _6587_/D VGND VGND VPWR VPWR _6587_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_11_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5607_ _7157_/Q _5615_/D VGND VGND VPWR VPWR _5609_/B sky130_fd_sc_hd__nand2_1
X_3799_ _6486_/Q _3801_/B VGND VGND VPWR VPWR _3802_/A sky130_fd_sc_hd__nand2_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5538_ _5583_/A0 hold708/X _5539_/S VGND VGND VPWR VPWR _5538_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7208_ _7208_/CLK _7208_/D VGND VGND VPWR VPWR _7208_/Q sky130_fd_sc_hd__dfxtp_4
X_5469_ _5541_/A0 _5469_/A1 _5476_/S VGND VGND VPWR VPWR _7037_/D sky130_fd_sc_hd__mux2_1
XFILLER_78_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout365 _5486_/B VGND VGND VPWR VPWR _5558_/B sky130_fd_sc_hd__buf_8
X_7139_ _7139_/CLK _7139_/D fanout435/X VGND VGND VPWR VPWR _7139_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout376 hold78/X VGND VGND VPWR VPWR _5600_/A0 sky130_fd_sc_hd__buf_8
Xfanout398 hold67/X VGND VGND VPWR VPWR _5596_/A0 sky130_fd_sc_hd__buf_8
Xfanout387 hold135/X VGND VGND VPWR VPWR hold71/A sky130_fd_sc_hd__buf_8
XFILLER_101_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput18 mask_rev_in[22] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__clkbuf_4
Xinput29 mask_rev_in[3] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__clkbuf_4
XFILLER_155_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_270 wb_adr_i[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4840_ _4840_/A _4957_/A VGND VGND VPWR VPWR _5046_/A sky130_fd_sc_hd__or2_2
XANTENNA_281 wb_dat_i[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_292 input97/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4771_ _4986_/B _5031_/B VGND VGND VPWR VPWR _4806_/B sky130_fd_sc_hd__nor2_1
X_6510_ _6976_/CLK _6510_/D fanout450/X VGND VGND VPWR VPWR _6510_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3722_ _7030_/Q _5459_/A _5423_/A _6998_/Q _3721_/X VGND VGND VPWR VPWR _3725_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6441_ _6446_/A _6446_/B VGND VGND VPWR VPWR _6441_/X sky130_fd_sc_hd__and2_1
X_3653_ _7087_/Q hold54/A _3978_/A _6490_/Q _3652_/X VGND VGND VPWR VPWR _3654_/D
+ sky130_fd_sc_hd__a221o_1
X_6372_ _6372_/A _6372_/B VGND VGND VPWR VPWR _6372_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5323_ _5602_/A0 hold529/X _5323_/S VGND VGND VPWR VPWR _5323_/X sky130_fd_sc_hd__mux2_1
X_3584_ input55/X _4025_/A _4154_/A _6627_/Q _3583_/X VGND VGND VPWR VPWR _3587_/C
+ sky130_fd_sc_hd__a221o_4
XFILLER_127_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5254_ _5254_/A0 hold912/X _5260_/S VGND VGND VPWR VPWR _5254_/X sky130_fd_sc_hd__mux2_1
X_4205_ hold317/X _5596_/A0 _4217_/S VGND VGND VPWR VPWR _4205_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5185_ _5185_/A _6406_/B VGND VGND VPWR VPWR _5190_/S sky130_fd_sc_hd__nand2_4
X_4136_ _4136_/A _5558_/B VGND VGND VPWR VPWR _4141_/S sky130_fd_sc_hd__nand2_4
Xclkbuf_3_6_0_csclk clkbuf_3_7_0_csclk/A VGND VGND VPWR VPWR _7137_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_3_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4067_ _4067_/A _5558_/B VGND VGND VPWR VPWR _4072_/S sky130_fd_sc_hd__nand2_4
XFILLER_37_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4969_ _4949_/B _4571_/Y _4959_/A _4905_/B VGND VGND VPWR VPWR _4973_/C sky130_fd_sc_hd__a31o_2
XFILLER_51_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6708_ _6717_/CLK _6708_/D fanout426/X VGND VGND VPWR VPWR _6708_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6639_ _6786_/CLK _6639_/D fanout417/X VGND VGND VPWR VPWR _6639_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6990_ _7136_/CLK _6990_/D fanout436/X VGND VGND VPWR VPWR _6990_/Q sky130_fd_sc_hd__dfstp_2
X_5941_ _6592_/Q _5680_/X _5700_/X _6538_/Q VGND VGND VPWR VPWR _5941_/X sky130_fd_sc_hd__a22o_1
X_5872_ _6860_/Q _5722_/B _5861_/X _5871_/X _6308_/S VGND VGND VPWR VPWR _5872_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4823_ _5164_/B _5017_/A _4756_/B _4898_/B VGND VGND VPWR VPWR _4823_/X sky130_fd_sc_hd__o22a_1
X_4754_ _4898_/B _4754_/B VGND VGND VPWR VPWR _4950_/B sky130_fd_sc_hd__nor2_4
XFILLER_146_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3705_ _6894_/Q _5306_/A _4136_/A _6610_/Q _3704_/X VGND VGND VPWR VPWR _3709_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4685_ _4685_/A _4746_/B VGND VGND VPWR VPWR _5017_/A sky130_fd_sc_hd__or2_4
XFILLER_146_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3636_ _3636_/A _3636_/B _3636_/C _3636_/D VGND VGND VPWR VPWR _3665_/A sky130_fd_sc_hd__or4_4
X_6424_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6424_/X sky130_fd_sc_hd__and2_1
XFILLER_127_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3567_ _6912_/Q _5324_/A _5387_/A _6968_/Q _3554_/X VGND VGND VPWR VPWR _3567_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_115_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6355_ _6355_/A _6355_/B _6355_/C _6355_/D VGND VGND VPWR VPWR _6356_/D sky130_fd_sc_hd__or4_2
X_5306_ _5306_/A _5558_/B VGND VGND VPWR VPWR _5314_/S sky130_fd_sc_hd__nand2_8
X_6286_ _6616_/Q _6022_/A _6025_/C _6601_/Q VGND VGND VPWR VPWR _6286_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5237_ _5289_/A0 _5237_/A1 _5237_/S VGND VGND VPWR VPWR _5237_/X sky130_fd_sc_hd__mux2_1
X_3498_ _6993_/Q _3299_/Y _6406_/A _7225_/Q VGND VGND VPWR VPWR _3498_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5168_ _6783_/Q _6376_/A _5155_/X _5158_/Y _5167_/X VGND VGND VPWR VPWR _5169_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5099_ _5099_/A _5099_/B _5099_/C VGND VGND VPWR VPWR _5101_/C sky130_fd_sc_hd__or3_1
XFILLER_84_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4119_ _4119_/A0 _6407_/A0 _4123_/S VGND VGND VPWR VPWR _4119_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold7 hold7/A VGND VGND VPWR VPWR hold7/X sky130_fd_sc_hd__bufbuf_16
XFILLER_121_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4470_ _4740_/A _4470_/B VGND VGND VPWR VPWR _5005_/A sky130_fd_sc_hd__nand2_1
XFILLER_156_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold407 _5467_/X VGND VGND VPWR VPWR _7036_/D sky130_fd_sc_hd__bufbuf_16
Xhold418 _7100_/Q VGND VGND VPWR VPWR hold418/X sky130_fd_sc_hd__bufbuf_16
XFILLER_143_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3421_ _3421_/A _3421_/B _3421_/C VGND VGND VPWR VPWR _3543_/B sky130_fd_sc_hd__or3_4
Xhold429 _6852_/Q VGND VGND VPWR VPWR hold429/X sky130_fd_sc_hd__bufbuf_16
XFILLER_171_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6140_ _7001_/Q _5987_/Y _6022_/D _6921_/Q VGND VGND VPWR VPWR _6140_/X sky130_fd_sc_hd__a22o_1
XFILLER_98_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3352_ _3673_/B _3543_/A VGND VGND VPWR VPWR _5306_/A sky130_fd_sc_hd__nor2_8
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xload_slew354 _3457_/A VGND VGND VPWR VPWR _3540_/A sky130_fd_sc_hd__buf_8
XFILLER_58_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3283_ _5225_/A _3534_/A VGND VGND VPWR VPWR _3283_/Y sky130_fd_sc_hd__nor2_8
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _6071_/A _6071_/B _6071_/C _6071_/D VGND VGND VPWR VPWR _6071_/X sky130_fd_sc_hd__or4_1
Xhold1118 _6552_/Q VGND VGND VPWR VPWR _4070_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1129 _6599_/Q VGND VGND VPWR VPWR _4125_/A0 sky130_fd_sc_hd__bufbuf_16
X_5022_ _5022_/A _5022_/B _5022_/C _5022_/D VGND VGND VPWR VPWR _5180_/C sky130_fd_sc_hd__or4_2
XFILLER_100_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1107 _7105_/Q VGND VGND VPWR VPWR _5545_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_65_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6973_ _7133_/CLK _6973_/D fanout443/X VGND VGND VPWR VPWR _6973_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_53_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5924_ _6596_/Q _5681_/X _5923_/X VGND VGND VPWR VPWR _5927_/C sky130_fd_sc_hd__a21o_1
XFILLER_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5855_ _7020_/Q _5682_/X _5688_/X _7036_/Q VGND VGND VPWR VPWR _5855_/X sky130_fd_sc_hd__a22o_1
X_4806_ _5142_/A _4806_/B _5099_/B _4806_/D VGND VGND VPWR VPWR _4806_/X sky130_fd_sc_hd__or4_1
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5786_ _5663_/A _7178_/Q _6358_/B1 VGND VGND VPWR VPWR _5786_/X sky130_fd_sc_hd__a21o_1
X_4737_ _4898_/B _5062_/C VGND VGND VPWR VPWR _4737_/Y sky130_fd_sc_hd__nor2_4
XFILLER_135_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4668_ _4758_/B _4668_/B VGND VGND VPWR VPWR _4886_/B sky130_fd_sc_hd__nand2_8
XFILLER_147_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3619_ _6967_/Q _5387_/A _5360_/A _6943_/Q VGND VGND VPWR VPWR _3619_/X sky130_fd_sc_hd__a22o_2
XFILLER_107_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold930 _6686_/Q VGND VGND VPWR VPWR hold930/X sky130_fd_sc_hd__bufbuf_16
X_6407_ _6407_/A0 _6407_/A1 _6411_/S VGND VGND VPWR VPWR _6407_/X sky130_fd_sc_hd__mux2_1
XFILLER_162_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold952 _6591_/Q VGND VGND VPWR VPWR hold952/X sky130_fd_sc_hd__bufbuf_16
X_4599_ _4622_/B _4868_/A VGND VGND VPWR VPWR _4893_/A sky130_fd_sc_hd__nand2_4
Xhold963 _6845_/Q VGND VGND VPWR VPWR hold963/X sky130_fd_sc_hd__bufbuf_16
Xhold941 _4198_/X VGND VGND VPWR VPWR _6660_/D sky130_fd_sc_hd__bufbuf_16
Xhold985 _6861_/Q VGND VGND VPWR VPWR hold985/X sky130_fd_sc_hd__bufbuf_16
Xhold974 _6869_/Q VGND VGND VPWR VPWR hold974/X sky130_fd_sc_hd__bufbuf_16
XFILLER_143_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold996 _6787_/Q VGND VGND VPWR VPWR hold996/X sky130_fd_sc_hd__bufbuf_16
X_6338_ _6658_/Q _6311_/B _6036_/Y _6752_/Q _6335_/X VGND VGND VPWR VPWR _6343_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6269_ _6269_/A _6269_/B _6269_/C _6269_/D VGND VGND VPWR VPWR _6269_/X sky130_fd_sc_hd__or4_2
XFILLER_130_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_3_0_csclk clkbuf_2_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_7_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_69_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3970_ _3970_/A _3970_/B VGND VGND VPWR VPWR _3970_/X sky130_fd_sc_hd__and2_2
XFILLER_149_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5640_ _7167_/Q _7166_/Q VGND VGND VPWR VPWR _6032_/A sky130_fd_sc_hd__and2b_4
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5571_ _5571_/A0 hold601/X _5575_/S VGND VGND VPWR VPWR _5571_/X sky130_fd_sc_hd__mux2_1
X_4522_ _5023_/A _4871_/A _4617_/A VGND VGND VPWR VPWR _5022_/A sky130_fd_sc_hd__a21oi_2
Xhold204 _6465_/Q VGND VGND VPWR VPWR hold204/X sky130_fd_sc_hd__bufbuf_16
X_4453_ _4584_/A _4663_/B VGND VGND VPWR VPWR _4453_/Y sky130_fd_sc_hd__nor2_8
XFILLER_144_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold215 hold812/X VGND VGND VPWR VPWR _5252_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold226 _3344_/Y VGND VGND VPWR VPWR _3995_/A sky130_fd_sc_hd__bufbuf_16
XFILLER_172_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3404_ _7115_/Q hold85/A _5594_/A _7155_/Q VGND VGND VPWR VPWR _3404_/X sky130_fd_sc_hd__a22o_4
XFILLER_144_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold248 _7073_/Q VGND VGND VPWR VPWR hold248/X sky130_fd_sc_hd__bufbuf_16
Xhold237 _6945_/Q VGND VGND VPWR VPWR hold237/X sky130_fd_sc_hd__bufbuf_16
Xhold259 _5436_/X VGND VGND VPWR VPWR _7008_/D sky130_fd_sc_hd__bufbuf_16
X_4384_ _5031_/A _4584_/A VGND VGND VPWR VPWR _4871_/A sky130_fd_sc_hd__or2_4
XFILLER_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7172_ _7196_/CLK _7172_/D fanout433/X VGND VGND VPWR VPWR _7172_/Q sky130_fd_sc_hd__dfrtp_1
X_6123_ _6888_/Q _6020_/A _6021_/D _7144_/Q _6122_/X VGND VGND VPWR VPWR _6123_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_131_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3335_ _5225_/A hold84/X VGND VGND VPWR VPWR _3978_/A sky130_fd_sc_hd__nor2_8
XFILLER_140_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6054_ _6925_/Q _6025_/C _6010_/Y _7021_/Q _6053_/X VGND VGND VPWR VPWR _6057_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3266_ _3991_/S hold88/X hold113/X VGND VGND VPWR VPWR hold89/A sky130_fd_sc_hd__a21oi_4
X_5005_ _5005_/A _5062_/A _5005_/C VGND VGND VPWR VPWR _5050_/C sky130_fd_sc_hd__and3_4
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3197_ _5663_/A VGND VGND VPWR VPWR _3197_/Y sky130_fd_sc_hd__inv_8
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6956_ _6964_/CLK _6956_/D fanout443/X VGND VGND VPWR VPWR _6956_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5907_ _6635_/Q _5675_/X _5684_/X _6724_/Q _5906_/X VGND VGND VPWR VPWR _5910_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_53_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6887_ _7153_/CLK _6887_/D fanout444/X VGND VGND VPWR VPWR _6887_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_14_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5838_ _6963_/Q _5673_/X _5699_/X _6931_/Q _5837_/X VGND VGND VPWR VPWR _5839_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5769_ _7000_/Q _5667_/X _5687_/X _7048_/Q VGND VGND VPWR VPWR _5769_/X sky130_fd_sc_hd__a22o_1
XFILLER_163_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold771 _4018_/X VGND VGND VPWR VPWR _6510_/D sky130_fd_sc_hd__bufbuf_16
Xhold782 _6976_/Q VGND VGND VPWR VPWR hold782/X sky130_fd_sc_hd__bufbuf_16
Xhold760 _4035_/X VGND VGND VPWR VPWR _6522_/D sky130_fd_sc_hd__bufbuf_16
Xhold793 _6936_/Q VGND VGND VPWR VPWR hold793/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput309 _3385_/X VGND VGND VPWR VPWR serial_data_2 sky130_fd_sc_hd__buf_8
XFILLER_113_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6810_ _6810_/CLK _6810_/D fanout419/X VGND VGND VPWR VPWR _6810_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6741_ _6759_/CLK _6741_/D fanout419/X VGND VGND VPWR VPWR _6741_/Q sky130_fd_sc_hd__dfrtp_2
X_3953_ _3991_/S _3953_/B VGND VGND VPWR VPWR _3953_/Y sky130_fd_sc_hd__nor2_2
X_6672_ _6672_/CLK _6672_/D fanout453/X VGND VGND VPWR VPWR _6672_/Q sky130_fd_sc_hd__dfrtp_2
X_3884_ _6472_/Q _6456_/Q _6454_/B VGND VGND VPWR VPWR _3974_/B sky130_fd_sc_hd__o21ai_4
X_5623_ _7162_/Q _7161_/Q VGND VGND VPWR VPWR _5702_/B sky130_fd_sc_hd__nor2_8
X_5554_ hold819/X _5599_/A0 hold86/X VGND VGND VPWR VPWR _5554_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4505_ _4812_/A _4687_/A VGND VGND VPWR VPWR _4505_/X sky130_fd_sc_hd__or2_4
XFILLER_172_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5485_ hold505/X _5584_/A0 _5485_/S VGND VGND VPWR VPWR _5485_/X sky130_fd_sc_hd__mux2_1
X_4436_ _4696_/A _4436_/B _4446_/B VGND VGND VPWR VPWR _4529_/C sky130_fd_sc_hd__and3_4
XFILLER_116_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7224_ _7225_/CLK _7224_/D fanout420/X VGND VGND VPWR VPWR _7224_/Q sky130_fd_sc_hd__dfrtp_2
X_7155_ _7156_/CLK _7155_/D fanout452/X VGND VGND VPWR VPWR _7155_/Q sky130_fd_sc_hd__dfrtp_2
X_4367_ _4728_/A _4478_/B _4986_/A _6705_/Q VGND VGND VPWR VPWR _4367_/X sky130_fd_sc_hd__o31a_2
XFILLER_132_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6106_ _6106_/A _6106_/B _6106_/C _6106_/D VGND VGND VPWR VPWR _6107_/C sky130_fd_sc_hd__or4_1
XFILLER_113_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3318_ _6860_/Q _3315_/Y _3317_/Y _7068_/Q VGND VGND VPWR VPWR _3318_/X sky130_fd_sc_hd__a22o_1
XFILLER_112_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4298_ _4298_/A _6406_/B VGND VGND VPWR VPWR _4303_/S sky130_fd_sc_hd__nand2_4
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7086_ _7129_/CLK _7086_/D fanout428/X VGND VGND VPWR VPWR _7086_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_132_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6037_ _6037_/A _6037_/B _6037_/C VGND VGND VPWR VPWR _6335_/B sky130_fd_sc_hd__and3_4
XFILLER_100_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3249_ _3845_/A _3249_/B VGND VGND VPWR VPWR _3249_/Y sky130_fd_sc_hd__nand2b_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6939_ _6939_/CLK _6939_/D fanout454/X VGND VGND VPWR VPWR _6939_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_csclk _3954_/X VGND VGND VPWR VPWR clkbuf_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_173_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold590 _5340_/X VGND VGND VPWR VPWR _6923_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_0_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_1_0_1_csclk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_441 hold319/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_452 _3802_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_430 _5561_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_474 _6693_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_463 _5602_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5270_ hold28/X _5594_/B VGND VGND VPWR VPWR hold29/A sky130_fd_sc_hd__nand2_8
XFILLER_114_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4221_ _4221_/A0 _4220_/X _4235_/S VGND VGND VPWR VPWR _4221_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4152_ hold817/X _4326_/A0 _4153_/S VGND VGND VPWR VPWR _4152_/X sky130_fd_sc_hd__mux2_1
X_4083_ _4083_/A0 _5289_/A0 _4087_/S VGND VGND VPWR VPWR _4083_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4985_ _4507_/A _5004_/B _4842_/X VGND VGND VPWR VPWR _4985_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_23_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6724_ _6747_/CLK _6724_/D fanout427/X VGND VGND VPWR VPWR _6724_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3936_ _6842_/Q input81/X _3970_/B VGND VGND VPWR VPWR _3936_/X sky130_fd_sc_hd__mux2_8
XFILLER_51_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_2_0_csclk clkbuf_3_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_2_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_137_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6655_ _7225_/CLK _6655_/D fanout422/X VGND VGND VPWR VPWR _6655_/Q sky130_fd_sc_hd__dfrtp_2
X_3867_ _3875_/B _3864_/B _3861_/B _6467_/Q _3866_/X VGND VGND VPWR VPWR _6467_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6586_ _7220_/CLK _6586_/D VGND VGND VPWR VPWR _6586_/Q sky130_fd_sc_hd__dfxtp_2
X_3798_ _6664_/Q _3797_/X _6485_/Q VGND VGND VPWR VPWR _3801_/B sky130_fd_sc_hd__o21a_1
X_5606_ _6680_/Q _5606_/B _5665_/B VGND VGND VPWR VPWR _5617_/A sky130_fd_sc_hd__or3_2
XFILLER_192_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5537_ _5582_/A0 hold634/X _5539_/S VGND VGND VPWR VPWR _5537_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7207_ _7209_/CLK _7207_/D VGND VGND VPWR VPWR _7207_/Q sky130_fd_sc_hd__dfxtp_4
X_5468_ _5468_/A _5576_/B VGND VGND VPWR VPWR _5476_/S sky130_fd_sc_hd__nand2_8
XFILLER_160_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4419_ _4707_/B _4773_/A VGND VGND VPWR VPWR _4426_/A sky130_fd_sc_hd__nand2_2
X_5399_ hold784/X _5597_/A0 _5404_/S VGND VGND VPWR VPWR _5399_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout366 _5486_/B VGND VGND VPWR VPWR _5594_/B sky130_fd_sc_hd__bufbuf_16
XFILLER_86_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7138_ _7138_/CLK _7138_/D fanout456/X VGND VGND VPWR VPWR _7138_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout377 hold76/X VGND VGND VPWR VPWR hold77/A sky130_fd_sc_hd__buf_8
XFILLER_143_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout388 _5561_/A0 VGND VGND VPWR VPWR _6409_/A0 sky130_fd_sc_hd__buf_8
XFILLER_59_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7069_ _7136_/CLK _7069_/D fanout436/X VGND VGND VPWR VPWR _7069_/Q sky130_fd_sc_hd__dfstp_4
Xfanout399 _6407_/A0 VGND VGND VPWR VPWR _5234_/C sky130_fd_sc_hd__buf_8
XFILLER_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput19 mask_rev_in[23] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__clkbuf_4
XFILLER_182_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_260 spi_sdoenb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_271 wb_adr_i[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_282 wb_dat_i[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_293 input96/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4770_ _5087_/A _5087_/C _5165_/A VGND VGND VPWR VPWR _5035_/B sky130_fd_sc_hd__o21a_2
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3721_ _6497_/Q _3344_/Y _4262_/A _6719_/Q VGND VGND VPWR VPWR _3721_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3652_ _7103_/Q hold21/A _3551_/Y input97/X VGND VGND VPWR VPWR _3652_/X sky130_fd_sc_hd__a22o_2
X_6440_ _6446_/A _6446_/B VGND VGND VPWR VPWR _6440_/X sky130_fd_sc_hd__and2_1
X_6371_ _6372_/A _6371_/B VGND VGND VPWR VPWR _6371_/Y sky130_fd_sc_hd__nand2_1
X_3583_ _7128_/Q _5567_/A _4160_/A _6632_/Q VGND VGND VPWR VPWR _3583_/X sky130_fd_sc_hd__a22o_1
XFILLER_127_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5322_ _5601_/A0 hold737/X _5323_/S VGND VGND VPWR VPWR _5322_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5253_ _5234_/C hold963/X _5260_/S VGND VGND VPWR VPWR _5253_/X sky130_fd_sc_hd__mux2_1
X_4204_ hold953/X _4203_/X _4218_/S VGND VGND VPWR VPWR _4204_/X sky130_fd_sc_hd__mux2_1
X_5184_ _5184_/A _5184_/B VGND VGND VPWR VPWR _6784_/D sky130_fd_sc_hd__or2_2
X_4135_ _5545_/A0 _4135_/A1 _4135_/S VGND VGND VPWR VPWR _4135_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_63_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7136_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_83_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4066_ _5545_/A0 _4066_/A1 _4066_/S VGND VGND VPWR VPWR _4066_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_78_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6845_/CLK sky130_fd_sc_hd__clkbuf_8
X_4968_ _4537_/X _4959_/A _4959_/B _4906_/B VGND VGND VPWR VPWR _5071_/D sky130_fd_sc_hd__a31o_4
XFILLER_165_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4899_ _4965_/A _4899_/B VGND VGND VPWR VPWR _4976_/A sky130_fd_sc_hd__nor2_1
X_6707_ _7209_/CLK _6707_/D _6362_/B VGND VGND VPWR VPWR _6707_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3919_ _6832_/Q _5626_/A _3918_/X VGND VGND VPWR VPWR _6677_/D sky130_fd_sc_hd__o21ai_1
XFILLER_165_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6638_ _6786_/CLK _6638_/D fanout417/X VGND VGND VPWR VPWR _6638_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_106_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6569_ _7220_/CLK _6569_/D VGND VGND VPWR VPWR _6569_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_16_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _6745_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_133_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5940_ _7186_/Q _6309_/S _5938_/X _5939_/X VGND VGND VPWR VPWR _7186_/D sky130_fd_sc_hd__o22a_1
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5871_ _5871_/A _5871_/B _5871_/C _5871_/D VGND VGND VPWR VPWR _5871_/X sky130_fd_sc_hd__or4_2
XFILLER_34_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4822_ _4956_/C _4684_/Y _4653_/Y VGND VGND VPWR VPWR _5047_/C sky130_fd_sc_hd__a21o_2
XFILLER_61_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4753_ _4753_/A _4753_/B _4753_/C _4753_/D VGND VGND VPWR VPWR _4753_/X sky130_fd_sc_hd__and4_1
XFILLER_146_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3704_ _6878_/Q _5288_/A _4148_/A _6620_/Q VGND VGND VPWR VPWR _3704_/X sky130_fd_sc_hd__a22o_1
X_4684_ _4685_/A _4746_/B VGND VGND VPWR VPWR _4684_/Y sky130_fd_sc_hd__nor2_4
X_6423_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6423_/X sky130_fd_sc_hd__and2_1
X_3635_ _3635_/A _3635_/B _3635_/C _3635_/D VGND VGND VPWR VPWR _3636_/D sky130_fd_sc_hd__or4_1
XFILLER_134_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3566_ _6936_/Q _5351_/A _4256_/A _6716_/Q VGND VGND VPWR VPWR _3588_/A sky130_fd_sc_hd__a22o_1
X_6354_ _6717_/Q _6023_/B _6021_/C _6549_/Q _6353_/X VGND VGND VPWR VPWR _6355_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5305_ _5602_/A0 hold366/X _5305_/S VGND VGND VPWR VPWR _5305_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6285_ _7198_/Q _6309_/S _6284_/X VGND VGND VPWR VPWR _7198_/D sky130_fd_sc_hd__o21a_1
X_3497_ hold53/X _5234_/B VGND VGND VPWR VPWR _6406_/A sky130_fd_sc_hd__nor2_8
X_5236_ _5236_/A _5558_/B VGND VGND VPWR VPWR _5237_/S sky130_fd_sc_hd__nand2_1
XFILLER_115_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5167_ _5101_/B _5163_/X _5166_/X _5161_/X VGND VGND VPWR VPWR _5167_/X sky130_fd_sc_hd__o31a_1
XFILLER_130_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5098_ _5098_/A _5098_/B _5098_/C VGND VGND VPWR VPWR _5101_/B sky130_fd_sc_hd__or3_2
X_4118_ _4118_/A hold47/X VGND VGND VPWR VPWR _4123_/S sky130_fd_sc_hd__and2_4
XFILLER_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4049_ _4049_/A _6406_/B VGND VGND VPWR VPWR _4054_/S sky130_fd_sc_hd__and2_4
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold8 hold8/A VGND VGND VPWR VPWR hold8/X sky130_fd_sc_hd__bufbuf_16
XFILLER_181_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold408 _6495_/Q VGND VGND VPWR VPWR hold408/X sky130_fd_sc_hd__bufbuf_16
X_3420_ _4241_/A _3732_/B VGND VGND VPWR VPWR _5245_/A sky130_fd_sc_hd__nor2_8
XFILLER_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold419 _5539_/X VGND VGND VPWR VPWR _7100_/D sky130_fd_sc_hd__bufbuf_16
X_3351_ _7004_/Q _5423_/A _5594_/A _7156_/Q _3348_/X VGND VGND VPWR VPWR _3378_/C
+ sky130_fd_sc_hd__a221o_4
XFILLER_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6070_ _6982_/Q _6028_/X _6034_/Y _6990_/Q _6069_/X VGND VGND VPWR VPWR _6071_/D
+ sky130_fd_sc_hd__a221o_2
Xload_slew355 _3473_/A VGND VGND VPWR VPWR _3543_/A sky130_fd_sc_hd__buf_8
X_3282_ hold90/X _3383_/C VGND VGND VPWR VPWR _3534_/A sky130_fd_sc_hd__or2_4
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1119 _6743_/Q VGND VGND VPWR VPWR _4293_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_112_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5021_ _6780_/Q _4239_/X _4979_/X _5020_/X VGND VGND VPWR VPWR _6780_/D sky130_fd_sc_hd__o22a_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1108 _5545_/X VGND VGND VPWR VPWR _7105_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_66_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6972_ _7156_/CLK _6972_/D fanout451/X VGND VGND VPWR VPWR _6972_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5923_ _6591_/Q _5680_/X _5687_/X _6641_/Q VGND VGND VPWR VPWR _5923_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5854_ _6964_/Q _5673_/X _5676_/X _6980_/Q _5853_/X VGND VGND VPWR VPWR _5861_/A
+ sky130_fd_sc_hd__a221o_4
XFILLER_179_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4805_ _4805_/A _4805_/B _4805_/C _4638_/X VGND VGND VPWR VPWR _4806_/D sky130_fd_sc_hd__or4b_1
XFILLER_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5785_ _6856_/Q _5722_/B _5777_/X _5784_/X _3197_/Y VGND VGND VPWR VPWR _5785_/X
+ sky130_fd_sc_hd__o221a_1
X_4736_ _4748_/A _4736_/B VGND VGND VPWR VPWR _5147_/C sky130_fd_sc_hd__nor2_2
XFILLER_119_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4667_ _5050_/A _4714_/B VGND VGND VPWR VPWR _5147_/B sky130_fd_sc_hd__or2_4
XFILLER_135_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3618_ _6606_/Q _4130_/A _4082_/A _6565_/Q VGND VGND VPWR VPWR _3618_/X sky130_fd_sc_hd__a22o_1
Xhold931 _4231_/X VGND VGND VPWR VPWR _6686_/D sky130_fd_sc_hd__bufbuf_16
Xhold920 _6489_/Q VGND VGND VPWR VPWR hold920/X sky130_fd_sc_hd__bufbuf_16
X_6406_ _6406_/A _6406_/B VGND VGND VPWR VPWR _6411_/S sky130_fd_sc_hd__nand2_4
Xhold942 _6725_/Q VGND VGND VPWR VPWR hold942/X sky130_fd_sc_hd__bufbuf_16
XFILLER_143_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold953 _6669_/Q VGND VGND VPWR VPWR hold953/X sky130_fd_sc_hd__bufbuf_16
XFILLER_134_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4598_ _4997_/A _4749_/C VGND VGND VPWR VPWR _4846_/B sky130_fd_sc_hd__nor2_4
XFILLER_115_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6337_ _6762_/Q _6010_/Y _6031_/X _6648_/Q _6336_/X VGND VGND VPWR VPWR _6343_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold964 _5253_/X VGND VGND VPWR VPWR _6845_/D sky130_fd_sc_hd__bufbuf_16
Xhold975 _6981_/Q VGND VGND VPWR VPWR hold975/X sky130_fd_sc_hd__bufbuf_16
XFILLER_142_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold986 _6565_/Q VGND VGND VPWR VPWR hold986/X sky130_fd_sc_hd__bufbuf_16
Xhold997 _6490_/Q VGND VGND VPWR VPWR hold997/X sky130_fd_sc_hd__bufbuf_16
XFILLER_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3549_ _4108_/A1 _6793_/Q _3857_/C VGND VGND VPWR VPWR _3549_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6268_ _6625_/Q _6028_/X _6034_/Y _6724_/Q _6267_/X VGND VGND VPWR VPWR _6269_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6199_ _6907_/Q _6021_/A _6025_/A _6939_/Q _6198_/X VGND VGND VPWR VPWR _6206_/A
+ sky130_fd_sc_hd__a221o_1
X_5219_ _5219_/A0 _5541_/A0 _5222_/S VGND VGND VPWR VPWR _5219_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5570_ _5597_/A0 hold437/X _5575_/S VGND VGND VPWR VPWR _5570_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4521_ _4871_/A _4617_/A VGND VGND VPWR VPWR _4798_/A sky130_fd_sc_hd__nor2_1
Xhold205 hold205/A VGND VGND VPWR VPWR hold205/X sky130_fd_sc_hd__bufbuf_16
XFILLER_172_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4452_ _4694_/A VGND VGND VPWR VPWR _4452_/Y sky130_fd_sc_hd__inv_2
Xhold216 _5252_/X VGND VGND VPWR VPWR _5260_/S sky130_fd_sc_hd__bufbuf_16
XFILLER_132_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold249 _5509_/X VGND VGND VPWR VPWR _7073_/D sky130_fd_sc_hd__bufbuf_16
X_3403_ _7131_/Q _5567_/A _5279_/A _6875_/Q VGND VGND VPWR VPWR _3403_/X sky130_fd_sc_hd__a22o_1
Xhold227 _4002_/X VGND VGND VPWR VPWR _6502_/D sky130_fd_sc_hd__bufbuf_16
Xhold238 _5365_/X VGND VGND VPWR VPWR _6945_/D sky130_fd_sc_hd__bufbuf_16
X_4383_ _5031_/A _4584_/A VGND VGND VPWR VPWR _4500_/A sky130_fd_sc_hd__nor2_8
XFILLER_125_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7171_ _7193_/CLK _7171_/D fanout456/X VGND VGND VPWR VPWR _7171_/Q sky130_fd_sc_hd__dfrtp_2
X_6122_ _7112_/Q _6027_/B _6021_/B _7152_/Q VGND VGND VPWR VPWR _6122_/X sky130_fd_sc_hd__a22o_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3334_ _3506_/A hold20/X VGND VGND VPWR VPWR _3334_/Y sky130_fd_sc_hd__nor2_8
XFILLER_105_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6053_ _6949_/Q _6022_/A _6009_/X _7069_/Q VGND VGND VPWR VPWR _6053_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_0__1132_ _3548_/X VGND VGND VPWR VPWR clkbuf_0__1132_/X sky130_fd_sc_hd__clkbuf_8
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ _3991_/S hold286/X hold113/X VGND VGND VPWR VPWR _3265_/X sky130_fd_sc_hd__a21o_4
X_5004_ _5004_/A _5004_/B VGND VGND VPWR VPWR _5037_/B sky130_fd_sc_hd__and2_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3196_ _6666_/Q VGND VGND VPWR VPWR _3196_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6955_ _6976_/CLK _6955_/D fanout450/X VGND VGND VPWR VPWR _6955_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_121_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5906_ _6546_/Q _5674_/X _5688_/X _6769_/Q VGND VGND VPWR VPWR _5906_/X sky130_fd_sc_hd__a22o_1
X_6886_ _7111_/CLK _6886_/D fanout444/X VGND VGND VPWR VPWR _6886_/Q sky130_fd_sc_hd__dfstp_4
X_5837_ _7003_/Q _5667_/X _5681_/X _6923_/Q VGND VGND VPWR VPWR _5837_/X sky130_fd_sc_hd__a22o_1
XFILLER_167_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5768_ _7088_/Q _5685_/X _5699_/X _6928_/Q VGND VGND VPWR VPWR _5768_/X sky130_fd_sc_hd__a22o_1
XFILLER_182_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4719_ _4690_/A _4719_/B _4719_/C VGND VGND VPWR VPWR _4719_/X sky130_fd_sc_hd__and3b_4
XFILLER_154_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5699_ _5864_/B _5706_/B _5707_/B VGND VGND VPWR VPWR _5699_/X sky130_fd_sc_hd__and3_4
XFILLER_107_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold772 _6711_/Q VGND VGND VPWR VPWR hold772/X sky130_fd_sc_hd__bufbuf_16
Xhold761 _6597_/Q VGND VGND VPWR VPWR hold761/X sky130_fd_sc_hd__bufbuf_16
Xhold750 _7225_/Q VGND VGND VPWR VPWR hold750/X sky130_fd_sc_hd__bufbuf_16
Xhold794 _6613_/Q VGND VGND VPWR VPWR hold794/X sky130_fd_sc_hd__bufbuf_16
Xhold783 _5400_/X VGND VGND VPWR VPWR _6976_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_131_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6740_ _6759_/CLK _6740_/D fanout421/X VGND VGND VPWR VPWR _6740_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_23_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3952_ _7174_/Q _6827_/Q _6831_/Q VGND VGND VPWR VPWR _3952_/X sky130_fd_sc_hd__mux2_2
XFILLER_188_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6671_ _6672_/CLK _6671_/D fanout453/X VGND VGND VPWR VPWR _6671_/Q sky130_fd_sc_hd__dfrtp_2
X_3883_ _6472_/Q _6456_/Q _6454_/B VGND VGND VPWR VPWR _3883_/X sky130_fd_sc_hd__o21a_4
XFILLER_188_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5622_ _6679_/Q _5620_/Y _7161_/Q VGND VGND VPWR VPWR _7161_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5553_ hold584/X _5571_/A0 hold86/X VGND VGND VPWR VPWR _7112_/D sky130_fd_sc_hd__mux2_1
XFILLER_136_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4504_ _4812_/A _5164_/B VGND VGND VPWR VPWR _5087_/B sky130_fd_sc_hd__nor2_2
XFILLER_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5484_ hold721/X _5583_/A0 _5485_/S VGND VGND VPWR VPWR _5484_/X sky130_fd_sc_hd__mux2_1
X_4435_ _4696_/A _4446_/B VGND VGND VPWR VPWR _4440_/B sky130_fd_sc_hd__nand2_4
XFILLER_105_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7223_ _7225_/CLK _7223_/D fanout422/X VGND VGND VPWR VPWR _7223_/Q sky130_fd_sc_hd__dfstp_4
X_7154_ _7154_/CLK _7154_/D fanout451/X VGND VGND VPWR VPWR _7154_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_160_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4366_ _4364_/A _4364_/B _4388_/B VGND VGND VPWR VPWR _4553_/B sky130_fd_sc_hd__o21bai_4
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6105_ _6863_/Q _6025_/D _6029_/X _7047_/Q _6104_/X VGND VGND VPWR VPWR _6106_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_113_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3317_ _3501_/A _3515_/B VGND VGND VPWR VPWR _3317_/Y sky130_fd_sc_hd__nor2_8
XFILLER_86_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4297_ _5545_/A0 _4297_/A1 _4297_/S VGND VGND VPWR VPWR _4297_/X sky130_fd_sc_hd__mux2_1
X_7085_ _7132_/CLK _7085_/D fanout428/X VGND VGND VPWR VPWR _7085_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_100_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6036_ _6036_/A _6036_/B VGND VGND VPWR VPWR _6036_/Y sky130_fd_sc_hd__nor2_8
X_3248_ _6487_/Q _6486_/Q _6485_/Q VGND VGND VPWR VPWR _3857_/C sky130_fd_sc_hd__or3_4
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6938_ _7154_/CLK _6938_/D fanout451/X VGND VGND VPWR VPWR _6938_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6869_ _7151_/CLK _6869_/D fanout447/X VGND VGND VPWR VPWR _6869_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_22_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold580 _5384_/X VGND VGND VPWR VPWR _6962_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold591 _6928_/Q VGND VGND VPWR VPWR hold591/X sky130_fd_sc_hd__bufbuf_16
XFILLER_77_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_442 hold337/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_453 _3924_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_431 _5578_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_420 input1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_475 _4029_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_464 _6411_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4220_ hold963/X _5234_/C _4234_/S VGND VGND VPWR VPWR _4220_/X sky130_fd_sc_hd__mux2_1
X_4151_ hold950/X _5300_/A0 _4153_/S VGND VGND VPWR VPWR _4151_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4082_ _4082_/A _5558_/B VGND VGND VPWR VPWR _4087_/S sky130_fd_sc_hd__and2_4
XFILLER_110_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4984_ _4871_/A _4749_/C _4812_/A VGND VGND VPWR VPWR _5004_/B sky130_fd_sc_hd__a21oi_4
XFILLER_51_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6723_ _6725_/CLK _6723_/D fanout442/X VGND VGND VPWR VPWR _6723_/Q sky130_fd_sc_hd__dfrtp_2
X_3935_ _6840_/Q input78/X _3970_/B VGND VGND VPWR VPWR _3935_/X sky130_fd_sc_hd__mux2_8
XFILLER_177_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6654_ _7225_/CLK _6654_/D fanout422/X VGND VGND VPWR VPWR _6654_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_176_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5605_ _5615_/D VGND VGND VPWR VPWR _5605_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3866_ _6664_/Q _3866_/B VGND VGND VPWR VPWR _3866_/X sky130_fd_sc_hd__and2b_1
XFILLER_176_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6585_ _7220_/CLK _6585_/D VGND VGND VPWR VPWR _6585_/Q sky130_fd_sc_hd__dfxtp_2
X_3797_ _6667_/Q _6666_/Q VGND VGND VPWR VPWR _3797_/X sky130_fd_sc_hd__or2_4
XFILLER_127_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5536_ hold185/A hold269/X _5539_/S VGND VGND VPWR VPWR _5536_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5467_ _5584_/A0 hold406/X _5467_/S VGND VGND VPWR VPWR _5467_/X sky130_fd_sc_hd__mux2_1
X_4418_ _5050_/A _4711_/A VGND VGND VPWR VPWR _4773_/A sky130_fd_sc_hd__xor2_4
XFILLER_132_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7206_ _7208_/CLK _7206_/D VGND VGND VPWR VPWR _7206_/Q sky130_fd_sc_hd__dfxtp_4
X_5398_ hold508/X _5587_/A0 _5404_/S VGND VGND VPWR VPWR _6974_/D sky130_fd_sc_hd__mux2_1
X_4349_ _4349_/A _4349_/B _4349_/C _4349_/D VGND VGND VPWR VPWR _4352_/A sky130_fd_sc_hd__and4_1
X_7137_ _7137_/CLK _7137_/D fanout443/X VGND VGND VPWR VPWR _7137_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout367 _4719_/C VGND VGND VPWR VPWR _4758_/B sky130_fd_sc_hd__buf_8
X_7068_ _7122_/CLK _7068_/D fanout443/X VGND VGND VPWR VPWR _7068_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_101_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout378 _6411_/A0 VGND VGND VPWR VPWR _5545_/A0 sky130_fd_sc_hd__buf_8
XFILLER_86_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout389 hold43/A VGND VGND VPWR VPWR _5561_/A0 sky130_fd_sc_hd__buf_8
XFILLER_100_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6019_ _6019_/A _6036_/B VGND VGND VPWR VPWR _6021_/D sky130_fd_sc_hd__nor2_8
XFILLER_74_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_261 spimemio_flash_io3_do VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_250 mask_rev_in[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_283 wb_dat_i[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_272 wb_adr_i[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_294 input93/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3720_ _6990_/Q _3299_/Y _3368_/Y input12/X _3679_/X VGND VGND VPWR VPWR _3725_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3651_ _6532_/Q _4043_/A _4166_/A _6636_/Q _3650_/X VGND VGND VPWR VPWR _3654_/C
+ sky130_fd_sc_hd__a221o_4
XFILLER_146_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3582_ _6920_/Q _5333_/A _5306_/A _6896_/Q _3581_/X VGND VGND VPWR VPWR _3587_/B
+ sky130_fd_sc_hd__a221o_1
X_6370_ _7210_/Q _3379_/X _6370_/S VGND VGND VPWR VPWR _7210_/D sky130_fd_sc_hd__mux2_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5321_ _5600_/A0 hold581/X _5323_/S VGND VGND VPWR VPWR _5321_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5252_ _5252_/A _5252_/B _6454_/B _5252_/D VGND VGND VPWR VPWR _5252_/X sky130_fd_sc_hd__or4_4
X_5183_ _5143_/Y _5146_/Y _5175_/X _5182_/X VGND VGND VPWR VPWR _5184_/B sky130_fd_sc_hd__a31o_1
X_4203_ hold956/X hold885/X _4217_/S VGND VGND VPWR VPWR _4203_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4134_ _4326_/A0 _4134_/A1 _4135_/S VGND VGND VPWR VPWR _4134_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4065_ _4326_/A0 hold786/X _4066_/S VGND VGND VPWR VPWR _6548_/D sky130_fd_sc_hd__mux2_1
XFILLER_64_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4967_ _4956_/C _4719_/X _4959_/X _4571_/Y _4628_/Y VGND VGND VPWR VPWR _5073_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_51_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4898_ _4965_/A _4898_/B VGND VGND VPWR VPWR _4911_/B sky130_fd_sc_hd__nor2_1
X_6706_ _7220_/CLK _6706_/D _6362_/B VGND VGND VPWR VPWR _6706_/Q sky130_fd_sc_hd__dfrtp_2
X_3918_ _5659_/C _3918_/B VGND VGND VPWR VPWR _3918_/X sky130_fd_sc_hd__or2_1
XFILLER_192_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3849_ _3196_/Y _6668_/Q _3859_/B _6473_/Q VGND VGND VPWR VPWR _6473_/D sky130_fd_sc_hd__a31o_1
X_6637_ _6786_/CLK _6637_/D fanout418/X VGND VGND VPWR VPWR _6637_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_137_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6568_ _7209_/CLK _6568_/D VGND VGND VPWR VPWR _6568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5519_ _5582_/A0 hold670/X _5521_/S VGND VGND VPWR VPWR _5519_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6499_ _6810_/CLK _6499_/D fanout419/X VGND VGND VPWR VPWR _6499_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_160_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5870_ _6972_/Q _5691_/X _5699_/X _6932_/Q _5869_/X VGND VGND VPWR VPWR _5871_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4821_ _5119_/A _5135_/A VGND VGND VPWR VPWR _5013_/B sky130_fd_sc_hd__or2_2
XFILLER_73_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4752_ _4947_/B _5147_/C _4756_/B VGND VGND VPWR VPWR _4753_/D sky130_fd_sc_hd__a21o_1
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4683_ _4745_/A _4832_/B VGND VGND VPWR VPWR _5151_/A sky130_fd_sc_hd__nor2_2
X_3703_ _6926_/Q _5342_/A _5396_/A _6974_/Q _3702_/X VGND VGND VPWR VPWR _3709_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3634_ _6863_/Q hold28/A _5306_/A _6895_/Q _3633_/X VGND VGND VPWR VPWR _3635_/D
+ sky130_fd_sc_hd__a221o_1
X_6422_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6422_/X sky130_fd_sc_hd__and2_1
XFILLER_146_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6353_ _6663_/Q _5996_/X _6020_/C _6593_/Q VGND VGND VPWR VPWR _6353_/X sky130_fd_sc_hd__a22o_1
X_3565_ _7016_/Q _3359_/Y _4274_/A _6731_/Q VGND VGND VPWR VPWR _3565_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5304_ _5601_/A0 hold539/X _5305_/S VGND VGND VPWR VPWR _5304_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6284_ _5611_/A _7197_/Q _6358_/B1 _6283_/X VGND VGND VPWR VPWR _6284_/X sky130_fd_sc_hd__a211o_1
X_3496_ input24/X _3302_/Y _5360_/A _6945_/Q _3495_/X VGND VGND VPWR VPWR _3504_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5235_ _5235_/A1 _5227_/A _5576_/B _5234_/X VGND VGND VPWR VPWR _5235_/X sky130_fd_sc_hd__o211a_1
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5166_ _5166_/A _5166_/B _5166_/C _4935_/C VGND VGND VPWR VPWR _5166_/X sky130_fd_sc_hd__or4b_2
XFILLER_69_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5097_ _5164_/A _4995_/A _5096_/X VGND VGND VPWR VPWR _5098_/C sky130_fd_sc_hd__o21ai_1
XFILLER_110_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4117_ _5545_/A0 _4117_/A1 _4117_/S VGND VGND VPWR VPWR _4117_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4048_ _4048_/A0 _5545_/A0 _4048_/S VGND VGND VPWR VPWR _6534_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5999_ _6019_/A _6004_/A VGND VGND VPWR VPWR _6023_/A sky130_fd_sc_hd__nor2_8
XFILLER_24_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput290 _6818_/Q VGND VGND VPWR VPWR pll_trim[23] sky130_fd_sc_hd__buf_8
XFILLER_181_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold9 hold9/A VGND VGND VPWR VPWR hold9/X sky130_fd_sc_hd__bufbuf_16
XFILLER_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire351 _6232_/A VGND VGND VPWR VPWR _6306_/A sky130_fd_sc_hd__buf_6
Xhold409 _6986_/Q VGND VGND VPWR VPWR hold409/X sky130_fd_sc_hd__bufbuf_16
XFILLER_143_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_62_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7101_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_128_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3350_ _3673_/B _4241_/A VGND VGND VPWR VPWR _5594_/A sky130_fd_sc_hd__nor2_8
XFILLER_124_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_77_csclk clkbuf_opt_2_0_csclk/X VGND VGND VPWR VPWR _6824_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_3_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5020_ _5102_/C _4946_/X _5002_/X _5019_/X VGND VGND VPWR VPWR _5020_/X sky130_fd_sc_hd__a211o_4
XFILLER_98_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3281_ hold18/X hold82/X VGND VGND VPWR VPWR _3383_/C sky130_fd_sc_hd__nand2_2
XFILLER_2_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xload_slew356 _3476_/A VGND VGND VPWR VPWR _5225_/A sky130_fd_sc_hd__buf_8
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1109 _6609_/Q VGND VGND VPWR VPWR _4137_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_85_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6971_ _6971_/CLK _6971_/D fanout451/X VGND VGND VPWR VPWR _6971_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_81_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5922_ _6715_/Q _5676_/X _5682_/X _6750_/Q _5921_/X VGND VGND VPWR VPWR _5927_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_15_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _6725_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5853_ _6924_/Q _5681_/X _5707_/X _7028_/Q VGND VGND VPWR VPWR _5853_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4804_ _4654_/A _4958_/A _4702_/A _4711_/C _4803_/X VGND VGND VPWR VPWR _4805_/C
+ sky130_fd_sc_hd__a41o_1
X_5784_ _5784_/A _5784_/B _5784_/C VGND VGND VPWR VPWR _5784_/X sky130_fd_sc_hd__or3_4
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4735_ _4818_/A _4735_/B _4566_/A VGND VGND VPWR VPWR _4735_/X sky130_fd_sc_hd__or3b_2
XFILLER_159_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4666_ _5050_/A _4714_/B VGND VGND VPWR VPWR _4668_/B sky130_fd_sc_hd__nor2_8
XFILLER_119_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3617_ _6887_/Q _5297_/A _5288_/A _6879_/Q VGND VGND VPWR VPWR _3617_/X sky130_fd_sc_hd__a22o_1
X_4597_ _4648_/B _4947_/B VGND VGND VPWR VPWR _4957_/A sky130_fd_sc_hd__nor2_4
XFILLER_134_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6405_ _7220_/Q _6704_/Q _4239_/X _6404_/X VGND VGND VPWR VPWR _7220_/D sky130_fd_sc_hd__o31a_1
Xhold910 _6640_/Q VGND VGND VPWR VPWR hold910/X sky130_fd_sc_hd__bufbuf_16
Xhold921 _6683_/Q VGND VGND VPWR VPWR hold921/X sky130_fd_sc_hd__bufbuf_16
Xhold943 _6509_/Q VGND VGND VPWR VPWR hold943/X sky130_fd_sc_hd__bufbuf_16
Xhold954 _4204_/X VGND VGND VPWR VPWR _6669_/D sky130_fd_sc_hd__bufbuf_16
X_3548_ _3548_/A _3548_/B _3548_/C VGND VGND VPWR VPWR _3548_/X sky130_fd_sc_hd__or3_2
X_6336_ _6737_/Q _6020_/B _6011_/X _6789_/Q VGND VGND VPWR VPWR _6336_/X sky130_fd_sc_hd__a22o_1
Xhold932 _6801_/Q VGND VGND VPWR VPWR hold932/X sky130_fd_sc_hd__bufbuf_16
Xhold965 _6893_/Q VGND VGND VPWR VPWR hold965/X sky130_fd_sc_hd__bufbuf_16
Xhold976 _7109_/Q VGND VGND VPWR VPWR hold976/X sky130_fd_sc_hd__bufbuf_16
Xhold987 _4085_/X VGND VGND VPWR VPWR _6565_/D sky130_fd_sc_hd__bufbuf_16
Xhold998 _6532_/Q VGND VGND VPWR VPWR hold998/X sky130_fd_sc_hd__bufbuf_16
XFILLER_142_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3479_ _6873_/Q _5279_/A _4148_/A _6623_/Q _3477_/X VGND VGND VPWR VPWR _3488_/B
+ sky130_fd_sc_hd__a221o_1
X_6267_ _7222_/Q _6009_/X _6020_/D _6709_/Q VGND VGND VPWR VPWR _6267_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6198_ _6955_/Q _6022_/A _6025_/C _6931_/Q VGND VGND VPWR VPWR _6198_/X sky130_fd_sc_hd__a22o_1
XFILLER_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5218_ _5218_/A _5576_/B VGND VGND VPWR VPWR _5222_/S sky130_fd_sc_hd__and2_4
XFILLER_130_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5149_ _5146_/A _5146_/B _5175_/C _5143_/Y VGND VGND VPWR VPWR _5169_/B sky130_fd_sc_hd__o31a_1
XFILLER_72_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4520_ _4370_/Y _4503_/Y _4506_/X _4484_/B _4533_/A VGND VGND VPWR VPWR _4520_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_144_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold206 _3991_/X VGND VGND VPWR VPWR hold206/X sky130_fd_sc_hd__bufbuf_16
X_4451_ _4525_/A _4590_/A VGND VGND VPWR VPWR _4694_/A sky130_fd_sc_hd__or2_4
Xhold217 _5256_/X VGND VGND VPWR VPWR _6848_/D sky130_fd_sc_hd__bufbuf_16
X_7170_ _7193_/CLK _7170_/D fanout455/X VGND VGND VPWR VPWR _7170_/Q sky130_fd_sc_hd__dfstp_4
Xhold239 _7072_/Q VGND VGND VPWR VPWR hold239/X sky130_fd_sc_hd__bufbuf_16
X_3402_ _6883_/Q _5288_/A _5360_/A _6947_/Q _3401_/X VGND VGND VPWR VPWR _3415_/B
+ sky130_fd_sc_hd__a221o_4
Xhold228 _7024_/Q VGND VGND VPWR VPWR hold228/X sky130_fd_sc_hd__bufbuf_16
X_4382_ _4469_/A _4819_/A VGND VGND VPWR VPWR _4584_/A sky130_fd_sc_hd__nand2_8
XFILLER_125_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6121_ _6121_/A _6121_/B _6121_/C _6121_/D VGND VGND VPWR VPWR _6121_/X sky130_fd_sc_hd__or4_4
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _3476_/A _3733_/B VGND VGND VPWR VPWR _5207_/A sky130_fd_sc_hd__nor2_8
X_6052_ _6901_/Q _6021_/A _6021_/B _7149_/Q _6051_/X VGND VGND VPWR VPWR _6057_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ _3991_/S _3264_/B VGND VGND VPWR VPWR _3264_/X sky130_fd_sc_hd__and2b_4
X_5003_ _5003_/A _5003_/B _5003_/C VGND VGND VPWR VPWR _5003_/X sky130_fd_sc_hd__and3_1
XFILLER_140_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3195_ _6704_/Q VGND VGND VPWR VPWR _3916_/A sky130_fd_sc_hd__clkinv_8
XFILLER_66_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6954_ _6971_/CLK _6954_/D fanout451/X VGND VGND VPWR VPWR _6954_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_121_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5905_ _6620_/Q _5673_/X _5681_/X _6595_/Q _5904_/X VGND VGND VPWR VPWR _5910_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_81_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6885_ _7054_/CLK _6885_/D fanout444/X VGND VGND VPWR VPWR _6885_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5836_ _6971_/Q _5691_/X _5835_/X VGND VGND VPWR VPWR _5839_/C sky130_fd_sc_hd__a21o_1
X_5767_ _6896_/Q _5694_/X _5706_/X _7056_/Q VGND VGND VPWR VPWR _5767_/X sky130_fd_sc_hd__a22o_1
XFILLER_182_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4718_ _4745_/A _4757_/B VGND VGND VPWR VPWR _5178_/A sky130_fd_sc_hd__nor2_4
X_5698_ _5864_/B _5698_/B VGND VGND VPWR VPWR _5722_/B sky130_fd_sc_hd__nand2_8
XFILLER_190_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4649_ _4722_/B _4650_/B VGND VGND VPWR VPWR _4719_/C sky130_fd_sc_hd__nor2_8
XFILLER_135_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold773 _4254_/X VGND VGND VPWR VPWR _6711_/D sky130_fd_sc_hd__bufbuf_16
Xhold740 _4291_/X VGND VGND VPWR VPWR _6742_/D sky130_fd_sc_hd__bufbuf_16
Xhold751 _6411_/X VGND VGND VPWR VPWR _7225_/D sky130_fd_sc_hd__bufbuf_16
Xhold762 _4122_/X VGND VGND VPWR VPWR _6597_/D sky130_fd_sc_hd__bufbuf_16
Xhold795 _4141_/X VGND VGND VPWR VPWR _6613_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_150_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold784 _6975_/Q VGND VGND VPWR VPWR hold784/X sky130_fd_sc_hd__bufbuf_16
XFILLER_115_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6319_ _7224_/Q _6009_/X _6020_/D _6711_/Q VGND VGND VPWR VPWR _6319_/X sky130_fd_sc_hd__a22o_1
XFILLER_162_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3951_ _7172_/Q _6828_/Q _6831_/Q VGND VGND VPWR VPWR _3951_/X sky130_fd_sc_hd__mux2_4
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6670_ _6672_/CLK _6670_/D fanout453/X VGND VGND VPWR VPWR _6670_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3882_ _7173_/Q _6826_/Q _6831_/Q VGND VGND VPWR VPWR _3920_/B sky130_fd_sc_hd__mux2_8
X_5621_ _6677_/Q _6679_/Q VGND VGND VPWR VPWR _5621_/X sky130_fd_sc_hd__or2_2
X_5552_ hold543/X _5597_/A0 hold86/X VGND VGND VPWR VPWR _5552_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4503_ _5087_/A VGND VGND VPWR VPWR _4503_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5483_ hold655/X _5582_/A0 _5485_/S VGND VGND VPWR VPWR _5483_/X sky130_fd_sc_hd__mux2_1
X_4434_ _4818_/A _4672_/A _4469_/A _4395_/D VGND VGND VPWR VPWR _4446_/B sky130_fd_sc_hd__o211a_4
XFILLER_144_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7222_ _7222_/CLK _7222_/D fanout422/X VGND VGND VPWR VPWR _7222_/Q sky130_fd_sc_hd__dfrtp_2
X_7153_ _7153_/CLK _7153_/D fanout444/X VGND VGND VPWR VPWR _7153_/Q sky130_fd_sc_hd__dfrtp_2
X_4365_ _4707_/B _4364_/B _4340_/B VGND VGND VPWR VPWR _4388_/B sky130_fd_sc_hd__o21a_1
XFILLER_113_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6104_ _7103_/Q _5653_/X _6022_/B _6943_/Q VGND VGND VPWR VPWR _6104_/X sky130_fd_sc_hd__a22o_1
XFILLER_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3316_ _3421_/A _3421_/B hold83/X VGND VGND VPWR VPWR _3386_/B sky130_fd_sc_hd__or3_4
X_7084_ _7140_/CLK _7084_/D fanout430/X VGND VGND VPWR VPWR _7084_/Q sky130_fd_sc_hd__dfrtp_2
X_6035_ _6035_/A _6037_/C _6035_/C VGND VGND VPWR VPWR _6311_/B sky130_fd_sc_hd__and3_4
X_4296_ _4326_/A0 hold835/X _4297_/S VGND VGND VPWR VPWR _4296_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3247_ _4707_/B VGND VGND VPWR VPWR _4655_/A sky130_fd_sc_hd__inv_4
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6937_ _7121_/CLK _6937_/D fanout442/X VGND VGND VPWR VPWR _6937_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_81_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6868_ _7124_/CLK hold30/X fanout437/X VGND VGND VPWR VPWR _6868_/Q sky130_fd_sc_hd__dfrtp_2
X_5819_ _7042_/Q _5683_/X _5704_/X _6938_/Q _5810_/X VGND VGND VPWR VPWR _5826_/A
+ sky130_fd_sc_hd__a221o_1
X_6799_ _6804_/CLK _6799_/D _6439_/A VGND VGND VPWR VPWR _6799_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold581 _6906_/Q VGND VGND VPWR VPWR hold581/X sky130_fd_sc_hd__bufbuf_16
XFILLER_123_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold570 _7002_/Q VGND VGND VPWR VPWR hold570/X sky130_fd_sc_hd__bufbuf_16
XFILLER_173_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold592 _5346_/X VGND VGND VPWR VPWR _6928_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_106_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_410 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_432 _5596_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_443 hold411/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_421 _6356_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_454 _5341_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_465 _5581_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_476 _4235_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4150_ hold637/X _5587_/A0 _4153_/S VGND VGND VPWR VPWR _4150_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4081_ _6562_/Q _3379_/X _4081_/S VGND VGND VPWR VPWR _6562_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4983_ _5013_/A _4983_/B VGND VGND VPWR VPWR _5135_/B sky130_fd_sc_hd__or2_2
XFILLER_63_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6722_ _6722_/CLK _6722_/D fanout427/X VGND VGND VPWR VPWR _6722_/Q sky130_fd_sc_hd__dfstp_1
X_3934_ _6839_/Q input80/X _3970_/B VGND VGND VPWR VPWR _3934_/X sky130_fd_sc_hd__mux2_8
X_3865_ _3866_/B _3865_/B VGND VGND VPWR VPWR _6468_/D sky130_fd_sc_hd__xnor2_1
X_6653_ _6777_/CLK _6653_/D fanout424/X VGND VGND VPWR VPWR _6653_/Q sky130_fd_sc_hd__dfrtp_2
X_5604_ _5663_/A _6680_/Q _6679_/Q _3920_/Y VGND VGND VPWR VPWR _5615_/D sky130_fd_sc_hd__o31a_4
XFILLER_191_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6584_ _7220_/CLK _6584_/D VGND VGND VPWR VPWR _6584_/Q sky130_fd_sc_hd__dfxtp_2
X_3796_ _6790_/Q _3928_/A _3794_/X _3795_/Y VGND VGND VPWR VPWR _6790_/D sky130_fd_sc_hd__a22o_1
XFILLER_164_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5535_ hold136/X hold221/X _5539_/S VGND VGND VPWR VPWR _7096_/D sky130_fd_sc_hd__mux2_1
XFILLER_191_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5466_ _5583_/A0 hold653/X _5467_/S VGND VGND VPWR VPWR _5466_/X sky130_fd_sc_hd__mux2_1
X_4417_ _4650_/B _4416_/B _4415_/X VGND VGND VPWR VPWR _5165_/A sky130_fd_sc_hd__a21oi_4
XFILLER_160_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7205_ _7209_/CLK _7205_/D VGND VGND VPWR VPWR _7205_/Q sky130_fd_sc_hd__dfxtp_4
X_5397_ hold918/X hold885/X _5404_/S VGND VGND VPWR VPWR _6973_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4348_ _4368_/A _4722_/B VGND VGND VPWR VPWR _4774_/A sky130_fd_sc_hd__or2_4
XFILLER_113_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7136_ _7136_/CLK _7136_/D fanout437/X VGND VGND VPWR VPWR _7136_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout368 _4687_/A VGND VGND VPWR VPWR _5164_/B sky130_fd_sc_hd__buf_8
XFILLER_100_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout379 hold185/A VGND VGND VPWR VPWR _6411_/A0 sky130_fd_sc_hd__buf_8
XFILLER_74_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7067_ _7131_/CLK _7067_/D fanout432/X VGND VGND VPWR VPWR _7067_/Q sky130_fd_sc_hd__dfrtp_2
X_4279_ _6411_/A0 hold788/X _4279_/S VGND VGND VPWR VPWR _4279_/X sky130_fd_sc_hd__mux2_1
X_6018_ _6018_/A _6035_/C _6032_/C VGND VGND VPWR VPWR _6022_/D sky130_fd_sc_hd__and3_4
XFILLER_86_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_251 _6512_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_240 mask_rev_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_284 wb_dat_i[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_273 wb_adr_i[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_262 spimemio_flash_io3_oeb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_295 _7227_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3650_ input13/X _3368_/Y _5238_/A _6834_/Q VGND VGND VPWR VPWR _3650_/X sky130_fd_sc_hd__a22o_4
XFILLER_127_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3581_ _6904_/Q _5315_/A _4097_/A _6579_/Q VGND VGND VPWR VPWR _3581_/X sky130_fd_sc_hd__a22o_1
X_5320_ _5581_/A0 hold444/X _5323_/S VGND VGND VPWR VPWR _5320_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5251_ hold78/X hold95/X _5251_/S VGND VGND VPWR VPWR hold96/A sky130_fd_sc_hd__mux2_1
XFILLER_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4202_ _4241_/B _6421_/B _4007_/X _4217_/S _5594_/B VGND VGND VPWR VPWR _4218_/S
+ sky130_fd_sc_hd__o221a_4
XFILLER_130_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5182_ _6784_/Q _6376_/A _5158_/Y _5178_/X _5181_/X VGND VGND VPWR VPWR _5182_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_87_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4133_ _5300_/A0 hold955/X _4135_/S VGND VGND VPWR VPWR _6606_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4064_ _5300_/A0 hold958/X _4066_/S VGND VGND VPWR VPWR _4064_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4966_ _4443_/X _4536_/B _4959_/A _4909_/B VGND VGND VPWR VPWR _5145_/B sky130_fd_sc_hd__a31o_1
X_6705_ _7220_/CLK _6705_/D _6362_/B VGND VGND VPWR VPWR _6705_/Q sky130_fd_sc_hd__dfrtp_2
X_4897_ _5003_/A _4897_/B VGND VGND VPWR VPWR _4913_/B sky130_fd_sc_hd__nand2_1
X_3917_ _6457_/Q _3192_/Y _6664_/Q _3843_/B _6665_/Q VGND VGND VPWR VPWR _6665_/D
+ sky130_fd_sc_hd__a41o_1
XFILLER_125_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3848_ _6474_/Q _6459_/Q _3848_/S VGND VGND VPWR VPWR _6474_/D sky130_fd_sc_hd__mux2_1
XFILLER_22_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6636_ _6786_/CLK _6636_/D fanout418/X VGND VGND VPWR VPWR _6636_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_118_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6567_ _6715_/CLK _6567_/D fanout439/X VGND VGND VPWR VPWR _6567_/Q sky130_fd_sc_hd__dfrtp_2
X_3779_ _7175_/Q _5227_/A _6406_/A _7221_/Q VGND VGND VPWR VPWR _3779_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5518_ hold185/X hold299/X _5521_/S VGND VGND VPWR VPWR _5518_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6498_ _6810_/CLK _6498_/D fanout419/X VGND VGND VPWR VPWR _6498_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_78_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5449_ _5584_/A0 hold421/X _5449_/S VGND VGND VPWR VPWR _5449_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7119_ _7119_/CLK _7119_/D fanout437/X VGND VGND VPWR VPWR _7119_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_86_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _6401_/A1 sky130_fd_sc_hd__clkbuf_8
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4820_ _5003_/C _4820_/B VGND VGND VPWR VPWR _4827_/A sky130_fd_sc_hd__nand2_1
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4751_ _4754_/B _4735_/X _5123_/B _4935_/D _5144_/B VGND VGND VPWR VPWR _4753_/C
+ sky130_fd_sc_hd__o2111a_1
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4682_ _4697_/A _4832_/B VGND VGND VPWR VPWR _4682_/Y sky130_fd_sc_hd__nor2_1
X_3702_ _6902_/Q _5315_/A _4061_/A _6546_/Q VGND VGND VPWR VPWR _3702_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6421_ _6421_/A _6421_/B VGND VGND VPWR VPWR _6421_/X sky130_fd_sc_hd__and2_1
X_3633_ _7127_/Q _5567_/A hold61/A _7135_/Q VGND VGND VPWR VPWR _3633_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6352_ _6539_/Q _6025_/D _6029_/X _6643_/Q _6351_/X VGND VGND VPWR VPWR _6355_/C
+ sky130_fd_sc_hd__a221o_1
X_3564_ _7000_/Q _5423_/A _4310_/A _6761_/Q VGND VGND VPWR VPWR _3564_/X sky130_fd_sc_hd__a22o_1
X_5303_ _5600_/A0 hold468/X _5305_/S VGND VGND VPWR VPWR _5303_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3495_ _6732_/Q _4274_/A _4196_/A _6663_/Q VGND VGND VPWR VPWR _3495_/X sky130_fd_sc_hd__a22o_1
X_6283_ _6531_/Q _6060_/B _6269_/X _6282_/X _6308_/S VGND VGND VPWR VPWR _6283_/X
+ sky130_fd_sc_hd__o221a_2
X_5234_ _5234_/A _5234_/B _5234_/C VGND VGND VPWR VPWR _5234_/X sky130_fd_sc_hd__or3_4
X_5165_ _5165_/A _5165_/B _5165_/C VGND VGND VPWR VPWR _5166_/B sky130_fd_sc_hd__and3_1
XFILLER_130_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4116_ _4326_/A0 hold829/X _4117_/S VGND VGND VPWR VPWR _4116_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5096_ _5164_/B _5017_/A _4756_/B _4724_/B VGND VGND VPWR VPWR _5096_/X sky130_fd_sc_hd__o22a_1
XFILLER_110_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4047_ hold792/X _4326_/A0 _4048_/S VGND VGND VPWR VPWR _6533_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5998_ _6019_/A _6037_/B _6033_/C VGND VGND VPWR VPWR _6020_/B sky130_fd_sc_hd__and3b_4
XFILLER_12_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4949_ _4949_/A _4949_/B _4949_/C _4959_/A VGND VGND VPWR VPWR _4950_/C sky130_fd_sc_hd__and4_1
XFILLER_178_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6619_ _6649_/CLK _6619_/D fanout439/X VGND VGND VPWR VPWR _6619_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_153_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput280 _6494_/Q VGND VGND VPWR VPWR pll_trim[14] sky130_fd_sc_hd__buf_8
XFILLER_121_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput291 _6504_/Q VGND VGND VPWR VPWR pll_trim[24] sky130_fd_sc_hd__buf_8
XFILLER_75_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3280_ _3476_/A VGND VGND VPWR VPWR _3280_/Y sky130_fd_sc_hd__inv_2
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew357 hold53/X VGND VGND VPWR VPWR _3501_/A sky130_fd_sc_hd__buf_8
XFILLER_66_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6970_ _7154_/CLK _6970_/D fanout451/X VGND VGND VPWR VPWR _6970_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5921_ _6661_/Q _5669_/X _5684_/X _6725_/Q VGND VGND VPWR VPWR _5921_/X sky130_fd_sc_hd__a22o_1
XFILLER_81_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5852_ _7182_/Q _6309_/S _5850_/X _5851_/X VGND VGND VPWR VPWR _7182_/D sky130_fd_sc_hd__o22a_1
XFILLER_179_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4803_ _4654_/A _4958_/A _5165_/A _4702_/A _4704_/X VGND VGND VPWR VPWR _4803_/X
+ sky130_fd_sc_hd__a41o_1
X_5783_ _6944_/Q _5705_/X _5707_/X _7024_/Q _5782_/X VGND VGND VPWR VPWR _5784_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4734_ _4724_/A _4724_/B _4503_/Y VGND VGND VPWR VPWR _4734_/X sky130_fd_sc_hd__o21a_1
XFILLER_147_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4665_ _4707_/B _4696_/B VGND VGND VPWR VPWR _4714_/B sky130_fd_sc_hd__nand2_8
XFILLER_135_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6404_ _3916_/A _4238_/B _6374_/X _6403_/X _6372_/A VGND VGND VPWR VPWR _6404_/X
+ sky130_fd_sc_hd__a32o_4
X_4596_ _4745_/B _4947_/B VGND VGND VPWR VPWR _5135_/A sky130_fd_sc_hd__nor2_8
X_3616_ _6959_/Q _5378_/A _5396_/A _6975_/Q VGND VGND VPWR VPWR _3616_/X sky130_fd_sc_hd__a22o_1
XFILLER_135_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold911 _4174_/X VGND VGND VPWR VPWR _6640_/D sky130_fd_sc_hd__bufbuf_16
Xhold922 _4225_/X VGND VGND VPWR VPWR _6683_/D sky130_fd_sc_hd__bufbuf_16
Xhold900 _4045_/X VGND VGND VPWR VPWR _6531_/D sky130_fd_sc_hd__bufbuf_16
Xhold944 _4016_/X VGND VGND VPWR VPWR _6509_/D sky130_fd_sc_hd__bufbuf_16
Xhold955 _6606_/Q VGND VGND VPWR VPWR hold955/X sky130_fd_sc_hd__bufbuf_16
X_3547_ _3547_/A _3547_/B _3547_/C _3547_/D VGND VGND VPWR VPWR _3548_/C sky130_fd_sc_hd__or4_2
X_6335_ _6777_/Q _6335_/B VGND VGND VPWR VPWR _6335_/X sky130_fd_sc_hd__and2_1
Xhold933 _5196_/X VGND VGND VPWR VPWR _6801_/D sky130_fd_sc_hd__bufbuf_16
Xhold988 _7141_/Q VGND VGND VPWR VPWR hold988/X sky130_fd_sc_hd__bufbuf_16
XFILLER_89_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold977 _7224_/Q VGND VGND VPWR VPWR hold977/X sky130_fd_sc_hd__bufbuf_16
Xhold966 _6637_/Q VGND VGND VPWR VPWR hold966/X sky130_fd_sc_hd__bufbuf_16
X_3478_ _3534_/A _3540_/A VGND VGND VPWR VPWR _4148_/A sky130_fd_sc_hd__nor2_8
Xhold999 _4046_/X VGND VGND VPWR VPWR _6532_/D sky130_fd_sc_hd__bufbuf_16
X_6266_ _6754_/Q _6023_/D _6030_/Y _6769_/Q _6265_/X VGND VGND VPWR VPWR _6269_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_57_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6197_ _7131_/Q _6023_/A _6033_/X _7011_/Q _6196_/X VGND VGND VPWR VPWR _6207_/C
+ sky130_fd_sc_hd__a221o_1
X_5217_ _5541_/A0 _5217_/A1 _5217_/S VGND VGND VPWR VPWR _6819_/D sky130_fd_sc_hd__mux2_1
X_5148_ _5148_/A _5148_/B _5066_/A _4612_/A VGND VGND VPWR VPWR _5175_/C sky130_fd_sc_hd__or4bb_4
XFILLER_151_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5079_ _5079_/A _5079_/B _5079_/C VGND VGND VPWR VPWR _5137_/A sky130_fd_sc_hd__or3_1
XFILLER_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold207 hold207/A VGND VGND VPWR VPWR hold207/X sky130_fd_sc_hd__bufbuf_16
X_4450_ _4572_/A _4572_/B VGND VGND VPWR VPWR _4590_/A sky130_fd_sc_hd__or2_2
XFILLER_171_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4381_ _4395_/D _4987_/B VGND VGND VPWR VPWR _5023_/A sky130_fd_sc_hd__nand2_8
Xhold218 _7129_/Q VGND VGND VPWR VPWR hold218/X sky130_fd_sc_hd__bufbuf_16
Xhold229 _5454_/X VGND VGND VPWR VPWR _7024_/D sky130_fd_sc_hd__bufbuf_16
X_3401_ _6979_/Q _5396_/A _3399_/X _3400_/X VGND VGND VPWR VPWR _3401_/X sky130_fd_sc_hd__a211o_1
X_6120_ _6984_/Q _6028_/X _6034_/Y _6992_/Q _6119_/X VGND VGND VPWR VPWR _6121_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_112_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3332_ _3383_/C _3343_/A VGND VGND VPWR VPWR _3733_/B sky130_fd_sc_hd__or2_4
XFILLER_140_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ _7125_/Q _6023_/A _6020_/D _6965_/Q VGND VGND VPWR VPWR _6051_/X sky130_fd_sc_hd__a22o_1
XFILLER_112_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ hold111/X hold24/X _3845_/A VGND VGND VPWR VPWR _3263_/X sky130_fd_sc_hd__mux2_1
X_5002_ _5084_/B _5001_/X _5121_/A VGND VGND VPWR VPWR _5002_/X sky130_fd_sc_hd__o21ba_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3194_ _6880_/Q VGND VGND VPWR VPWR _3194_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6953_ _7153_/CLK _6953_/D fanout442/X VGND VGND VPWR VPWR _6953_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_53_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6884_ _7156_/CLK _6884_/D fanout447/X VGND VGND VPWR VPWR _6884_/Q sky130_fd_sc_hd__dfrtp_2
X_5904_ _6709_/Q _5691_/X _5701_/X _6615_/Q VGND VGND VPWR VPWR _5904_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5835_ _7091_/Q _5685_/X _5689_/X _6907_/Q VGND VGND VPWR VPWR _5835_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5766_ _7178_/Q _6309_/S _5764_/X _5765_/X VGND VGND VPWR VPWR _7178_/D sky130_fd_sc_hd__o22a_1
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5697_ _5864_/B _5702_/B _5703_/B VGND VGND VPWR VPWR _5697_/X sky130_fd_sc_hd__and3_4
XFILLER_148_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4717_ _5164_/B _4717_/B VGND VGND VPWR VPWR _5022_/C sky130_fd_sc_hd__nor2_1
X_4648_ _4671_/A _4648_/B VGND VGND VPWR VPWR _4708_/B sky130_fd_sc_hd__nor2_1
XFILLER_135_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold730 _5457_/X VGND VGND VPWR VPWR _7027_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_190_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4579_ _4818_/C _5062_/A VGND VGND VPWR VPWR _4874_/B sky130_fd_sc_hd__or2_4
Xhold752 _6955_/Q VGND VGND VPWR VPWR hold752/X sky130_fd_sc_hd__bufbuf_16
Xhold741 _6902_/Q VGND VGND VPWR VPWR hold741/X sky130_fd_sc_hd__bufbuf_16
Xhold763 _6762_/Q VGND VGND VPWR VPWR hold763/X sky130_fd_sc_hd__bufbuf_16
Xhold796 _6952_/Q VGND VGND VPWR VPWR hold796/X sky130_fd_sc_hd__bufbuf_16
Xhold785 _5399_/X VGND VGND VPWR VPWR _6975_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_115_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold774 _6995_/Q VGND VGND VPWR VPWR hold774/X sky130_fd_sc_hd__bufbuf_16
X_6318_ _6731_/Q _5987_/Y _6022_/D _6597_/Q _6317_/X VGND VGND VPWR VPWR _6321_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6249_ _6733_/Q _6020_/B _6025_/C _6599_/Q VGND VGND VPWR VPWR _6249_/X sky130_fd_sc_hd__a22o_1
XFILLER_77_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_61_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7078_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_76_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6804_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_40_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_14_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _6843_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_134_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_29_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7127_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_82_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold90 hold90/A VGND VGND VPWR VPWR hold90/X sky130_fd_sc_hd__bufbuf_16
XFILLER_48_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3950_ _6511_/Q input93/X _6836_/Q VGND VGND VPWR VPWR _3950_/X sky130_fd_sc_hd__mux2_8
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3881_ _6471_/Q _6456_/Q _6666_/Q _3843_/B VGND VGND VPWR VPWR _6456_/D sky130_fd_sc_hd__o211a_1
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5620_ _6677_/Q _6679_/Q VGND VGND VPWR VPWR _5620_/Y sky130_fd_sc_hd__nor2_2
X_5551_ hold547/X _5587_/A0 hold86/X VGND VGND VPWR VPWR _7110_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4502_ _4986_/A _4812_/A VGND VGND VPWR VPWR _5087_/A sky130_fd_sc_hd__nor2_4
XFILLER_144_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7221_ _7222_/CLK _7221_/D fanout420/X VGND VGND VPWR VPWR _7221_/Q sky130_fd_sc_hd__dfrtp_2
X_5482_ hold271/X hold185/X _5485_/S VGND VGND VPWR VPWR _5482_/X sky130_fd_sc_hd__mux2_1
X_4433_ _4818_/A _4672_/A VGND VGND VPWR VPWR _4663_/B sky130_fd_sc_hd__or2_4
XFILLER_172_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7152_ _7152_/CLK _7152_/D fanout452/X VGND VGND VPWR VPWR _7152_/Q sky130_fd_sc_hd__dfrtp_2
X_4364_ _4364_/A _4364_/B VGND VGND VPWR VPWR _4478_/C sky130_fd_sc_hd__or2_4
XFILLER_116_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4295_ _5588_/A0 _4295_/A1 _4297_/S VGND VGND VPWR VPWR _6745_/D sky130_fd_sc_hd__mux2_1
X_6103_ _6871_/Q _6023_/C _6025_/B _6895_/Q _6102_/X VGND VGND VPWR VPWR _6106_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_113_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3315_ hold84/X _5234_/A VGND VGND VPWR VPWR _3315_/Y sky130_fd_sc_hd__nor2_8
X_7083_ _7139_/CLK _7083_/D fanout435/X VGND VGND VPWR VPWR _7083_/Q sky130_fd_sc_hd__dfrtp_2
X_3246_ _4958_/A VGND VGND VPWR VPWR _4654_/B sky130_fd_sc_hd__inv_6
XFILLER_140_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6034_ _6036_/A _6034_/B VGND VGND VPWR VPWR _6034_/Y sky130_fd_sc_hd__nor2_8
XFILLER_132_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6936_ _6976_/CLK _6936_/D fanout450/X VGND VGND VPWR VPWR _6936_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6867_ _7090_/CLK _6867_/D fanout438/X VGND VGND VPWR VPWR _6867_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5818_ _6946_/Q _5705_/X _5707_/X _7026_/Q _5817_/X VGND VGND VPWR VPWR _5827_/C
+ sky130_fd_sc_hd__a221o_1
X_6798_ _6824_/CLK _6798_/D _6439_/A VGND VGND VPWR VPWR _6798_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5749_ _6935_/Q _5704_/X _5706_/X _7055_/Q VGND VGND VPWR VPWR _5749_/X sky130_fd_sc_hd__a22o_1
XFILLER_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold560 _6987_/Q VGND VGND VPWR VPWR hold560/X sky130_fd_sc_hd__bufbuf_16
Xhold571 _5429_/X VGND VGND VPWR VPWR _7002_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_173_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold582 _5321_/X VGND VGND VPWR VPWR _6906_/D sky130_fd_sc_hd__bufbuf_16
Xhold593 _6940_/Q VGND VGND VPWR VPWR hold593/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1260 _6999_/Q VGND VGND VPWR VPWR _5426_/A1 sky130_fd_sc_hd__bufbuf_16
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_400 _6610_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_411 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_444 hold537/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_433 _5541_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_422 _6309_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_466 _5581_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_455 _5694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_477 _3875_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4080_ _6561_/Q _3415_/X _4081_/S VGND VGND VPWR VPWR _6561_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4982_ _4758_/A _4634_/B _4554_/A _4863_/B _4766_/A VGND VGND VPWR VPWR _5084_/B
+ sky130_fd_sc_hd__a311o_2
X_6721_ _6746_/CLK _6721_/D fanout427/X VGND VGND VPWR VPWR _6721_/Q sky130_fd_sc_hd__dfstp_2
X_3933_ _3205_/Y input82/X _3970_/B VGND VGND VPWR VPWR _3933_/X sky130_fd_sc_hd__mux2_8
XFILLER_177_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3864_ _6468_/Q _3864_/B VGND VGND VPWR VPWR _3865_/B sky130_fd_sc_hd__nor2_1
X_6652_ _6777_/CLK _6652_/D fanout424/X VGND VGND VPWR VPWR _6652_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5603_ _5663_/A _6679_/Q VGND VGND VPWR VPWR _5665_/B sky130_fd_sc_hd__nor2_4
XFILLER_164_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6583_ _7220_/CLK _6583_/D VGND VGND VPWR VPWR _6583_/Q sky130_fd_sc_hd__dfxtp_1
X_3795_ _3857_/C _3928_/A VGND VGND VPWR VPWR _3795_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5534_ hold43/X _5534_/A1 _5539_/S VGND VGND VPWR VPWR _5534_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5465_ _5582_/A0 hold615/X _5467_/S VGND VGND VPWR VPWR _5465_/X sky130_fd_sc_hd__mux2_1
X_4416_ _4722_/A _4416_/B VGND VGND VPWR VPWR _4774_/C sky130_fd_sc_hd__xor2_4
X_7204_ _7220_/CLK _7204_/D VGND VGND VPWR VPWR _7204_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_160_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5396_ _5396_/A _5594_/B VGND VGND VPWR VPWR _5404_/S sky130_fd_sc_hd__and2_4
XFILLER_99_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7135_ _7135_/CLK hold63/X fanout430/X VGND VGND VPWR VPWR _7135_/Q sky130_fd_sc_hd__dfrtp_2
X_4347_ _4368_/A _4722_/B VGND VGND VPWR VPWR _4467_/B sky130_fd_sc_hd__nor2_4
XFILLER_160_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7066_ _7130_/CLK _7066_/D fanout454/X VGND VGND VPWR VPWR _7066_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout369 hold3/X VGND VGND VPWR VPWR _5584_/A0 sky130_fd_sc_hd__buf_8
X_4278_ _6410_/A0 _4278_/A1 _4279_/S VGND VGND VPWR VPWR _4278_/X sky130_fd_sc_hd__mux2_1
X_3229_ _6944_/Q VGND VGND VPWR VPWR _3229_/Y sky130_fd_sc_hd__inv_2
X_6017_ _6019_/A _6034_/B VGND VGND VPWR VPWR _6023_/D sky130_fd_sc_hd__nor2_8
XFILLER_86_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _3954_/A2 sky130_fd_sc_hd__clkbuf_8
X_6919_ _7121_/CLK _6919_/D fanout442/X VGND VGND VPWR VPWR _6919_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold390 _7156_/Q VGND VGND VPWR VPWR hold390/X sky130_fd_sc_hd__bufbuf_16
XFILLER_151_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1090 _6755_/Q VGND VGND VPWR VPWR _4307_/A0 sky130_fd_sc_hd__bufbuf_16
XFILLER_46_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_230 _6476_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_252 mgmt_gpio_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_241 mask_rev_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_274 wb_adr_i[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_285 wb_dat_i[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_263 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_296 _7227_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3580_ _6864_/Q hold28/A _4055_/A _6543_/Q _3579_/X VGND VGND VPWR VPWR _3587_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_173_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5250_ _5599_/A0 hold880/X _5251_/S VGND VGND VPWR VPWR _5250_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4201_ _6411_/A0 hold821/X _4201_/S VGND VGND VPWR VPWR _4201_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5181_ _5095_/X _5166_/X _5180_/X _5161_/X VGND VGND VPWR VPWR _5181_/X sky130_fd_sc_hd__o31a_1
XFILLER_68_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4132_ _6408_/A0 hold503/X _4135_/S VGND VGND VPWR VPWR _4132_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4063_ _5587_/A0 hold323/X _4066_/S VGND VGND VPWR VPWR _4063_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4965_ _4965_/A _5062_/A VGND VGND VPWR VPWR _5069_/D sky130_fd_sc_hd__nor2_1
XFILLER_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3916_ _3916_/A _3916_/B VGND VGND VPWR VPWR _6698_/D sky130_fd_sc_hd__nand2_1
X_6704_ _7220_/CLK _6704_/D _6362_/B VGND VGND VPWR VPWR _6704_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4896_ _4987_/A _4586_/B _4736_/B _4689_/Y VGND VGND VPWR VPWR _4905_/C sky130_fd_sc_hd__a22o_4
XFILLER_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3847_ _6485_/Q _3847_/B VGND VGND VPWR VPWR _3848_/S sky130_fd_sc_hd__nor2_2
X_6635_ _6786_/CLK _6635_/D fanout418/X VGND VGND VPWR VPWR _6635_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6566_ _6715_/CLK hold72/X fanout439/X VGND VGND VPWR VPWR _6566_/Q sky130_fd_sc_hd__dfrtp_2
X_3778_ _6530_/Q _4043_/A _4304_/A _6753_/Q _3777_/X VGND VGND VPWR VPWR _3785_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5517_ hold136/X hold235/X _5521_/S VGND VGND VPWR VPWR _5517_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6497_ _6759_/CLK _6497_/D fanout419/X VGND VGND VPWR VPWR _6497_/Q sky130_fd_sc_hd__dfstp_4
X_5448_ _5583_/A0 hold685/X _5449_/S VGND VGND VPWR VPWR _5448_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5379_ hold885/X _6957_/Q _5386_/S VGND VGND VPWR VPWR _5379_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7118_ _7118_/CLK hold37/X fanout436/X VGND VGND VPWR VPWR _7118_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_101_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7049_ _7078_/CLK _7049_/D fanout431/X VGND VGND VPWR VPWR _7049_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_170_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4750_ _5062_/A _4832_/B VGND VGND VPWR VPWR _5144_/B sky130_fd_sc_hd__or2_4
XFILLER_159_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4681_ _4697_/A _4886_/B VGND VGND VPWR VPWR _5033_/B sky130_fd_sc_hd__nor2_1
XFILLER_119_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3701_ _7046_/Q _5477_/A _4043_/A _6531_/Q _3700_/X VGND VGND VPWR VPWR _3701_/X
+ sky130_fd_sc_hd__a221o_1
X_6420_ _6421_/A _6421_/B VGND VGND VPWR VPWR _6420_/X sky130_fd_sc_hd__and2_1
X_3632_ _6626_/Q _4154_/A _4097_/A _6578_/Q _3612_/X VGND VGND VPWR VPWR _3635_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6351_ _6638_/Q _5653_/X _6022_/B _6613_/Q VGND VGND VPWR VPWR _6351_/X sky130_fd_sc_hd__a22o_1
X_5302_ _5599_/A0 hold851/X _5305_/S VGND VGND VPWR VPWR _5302_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3563_ _6856_/Q _3315_/Y _4196_/A _6662_/Q VGND VGND VPWR VPWR _3563_/X sky130_fd_sc_hd__a22o_1
X_6282_ _6356_/A _6282_/B _6282_/C VGND VGND VPWR VPWR _6282_/X sky130_fd_sc_hd__or3_2
X_3494_ hold53/X _3543_/B VGND VGND VPWR VPWR _4196_/A sky130_fd_sc_hd__nor2_8
XFILLER_170_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5233_ _5578_/A0 _6831_/Q _5233_/S VGND VGND VPWR VPWR _5233_/X sky130_fd_sc_hd__mux2_1
X_5164_ _5164_/A _5164_/B VGND VGND VPWR VPWR _5165_/C sky130_fd_sc_hd__nand2_1
XFILLER_130_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_opt_3_0_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7119_/CLK sky130_fd_sc_hd__clkbuf_8
X_4115_ _5300_/A0 hold952/X _4117_/S VGND VGND VPWR VPWR _6591_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5095_ _5095_/A _5095_/B _5095_/C _5095_/D VGND VGND VPWR VPWR _5095_/X sky130_fd_sc_hd__or4_2
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4046_ hold998/X _6409_/A0 _4048_/S VGND VGND VPWR VPWR _4046_/X sky130_fd_sc_hd__mux2_1
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5997_ _6012_/A _6018_/A _6032_/C VGND VGND VPWR VPWR _6025_/A sky130_fd_sc_hd__and3_4
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4948_ _4949_/B _4537_/X _4959_/A _5130_/A VGND VGND VPWR VPWR _5065_/A sky130_fd_sc_hd__a31o_2
XFILLER_165_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4879_ _5005_/C _4832_/B _4633_/X VGND VGND VPWR VPWR _5145_/A sky130_fd_sc_hd__o21ai_2
XFILLER_193_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6618_ _6713_/CLK _6618_/D fanout427/X VGND VGND VPWR VPWR _6618_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6549_ _6840_/CLK _6549_/D fanout424/X VGND VGND VPWR VPWR _6549_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_4_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput270 _6804_/Q VGND VGND VPWR VPWR pll_div[4] sky130_fd_sc_hd__buf_8
XFILLER_160_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput281 _6495_/Q VGND VGND VPWR VPWR pll_trim[15] sky130_fd_sc_hd__buf_8
Xoutput292 _6505_/Q VGND VGND VPWR VPWR pll_trim[25] sky130_fd_sc_hd__buf_8
XFILLER_181_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew358 _5252_/A VGND VGND VPWR VPWR _4241_/A sky130_fd_sc_hd__buf_8
XFILLER_93_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5920_ _6578_/Q _5689_/X _5694_/X _6565_/Q _5919_/X VGND VGND VPWR VPWR _5927_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5851_ _5663_/A _7181_/Q _6358_/B1 VGND VGND VPWR VPWR _5851_/X sky130_fd_sc_hd__a21o_1
X_4802_ _4802_/A _4802_/B _4802_/C _4802_/D VGND VGND VPWR VPWR _4805_/B sky130_fd_sc_hd__or4_2
X_5782_ _7008_/Q _5678_/X _5692_/X _7072_/Q VGND VGND VPWR VPWR _5782_/X sky130_fd_sc_hd__a22o_1
X_4733_ _4672_/A _4566_/A _4648_/B _4732_/X VGND VGND VPWR VPWR _4733_/X sky130_fd_sc_hd__o31a_1
XFILLER_147_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6403_ _6706_/Q _6371_/B _6402_/X VGND VGND VPWR VPWR _6403_/X sky130_fd_sc_hd__a21o_1
X_4664_ _5164_/B _4832_/B _4724_/B _4832_/A VGND VGND VPWR VPWR _4664_/X sky130_fd_sc_hd__o22a_1
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4595_ _4949_/C _4595_/B VGND VGND VPWR VPWR _4612_/C sky130_fd_sc_hd__nand2_1
X_3615_ _6935_/Q _5351_/A _3511_/Y _6616_/Q VGND VGND VPWR VPWR _3615_/X sky130_fd_sc_hd__a22o_1
Xhold912 _6846_/Q VGND VGND VPWR VPWR hold912/X sky130_fd_sc_hd__bufbuf_16
Xhold901 _6786_/Q VGND VGND VPWR VPWR hold901/X sky130_fd_sc_hd__bufbuf_16
XFILLER_190_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold945 _6887_/Q VGND VGND VPWR VPWR hold945/X sky130_fd_sc_hd__bufbuf_16
XFILLER_143_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold923 _7133_/Q VGND VGND VPWR VPWR hold923/X sky130_fd_sc_hd__bufbuf_16
X_3546_ _3546_/A _3546_/B _3546_/C _3546_/D VGND VGND VPWR VPWR _3547_/D sky130_fd_sc_hd__or4_2
Xhold934 _6729_/Q VGND VGND VPWR VPWR hold934/X sky130_fd_sc_hd__bufbuf_16
X_6334_ _7200_/Q _6309_/S _6333_/X VGND VGND VPWR VPWR _7200_/D sky130_fd_sc_hd__o21a_1
XFILLER_143_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold956 _6690_/Q VGND VGND VPWR VPWR hold956/X sky130_fd_sc_hd__bufbuf_16
XFILLER_135_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold978 _6410_/X VGND VGND VPWR VPWR _7224_/D sky130_fd_sc_hd__bufbuf_16
Xhold989 _6538_/Q VGND VGND VPWR VPWR hold989/X sky130_fd_sc_hd__bufbuf_16
Xhold967 _4170_/X VGND VGND VPWR VPWR _6637_/D sky130_fd_sc_hd__bufbuf_16
X_6265_ _6729_/Q _5987_/Y _6022_/D _6595_/Q VGND VGND VPWR VPWR _6265_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3477_ _3973_/B _4023_/S _3726_/A _3476_/Y VGND VGND VPWR VPWR _3477_/X sky130_fd_sc_hd__a211o_4
X_5216_ _5216_/A _5576_/B VGND VGND VPWR VPWR _5217_/S sky130_fd_sc_hd__nand2_1
X_6196_ _6891_/Q _6020_/A _6021_/D _7147_/Q _6195_/X VGND VGND VPWR VPWR _6196_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_97_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5147_ _5147_/A _5147_/B _5147_/C VGND VGND VPWR VPWR _5148_/B sky130_fd_sc_hd__nor3_1
XFILLER_84_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5078_ _5078_/A _5078_/B _5078_/C VGND VGND VPWR VPWR _5079_/C sky130_fd_sc_hd__or3_1
X_4029_ hold71/X hold165/X _4033_/S VGND VGND VPWR VPWR _4029_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold208 hold208/A VGND VGND VPWR VPWR hold208/X sky130_fd_sc_hd__bufbuf_16
XFILLER_144_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4380_ _4740_/A _4395_/D VGND VGND VPWR VPWR _4818_/B sky130_fd_sc_hd__nand2_8
XFILLER_172_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold219 _5572_/X VGND VGND VPWR VPWR _7129_/D sky130_fd_sc_hd__bufbuf_16
X_3400_ _7067_/Q _3317_/Y _5207_/A _6817_/Q _3389_/X VGND VGND VPWR VPWR _3400_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_171_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3331_ _3331_/A _3331_/B _3331_/C _3331_/D VGND VGND VPWR VPWR _3379_/B sky130_fd_sc_hd__or4_1
XFILLER_98_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _7133_/Q _6020_/B _6023_/B _6973_/Q _6049_/X VGND VGND VPWR VPWR _6057_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ hold25/X hold121/X _3991_/S VGND VGND VPWR VPWR _3262_/X sky130_fd_sc_hd__mux2_8
XFILLER_39_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5001_ _5135_/B _5001_/B _5001_/C _5001_/D VGND VGND VPWR VPWR _5001_/X sky130_fd_sc_hd__or4_1
XFILLER_112_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3193_ _6698_/Q VGND VGND VPWR VPWR _6360_/A sky130_fd_sc_hd__inv_2
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6952_ _6976_/CLK _6952_/D fanout450/X VGND VGND VPWR VPWR _6952_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_81_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6883_ _6939_/CLK _6883_/D fanout453/X VGND VGND VPWR VPWR _6883_/Q sky130_fd_sc_hd__dfrtp_2
X_5903_ _6774_/Q _5683_/X _5704_/X _6605_/Q _5902_/X VGND VGND VPWR VPWR _5910_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5834_ _6955_/Q _5701_/X _5707_/X _7027_/Q _5833_/X VGND VGND VPWR VPWR _5839_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5765_ _5663_/A _7177_/Q _6358_/B1 VGND VGND VPWR VPWR _5765_/X sky130_fd_sc_hd__a21o_1
XFILLER_148_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5696_ _5702_/B _5703_/B VGND VGND VPWR VPWR _5698_/B sky130_fd_sc_hd__and2_4
X_4716_ _4754_/B _4724_/B VGND VGND VPWR VPWR _4797_/C sky130_fd_sc_hd__nor2_1
X_4647_ _4654_/B _4422_/Y _4707_/A _6706_/Q VGND VGND VPWR VPWR _4917_/B sky130_fd_sc_hd__o31a_4
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold720 _4012_/X VGND VGND VPWR VPWR _6507_/D sky130_fd_sc_hd__bufbuf_16
X_4578_ _4818_/B _4740_/B VGND VGND VPWR VPWR _5062_/A sky130_fd_sc_hd__or2_4
Xhold753 _5376_/X VGND VGND VPWR VPWR _6955_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_122_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold742 _6716_/Q VGND VGND VPWR VPWR hold742/X sky130_fd_sc_hd__bufbuf_16
Xhold764 _4315_/X VGND VGND VPWR VPWR _6762_/D sky130_fd_sc_hd__bufbuf_16
Xhold731 _6658_/Q VGND VGND VPWR VPWR hold731/X sky130_fd_sc_hd__bufbuf_16
X_6317_ _6756_/Q _6023_/D _6030_/Y _6771_/Q VGND VGND VPWR VPWR _6317_/X sky130_fd_sc_hd__a22o_1
Xhold797 _5373_/X VGND VGND VPWR VPWR _6952_/D sky130_fd_sc_hd__bufbuf_16
X_3529_ _3543_/A _4241_/B VGND VGND VPWR VPWR _4112_/A sky130_fd_sc_hd__nor2_8
Xhold786 _6548_/Q VGND VGND VPWR VPWR hold786/X sky130_fd_sc_hd__bufbuf_16
Xhold775 _5421_/X VGND VGND VPWR VPWR _6995_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_130_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6248_ _6248_/A _6248_/B _6248_/C VGND VGND VPWR VPWR _6248_/X sky130_fd_sc_hd__or3_2
XFILLER_77_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6179_ _6866_/Q _6025_/D _6029_/X _7050_/Q _6178_/X VGND VGND VPWR VPWR _6181_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold80 hold80/A VGND VGND VPWR VPWR hold80/X sky130_fd_sc_hd__bufbuf_16
Xhold91 hold91/A VGND VGND VPWR VPWR hold91/X sky130_fd_sc_hd__bufbuf_16
XFILLER_63_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3880_ _3875_/B _3848_/S _3879_/X _6457_/Q VGND VGND VPWR VPWR _6457_/D sky130_fd_sc_hd__a22o_1
XFILLER_43_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5550_ hold976/X _5595_/A0 hold86/X VGND VGND VPWR VPWR _7109_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4501_ _4501_/A _4812_/A VGND VGND VPWR VPWR _4672_/B sky130_fd_sc_hd__nor2_2
XFILLER_157_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5481_ hold266/X hold136/X _5485_/S VGND VGND VPWR VPWR _7048_/D sky130_fd_sc_hd__mux2_1
X_4432_ _4818_/A _4672_/A VGND VGND VPWR VPWR _4470_/B sky130_fd_sc_hd__nor2_4
X_7220_ _7220_/CLK _7220_/D _6362_/B VGND VGND VPWR VPWR _7220_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_132_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7151_ _7151_/CLK _7151_/D fanout446/X VGND VGND VPWR VPWR _7151_/Q sky130_fd_sc_hd__dfrtp_2
X_4363_ _5050_/A _4413_/C VGND VGND VPWR VPWR _4364_/B sky130_fd_sc_hd__and2_2
XFILLER_140_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6102_ _6959_/Q _6022_/C _6032_/X _7055_/Q VGND VGND VPWR VPWR _6102_/X sky130_fd_sc_hd__a22o_1
XFILLER_113_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4294_ _6408_/A0 hold568/X _4297_/S VGND VGND VPWR VPWR _4294_/X sky130_fd_sc_hd__mux2_1
X_3314_ _3314_/A _3314_/B VGND VGND VPWR VPWR _3551_/A sky130_fd_sc_hd__or2_4
X_7082_ _7139_/CLK _7082_/D fanout435/X VGND VGND VPWR VPWR _7082_/Q sky130_fd_sc_hd__dfrtp_2
X_3245_ _4395_/D VGND VGND VPWR VPWR _4819_/A sky130_fd_sc_hd__inv_6
X_6033_ _6037_/B _6037_/C _6033_/C VGND VGND VPWR VPWR _6033_/X sky130_fd_sc_hd__and3_4
XFILLER_58_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6935_ _7121_/CLK _6935_/D fanout442/X VGND VGND VPWR VPWR _6935_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6866_ _7154_/CLK hold79/X fanout452/X VGND VGND VPWR VPWR _6866_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5817_ _7010_/Q _5678_/X _5692_/X _7074_/Q VGND VGND VPWR VPWR _5817_/X sky130_fd_sc_hd__a22o_1
XFILLER_10_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6797_ _3545_/A1 _6797_/D _6455_/X VGND VGND VPWR VPWR _6797_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_157_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5748_ _7015_/Q _5682_/X _5685_/X _7087_/Q _5747_/X VGND VGND VPWR VPWR _5753_/B
+ sky130_fd_sc_hd__a221o_4
XFILLER_41_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5679_ _7164_/Q _7163_/Q VGND VGND VPWR VPWR _5707_/C sky130_fd_sc_hd__and2b_4
XFILLER_136_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold561 _5412_/X VGND VGND VPWR VPWR _6987_/D sky130_fd_sc_hd__bufbuf_16
Xhold572 _6888_/Q VGND VGND VPWR VPWR hold572/X sky130_fd_sc_hd__bufbuf_16
Xhold550 _6967_/Q VGND VGND VPWR VPWR hold550/X sky130_fd_sc_hd__bufbuf_16
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold583 _6896_/Q VGND VGND VPWR VPWR hold583/X sky130_fd_sc_hd__bufbuf_16
Xhold594 _5359_/X VGND VGND VPWR VPWR _6940_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_89_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1250 _7071_/Q VGND VGND VPWR VPWR _5507_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1261 _6823_/Q VGND VGND VPWR VPWR _5222_/A0 sky130_fd_sc_hd__bufbuf_16
XANTENNA_401 _6861_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_434 hold7/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_412 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_423 _5582_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_445 hold601/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_456 _6025_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_467 _5561_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_478 _6407_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput170 wb_we_i VGND VGND VPWR VPWR _6372_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4981_ _5003_/A _5102_/D VGND VGND VPWR VPWR _5121_/B sky130_fd_sc_hd__nand2_2
XFILLER_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3932_ _3204_/Y input90/X _3932_/S VGND VGND VPWR VPWR _3932_/X sky130_fd_sc_hd__mux2_8
XFILLER_149_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6720_ _6951_/CLK _6720_/D fanout442/X VGND VGND VPWR VPWR _6720_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_32_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3863_ _6469_/Q _3864_/B _3862_/Y _6468_/Q VGND VGND VPWR VPWR _6469_/D sky130_fd_sc_hd__o22a_1
X_6651_ _6777_/CLK _6651_/D fanout424/X VGND VGND VPWR VPWR _6651_/Q sky130_fd_sc_hd__dfstp_4
X_5602_ _5602_/A0 hold390/X _5602_/S VGND VGND VPWR VPWR _5602_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6582_ _7201_/CLK _6582_/D VGND VGND VPWR VPWR _6582_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_118_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3794_ _3794_/A _3794_/B _3794_/C _3794_/D VGND VGND VPWR VPWR _3794_/X sky130_fd_sc_hd__or4_4
X_5533_ _5578_/A0 hold360/X _5539_/S VGND VGND VPWR VPWR _7094_/D sky130_fd_sc_hd__mux2_1
XFILLER_157_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5464_ _6411_/A0 hold857/X _5467_/S VGND VGND VPWR VPWR _5464_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_60_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7135_/CLK sky130_fd_sc_hd__clkbuf_8
X_4415_ _4529_/A _4529_/B _4414_/B _4533_/A VGND VGND VPWR VPWR _4415_/X sky130_fd_sc_hd__a31o_2
X_5395_ _5602_/A0 hold368/X _5395_/S VGND VGND VPWR VPWR _5395_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7203_ _7208_/CLK _7203_/D VGND VGND VPWR VPWR _7203_/Q sky130_fd_sc_hd__dfxtp_4
X_4346_ _4722_/B _4345_/Y _4346_/S VGND VGND VPWR VPWR _4533_/A sky130_fd_sc_hd__mux2_8
XFILLER_99_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7134_ _7134_/CLK _7134_/D fanout428/X VGND VGND VPWR VPWR _7134_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_99_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7065_ _7133_/CLK _7065_/D fanout443/X VGND VGND VPWR VPWR _7065_/Q sky130_fd_sc_hd__dfrtp_2
Xclkbuf_leaf_75_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6810_/CLK sky130_fd_sc_hd__clkbuf_8
X_4277_ _6409_/A0 _4277_/A1 _4279_/S VGND VGND VPWR VPWR _6730_/D sky130_fd_sc_hd__mux2_1
X_3228_ _6952_/Q VGND VGND VPWR VPWR _3228_/Y sky130_fd_sc_hd__inv_2
X_6016_ _6032_/A _6035_/A _6018_/A VGND VGND VPWR VPWR _6022_/C sky130_fd_sc_hd__and3_4
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6918_ _7121_/CLK _6918_/D fanout442/X VGND VGND VPWR VPWR _6918_/Q sky130_fd_sc_hd__dfstp_4
Xclkbuf_leaf_13_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _6616_/CLK sky130_fd_sc_hd__clkbuf_8
X_6849_ _7106_/CLK _6849_/D fanout438/X VGND VGND VPWR VPWR _6849_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_10_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_28_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7151_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_151_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold380 _7004_/Q VGND VGND VPWR VPWR hold380/X sky130_fd_sc_hd__bufbuf_16
XFILLER_77_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold391 _5602_/X VGND VGND VPWR VPWR _7156_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_77_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1080 _7013_/Q VGND VGND VPWR VPWR _5442_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1091 _4307_/X VGND VGND VPWR VPWR _6755_/D sky130_fd_sc_hd__bufbuf_16
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_220 _6918_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_231 _6476_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_242 mask_rev_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_286 wb_dat_i[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_275 wb_adr_i[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_264 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_253 _7164_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_297 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4200_ _6410_/A0 _4200_/A1 _4201_/S VGND VGND VPWR VPWR _4200_/X sky130_fd_sc_hd__mux2_1
X_5180_ _5180_/A _5180_/B _5180_/C _5179_/X VGND VGND VPWR VPWR _5180_/X sky130_fd_sc_hd__or4b_2
X_4131_ _5289_/A0 _4131_/A1 _4135_/S VGND VGND VPWR VPWR _4131_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4062_ _5289_/A0 _4062_/A1 _4066_/S VGND VGND VPWR VPWR _4062_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4964_ _4536_/B _4959_/X _4906_/C VGND VGND VPWR VPWR _5174_/D sky130_fd_sc_hd__a21o_2
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6703_ _7220_/CLK _6703_/D _6362_/B VGND VGND VPWR VPWR _6703_/Q sky130_fd_sc_hd__dfrtp_2
X_3915_ _6360_/A _3915_/B VGND VGND VPWR VPWR _3916_/B sky130_fd_sc_hd__or2_1
XFILLER_177_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4895_ _4987_/A _4409_/Y _4736_/B _4748_/B VGND VGND VPWR VPWR _5129_/A sky130_fd_sc_hd__a22o_2
XFILLER_149_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6634_ _6786_/CLK _6634_/D fanout417/X VGND VGND VPWR VPWR _6634_/Q sky130_fd_sc_hd__dfrtp_2
X_3846_ _3196_/Y _6665_/Q _3201_/Y _3859_/B _6475_/Q VGND VGND VPWR VPWR _6475_/D
+ sky130_fd_sc_hd__a41o_1
XFILLER_164_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6565_ _6616_/CLK _6565_/D fanout439/X VGND VGND VPWR VPWR _6565_/Q sky130_fd_sc_hd__dfstp_2
X_3777_ _7077_/Q _5513_/A _4178_/A _6644_/Q VGND VGND VPWR VPWR _3777_/X sky130_fd_sc_hd__a22o_2
X_5516_ hold43/X hold157/X _5521_/S VGND VGND VPWR VPWR _5516_/X sky130_fd_sc_hd__mux2_1
X_6496_ _6810_/CLK _6496_/D fanout419/X VGND VGND VPWR VPWR _6496_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_145_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5447_ _5582_/A0 hold632/X _5449_/S VGND VGND VPWR VPWR _5447_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5378_ _5378_/A _5594_/B VGND VGND VPWR VPWR _5378_/Y sky130_fd_sc_hd__nand2_8
X_7117_ _7141_/CLK _7117_/D fanout447/X VGND VGND VPWR VPWR _7117_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_113_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4329_ _5234_/C _4329_/A1 _4333_/S VGND VGND VPWR VPWR _4329_/X sky130_fd_sc_hd__mux2_1
X_7048_ _7123_/CLK _7048_/D fanout434/X VGND VGND VPWR VPWR _7048_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_101_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3700_ _6551_/Q _4067_/A _4196_/A _6660_/Q VGND VGND VPWR VPWR _3700_/X sky130_fd_sc_hd__a22o_1
X_4680_ _5099_/A _5024_/A _4680_/C _4670_/X VGND VGND VPWR VPWR _4708_/D sky130_fd_sc_hd__or4b_1
XFILLER_41_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3631_ _6903_/Q _5315_/A _5279_/A _6871_/Q _3611_/X VGND VGND VPWR VPWR _3635_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6350_ _6544_/Q _6023_/C _6025_/B _6567_/Q _6349_/X VGND VGND VPWR VPWR _6355_/B
+ sky130_fd_sc_hd__a221o_1
X_3562_ _6652_/Q _4184_/A _4286_/A _6741_/Q VGND VGND VPWR VPWR _3562_/X sky130_fd_sc_hd__a22o_4
X_5301_ _5571_/A0 hold572/X _5305_/S VGND VGND VPWR VPWR _6888_/D sky130_fd_sc_hd__mux2_1
X_6281_ _6281_/A _6281_/B _6281_/C _6281_/D VGND VGND VPWR VPWR _6282_/C sky130_fd_sc_hd__or4_1
X_3493_ _3506_/A _3543_/B VGND VGND VPWR VPWR _4274_/A sky130_fd_sc_hd__nor2_8
XFILLER_142_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5232_ _5583_/A0 hold672/X _5233_/S VGND VGND VPWR VPWR _5232_/X sky130_fd_sc_hd__mux2_1
X_5163_ _5163_/A _5163_/B _5163_/C VGND VGND VPWR VPWR _5163_/X sky130_fd_sc_hd__or3_1
XFILLER_111_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4114_ _6408_/A0 hold557/X _4117_/S VGND VGND VPWR VPWR _4114_/X sky130_fd_sc_hd__mux2_1
X_5094_ _4395_/D _4987_/B _4586_/B _5116_/A _4797_/C VGND VGND VPWR VPWR _5095_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4045_ hold899/X _5254_/A0 _4048_/S VGND VGND VPWR VPWR _4045_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5996_ _6012_/A _6037_/C _6032_/C VGND VGND VPWR VPWR _5996_/X sky130_fd_sc_hd__and3_4
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4947_ _4986_/C _4947_/B VGND VGND VPWR VPWR _4959_/A sky130_fd_sc_hd__nand2_8
X_4878_ _4878_/A VGND VGND VPWR VPWR _5130_/A sky130_fd_sc_hd__inv_2
XFILLER_137_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6617_ _6713_/CLK _6617_/D fanout427/X VGND VGND VPWR VPWR _6617_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3829_ _3828_/X _6481_/Q _3840_/S VGND VGND VPWR VPWR _6481_/D sky130_fd_sc_hd__mux2_1
XFILLER_165_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6548_ _6840_/CLK _6548_/D fanout424/X VGND VGND VPWR VPWR _6548_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_180_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6479_ _6668_/CLK _6479_/D _6434_/X VGND VGND VPWR VPWR hold24/A sky130_fd_sc_hd__dfrtp_2
XFILLER_133_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput260 _3962_/A VGND VGND VPWR VPWR pad_flash_io1_oeb sky130_fd_sc_hd__buf_8
Xoutput271 _6798_/Q VGND VGND VPWR VPWR pll_ena sky130_fd_sc_hd__buf_8
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput293 _6498_/Q VGND VGND VPWR VPWR pll_trim[2] sky130_fd_sc_hd__buf_8
Xoutput282 _6811_/Q VGND VGND VPWR VPWR pll_trim[16] sky130_fd_sc_hd__buf_8
XFILLER_87_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5850_ _6859_/Q _5722_/B _5839_/X _5849_/X _6308_/S VGND VGND VPWR VPWR _5850_/X
+ sky130_fd_sc_hd__o221a_2
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4801_ _4758_/C _4719_/X _4789_/X _4800_/X _5078_/A VGND VGND VPWR VPWR _4802_/D
+ sky130_fd_sc_hd__a2111o_1
X_5781_ _7096_/Q _5690_/X _5693_/X _7080_/Q _5780_/X VGND VGND VPWR VPWR _5784_/B
+ sky130_fd_sc_hd__a221o_1
X_4732_ _4562_/B _4812_/C _4723_/X _4727_/Y _4731_/X VGND VGND VPWR VPWR _4732_/X
+ sky130_fd_sc_hd__o2111a_1
X_4663_ _4663_/A _4663_/B VGND VGND VPWR VPWR _4724_/B sky130_fd_sc_hd__or2_4
XFILLER_30_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6402_ _6707_/Q _6402_/A2 _6372_/B _6705_/Q VGND VGND VPWR VPWR _6402_/X sky130_fd_sc_hd__a22o_1
X_3614_ _7151_/Q _5594_/A _3552_/Y _6822_/Q VGND VGND VPWR VPWR _3614_/X sky130_fd_sc_hd__a22o_2
XFILLER_174_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4594_ _4871_/A _4947_/B _4812_/A VGND VGND VPWR VPWR _4595_/B sky130_fd_sc_hd__a21oi_4
XFILLER_134_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold913 _5254_/X VGND VGND VPWR VPWR _6846_/D sky130_fd_sc_hd__bufbuf_16
Xhold902 _5187_/X VGND VGND VPWR VPWR _6786_/D sky130_fd_sc_hd__bufbuf_16
Xhold924 _7053_/Q VGND VGND VPWR VPWR hold924/X sky130_fd_sc_hd__bufbuf_16
XFILLER_162_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold946 _5300_/X VGND VGND VPWR VPWR _6887_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_127_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3545_ _3545_/A1 _4234_/S _4055_/A _6544_/Q _3544_/X VGND VGND VPWR VPWR _3546_/D
+ sky130_fd_sc_hd__a221o_2
Xhold935 _4276_/X VGND VGND VPWR VPWR _6729_/D sky130_fd_sc_hd__bufbuf_16
X_6333_ _5611_/A _7199_/Q _6358_/B1 _6332_/X VGND VGND VPWR VPWR _6333_/X sky130_fd_sc_hd__a211o_1
Xhold957 _4242_/X VGND VGND VPWR VPWR _6690_/D sky130_fd_sc_hd__bufbuf_16
Xhold979 _6616_/Q VGND VGND VPWR VPWR hold979/X sky130_fd_sc_hd__bufbuf_16
Xhold968 _6631_/Q VGND VGND VPWR VPWR hold968/X sky130_fd_sc_hd__bufbuf_16
XFILLER_135_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6264_ _6749_/Q _6036_/Y _6335_/B _6774_/Q _6261_/X VGND VGND VPWR VPWR _6269_/B
+ sky130_fd_sc_hd__a221o_1
X_3476_ _3476_/A _5234_/B VGND VGND VPWR VPWR _3476_/Y sky130_fd_sc_hd__nor2_4
XFILLER_130_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5215_ hold417/X _5584_/A0 _5215_/S VGND VGND VPWR VPWR _6818_/D sky130_fd_sc_hd__mux2_1
X_6195_ _7115_/Q _6027_/B _6021_/B _7155_/Q VGND VGND VPWR VPWR _6195_/X sky130_fd_sc_hd__a22o_1
X_5146_ _5146_/A _5146_/B VGND VGND VPWR VPWR _5146_/Y sky130_fd_sc_hd__nor2_1
XFILLER_151_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5077_ _5121_/A _5121_/B VGND VGND VPWR VPWR _5077_/Y sky130_fd_sc_hd__nor2_1
XFILLER_84_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4028_ _5597_/A0 hold509/X _4033_/S VGND VGND VPWR VPWR _4028_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5979_ _6752_/Q _5682_/X _5703_/X _6544_/Q VGND VGND VPWR VPWR _5979_/X sky130_fd_sc_hd__a22o_1
XFILLER_100_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold209 hold209/A VGND VGND VPWR VPWR hold209/X sky130_fd_sc_hd__bufbuf_16
XFILLER_125_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3330_ _6972_/Q _5387_/A _4217_/S input51/X _3326_/X VGND VGND VPWR VPWR _3331_/D
+ sky130_fd_sc_hd__a221o_4
XFILLER_140_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _5121_/B _5081_/C _5000_/C _5136_/D VGND VGND VPWR VPWR _5001_/D sky130_fd_sc_hd__or4_1
XFILLER_112_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3261_ hold24/X hold16/X _3845_/A VGND VGND VPWR VPWR hold25/A sky130_fd_sc_hd__mux2_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3192_ _6459_/Q VGND VGND VPWR VPWR _3192_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6951_ _6951_/CLK _6951_/D fanout442/X VGND VGND VPWR VPWR _6951_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_19_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6882_ _7130_/CLK _6882_/D fanout453/X VGND VGND VPWR VPWR _6882_/Q sky130_fd_sc_hd__dfrtp_2
X_5902_ _6729_/Q _5667_/X _5687_/X _6640_/Q VGND VGND VPWR VPWR _5902_/X sky130_fd_sc_hd__a22o_1
X_5833_ _6915_/Q _5680_/X _5700_/X _6867_/Q VGND VGND VPWR VPWR _5833_/X sky130_fd_sc_hd__a22o_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5764_ _6855_/Q _5722_/B _5753_/X _5763_/X _6308_/S VGND VGND VPWR VPWR _5764_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_187_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4715_ _4453_/Y _4758_/B _4695_/X _5166_/A VGND VGND VPWR VPWR _4797_/B sky130_fd_sc_hd__a31o_1
X_5695_ _7077_/Q _5693_/X _5694_/X _6893_/Q VGND VGND VPWR VPWR _5695_/X sky130_fd_sc_hd__a22o_1
X_4646_ _4774_/A _4774_/C VGND VGND VPWR VPWR _4707_/A sky130_fd_sc_hd__or2_2
XFILLER_190_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4577_ _4818_/B _4740_/B VGND VGND VPWR VPWR _4748_/A sky130_fd_sc_hd__nor2_8
XFILLER_163_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold710 _6946_/Q VGND VGND VPWR VPWR hold710/X sky130_fd_sc_hd__bufbuf_16
Xhold721 _7051_/Q VGND VGND VPWR VPWR hold721/X sky130_fd_sc_hd__bufbuf_16
Xhold743 _4260_/X VGND VGND VPWR VPWR _6716_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold732 _4195_/X VGND VGND VPWR VPWR _6658_/D sky130_fd_sc_hd__bufbuf_16
Xhold754 _6638_/Q VGND VGND VPWR VPWR hold754/X sky130_fd_sc_hd__bufbuf_16
X_6316_ _6751_/Q _6036_/Y _6335_/B _6776_/Q _6311_/X VGND VGND VPWR VPWR _6321_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold776 _7031_/Q VGND VGND VPWR VPWR hold776/X sky130_fd_sc_hd__bufbuf_16
Xhold765 _7074_/Q VGND VGND VPWR VPWR hold765/X sky130_fd_sc_hd__bufbuf_16
X_3528_ _5252_/A _3528_/B VGND VGND VPWR VPWR _4160_/A sky130_fd_sc_hd__nor2_8
Xhold787 _6809_/Q VGND VGND VPWR VPWR hold787/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6247_ _6247_/A _6247_/B _6247_/C _6247_/D VGND VGND VPWR VPWR _6248_/C sky130_fd_sc_hd__or4_1
XFILLER_103_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold798 _6761_/Q VGND VGND VPWR VPWR hold798/X sky130_fd_sc_hd__bufbuf_16
X_3459_ _3501_/A _5252_/B VGND VGND VPWR VPWR _4316_/A sky130_fd_sc_hd__nor2_8
X_6178_ _7106_/Q _5653_/X _6022_/B _6946_/Q VGND VGND VPWR VPWR _6178_/X sky130_fd_sc_hd__a22o_4
X_5129_ _5129_/A _5129_/B _5123_/C _5123_/B VGND VGND VPWR VPWR _5130_/C sky130_fd_sc_hd__or4bb_1
XFILLER_85_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold70 hold70/A VGND VGND VPWR VPWR hold70/X sky130_fd_sc_hd__bufbuf_16
XFILLER_76_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold81 hold81/A VGND VGND VPWR VPWR hold81/X sky130_fd_sc_hd__bufbuf_16
XFILLER_36_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold92 hold92/A VGND VGND VPWR VPWR hold92/X sky130_fd_sc_hd__bufbuf_16
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4500_ _4500_/A _4586_/B VGND VGND VPWR VPWR _5116_/A sky130_fd_sc_hd__and2_2
X_5480_ hold702/X _5561_/A0 _5485_/S VGND VGND VPWR VPWR _5480_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4431_ _4992_/A _4851_/B _4499_/C _4507_/A VGND VGND VPWR VPWR _4539_/D sky130_fd_sc_hd__o211a_2
XFILLER_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1 _6482_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7150_ _7150_/CLK _7150_/D fanout444/X VGND VGND VPWR VPWR _7150_/Q sky130_fd_sc_hd__dfstp_2
X_4362_ _5050_/A _4413_/C VGND VGND VPWR VPWR _4364_/A sky130_fd_sc_hd__nor2_2
XFILLER_125_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4293_ _5289_/A0 _4293_/A1 _4297_/S VGND VGND VPWR VPWR _4293_/X sky130_fd_sc_hd__mux2_1
X_3313_ _6964_/Q _5378_/A _5342_/A _6932_/Q _3312_/X VGND VGND VPWR VPWR _3331_/B
+ sky130_fd_sc_hd__a221o_4
X_6101_ _6903_/Q _6021_/A _6025_/A _6935_/Q _6100_/X VGND VGND VPWR VPWR _6106_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_140_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7081_ _7081_/CLK _7081_/D fanout437/X VGND VGND VPWR VPWR _7081_/Q sky130_fd_sc_hd__dfrtp_2
X_3244_ _4469_/A VGND VGND VPWR VPWR _4740_/A sky130_fd_sc_hd__inv_8
X_6032_ _6032_/A _6037_/C _6032_/C VGND VGND VPWR VPWR _6032_/X sky130_fd_sc_hd__and3_4
XFILLER_98_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6934_ _7151_/CLK _6934_/D fanout447/X VGND VGND VPWR VPWR _6934_/Q sky130_fd_sc_hd__dfstp_4
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6865_ _7127_/CLK _6865_/D fanout449/X VGND VGND VPWR VPWR _6865_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5816_ _7098_/Q _5690_/X _5693_/X _7082_/Q _5815_/X VGND VGND VPWR VPWR _5827_/B
+ sky130_fd_sc_hd__a221o_2
X_6796_ _3545_/A1 _6796_/D _6454_/X VGND VGND VPWR VPWR _6796_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_148_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5747_ _6991_/Q _5684_/X _5692_/X _7071_/Q VGND VGND VPWR VPWR _5747_/X sky130_fd_sc_hd__a22o_1
XFILLER_157_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5678_ _7165_/Q _5705_/B _5703_/B VGND VGND VPWR VPWR _5678_/X sky130_fd_sc_hd__and3_4
XFILLER_135_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4629_ _4996_/A _4749_/C VGND VGND VPWR VPWR _5079_/B sky130_fd_sc_hd__nor2_2
Xhold540 _5304_/X VGND VGND VPWR VPWR _6891_/D sky130_fd_sc_hd__bufbuf_16
Xhold551 _5390_/X VGND VGND VPWR VPWR _6967_/D sky130_fd_sc_hd__bufbuf_16
Xhold562 _6954_/Q VGND VGND VPWR VPWR hold562/X sky130_fd_sc_hd__bufbuf_16
XFILLER_116_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold584 _7112_/Q VGND VGND VPWR VPWR hold584/X sky130_fd_sc_hd__bufbuf_16
Xhold573 _6912_/Q VGND VGND VPWR VPWR hold573/X sky130_fd_sc_hd__bufbuf_16
XFILLER_143_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold595 _6630_/Q VGND VGND VPWR VPWR hold595/X sky130_fd_sc_hd__bufbuf_16
XFILLER_1_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1240 _6673_/Q VGND VGND VPWR VPWR _4212_/A0 sky130_fd_sc_hd__bufbuf_16
XFILLER_92_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1251 _7095_/Q VGND VGND VPWR VPWR _5534_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_66_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1262 _6943_/Q VGND VGND VPWR VPWR _5363_/A1 sky130_fd_sc_hd__bufbuf_16
XANTENNA_435 hold165/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_402 _6917_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_413 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_424 _5582_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_457 _6011_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_446 hold739/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_468 _5541_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_479 _6407_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput160 wb_dat_i[6] VGND VGND VPWR VPWR _6396_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4980_ _4980_/A _4980_/B _4980_/C _4367_/X VGND VGND VPWR VPWR _5121_/A sky130_fd_sc_hd__or4b_4
XFILLER_91_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3931_ _3203_/Y input92/X _3932_/S VGND VGND VPWR VPWR _3931_/X sky130_fd_sc_hd__mux2_8
XFILLER_32_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6650_ _6715_/CLK _6650_/D fanout439/X VGND VGND VPWR VPWR _6650_/Q sky130_fd_sc_hd__dfrtp_2
X_3862_ _6469_/Q _3866_/B _3864_/B VGND VGND VPWR VPWR _3862_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_32_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5601_ _5601_/A0 hold603/X _5602_/S VGND VGND VPWR VPWR _5601_/X sky130_fd_sc_hd__mux2_1
X_6581_ _7220_/CLK _6581_/D VGND VGND VPWR VPWR _6581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5532_ _5541_/A0 _5532_/A1 _5539_/S VGND VGND VPWR VPWR _7093_/D sky130_fd_sc_hd__mux2_1
X_3793_ _3793_/A _3793_/B _3793_/C _3793_/D VGND VGND VPWR VPWR _3794_/D sky130_fd_sc_hd__or4_4
XFILLER_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5463_ hold136/X hold240/X _5467_/S VGND VGND VPWR VPWR _5463_/X sky130_fd_sc_hd__mux2_1
X_4414_ _4529_/B _4414_/B VGND VGND VPWR VPWR _4416_/B sky130_fd_sc_hd__nand2_8
X_5394_ _5601_/A0 hold746/X _5395_/S VGND VGND VPWR VPWR _5394_/X sky130_fd_sc_hd__mux2_1
X_7202_ _7220_/CLK _7202_/D _6362_/B VGND VGND VPWR VPWR _7202_/Q sky130_fd_sc_hd__dfrtp_2
X_4345_ _4345_/A _4345_/B VGND VGND VPWR VPWR _4345_/Y sky130_fd_sc_hd__nand2_1
X_7133_ _7133_/CLK _7133_/D fanout443/X VGND VGND VPWR VPWR _7133_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_99_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7064_ _7152_/CLK _7064_/D fanout454/X VGND VGND VPWR VPWR _7064_/Q sky130_fd_sc_hd__dfrtp_2
X_4276_ _5254_/A0 hold934/X _4279_/S VGND VGND VPWR VPWR _4276_/X sky130_fd_sc_hd__mux2_1
X_3227_ _6960_/Q VGND VGND VPWR VPWR _3227_/Y sky130_fd_sc_hd__inv_2
X_6015_ _6037_/B _6018_/A _6032_/C VGND VGND VPWR VPWR _6022_/B sky130_fd_sc_hd__and3_4
XFILLER_86_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6917_ _7127_/CLK _6917_/D fanout447/X VGND VGND VPWR VPWR _6917_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_167_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6848_ _7107_/CLK _6848_/D fanout434/X VGND VGND VPWR VPWR _6848_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_52_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6779_ _7208_/CLK _6779_/D _6362_/B VGND VGND VPWR VPWR _6779_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_182_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold370 _6988_/Q VGND VGND VPWR VPWR hold370/X sky130_fd_sc_hd__bufbuf_16
Xhold381 _5431_/X VGND VGND VPWR VPWR _7004_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_151_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold392 _6862_/Q VGND VGND VPWR VPWR hold392/X sky130_fd_sc_hd__bufbuf_16
XFILLER_65_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1070 _4269_/X VGND VGND VPWR VPWR _6723_/D sky130_fd_sc_hd__bufbuf_16
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1092 _7101_/Q VGND VGND VPWR VPWR _5541_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1081 _6682_/Q VGND VGND VPWR VPWR _4223_/A0 sky130_fd_sc_hd__bufbuf_16
XFILLER_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_210 _7064_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_221 _6918_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_232 _6459_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_243 mask_rev_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_265 wb_adr_i[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_276 wb_adr_i[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_254 pad_flash_io0_di VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_287 wb_dat_i[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_298 _3972_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4130_ _4130_/A hold47/X VGND VGND VPWR VPWR _4135_/S sky130_fd_sc_hd__nand2_8
XFILLER_110_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4061_ _4061_/A _5558_/B VGND VGND VPWR VPWR _4066_/S sky130_fd_sc_hd__nand2_8
XFILLER_68_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4963_ _4971_/B VGND VGND VPWR VPWR _4963_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6702_ _7220_/CLK _6702_/D _6362_/B VGND VGND VPWR VPWR _6702_/Q sky130_fd_sc_hd__dfrtp_2
X_3914_ _6706_/Q _3883_/X _6701_/Q VGND VGND VPWR VPWR _6706_/D sky130_fd_sc_hd__a21o_1
XFILLER_149_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4894_ _4956_/C _4689_/Y _4617_/Y VGND VGND VPWR VPWR _4906_/C sky130_fd_sc_hd__a21o_1
X_6633_ _6746_/CLK _6633_/D fanout427/X VGND VGND VPWR VPWR _6633_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_177_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3845_ _3845_/A _6664_/Q VGND VGND VPWR VPWR _3859_/B sky130_fd_sc_hd__nor2_8
XFILLER_192_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6564_ _6715_/CLK _6564_/D fanout439/X VGND VGND VPWR VPWR _6564_/Q sky130_fd_sc_hd__dfrtp_2
X_3776_ _6800_/Q _5194_/A _3771_/X _3773_/X _3775_/X VGND VGND VPWR VPWR _3793_/B
+ sky130_fd_sc_hd__a2111o_1
X_6495_ _7129_/CLK _6495_/D fanout429/X VGND VGND VPWR VPWR _6495_/Q sky130_fd_sc_hd__dfstp_4
X_5515_ _5578_/A0 hold415/X _5521_/S VGND VGND VPWR VPWR _5515_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5446_ hold185/X hold189/X _5449_/S VGND VGND VPWR VPWR _5446_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5377_ _5602_/A0 hold499/X _5377_/S VGND VGND VPWR VPWR _5377_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7116_ _7152_/CLK hold15/X fanout447/X VGND VGND VPWR VPWR _7116_/Q sky130_fd_sc_hd__dfrtp_2
X_4328_ _4328_/A hold47/X VGND VGND VPWR VPWR _4333_/S sky130_fd_sc_hd__nand2_4
XFILLER_113_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4259_ hold867/X _5300_/A0 _4261_/S VGND VGND VPWR VPWR _6715_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7047_ _7135_/CLK _7047_/D fanout429/X VGND VGND VPWR VPWR _7047_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_101_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_74_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7225_/CLK sky130_fd_sc_hd__clkbuf_8
X_3630_ _6927_/Q _5342_/A _4136_/A _6611_/Q _3618_/X VGND VGND VPWR VPWR _3635_/A
+ sky130_fd_sc_hd__a221o_1
X_3561_ _6992_/Q _3299_/Y _3334_/Y _7040_/Q VGND VGND VPWR VPWR _3561_/X sky130_fd_sc_hd__a22o_1
X_5300_ _5300_/A0 hold945/X _5305_/S VGND VGND VPWR VPWR _5300_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3492_ _6889_/Q _5297_/A _5185_/A _6789_/Q _3490_/X VGND VGND VPWR VPWR _3504_/A
+ sky130_fd_sc_hd__a221o_4
X_6280_ _6714_/Q _6023_/B _6021_/C _6546_/Q _6279_/X VGND VGND VPWR VPWR _6281_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5231_ _5582_/A0 hold575/X _5233_/S VGND VGND VPWR VPWR _5231_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5162_ _5164_/A _4636_/A _4664_/X VGND VGND VPWR VPWR _5163_/C sky130_fd_sc_hd__o21ai_1
XFILLER_96_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5093_ _5061_/Y _5076_/X _5092_/X _5059_/X VGND VGND VPWR VPWR _6781_/D sky130_fd_sc_hd__a211o_1
X_4113_ _5289_/A0 _4113_/A1 _4117_/S VGND VGND VPWR VPWR _4113_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_12_csclk clkbuf_opt_4_0_csclk/X VGND VGND VPWR VPWR _6715_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_111_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4044_ _4044_/A0 _5234_/C _4048_/S VGND VGND VPWR VPWR _4044_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_27_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7111_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5995_ _7168_/Q _7169_/Q VGND VGND VPWR VPWR _6032_/C sky130_fd_sc_hd__and2b_4
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4946_ _4946_/A _4946_/B VGND VGND VPWR VPWR _4946_/X sky130_fd_sc_hd__or2_1
XFILLER_33_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4877_ _5147_/A _4877_/B VGND VGND VPWR VPWR _4878_/A sky130_fd_sc_hd__or2_2
X_6616_ _6616_/CLK _6616_/D fanout439/X VGND VGND VPWR VPWR _6616_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_138_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3828_ hold58/A _3249_/Y _3828_/S VGND VGND VPWR VPWR _3828_/X sky130_fd_sc_hd__mux2_1
X_6547_ _6649_/CLK _6547_/D fanout439/X VGND VGND VPWR VPWR _6547_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_165_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3759_ _3759_/A _3759_/B _3759_/C _3759_/D VGND VGND VPWR VPWR _3794_/B sky130_fd_sc_hd__or4_1
XFILLER_106_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6478_ _3957_/A1 _6478_/D _6433_/X VGND VGND VPWR VPWR hold16/A sky130_fd_sc_hd__dfrtp_2
XFILLER_160_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput250 _3938_/X VGND VGND VPWR VPWR mgmt_gpio_out[9] sky130_fd_sc_hd__clkbuf_4
Xoutput261 _6808_/Q VGND VGND VPWR VPWR pll90_sel[0] sky130_fd_sc_hd__buf_8
X_5429_ _5582_/A0 hold570/X hold48/X VGND VGND VPWR VPWR _5429_/X sky130_fd_sc_hd__mux2_1
Xoutput294 _6499_/Q VGND VGND VPWR VPWR pll_trim[3] sky130_fd_sc_hd__buf_8
Xoutput272 _6805_/Q VGND VGND VPWR VPWR pll_sel[0] sky130_fd_sc_hd__buf_8
Xoutput283 _6812_/Q VGND VGND VPWR VPWR pll_trim[17] sky130_fd_sc_hd__buf_8
XFILLER_102_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_1_wb_clk_i clkbuf_1_1_1_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_151_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4800_ _4800_/A _4800_/B _4800_/C _4800_/D VGND VGND VPWR VPWR _4800_/X sky130_fd_sc_hd__or4_1
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5780_ _7016_/Q _5682_/X _5703_/X _6872_/Q VGND VGND VPWR VPWR _5780_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4731_ _4898_/B _4756_/B _4728_/X _4947_/B _4730_/X VGND VGND VPWR VPWR _4731_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_187_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4662_ _4663_/A _4663_/B VGND VGND VPWR VPWR _4758_/C sky130_fd_sc_hd__nor2_8
X_3613_ _3875_/B _4234_/S _5558_/A _7119_/Q VGND VGND VPWR VPWR _3613_/X sky130_fd_sc_hd__a22o_4
X_6401_ _6401_/A1 _4237_/X _6376_/A _3916_/A VGND VGND VPWR VPWR _7219_/D sky130_fd_sc_hd__o211a_2
X_4593_ _4593_/A _4693_/B _5087_/C VGND VGND VPWR VPWR _4593_/Y sky130_fd_sc_hd__nand3_2
XFILLER_134_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold903 _6814_/Q VGND VGND VPWR VPWR hold903/X sky130_fd_sc_hd__bufbuf_16
XFILLER_127_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3544_ _6492_/Q _3978_/A _5594_/A _7153_/Q VGND VGND VPWR VPWR _3544_/X sky130_fd_sc_hd__a22o_1
Xhold925 _6737_/Q VGND VGND VPWR VPWR hold925/X sky130_fd_sc_hd__bufbuf_16
Xhold936 _6838_/Q VGND VGND VPWR VPWR hold936/X sky130_fd_sc_hd__bufbuf_16
Xhold914 _6764_/Q VGND VGND VPWR VPWR hold914/X sky130_fd_sc_hd__bufbuf_16
X_6332_ _6533_/Q _6060_/B _6321_/X _6331_/X _6308_/S VGND VGND VPWR VPWR _6332_/X
+ sky130_fd_sc_hd__o221a_2
Xhold947 _6735_/Q VGND VGND VPWR VPWR hold947/X sky130_fd_sc_hd__bufbuf_16
X_3475_ _6881_/Q _5288_/A _5405_/A _6985_/Q _3474_/X VGND VGND VPWR VPWR _3488_/A
+ sky130_fd_sc_hd__a221o_4
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold969 _4163_/X VGND VGND VPWR VPWR _6631_/D sky130_fd_sc_hd__bufbuf_16
Xhold958 _6547_/Q VGND VGND VPWR VPWR hold958/X sky130_fd_sc_hd__bufbuf_16
XFILLER_103_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6263_ _6759_/Q _6010_/Y _6031_/X _6645_/Q _6262_/X VGND VGND VPWR VPWR _6269_/A
+ sky130_fd_sc_hd__a221o_1
X_5214_ hold679/X _5583_/A0 _5215_/S VGND VGND VPWR VPWR _6817_/D sky130_fd_sc_hd__mux2_1
X_6194_ _6194_/A _6194_/B _6194_/C _6194_/D VGND VGND VPWR VPWR _6207_/B sky130_fd_sc_hd__or4_1
X_5145_ _5145_/A _5145_/B _5145_/C _5145_/D VGND VGND VPWR VPWR _5146_/B sky130_fd_sc_hd__or4_2
XFILLER_111_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5076_ _5142_/B _5076_/B _5076_/C _5076_/D VGND VGND VPWR VPWR _5076_/X sky130_fd_sc_hd__or4_2
XFILLER_84_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4027_ _5596_/A0 hold309/X _4033_/S VGND VGND VPWR VPWR _4027_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5978_ _6580_/Q _5689_/X _5967_/X _5977_/X VGND VGND VPWR VPWR _5981_/C sky130_fd_sc_hd__a211o_1
XFILLER_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4929_ _4500_/A _4758_/A _4711_/C _4682_/Y VGND VGND VPWR VPWR _4932_/B sky130_fd_sc_hd__a31o_1
XFILLER_100_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3260_ _3309_/A _3275_/B _3275_/C VGND VGND VPWR VPWR _3260_/X sky130_fd_sc_hd__or3_4
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3191_ hold80/A VGND VGND VPWR VPWR _3191_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6950_ _6951_/CLK _6950_/D fanout442/X VGND VGND VPWR VPWR _6950_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_19_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5901_ _6564_/Q _5694_/X _5706_/X _6650_/Q VGND VGND VPWR VPWR _5901_/X sky130_fd_sc_hd__a22o_2
XFILLER_81_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6881_ _7121_/CLK _6881_/D _6421_/A VGND VGND VPWR VPWR _6881_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_34_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5832_ _7083_/Q _5693_/X _5694_/X _6899_/Q _5831_/X VGND VGND VPWR VPWR _5839_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_62_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5763_ _5763_/A _5763_/B _5763_/C _5763_/D VGND VGND VPWR VPWR _5763_/X sky130_fd_sc_hd__or4_4
X_4714_ _5062_/B _4714_/B VGND VGND VPWR VPWR _5050_/B sky130_fd_sc_hd__or2_1
XFILLER_147_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5694_ _5864_/B _5707_/B _5707_/C VGND VGND VPWR VPWR _5694_/X sky130_fd_sc_hd__and3_4
XFILLER_163_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4645_ _4887_/B _4787_/B _4642_/X _4644_/Y _4567_/X VGND VGND VPWR VPWR _4645_/X
+ sky130_fd_sc_hd__o41a_4
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4576_ _4871_/A _4953_/A VGND VGND VPWR VPWR _4708_/A sky130_fd_sc_hd__nor2_1
XFILLER_146_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold700 _6850_/Q VGND VGND VPWR VPWR hold700/X sky130_fd_sc_hd__bufbuf_16
Xhold711 _5366_/X VGND VGND VPWR VPWR _6946_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_190_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3527_ input48/X _4217_/S _5585_/A _7145_/Q _3526_/X VGND VGND VPWR VPWR _3533_/B
+ sky130_fd_sc_hd__a221o_4
Xhold744 _6643_/Q VGND VGND VPWR VPWR hold744/X sky130_fd_sc_hd__bufbuf_16
Xhold722 _5484_/X VGND VGND VPWR VPWR _7051_/D sky130_fd_sc_hd__bufbuf_16
Xhold755 _4171_/X VGND VGND VPWR VPWR _6638_/D sky130_fd_sc_hd__bufbuf_16
Xhold733 _6789_/Q VGND VGND VPWR VPWR hold733/X sky130_fd_sc_hd__bufbuf_16
X_6315_ _6761_/Q _6010_/Y _6031_/X _6647_/Q _6312_/X VGND VGND VPWR VPWR _6321_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold777 _5462_/X VGND VGND VPWR VPWR _7031_/D sky130_fd_sc_hd__bufbuf_16
Xhold766 _5510_/X VGND VGND VPWR VPWR _7074_/D sky130_fd_sc_hd__bufbuf_16
Xhold788 _6732_/Q VGND VGND VPWR VPWR hold788/X sky130_fd_sc_hd__bufbuf_16
XFILLER_162_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6246_ _6545_/Q _6021_/C _6031_/X _6644_/Q _6245_/X VGND VGND VPWR VPWR _6247_/D
+ sky130_fd_sc_hd__a221o_1
X_3458_ _7001_/Q _5423_/A _4154_/A _6628_/Q _3456_/X VGND VGND VPWR VPWR _3472_/A
+ sky130_fd_sc_hd__a221o_1
Xhold799 _4314_/X VGND VGND VPWR VPWR _6761_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_190_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6177_ _6874_/Q _6023_/C _6025_/B _6898_/Q _6176_/X VGND VGND VPWR VPWR _6181_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_85_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3389_ input32/X _3283_/Y _5477_/A _7051_/Q VGND VGND VPWR VPWR _3389_/X sky130_fd_sc_hd__a22o_1
X_5128_ _5128_/A _5128_/B _5128_/C _5128_/D VGND VGND VPWR VPWR _5143_/A sky130_fd_sc_hd__or4_4
XFILLER_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5059_ _4935_/D _5102_/C _5102_/D _5036_/X _5058_/X VGND VGND VPWR VPWR _5059_/X
+ sky130_fd_sc_hd__a41o_1
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold71 hold71/A VGND VGND VPWR VPWR hold71/X sky130_fd_sc_hd__bufbuf_16
Xhold82 hold82/A VGND VGND VPWR VPWR hold82/X sky130_fd_sc_hd__bufbuf_16
Xhold60 hold60/A VGND VGND VPWR VPWR hold60/X sky130_fd_sc_hd__bufbuf_16
Xhold93 hold93/A VGND VGND VPWR VPWR hold93/X sky130_fd_sc_hd__bufbuf_16
XFILLER_188_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4430_ _4507_/A _4500_/A _4851_/B _4499_/C VGND VGND VPWR VPWR _5140_/B sky130_fd_sc_hd__and4_2
XANTENNA_2 _6483_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4361_ _4566_/A _4558_/B VGND VGND VPWR VPWR _4986_/A sky130_fd_sc_hd__or2_4
XFILLER_160_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6100_ _6951_/Q _6022_/A _6025_/C _6927_/Q VGND VGND VPWR VPWR _6100_/X sky130_fd_sc_hd__a22o_1
XFILLER_125_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4292_ _4292_/A _5558_/B VGND VGND VPWR VPWR _4297_/S sky130_fd_sc_hd__nand2_8
X_3312_ input42/X _4023_/S hold85/A _7116_/Q VGND VGND VPWR VPWR _3312_/X sky130_fd_sc_hd__a22o_1
XFILLER_112_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7080_ _7097_/CLK _7080_/D fanout437/X VGND VGND VPWR VPWR _7080_/Q sky130_fd_sc_hd__dfrtp_2
X_3243_ _4672_/A VGND VGND VPWR VPWR _4735_/B sky130_fd_sc_hd__clkinv_4
XFILLER_112_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6031_ _6032_/A _6035_/A _6037_/C VGND VGND VPWR VPWR _6031_/X sky130_fd_sc_hd__and3_4
XFILLER_100_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6933_ _7054_/CLK _6933_/D fanout445/X VGND VGND VPWR VPWR _6933_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6864_ _7152_/CLK _6864_/D fanout452/X VGND VGND VPWR VPWR _6864_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5815_ _7018_/Q _5682_/X _5703_/X _6874_/Q VGND VGND VPWR VPWR _5815_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6795_ _3545_/A1 _6795_/D _6453_/X VGND VGND VPWR VPWR _6795_/Q sky130_fd_sc_hd__dfrtn_1
X_5746_ _7103_/Q _5675_/X _5701_/X _6951_/Q _5745_/X VGND VGND VPWR VPWR _5753_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_41_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5677_ _7101_/Q _5675_/X _5676_/X _6973_/Q VGND VGND VPWR VPWR _5677_/X sky130_fd_sc_hd__a22o_1
XFILLER_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4628_ _4995_/A _4989_/A VGND VGND VPWR VPWR _4628_/Y sky130_fd_sc_hd__nor2_1
XFILLER_163_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold530 _5323_/X VGND VGND VPWR VPWR _6908_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_190_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold552 _6898_/Q VGND VGND VPWR VPWR hold552/X sky130_fd_sc_hd__bufbuf_16
X_4559_ _4808_/A _5013_/A _4559_/C _4558_/X VGND VGND VPWR VPWR _4559_/X sky130_fd_sc_hd__or4b_2
XFILLER_151_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold563 _5375_/X VGND VGND VPWR VPWR _6954_/D sky130_fd_sc_hd__bufbuf_16
Xhold541 _6841_/Q VGND VGND VPWR VPWR hold541/X sky130_fd_sc_hd__bufbuf_16
XFILLER_116_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold574 _5328_/X VGND VGND VPWR VPWR _6912_/D sky130_fd_sc_hd__bufbuf_16
Xhold585 _6915_/Q VGND VGND VPWR VPWR hold585/X sky130_fd_sc_hd__bufbuf_16
XFILLER_104_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold596 _4162_/X VGND VGND VPWR VPWR _6630_/D sky130_fd_sc_hd__bufbuf_16
X_6229_ _7068_/Q _5996_/X _6020_/C _6916_/Q VGND VGND VPWR VPWR _6229_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1252 _6964_/Q VGND VGND VPWR VPWR _5386_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1241 _7108_/Q VGND VGND VPWR VPWR _5548_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_58_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1230 _6530_/Q VGND VGND VPWR VPWR _4044_/A0 sky130_fd_sc_hd__bufbuf_16
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1263 _7023_/Q VGND VGND VPWR VPWR _5453_/A1 sky130_fd_sc_hd__bufbuf_16
XANTENNA_425 _5600_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_414 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_403 _6482_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_447 hold874/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_458 _6022_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_436 hold185/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_469 _5611_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput150 wb_dat_i[26] VGND VGND VPWR VPWR _6384_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput161 wb_dat_i[7] VGND VGND VPWR VPWR _6399_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3930_ _6843_/Q input89/X _3932_/S VGND VGND VPWR VPWR _3930_/X sky130_fd_sc_hd__mux2_8
XFILLER_91_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3861_ _6467_/Q _3861_/B VGND VGND VPWR VPWR _3866_/B sky130_fd_sc_hd__nor2_2
XFILLER_176_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5600_ _5600_/A0 hold464/X _5602_/S VGND VGND VPWR VPWR _5600_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6580_ _6717_/CLK _6580_/D fanout426/X VGND VGND VPWR VPWR _6580_/Q sky130_fd_sc_hd__dfrtp_2
X_3792_ _3792_/A _3792_/B _3792_/C _3792_/D VGND VGND VPWR VPWR _3793_/D sky130_fd_sc_hd__or4_1
XFILLER_191_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5531_ _5531_/A _5576_/B VGND VGND VPWR VPWR _5539_/S sky130_fd_sc_hd__nand2_8
XFILLER_191_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5462_ _5561_/A0 hold776/X _5467_/S VGND VGND VPWR VPWR _5462_/X sky130_fd_sc_hd__mux2_1
X_7201_ _7201_/CLK _7201_/D fanout419/X VGND VGND VPWR VPWR _7201_/Q sky130_fd_sc_hd__dfrtp_2
X_4413_ _4672_/A _4696_/A _4413_/C _4436_/B VGND VGND VPWR VPWR _4414_/B sky130_fd_sc_hd__and4_4
X_5393_ _5600_/A0 hold476/X _5395_/S VGND VGND VPWR VPWR _5393_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4344_ _4408_/B _4408_/A VGND VGND VPWR VPWR _4553_/A sky130_fd_sc_hd__nand2b_4
XFILLER_141_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7132_ _7132_/CLK _7132_/D fanout432/X VGND VGND VPWR VPWR _7132_/Q sky130_fd_sc_hd__dfrtp_2
X_7063_ _7127_/CLK _7063_/D fanout449/X VGND VGND VPWR VPWR _7063_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_140_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6014_ _6014_/A _6034_/B VGND VGND VPWR VPWR _6025_/D sky130_fd_sc_hd__nor2_8
X_4275_ _5234_/C _4275_/A1 _4279_/S VGND VGND VPWR VPWR _4275_/X sky130_fd_sc_hd__mux2_1
X_3226_ _6968_/Q VGND VGND VPWR VPWR _3226_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6916_ _7156_/CLK _6916_/D fanout447/X VGND VGND VPWR VPWR _6916_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_42_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6847_ _7107_/CLK _6847_/D fanout434/X VGND VGND VPWR VPWR _6847_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6778_ _7208_/CLK _6778_/D _6362_/B VGND VGND VPWR VPWR _6778_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5729_ _6958_/Q _5673_/X _5681_/X _6918_/Q _5728_/X VGND VGND VPWR VPWR _5734_/B
+ sky130_fd_sc_hd__a221o_4
XFILLER_136_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold371 _5413_/X VGND VGND VPWR VPWR _6988_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_163_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold360 _7094_/Q VGND VGND VPWR VPWR hold360/X sky130_fd_sc_hd__bufbuf_16
Xhold393 _6882_/Q VGND VGND VPWR VPWR hold393/X sky130_fd_sc_hd__bufbuf_16
Xhold382 _6958_/Q VGND VGND VPWR VPWR hold382/X sky130_fd_sc_hd__bufbuf_16
XFILLER_117_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1060 _6802_/Q VGND VGND VPWR VPWR _5197_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1093 _6624_/Q VGND VGND VPWR VPWR _4155_/A0 sky130_fd_sc_hd__bufbuf_16
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_200 _6750_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1071 _6997_/Q VGND VGND VPWR VPWR _5424_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1082 _4223_/X VGND VGND VPWR VPWR _6682_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_211 _6658_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_222 hold80/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_233 mask_rev_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_266 wb_adr_i[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_277 wb_clk_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_255 pad_flash_io1_di VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_244 mask_rev_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_299 _7229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_288 wb_dat_i[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4060_ _5545_/A0 _4060_/A1 _4060_/S VGND VGND VPWR VPWR _4060_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4962_ _4962_/A _4962_/B VGND VGND VPWR VPWR _4971_/B sky130_fd_sc_hd__or2_2
X_4893_ _4893_/A _4893_/B VGND VGND VPWR VPWR _4906_/B sky130_fd_sc_hd__nand2_4
X_6701_ _7220_/CLK _6701_/D _6362_/B VGND VGND VPWR VPWR _6701_/Q sky130_fd_sc_hd__dfrtp_2
X_3913_ _6705_/Q _3883_/X _6700_/Q VGND VGND VPWR VPWR _6705_/D sky130_fd_sc_hd__a21o_1
X_6632_ _6833_/CLK _6632_/D fanout456/X VGND VGND VPWR VPWR _6632_/Q sky130_fd_sc_hd__dfstp_4
X_3844_ _6457_/Q _6476_/Q _3924_/C VGND VGND VPWR VPWR _6476_/D sky130_fd_sc_hd__mux2_1
XFILLER_149_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6563_ _6629_/CLK _6563_/D fanout439/X VGND VGND VPWR VPWR _6563_/Q sky130_fd_sc_hd__dfrtp_2
X_3775_ _7069_/Q hold92/A _4190_/A _6654_/Q _3774_/X VGND VGND VPWR VPWR _3775_/X
+ sky130_fd_sc_hd__a221o_4
X_5514_ _5541_/A0 _5514_/A1 _5521_/S VGND VGND VPWR VPWR _7077_/D sky130_fd_sc_hd__mux2_1
X_6494_ _7129_/CLK _6494_/D fanout428/X VGND VGND VPWR VPWR _6494_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_173_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5445_ hold136/X _7016_/Q _5449_/S VGND VGND VPWR VPWR _5445_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7115_ _7154_/CLK _7115_/D fanout451/X VGND VGND VPWR VPWR _7115_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_154_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5376_ _5601_/A0 hold752/X _5377_/S VGND VGND VPWR VPWR _5376_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4327_ _6411_/A0 hold790/X _4327_/S VGND VGND VPWR VPWR _4327_/X sky130_fd_sc_hd__mux2_1
X_4258_ hold527/X _6408_/A0 _4261_/S VGND VGND VPWR VPWR _4258_/X sky130_fd_sc_hd__mux2_1
X_7046_ _7078_/CLK _7046_/D fanout431/X VGND VGND VPWR VPWR _7046_/Q sky130_fd_sc_hd__dfstp_4
X_3209_ _7104_/Q VGND VGND VPWR VPWR _3209_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4189_ _4189_/A0 _5545_/A0 _4189_/S VGND VGND VPWR VPWR _4189_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold190 _5446_/X VGND VGND VPWR VPWR _7017_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_120_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_8_csclk _6722_/CLK VGND VGND VPWR VPWR _6746_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_160_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3560_ _7008_/Q _5432_/A _3368_/Y input14/X VGND VGND VPWR VPWR _3560_/X sky130_fd_sc_hd__a22o_2
XFILLER_161_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5230_ _5561_/A0 hold704/X _5233_/S VGND VGND VPWR VPWR _5230_/X sky130_fd_sc_hd__mux2_1
X_3491_ hold53/X _3732_/B VGND VGND VPWR VPWR _5185_/A sky130_fd_sc_hd__nor2_8
XFILLER_130_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5161_ _4940_/B _5101_/C _5161_/C _5161_/D VGND VGND VPWR VPWR _5161_/X sky130_fd_sc_hd__and4bb_2
XFILLER_123_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5092_ _5083_/X _5091_/X _5077_/Y VGND VGND VPWR VPWR _5092_/X sky130_fd_sc_hd__o21a_1
X_4112_ _4112_/A _5558_/B VGND VGND VPWR VPWR _4117_/S sky130_fd_sc_hd__nand2_8
XFILLER_96_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4043_ _4043_/A _6406_/B VGND VGND VPWR VPWR _4048_/S sky130_fd_sc_hd__and2_4
XFILLER_49_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5994_ _6030_/A _6014_/A VGND VGND VPWR VPWR _6021_/A sky130_fd_sc_hd__nor2_8
XFILLER_52_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4945_ _5095_/B _5022_/D _5180_/B _4945_/D VGND VGND VPWR VPWR _4946_/B sky130_fd_sc_hd__or4_1
XFILLER_178_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4876_ _4989_/A _4970_/B _4898_/B _5147_/B VGND VGND VPWR VPWR _4877_/B sky130_fd_sc_hd__o22a_1
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6615_ _6715_/CLK _6615_/D fanout439/X VGND VGND VPWR VPWR _6615_/Q sky130_fd_sc_hd__dfrtp_2
X_3827_ _3845_/A _3830_/B VGND VGND VPWR VPWR _3827_/Y sky130_fd_sc_hd__nor2_1
XFILLER_193_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3758_ _6957_/Q _5378_/A _4256_/A _6713_/Q _3740_/X VGND VGND VPWR VPWR _3759_/D
+ sky130_fd_sc_hd__a221o_2
X_6546_ _6715_/CLK _6546_/D fanout439/X VGND VGND VPWR VPWR _6546_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_180_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3689_ _6625_/Q _4154_/A _4250_/A _6709_/Q VGND VGND VPWR VPWR _3689_/X sky130_fd_sc_hd__a22o_4
X_6477_ _3957_/A1 _6477_/D _6432_/X VGND VGND VPWR VPWR hold80/A sky130_fd_sc_hd__dfrtp_2
Xoutput240 _6841_/Q VGND VGND VPWR VPWR mgmt_gpio_out[34] sky130_fd_sc_hd__buf_8
X_5428_ _5581_/A0 hold303/X hold48/X VGND VGND VPWR VPWR _5428_/X sky130_fd_sc_hd__mux2_1
Xoutput251 _3957_/X VGND VGND VPWR VPWR pad_flash_clk sky130_fd_sc_hd__clkbuf_4
Xoutput262 _6809_/Q VGND VGND VPWR VPWR pll90_sel[1] sky130_fd_sc_hd__buf_8
XFILLER_160_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5359_ _5602_/A0 hold593/X _5359_/S VGND VGND VPWR VPWR _5359_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput295 _6500_/Q VGND VGND VPWR VPWR pll_trim[4] sky130_fd_sc_hd__buf_8
Xoutput273 _6806_/Q VGND VGND VPWR VPWR pll_sel[1] sky130_fd_sc_hd__buf_8
Xoutput284 _6813_/Q VGND VGND VPWR VPWR pll_trim[18] sky130_fd_sc_hd__buf_8
XFILLER_160_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7029_ _7124_/CLK _7029_/D fanout436/X VGND VGND VPWR VPWR _7029_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_74_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4730_ _4740_/B _5017_/A _4729_/X VGND VGND VPWR VPWR _4730_/X sky130_fd_sc_hd__o21ba_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4661_ _4745_/A _4697_/A VGND VGND VPWR VPWR _4933_/B sky130_fd_sc_hd__nand2_2
XFILLER_119_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6400_ _6399_/X _7218_/Q _6400_/S VGND VGND VPWR VPWR _7218_/D sky130_fd_sc_hd__mux2_1
XFILLER_175_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3612_ _6552_/Q _4067_/A _4055_/A _6542_/Q VGND VGND VPWR VPWR _3612_/X sky130_fd_sc_hd__a22o_1
XFILLER_190_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4592_ _4812_/A _4947_/B VGND VGND VPWR VPWR _5087_/C sky130_fd_sc_hd__nor2_4
X_6331_ _6356_/A _6331_/B _6331_/C _6331_/D VGND VGND VPWR VPWR _6331_/X sky130_fd_sc_hd__or4_4
Xhold904 _5211_/X VGND VGND VPWR VPWR _6814_/D sky130_fd_sc_hd__bufbuf_16
X_3543_ _3543_/A _3543_/B VGND VGND VPWR VPWR _4055_/A sky130_fd_sc_hd__nor2_8
Xhold926 _4285_/X VGND VGND VPWR VPWR _6737_/D sky130_fd_sc_hd__bufbuf_16
Xhold937 _5244_/X VGND VGND VPWR VPWR _6838_/D sky130_fd_sc_hd__bufbuf_16
Xhold915 _4318_/X VGND VGND VPWR VPWR _6764_/D sky130_fd_sc_hd__bufbuf_16
X_3474_ _6921_/Q _5333_/A _4067_/A _6554_/Q VGND VGND VPWR VPWR _3474_/X sky130_fd_sc_hd__a22o_1
Xhold948 _6506_/Q VGND VGND VPWR VPWR hold948/X sky130_fd_sc_hd__bufbuf_16
Xhold959 _4064_/X VGND VGND VPWR VPWR _6547_/D sky130_fd_sc_hd__bufbuf_16
X_6262_ _6734_/Q _6020_/B _6011_/X _6786_/Q VGND VGND VPWR VPWR _6262_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6193_ _6987_/Q _6028_/X _6034_/Y _6995_/Q _6192_/X VGND VGND VPWR VPWR _6194_/D
+ sky130_fd_sc_hd__a221o_2
X_5213_ hold614/X _5582_/A0 _5215_/S VGND VGND VPWR VPWR _6816_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5144_ _5144_/A _5144_/B VGND VGND VPWR VPWR _5145_/D sky130_fd_sc_hd__nand2_1
XFILLER_97_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5075_ _5075_/A _5075_/B _5075_/C _5075_/D VGND VGND VPWR VPWR _5076_/D sky130_fd_sc_hd__or4_1
X_4026_ _5595_/A0 hold982/X _4033_/S VGND VGND VPWR VPWR _4026_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5977_ _6593_/Q _5680_/X _5700_/X _6539_/Q _5964_/X VGND VGND VPWR VPWR _5977_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4928_ _4932_/A VGND VGND VPWR VPWR _4928_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4859_ _4624_/B _4845_/B _4858_/X _5114_/A _5114_/B VGND VGND VPWR VPWR _4859_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_181_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6529_ _7141_/CLK _6529_/D fanout447/X VGND VGND VPWR VPWR _6529_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_73_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7222_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_28_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_11_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _6649_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_26_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7054_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_180_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5900_ _6739_/Q _5678_/X _5692_/X _7222_/Q _5898_/X VGND VGND VPWR VPWR _5915_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6880_ _6939_/CLK _6880_/D fanout453/X VGND VGND VPWR VPWR _6880_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5831_ _7107_/Q _5675_/X _5687_/X _7051_/Q VGND VGND VPWR VPWR _5831_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5762_ _6911_/Q _5680_/X _5687_/X _7047_/Q _5761_/X VGND VGND VPWR VPWR _5763_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_62_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4713_ _4713_/A _4713_/B _4713_/C _4713_/D VGND VGND VPWR VPWR _4713_/X sky130_fd_sc_hd__or4_1
XFILLER_148_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5693_ _7165_/Q _5702_/B _5701_/C VGND VGND VPWR VPWR _5693_/X sky130_fd_sc_hd__and3_4
X_4644_ _4917_/A _4897_/B VGND VGND VPWR VPWR _4644_/Y sky130_fd_sc_hd__nand2_1
XFILLER_163_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4575_ _4987_/A _4575_/B VGND VGND VPWR VPWR _4575_/Y sky130_fd_sc_hd__nand2_1
Xhold701 _5258_/X VGND VGND VPWR VPWR _6850_/D sky130_fd_sc_hd__bufbuf_16
Xhold712 _6596_/Q VGND VGND VPWR VPWR hold712/X sky130_fd_sc_hd__bufbuf_16
XFILLER_115_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6314_ _6716_/Q _6023_/B _6020_/C _6592_/Q VGND VGND VPWR VPWR _6330_/B sky130_fd_sc_hd__a22o_1
XFILLER_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3526_ _6815_/Q _5207_/A _3344_/Y _6500_/Q VGND VGND VPWR VPWR _3526_/X sky130_fd_sc_hd__a22o_4
Xhold745 _4177_/X VGND VGND VPWR VPWR _6643_/D sky130_fd_sc_hd__bufbuf_16
Xhold734 _5190_/X VGND VGND VPWR VPWR _6789_/D sky130_fd_sc_hd__bufbuf_16
Xhold723 _7139_/Q VGND VGND VPWR VPWR hold723/X sky130_fd_sc_hd__bufbuf_16
Xhold778 _6904_/Q VGND VGND VPWR VPWR hold778/X sky130_fd_sc_hd__bufbuf_16
Xhold767 _6875_/Q VGND VGND VPWR VPWR hold767/X sky130_fd_sc_hd__bufbuf_16
XFILLER_143_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6245_ _6763_/Q _6027_/B _6335_/B _6773_/Q VGND VGND VPWR VPWR _6245_/X sky130_fd_sc_hd__a22o_1
Xhold756 _6855_/Q VGND VGND VPWR VPWR hold756/X sky130_fd_sc_hd__bufbuf_16
XFILLER_103_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3457_ _3457_/A _5252_/B VGND VGND VPWR VPWR _4154_/A sky130_fd_sc_hd__nor2_8
Xhold789 _4279_/X VGND VGND VPWR VPWR _6732_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_162_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6176_ _6962_/Q _6022_/C _6032_/X _7058_/Q VGND VGND VPWR VPWR _6176_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3388_ _7147_/Q _5585_/A _4234_/S input69/X VGND VGND VPWR VPWR _3388_/X sky130_fd_sc_hd__a22o_1
X_5127_ _5127_/A VGND VGND VPWR VPWR _5146_/A sky130_fd_sc_hd__inv_2
XFILLER_69_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5058_ _6781_/Q _6376_/A _5038_/Y _5057_/X VGND VGND VPWR VPWR _5058_/X sky130_fd_sc_hd__a22o_1
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4009_ _4035_/A1 hold885/X _4023_/S VGND VGND VPWR VPWR _4009_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold50 hold50/A VGND VGND VPWR VPWR hold50/X sky130_fd_sc_hd__bufbuf_16
XFILLER_152_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold72 hold72/A VGND VGND VPWR VPWR hold72/X sky130_fd_sc_hd__bufbuf_16
Xhold83 hold83/A VGND VGND VPWR VPWR hold83/X sky130_fd_sc_hd__bufbuf_16
Xhold61 hold61/A VGND VGND VPWR VPWR hold61/X sky130_fd_sc_hd__bufbuf_16
Xhold94 hold94/A VGND VGND VPWR VPWR hold94/X sky130_fd_sc_hd__bufbuf_16
XFILLER_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_mgmt_gpio_in[4] clkbuf_2_3_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _3545_/A1
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_71_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_3 _6484_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4360_ _4566_/A _4558_/B VGND VGND VPWR VPWR _4987_/A sky130_fd_sc_hd__nor2_8
X_3311_ _3501_/A hold84/X VGND VGND VPWR VPWR hold85/A sky130_fd_sc_hd__nor2_8
XFILLER_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4291_ _6411_/A0 hold739/X _4291_/S VGND VGND VPWR VPWR _4291_/X sky130_fd_sc_hd__mux2_1
X_3242_ _4818_/A VGND VGND VPWR VPWR _4564_/A sky130_fd_sc_hd__clkinv_4
X_6030_ _6030_/A _6036_/A VGND VGND VPWR VPWR _6030_/Y sky130_fd_sc_hd__nor2_8
XFILLER_39_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6932_ _7141_/CLK _6932_/D fanout448/X VGND VGND VPWR VPWR _6932_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_82_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6863_ _7127_/CLK _6863_/D fanout449/X VGND VGND VPWR VPWR _6863_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5814_ _6906_/Q _5689_/X _5812_/X _5813_/X VGND VGND VPWR VPWR _5827_/A sky130_fd_sc_hd__a211o_4
XFILLER_62_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6794_ _3545_/A1 _6794_/D _6452_/X VGND VGND VPWR VPWR _6794_/Q sky130_fd_sc_hd__dfrtn_1
X_5745_ _6975_/Q _5676_/X _5703_/X _6871_/Q VGND VGND VPWR VPWR _5745_/X sky130_fd_sc_hd__a22o_1
XFILLER_163_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5676_ _5864_/B _5705_/B _5701_/C VGND VGND VPWR VPWR _5676_/X sky130_fd_sc_hd__and3_4
XFILLER_163_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4627_ _4986_/C _4990_/A _4623_/X _4624_/Y _4626_/Y VGND VGND VPWR VPWR _4627_/X
+ sky130_fd_sc_hd__o2111a_2
XFILLER_190_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold520 _5287_/X VGND VGND VPWR VPWR _6876_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_190_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold542 _5248_/X VGND VGND VPWR VPWR _6841_/D sky130_fd_sc_hd__bufbuf_16
Xhold553 _5312_/X VGND VGND VPWR VPWR _6898_/D sky130_fd_sc_hd__bufbuf_16
Xhold531 _6600_/Q VGND VGND VPWR VPWR hold531/X sky130_fd_sc_hd__bufbuf_16
X_4558_ _4819_/A _4558_/B _4844_/B VGND VGND VPWR VPWR _4558_/X sky130_fd_sc_hd__or3_1
XFILLER_2_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4489_ _4651_/B _4746_/A VGND VGND VPWR VPWR _4659_/A sky130_fd_sc_hd__nor2_8
Xhold586 _5331_/X VGND VGND VPWR VPWR _6915_/D sky130_fd_sc_hd__bufbuf_16
Xhold597 _7059_/Q VGND VGND VPWR VPWR hold597/X sky130_fd_sc_hd__bufbuf_16
Xhold564 _7120_/Q VGND VGND VPWR VPWR hold564/X sky130_fd_sc_hd__bufbuf_16
XFILLER_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold575 _6829_/Q VGND VGND VPWR VPWR hold575/X sky130_fd_sc_hd__bufbuf_16
X_3509_ _6826_/Q _5227_/A _4304_/A _6757_/Q _3507_/X VGND VGND VPWR VPWR _3522_/A
+ sky130_fd_sc_hd__a221o_4
XFILLER_106_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6228_ _6868_/Q _6025_/D _6029_/X _7052_/Q _6227_/X VGND VGND VPWR VPWR _6231_/C
+ sky130_fd_sc_hd__a221o_4
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _5663_/A _7192_/Q _5664_/X _6158_/X VGND VGND VPWR VPWR _6159_/X sky130_fd_sc_hd__a211o_1
Xhold1242 _6868_/Q VGND VGND VPWR VPWR _5278_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_66_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1220 _6753_/Q VGND VGND VPWR VPWR _4305_/A0 sky130_fd_sc_hd__bufbuf_16
Xhold1231 _4044_/X VGND VGND VPWR VPWR _6530_/D sky130_fd_sc_hd__bufbuf_16
Xhold1264 _7056_/Q VGND VGND VPWR VPWR _5490_/A1 sky130_fd_sc_hd__bufbuf_16
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1253 _6994_/Q VGND VGND VPWR VPWR _5420_/A1 sky130_fd_sc_hd__bufbuf_16
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_426 _6411_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_415 _7159_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_404 _6485_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_437 _5260_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_448 hold897/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_459 _6766_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput140 wb_dat_i[17] VGND VGND VPWR VPWR _6381_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput151 wb_dat_i[27] VGND VGND VPWR VPWR _6386_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput162 wb_dat_i[8] VGND VGND VPWR VPWR _6377_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_163_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3860_ _3898_/A _3810_/B _3874_/S _3858_/Y VGND VGND VPWR VPWR _3861_/B sky130_fd_sc_hd__o31a_2
X_3791_ _7021_/Q _5450_/A _3735_/Y _6825_/Q _3743_/X VGND VGND VPWR VPWR _3792_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_188_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5530_ _5584_/A0 hold435/X hold55/X VGND VGND VPWR VPWR _5530_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5461_ _5578_/A0 hold373/X _5467_/S VGND VGND VPWR VPWR _7030_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4412_ _4671_/A _4997_/A VGND VGND VPWR VPWR _4412_/Y sky130_fd_sc_hd__nor2_2
X_7200_ _7201_/CLK _7200_/D _6439_/A VGND VGND VPWR VPWR _7200_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_172_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5392_ _5581_/A0 hold283/X _5395_/S VGND VGND VPWR VPWR _5392_/X sky130_fd_sc_hd__mux2_1
X_4343_ _4340_/B _4690_/A _4341_/X VGND VGND VPWR VPWR _4408_/B sky130_fd_sc_hd__o21ai_4
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7131_ _7131_/CLK _7131_/D fanout432/X VGND VGND VPWR VPWR _7131_/Q sky130_fd_sc_hd__dfrtp_2
X_7062_ _7127_/CLK _7062_/D fanout446/X VGND VGND VPWR VPWR _7062_/Q sky130_fd_sc_hd__dfstp_4
X_4274_ _4274_/A _6406_/B VGND VGND VPWR VPWR _4279_/S sky130_fd_sc_hd__nand2_4
X_3225_ _6976_/Q VGND VGND VPWR VPWR _3225_/Y sky130_fd_sc_hd__inv_2
X_6013_ _6032_/A _6033_/C VGND VGND VPWR VPWR _6034_/B sky130_fd_sc_hd__nand2_8
XFILLER_79_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6915_ _7154_/CLK _6915_/D fanout450/X VGND VGND VPWR VPWR _6915_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_70_728 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6846_ _6851_/CLK _6846_/D fanout423/X VGND VGND VPWR VPWR _6846_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6777_ _6777_/CLK _6777_/D fanout424/X VGND VGND VPWR VPWR _6777_/Q sky130_fd_sc_hd__dfrtp_2
X_3989_ hold74/X _7216_/Q _3991_/S VGND VGND VPWR VPWR hold75/A sky130_fd_sc_hd__mux2_4
X_5728_ _6966_/Q _5691_/X _5701_/X _6950_/Q VGND VGND VPWR VPWR _5728_/X sky130_fd_sc_hd__a22o_1
XFILLER_182_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5659_ _7159_/Q _7160_/Q _5659_/C _7157_/Q VGND VGND VPWR VPWR _5659_/X sky130_fd_sc_hd__or4b_1
XFILLER_184_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold350 _5593_/X VGND VGND VPWR VPWR _7148_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_117_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold361 _7014_/Q VGND VGND VPWR VPWR hold361/X sky130_fd_sc_hd__bufbuf_16
Xhold383 _7150_/Q VGND VGND VPWR VPWR hold383/X sky130_fd_sc_hd__bufbuf_16
Xhold394 _5294_/X VGND VGND VPWR VPWR _6882_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_77_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold372 _6812_/Q VGND VGND VPWR VPWR hold372/X sky130_fd_sc_hd__bufbuf_16
XFILLER_77_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1050 _6607_/Q VGND VGND VPWR VPWR _4134_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1094 _4155_/X VGND VGND VPWR VPWR _6624_/D sky130_fd_sc_hd__bufbuf_16
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1061 _6504_/Q VGND VGND VPWR VPWR _4005_/A1 sky130_fd_sc_hd__bufbuf_16
Xhold1072 _6941_/Q VGND VGND VPWR VPWR _5361_/A1 sky130_fd_sc_hd__bufbuf_16
XFILLER_18_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1083 _7005_/Q VGND VGND VPWR VPWR _5433_/A1 sky130_fd_sc_hd__bufbuf_16
XANTENNA_201 _7016_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_212 _6872_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_223 hold16/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_234 mask_rev_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_267 wb_adr_i[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_256 ser_tx VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_245 mask_rev_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_278 wb_dat_i[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_289 wb_dat_i[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__1132_ clkbuf_0__1132_/X VGND VGND VPWR VPWR _4108_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_123_752 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4961_ _4749_/C _5005_/C _4875_/A VGND VGND VPWR VPWR _4962_/B sky130_fd_sc_hd__a21oi_1
X_4892_ _5005_/C _4756_/B _4623_/D VGND VGND VPWR VPWR _5071_/C sky130_fd_sc_hd__o21ai_2
X_6700_ _7220_/CLK _6700_/D _6362_/B VGND VGND VPWR VPWR _6700_/Q sky130_fd_sc_hd__dfrtp_2
X_3912_ _3905_/X _3909_/Y _3918_/B _6680_/Q VGND VGND VPWR VPWR _6680_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_44_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6631_ _6833_/CLK _6631_/D fanout456/X VGND VGND VPWR VPWR _6631_/Q sky130_fd_sc_hd__dfrtp_2
X_3843_ _6664_/Q _3843_/B VGND VGND VPWR VPWR _3924_/C sky130_fd_sc_hd__nand2_1
XFILLER_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6562_ _7220_/CLK _6562_/D VGND VGND VPWR VPWR _6562_/Q sky130_fd_sc_hd__dfxtp_4
X_3774_ _6535_/Q _4049_/A _3551_/Y input98/X VGND VGND VPWR VPWR _3774_/X sky130_fd_sc_hd__a22o_1
X_6493_ _7129_/CLK _6493_/D fanout428/X VGND VGND VPWR VPWR _6493_/Q sky130_fd_sc_hd__dfstp_4
X_5513_ _5513_/A _5576_/B VGND VGND VPWR VPWR _5521_/S sky130_fd_sc_hd__nand2_8
XFILLER_133_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5444_ _5561_/A0 hold665/X _5449_/S VGND VGND VPWR VPWR _5444_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7114_ _7154_/CLK hold87/X fanout452/X VGND VGND VPWR VPWR _7114_/Q sky130_fd_sc_hd__dfrtp_2
X_5375_ _5600_/A0 hold562/X _5377_/S VGND VGND VPWR VPWR _5375_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4326_ _4326_/A0 hold800/X _4327_/S VGND VGND VPWR VPWR _4326_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4257_ _4257_/A0 _6407_/A0 _4261_/S VGND VGND VPWR VPWR _4257_/X sky130_fd_sc_hd__mux2_1
X_7045_ _7101_/CLK _7045_/D fanout430/X VGND VGND VPWR VPWR _7045_/Q sky130_fd_sc_hd__dfstp_4
X_3208_ _7112_/Q VGND VGND VPWR VPWR _3208_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4188_ hold804/X _4326_/A0 _4189_/S VGND VGND VPWR VPWR _4188_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6829_ _7035_/CLK _6829_/D fanout432/X VGND VGND VPWR VPWR _6829_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_155_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold180 _6463_/Q VGND VGND VPWR VPWR hold180/X sky130_fd_sc_hd__bufbuf_16
XFILLER_151_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold191 _6482_/Q VGND VGND VPWR VPWR hold191/X sky130_fd_sc_hd__bufbuf_16
XFILLER_144_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3490_ _7228_/A _5245_/A _4136_/A _6613_/Q VGND VGND VPWR VPWR _3490_/X sky130_fd_sc_hd__a22o_2
XFILLER_115_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5160_ _4414_/B _4711_/C _4802_/A _5159_/X VGND VGND VPWR VPWR _5161_/D sky130_fd_sc_hd__a211oi_2
X_5091_ _5135_/B _5119_/B _5091_/C VGND VGND VPWR VPWR _5091_/X sky130_fd_sc_hd__or3_1
XFILLER_96_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4111_ _6588_/Q _3379_/X _4111_/S VGND VGND VPWR VPWR _6588_/D sky130_fd_sc_hd__mux2_1
X_4042_ _5602_/A0 hold355/X _4042_/S VGND VGND VPWR VPWR _4042_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5993_ _6019_/A _6033_/C _6035_/C VGND VGND VPWR VPWR _6027_/B sky130_fd_sc_hd__and3b_4
XFILLER_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4944_ _4772_/A _4624_/B _5114_/A _4943_/Y VGND VGND VPWR VPWR _4945_/D sky130_fd_sc_hd__a211o_1
X_4875_ _4875_/A _4899_/B VGND VGND VPWR VPWR _4936_/C sky130_fd_sc_hd__nor2_4
XFILLER_149_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6614_ _6616_/CLK _6614_/D fanout439/X VGND VGND VPWR VPWR _6614_/Q sky130_fd_sc_hd__dfrtp_2
X_3826_ _3826_/A _3826_/B VGND VGND VPWR VPWR _6482_/D sky130_fd_sc_hd__xor2_1
XFILLER_193_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3757_ _6733_/Q _4280_/A _5236_/A _6833_/Q _3742_/X VGND VGND VPWR VPWR _3759_/C
+ sky130_fd_sc_hd__a221o_1
X_6545_ _6649_/CLK _6545_/D fanout439/X VGND VGND VPWR VPWR _6545_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3688_ _6942_/Q _5360_/A _4268_/A _6724_/Q _3670_/X VGND VGND VPWR VPWR _3693_/A
+ sky130_fd_sc_hd__a221o_1
X_6476_ _3957_/A1 _6476_/D _6431_/X VGND VGND VPWR VPWR _6476_/Q sky130_fd_sc_hd__dfrtp_2
Xoutput230 _6515_/Q VGND VGND VPWR VPWR mgmt_gpio_out[25] sky130_fd_sc_hd__buf_8
Xoutput241 _3936_/X VGND VGND VPWR VPWR mgmt_gpio_out[35] sky130_fd_sc_hd__buf_8
X_5427_ _5571_/A0 hold629/X hold48/X VGND VGND VPWR VPWR _7000_/D sky130_fd_sc_hd__mux2_1
Xoutput252 _3958_/Y VGND VGND VPWR VPWR pad_flash_clk_oeb sky130_fd_sc_hd__buf_8
X_5358_ _5601_/A0 hold624/X _5359_/S VGND VGND VPWR VPWR _5358_/X sky130_fd_sc_hd__mux2_1
Xoutput285 _6814_/Q VGND VGND VPWR VPWR pll_trim[19] sky130_fd_sc_hd__buf_8
Xoutput274 _6807_/Q VGND VGND VPWR VPWR pll_sel[2] sky130_fd_sc_hd__buf_8
Xoutput263 _6810_/Q VGND VGND VPWR VPWR pll90_sel[2] sky130_fd_sc_hd__buf_8
XFILLER_99_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput296 _6501_/Q VGND VGND VPWR VPWR pll_trim[5] sky130_fd_sc_hd__buf_8
X_4309_ hold831/X _6411_/A0 _4309_/S VGND VGND VPWR VPWR _4309_/X sky130_fd_sc_hd__mux2_1
X_5289_ _5289_/A0 _5289_/A1 _5296_/S VGND VGND VPWR VPWR _6877_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7028_ _7123_/CLK _7028_/D fanout434/X VGND VGND VPWR VPWR _7028_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4660_ _4745_/A _4697_/A VGND VGND VPWR VPWR _4660_/X sky130_fd_sc_hd__and2_4
XFILLER_30_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3611_ input37/X _4023_/S _4118_/A _6596_/Q VGND VGND VPWR VPWR _3611_/X sky130_fd_sc_hd__a22o_1
XFILLER_162_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4591_ _4898_/B _4591_/B VGND VGND VPWR VPWR _4591_/X sky130_fd_sc_hd__or2_1
XFILLER_127_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6330_ _6330_/A _6330_/B _6330_/C _6330_/D VGND VGND VPWR VPWR _6331_/D sky130_fd_sc_hd__or4_1
Xhold905 _6733_/Q VGND VGND VPWR VPWR hold905/X sky130_fd_sc_hd__bufbuf_16
Xhold916 _6672_/Q VGND VGND VPWR VPWR hold916/X sky130_fd_sc_hd__bufbuf_16
XFILLER_128_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3542_ _7025_/Q _5450_/A _5324_/A _6913_/Q _3541_/X VGND VGND VPWR VPWR _3546_/C
+ sky130_fd_sc_hd__a221o_1
Xhold927 _6799_/Q VGND VGND VPWR VPWR hold927/X sky130_fd_sc_hd__bufbuf_16
Xhold938 _7055_/Q VGND VGND VPWR VPWR hold938/X sky130_fd_sc_hd__bufbuf_16
Xhold949 _4010_/X VGND VGND VPWR VPWR _6506_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_142_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3473_ _3473_/A _3473_/B VGND VGND VPWR VPWR _4067_/A sky130_fd_sc_hd__nor2_8
X_6261_ _6655_/Q _6311_/B VGND VGND VPWR VPWR _6261_/X sky130_fd_sc_hd__and2_1
XFILLER_170_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6192_ _7075_/Q _6009_/X _6020_/D _6971_/Q VGND VGND VPWR VPWR _6192_/X sky130_fd_sc_hd__a22o_1
X_5212_ hold466/X _6411_/A0 _5215_/S VGND VGND VPWR VPWR _5212_/X sky130_fd_sc_hd__mux2_1
X_5143_ _5143_/A _5143_/B _5143_/C VGND VGND VPWR VPWR _5143_/Y sky130_fd_sc_hd__nor3_2
XFILLER_97_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5074_ _5074_/A _5126_/A _5175_/A _5145_/C VGND VGND VPWR VPWR _5075_/D sky130_fd_sc_hd__or4_1
XFILLER_111_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4025_ _4025_/A _5594_/B VGND VGND VPWR VPWR _4033_/S sky130_fd_sc_hd__nand2_8
XFILLER_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5976_ _5976_/A _5976_/B _5976_/C _5976_/D VGND VGND VPWR VPWR _5976_/X sky130_fd_sc_hd__or4_2
XFILLER_178_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4927_ _5023_/A _4927_/B VGND VGND VPWR VPWR _4932_/A sky130_fd_sc_hd__nor2_2
XFILLER_80_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4858_ _4399_/Y _4845_/B _5171_/A _4856_/X _4857_/X VGND VGND VPWR VPWR _4858_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_193_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3809_ _6469_/Q _6468_/Q VGND VGND VPWR VPWR _3810_/B sky130_fd_sc_hd__nor2_1
X_4789_ _4772_/A _4575_/B _4453_/Y _4719_/X VGND VGND VPWR VPWR _4789_/X sky130_fd_sc_hd__a22o_1
X_6528_ _6987_/CLK _6528_/D fanout450/X VGND VGND VPWR VPWR _6528_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_7_csclk _6722_/CLK VGND VGND VPWR VPWR _6747_/CLK sky130_fd_sc_hd__clkbuf_8
X_6459_ _3957_/A1 _6459_/D _6414_/X VGND VGND VPWR VPWR _6459_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5830_ _7181_/Q _6309_/S _5828_/X _5829_/X VGND VGND VPWR VPWR _7181_/D sky130_fd_sc_hd__o22a_1
X_5761_ _7063_/Q _5669_/X _5690_/X _7095_/Q VGND VGND VPWR VPWR _5761_/X sky130_fd_sc_hd__a22o_1
XFILLER_187_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4712_ _4922_/A _4712_/B _5069_/B _4936_/A VGND VGND VPWR VPWR _4713_/D sky130_fd_sc_hd__or4_1
XFILLER_187_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5692_ _7165_/Q _5705_/B _5706_/B VGND VGND VPWR VPWR _5692_/X sky130_fd_sc_hd__and3_4
XFILLER_30_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4643_ _4812_/A _4819_/B _5062_/A VGND VGND VPWR VPWR _4897_/B sky130_fd_sc_hd__or3_4
X_4574_ _5128_/A VGND VGND VPWR VPWR _4574_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold702 _7047_/Q VGND VGND VPWR VPWR hold702/X sky130_fd_sc_hd__bufbuf_16
Xhold735 _6913_/Q VGND VGND VPWR VPWR hold735/X sky130_fd_sc_hd__bufbuf_16
Xhold746 _6971_/Q VGND VGND VPWR VPWR hold746/X sky130_fd_sc_hd__bufbuf_16
X_6313_ _6662_/Q _5996_/X _6021_/C _6548_/Q VGND VGND VPWR VPWR _6330_/A sky130_fd_sc_hd__a22o_1
X_3525_ _7033_/Q _5459_/A _4292_/A _6747_/Q _3523_/X VGND VGND VPWR VPWR _3533_/A
+ sky130_fd_sc_hd__a221o_1
Xhold713 _7083_/Q VGND VGND VPWR VPWR hold713/X sky130_fd_sc_hd__bufbuf_16
Xhold724 _5583_/X VGND VGND VPWR VPWR _7139_/D sky130_fd_sc_hd__bufbuf_16
Xhold779 _5319_/X VGND VGND VPWR VPWR _6904_/D sky130_fd_sc_hd__bufbuf_16
Xhold768 _5286_/X VGND VGND VPWR VPWR _6875_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_143_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6244_ _6540_/Q _6023_/C _6032_/X _6649_/Q _6243_/X VGND VGND VPWR VPWR _6247_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold757 _5264_/X VGND VGND VPWR VPWR _6855_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_131_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3456_ input16/X _3368_/Y _4130_/A _6608_/Q VGND VGND VPWR VPWR _3456_/X sky130_fd_sc_hd__a22o_1
X_3387_ input41/X _4023_/S _5324_/A _6915_/Q VGND VGND VPWR VPWR _3387_/X sky130_fd_sc_hd__a22o_1
X_6175_ _6906_/Q _6021_/A _6025_/A _6938_/Q _6174_/X VGND VGND VPWR VPWR _6181_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5126_ _5126_/A _5126_/B VGND VGND VPWR VPWR _5127_/A sky130_fd_sc_hd__nor2_1
X_5057_ _5057_/A _5057_/B VGND VGND VPWR VPWR _5057_/X sky130_fd_sc_hd__or2_2
XFILLER_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4008_ hold20/X _6421_/B _4007_/X _4023_/S _5486_/B VGND VGND VPWR VPWR _4024_/S
+ sky130_fd_sc_hd__o221a_4
XFILLER_84_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5959_ _5959_/A _5959_/B _5959_/C _5959_/D VGND VGND VPWR VPWR _5959_/X sky130_fd_sc_hd__or4_1
XFILLER_25_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold40 hold40/A VGND VGND VPWR VPWR hold40/X sky130_fd_sc_hd__bufbuf_16
XFILLER_102_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold73 hold73/A VGND VGND VPWR VPWR hold5/A sky130_fd_sc_hd__bufbuf_16
Xhold51 hold51/A VGND VGND VPWR VPWR hold51/X sky130_fd_sc_hd__bufbuf_16
Xhold62 hold62/A VGND VGND VPWR VPWR hold62/X sky130_fd_sc_hd__bufbuf_16
XFILLER_48_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold95 hold95/A VGND VGND VPWR VPWR hold95/X sky130_fd_sc_hd__bufbuf_16
XFILLER_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold84 hold84/A VGND VGND VPWR VPWR hold84/X sky130_fd_sc_hd__bufbuf_16
XFILLER_90_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_4 _6497_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3310_ hold20/X _4241_/A VGND VGND VPWR VPWR _4023_/S sky130_fd_sc_hd__nor2_8
XFILLER_112_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4290_ _6410_/A0 hold990/X _4291_/S VGND VGND VPWR VPWR _4290_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3241_ _7165_/Q VGND VGND VPWR VPWR _5963_/B sky130_fd_sc_hd__inv_8
XFILLER_112_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6931_ _7130_/CLK _6931_/D fanout453/X VGND VGND VPWR VPWR _6931_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_81_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6862_ _7127_/CLK _6862_/D fanout446/X VGND VGND VPWR VPWR _6862_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_179_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5813_ _6914_/Q _5680_/X _5700_/X _6866_/Q _5811_/X VGND VGND VPWR VPWR _5813_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6793_ _3545_/A1 _6793_/D _6451_/X VGND VGND VPWR VPWR _6793_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_50_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5744_ _7177_/Q _6309_/S _5742_/X _5743_/X VGND VGND VPWR VPWR _7177_/D sky130_fd_sc_hd__o22a_1
XFILLER_187_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5675_ _7165_/Q _5705_/B _5701_/C VGND VGND VPWR VPWR _5675_/X sky130_fd_sc_hd__and3_4
Xclkbuf_leaf_72_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6759_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4626_ _5114_/B VGND VGND VPWR VPWR _4626_/Y sky130_fd_sc_hd__inv_2
Xhold510 _4028_/X VGND VGND VPWR VPWR _6516_/D sky130_fd_sc_hd__bufbuf_16
Xhold521 _6696_/Q VGND VGND VPWR VPWR hold521/X sky130_fd_sc_hd__bufbuf_16
Xhold543 _7111_/Q VGND VGND VPWR VPWR hold543/X sky130_fd_sc_hd__bufbuf_16
Xhold554 _6692_/Q VGND VGND VPWR VPWR hold554/X sky130_fd_sc_hd__bufbuf_16
Xhold532 _4126_/X VGND VGND VPWR VPWR _6600_/D sky130_fd_sc_hd__bufbuf_16
X_4557_ _4883_/A _5119_/A _4557_/C _4557_/D VGND VGND VPWR VPWR _4559_/C sky130_fd_sc_hd__or4_1
X_4488_ _4655_/A _4651_/B VGND VGND VPWR VPWR _4488_/X sky130_fd_sc_hd__or2_1
Xhold587 _6878_/Q VGND VGND VPWR VPWR hold587/X sky130_fd_sc_hd__bufbuf_16
Xhold565 _5562_/X VGND VGND VPWR VPWR _7120_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_104_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold576 _5231_/X VGND VGND VPWR VPWR _6829_/D sky130_fd_sc_hd__bufbuf_16
X_3508_ hold53/X _3733_/B VGND VGND VPWR VPWR _4304_/A sky130_fd_sc_hd__nor2_8
X_3439_ _6882_/Q _5288_/A _5405_/A _6986_/Q VGND VGND VPWR VPWR _3439_/X sky130_fd_sc_hd__a22o_4
Xhold598 _5493_/X VGND VGND VPWR VPWR _7059_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_103_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6227_ _7108_/Q _5653_/X _6022_/B _6948_/Q VGND VGND VPWR VPWR _6227_/X sky130_fd_sc_hd__a22o_1
XFILLER_58_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6158_ _6857_/Q _6060_/B _6144_/X _6157_/X _6308_/S VGND VGND VPWR VPWR _6158_/X
+ sky130_fd_sc_hd__o221a_4
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1243 _7116_/Q VGND VGND VPWR VPWR _5557_/A0 sky130_fd_sc_hd__bufbuf_16
X_5109_ _4748_/B _5041_/X _5056_/B _5104_/Y VGND VGND VPWR VPWR _5178_/B sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_10_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _6629_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1221 _4305_/X VGND VGND VPWR VPWR _6753_/D sky130_fd_sc_hd__bufbuf_16
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1232 _6763_/Q VGND VGND VPWR VPWR _4317_/A0 sky130_fd_sc_hd__bufbuf_16
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1210 _5246_/X VGND VGND VPWR VPWR _6839_/D sky130_fd_sc_hd__bufbuf_16
X_6089_ _6975_/Q _6023_/B _6021_/C _6879_/Q _6087_/X VGND VGND VPWR VPWR _6106_/A
+ sky130_fd_sc_hd__a221o_1
Xhold1265 _6693_/Q VGND VGND VPWR VPWR hold641/A sky130_fd_sc_hd__bufbuf_16
Xhold1254 _7135_/Q VGND VGND VPWR VPWR _5579_/A1 sky130_fd_sc_hd__bufbuf_16
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_416 _3972_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_405 mask_rev_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_csclk _7137_/CLK VGND VGND VPWR VPWR _6964_/CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA_427 _5581_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_438 _3995_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_449 hold907/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput152 wb_dat_i[28] VGND VGND VPWR VPWR _6390_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput130 wb_adr_i[9] VGND VGND VPWR VPWR _4351_/A sky130_fd_sc_hd__clkbuf_4
Xinput141 wb_dat_i[18] VGND VGND VPWR VPWR _6383_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput163 wb_dat_i[9] VGND VGND VPWR VPWR _6380_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_49_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3790_ _6997_/Q _5423_/A _4310_/A _6758_/Q _3789_/X VGND VGND VPWR VPWR _3792_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5460_ _5541_/A0 _5460_/A1 _5467_/S VGND VGND VPWR VPWR _7029_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4411_ _4871_/A _4997_/A VGND VGND VPWR VPWR _4411_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5391_ _5571_/A0 hold630/X _5395_/S VGND VGND VPWR VPWR _5391_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7130_ _7130_/CLK _7130_/D fanout454/X VGND VGND VPWR VPWR _7130_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_172_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4342_ _4654_/A _4654_/B VGND VGND VPWR VPWR _4690_/A sky130_fd_sc_hd__nand2_4
XFILLER_141_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4273_ hold872/X _6411_/A0 _4273_/S VGND VGND VPWR VPWR _4273_/X sky130_fd_sc_hd__mux2_1
X_7061_ _7129_/CLK _7061_/D fanout428/X VGND VGND VPWR VPWR _7061_/Q sky130_fd_sc_hd__dfstp_4
X_3224_ _6984_/Q VGND VGND VPWR VPWR _3224_/Y sky130_fd_sc_hd__inv_2
X_6012_ _6012_/A _6035_/A _6018_/A VGND VGND VPWR VPWR _6020_/D sky130_fd_sc_hd__and3_4
XFILLER_101_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
.ends

