magic
tech sky130A
timestamp 1534629073
<< checkpaint >>
rect -4974 13142 296936 347714
<< via3 >>
rect -4344 346852 -4072 347084
rect 296034 346852 296306 347084
rect -3864 346412 -3592 346644
rect 295554 346412 295826 346644
rect -2904 345972 -2632 346204
rect 294594 345972 294866 346204
rect -3384 345532 -3112 345764
rect 295074 345532 295346 345764
rect -2424 345092 -2152 345324
rect 294114 345092 294386 345324
rect -1944 344652 -1672 344884
rect 293634 344652 293906 344884
rect -1464 344212 -1192 344444
rect 293154 344212 293426 344444
rect -984 343772 -712 344004
rect 292674 343772 292946 344004
rect -4344 336852 -4072 337084
rect 296034 336852 296306 337084
rect -3864 336412 -3592 336644
rect 295554 336412 295826 336644
rect -2904 335972 -2632 336204
rect 294594 335972 294866 336204
rect 295074 335532 295346 335764
rect -2424 335092 -2152 335324
rect 294114 335092 294386 335324
rect -1944 334652 -1672 334884
rect 293634 334652 293906 334884
rect -1464 334212 -1192 334444
rect 293154 334212 293426 334444
rect -984 333772 -712 334004
rect 292674 333772 292946 334004
rect -4344 326852 -4072 327084
rect 296034 326852 296306 327084
rect -3864 326412 -3592 326644
rect 295554 326412 295826 326644
rect -2904 325972 -2632 326204
rect 294594 325972 294866 326204
rect -3384 325532 -3112 325764
rect 295074 325532 295346 325764
rect -2424 325092 -2152 325324
rect 294114 325092 294386 325324
rect -1944 324652 -1672 324884
rect 293634 324652 293906 324884
rect -1464 324212 -1192 324444
rect 293154 324212 293426 324444
rect -984 323772 -712 324004
rect 292674 323772 292946 324004
rect -4344 316852 -4072 317084
rect 296034 316852 296306 317084
rect -3864 316412 -3592 316644
rect 295554 316412 295826 316644
rect 294594 315972 294866 316204
rect -3384 315532 -3112 315764
rect 295074 315532 295346 315764
rect -2424 315092 -2152 315324
rect 294114 315092 294386 315324
rect -1944 314652 -1672 314884
rect 293634 314652 293906 314884
rect -1464 314212 -1192 314444
rect 293154 314212 293426 314444
rect -984 313772 -712 314004
rect 292674 313772 292946 314004
rect -4344 306852 -4072 307084
rect 296034 306852 296306 307084
rect -3864 306412 -3592 306644
rect 295554 306412 295826 306644
rect -2904 305972 -2632 306204
rect 294594 305972 294866 306204
rect -3384 305532 -3112 305764
rect 295074 305532 295346 305764
rect -2424 305092 -2152 305324
rect 294114 305092 294386 305324
rect -1944 304652 -1672 304884
rect 293634 304652 293906 304884
rect -1464 304212 -1192 304444
rect 293154 304212 293426 304444
rect -984 303772 -712 304004
rect 292674 303772 292946 304004
rect -4344 296852 -4072 297084
rect 296034 296852 296306 297084
rect 295554 296412 295826 296644
rect -2904 295972 -2632 296204
rect 294594 295972 294866 296204
rect -3384 295532 -3112 295764
rect 295074 295532 295346 295764
rect -2424 295092 -2152 295324
rect 294114 295092 294386 295324
rect -1944 294652 -1672 294884
rect 293634 294652 293906 294884
rect -1464 294212 -1192 294444
rect 293154 294212 293426 294444
rect -984 293772 -712 294004
rect 292674 293772 292946 294004
rect -4344 286852 -4072 287084
rect 296034 286852 296306 287084
rect -3864 286412 -3592 286644
rect 295554 286412 295826 286644
rect -2904 285972 -2632 286204
rect 294594 285972 294866 286204
rect -3384 285532 -3112 285764
rect 295074 285532 295346 285764
rect -2424 285092 -2152 285324
rect 294114 285092 294386 285324
rect -1944 284652 -1672 284884
rect 293634 284652 293906 284884
rect -1464 284212 -1192 284444
rect 293154 284212 293426 284444
rect -984 283772 -712 284004
rect 292674 283772 292946 284004
rect 296034 276852 296306 277084
rect -3864 276412 -3592 276644
rect 295554 276412 295826 276644
rect -2904 275972 -2632 276204
rect 294594 275972 294866 276204
rect -3384 275532 -3112 275764
rect 295074 275532 295346 275764
rect -2424 275092 -2152 275324
rect 294114 275092 294386 275324
rect -1944 274652 -1672 274884
rect 293634 274652 293906 274884
rect -1464 274212 -1192 274444
rect 293154 274212 293426 274444
rect -984 273772 -712 274004
rect 292674 273772 292946 274004
rect -4344 266852 -4072 267084
rect 296034 266852 296306 267084
rect -3864 266412 -3592 266644
rect 295554 266412 295826 266644
rect -2904 265972 -2632 266204
rect 294594 265972 294866 266204
rect -3384 265532 -3112 265764
rect 295074 265532 295346 265764
rect -2424 265092 -2152 265324
rect 294114 265092 294386 265324
rect -1944 264652 -1672 264884
rect 293634 264652 293906 264884
rect -1464 264212 -1192 264444
rect 293154 264212 293426 264444
rect 292674 263772 292946 264004
rect -4344 256852 -4072 257084
rect 296034 256852 296306 257084
rect -3864 256412 -3592 256644
rect 295554 256412 295826 256644
rect -2904 255972 -2632 256204
rect 294594 255972 294866 256204
rect -3384 255532 -3112 255764
rect 295074 255532 295346 255764
rect -2424 255092 -2152 255324
rect 294114 255092 294386 255324
rect -1944 254652 -1672 254884
rect 293634 254652 293906 254884
rect -1464 254212 -1192 254444
rect 293154 254212 293426 254444
rect -984 253772 -712 254004
rect 292674 253772 292946 254004
rect -4344 246852 -4072 247084
rect 296034 246852 296306 247084
rect -3864 246412 -3592 246644
rect 295554 246412 295826 246644
rect -2904 245972 -2632 246204
rect 294594 245972 294866 246204
rect -3384 245532 -3112 245764
rect 295074 245532 295346 245764
rect -2424 245092 -2152 245324
rect 294114 245092 294386 245324
rect -1944 244652 -1672 244884
rect 293634 244652 293906 244884
rect 293154 244212 293426 244444
rect -984 243772 -712 244004
rect 292674 243772 292946 244004
rect -4344 236852 -4072 237084
rect 296034 236852 296306 237084
rect -3864 236412 -3592 236644
rect 295554 236412 295826 236644
rect -2904 235972 -2632 236204
rect 294594 235972 294866 236204
rect -3384 235532 -3112 235764
rect 295074 235532 295346 235764
rect -2424 235092 -2152 235324
rect 294114 235092 294386 235324
rect -1944 234652 -1672 234884
rect 293634 234652 293906 234884
rect -1464 234212 -1192 234444
rect 293154 234212 293426 234444
rect -984 233772 -712 234004
rect 292674 233772 292946 234004
rect -4344 226852 -4072 227084
rect 296034 226852 296306 227084
rect -3864 226412 -3592 226644
rect 295554 226412 295826 226644
rect -2904 225972 -2632 226204
rect 294594 225972 294866 226204
rect -3384 225532 -3112 225764
rect 295074 225532 295346 225764
rect -2424 225092 -2152 225324
rect 294114 225092 294386 225324
rect 293634 224652 293906 224884
rect -1464 224212 -1192 224444
rect 293154 224212 293426 224444
rect -984 223772 -712 224004
rect 292674 223772 292946 224004
rect -4344 216852 -4072 217084
rect 296034 216852 296306 217084
rect -3864 216412 -3592 216644
rect 295554 216412 295826 216644
rect -2904 215972 -2632 216204
rect 294594 215972 294866 216204
rect -3384 215532 -3112 215764
rect 295074 215532 295346 215764
rect -2424 215092 -2152 215324
rect 294114 215092 294386 215324
rect -1944 214652 -1672 214884
rect 293634 214652 293906 214884
rect -1464 214212 -1192 214444
rect 293154 214212 293426 214444
rect -984 213772 -712 214004
rect 292674 213772 292946 214004
rect -4344 206852 -4072 207084
rect 296034 206852 296306 207084
rect -3864 206412 -3592 206644
rect 295554 206412 295826 206644
rect -2904 205972 -2632 206204
rect 294594 205972 294866 206204
rect -3384 205532 -3112 205764
rect 295074 205532 295346 205764
rect 294114 205092 294386 205324
rect -1944 204652 -1672 204884
rect 293634 204652 293906 204884
rect -1464 204212 -1192 204444
rect 293154 204212 293426 204444
rect -984 203772 -712 204004
rect 292674 203772 292946 204004
rect -4344 196852 -4072 197084
rect 296034 196852 296306 197084
rect -3864 196412 -3592 196644
rect 295554 196412 295826 196644
rect -2904 195972 -2632 196204
rect 294594 195972 294866 196204
rect -3384 195532 -3112 195764
rect 295074 195532 295346 195764
rect -2424 195092 -2152 195324
rect 294114 195092 294386 195324
rect -1944 194652 -1672 194884
rect 293634 194652 293906 194884
rect -1464 194212 -1192 194444
rect 293154 194212 293426 194444
rect -984 193772 -712 194004
rect 292674 193772 292946 194004
rect -4344 186852 -4072 187084
rect 296034 186852 296306 187084
rect -3864 186412 -3592 186644
rect 295554 186412 295826 186644
rect -2904 185972 -2632 186204
rect 294594 185972 294866 186204
rect 295074 185532 295346 185764
rect -2424 185092 -2152 185324
rect 294114 185092 294386 185324
rect -1944 184652 -1672 184884
rect 293634 184652 293906 184884
rect -1464 184212 -1192 184444
rect 293154 184212 293426 184444
rect -984 183772 -712 184004
rect 292674 183772 292946 184004
rect -4344 176852 -4072 177084
rect 296034 176852 296306 177084
rect -3864 176412 -3592 176644
rect 295554 176412 295826 176644
rect -2904 175972 -2632 176204
rect 294594 175972 294866 176204
rect -3384 175532 -3112 175764
rect 295074 175532 295346 175764
rect -2424 175092 -2152 175324
rect 294114 175092 294386 175324
rect -1944 174652 -1672 174884
rect 293634 174652 293906 174884
rect -1464 174212 -1192 174444
rect 293154 174212 293426 174444
rect -984 173772 -712 174004
rect 292674 173772 292946 174004
rect -4344 166852 -4072 167084
rect 296034 166852 296306 167084
rect -3864 166412 -3592 166644
rect 295554 166412 295826 166644
rect 294594 165972 294866 166204
rect -3384 165532 -3112 165764
rect 295074 165532 295346 165764
rect -2424 165092 -2152 165324
rect 294114 165092 294386 165324
rect -1944 164652 -1672 164884
rect 293634 164652 293906 164884
rect -1464 164212 -1192 164444
rect 293154 164212 293426 164444
rect -984 163772 -712 164004
rect 292674 163772 292946 164004
rect -4344 156852 -4072 157084
rect 296034 156852 296306 157084
rect -3864 156412 -3592 156644
rect 295554 156412 295826 156644
rect -2904 155972 -2632 156204
rect 294594 155972 294866 156204
rect -3384 155532 -3112 155764
rect 295074 155532 295346 155764
rect -2424 155092 -2152 155324
rect 294114 155092 294386 155324
rect -1944 154652 -1672 154884
rect 293634 154652 293906 154884
rect -1464 154212 -1192 154444
rect 293154 154212 293426 154444
rect -984 153772 -712 154004
rect 292674 153772 292946 154004
rect -4344 146852 -4072 147084
rect 296034 146852 296306 147084
rect 295554 146412 295826 146644
rect -2904 145972 -2632 146204
rect 294594 145972 294866 146204
rect -3384 145532 -3112 145764
rect 295074 145532 295346 145764
rect -2424 145092 -2152 145324
rect 294114 145092 294386 145324
rect -1944 144652 -1672 144884
rect 293634 144652 293906 144884
rect -1464 144212 -1192 144444
rect 293154 144212 293426 144444
rect -984 143772 -712 144004
rect 292674 143772 292946 144004
rect -4344 136852 -4072 137084
rect 296034 136852 296306 137084
rect -3864 136412 -3592 136644
rect 295554 136412 295826 136644
rect -2904 135972 -2632 136204
rect 294594 135972 294866 136204
rect -3384 135532 -3112 135764
rect 295074 135532 295346 135764
rect -2424 135092 -2152 135324
rect 294114 135092 294386 135324
rect -1944 134652 -1672 134884
rect 293634 134652 293906 134884
rect -1464 134212 -1192 134444
rect 293154 134212 293426 134444
rect -984 133772 -712 134004
rect 292674 133772 292946 134004
rect 296034 126852 296306 127084
rect -3864 126412 -3592 126644
rect 295554 126412 295826 126644
rect -2904 125972 -2632 126204
rect 294594 125972 294866 126204
rect -3384 125532 -3112 125764
rect 295074 125532 295346 125764
rect -2424 125092 -2152 125324
rect 294114 125092 294386 125324
rect -1944 124652 -1672 124884
rect 293634 124652 293906 124884
rect -1464 124212 -1192 124444
rect 293154 124212 293426 124444
rect -984 123772 -712 124004
rect 292674 123772 292946 124004
rect -4344 116852 -4072 117084
rect 296034 116852 296306 117084
rect -3864 116412 -3592 116644
rect 295554 116412 295826 116644
rect -2904 115972 -2632 116204
rect 294594 115972 294866 116204
rect -3384 115532 -3112 115764
rect 295074 115532 295346 115764
rect -2424 115092 -2152 115324
rect 294114 115092 294386 115324
rect -1944 114652 -1672 114884
rect 293634 114652 293906 114884
rect -1464 114212 -1192 114444
rect 293154 114212 293426 114444
rect 292674 113772 292946 114004
rect -4344 106852 -4072 107084
rect 296034 106852 296306 107084
rect -3864 106412 -3592 106644
rect 295554 106412 295826 106644
rect -2904 105972 -2632 106204
rect 294594 105972 294866 106204
rect -3384 105532 -3112 105764
rect 295074 105532 295346 105764
rect -2424 105092 -2152 105324
rect 294114 105092 294386 105324
rect -1944 104652 -1672 104884
rect 293634 104652 293906 104884
rect -1464 104212 -1192 104444
rect 293154 104212 293426 104444
rect -984 103772 -712 104004
rect 292674 103772 292946 104004
rect -4344 96852 -4072 97084
rect 296034 96852 296306 97084
rect -3864 96412 -3592 96644
rect 295554 96412 295826 96644
rect -2904 95972 -2632 96204
rect 294594 95972 294866 96204
rect -3384 95532 -3112 95764
rect 295074 95532 295346 95764
rect -2424 95092 -2152 95324
rect 294114 95092 294386 95324
rect -1944 94652 -1672 94884
rect 293634 94652 293906 94884
rect 293154 94212 293426 94444
rect -984 93772 -712 94004
rect 292674 93772 292946 94004
rect -4344 86852 -4072 87084
rect 296034 86852 296306 87084
rect -3864 86412 -3592 86644
rect 295554 86412 295826 86644
rect -2904 85972 -2632 86204
rect 294594 85972 294866 86204
rect -3384 85532 -3112 85764
rect 295074 85532 295346 85764
rect -2424 85092 -2152 85324
rect 294114 85092 294386 85324
rect -1944 84652 -1672 84884
rect 293634 84652 293906 84884
rect -1464 84212 -1192 84444
rect 293154 84212 293426 84444
rect -984 83772 -712 84004
rect 292674 83772 292946 84004
rect -4344 76852 -4072 77084
rect 296034 76852 296306 77084
rect -3864 76412 -3592 76644
rect 295554 76412 295826 76644
rect -2904 75972 -2632 76204
rect 294594 75972 294866 76204
rect -3384 75532 -3112 75764
rect 295074 75532 295346 75764
rect -2424 75092 -2152 75324
rect 294114 75092 294386 75324
rect 293634 74652 293906 74884
rect -1464 74212 -1192 74444
rect 293154 74212 293426 74444
rect -984 73772 -712 74004
rect 292674 73772 292946 74004
rect -4344 66852 -4072 67084
rect 296034 66852 296306 67084
rect -3864 66412 -3592 66644
rect 295554 66412 295826 66644
rect -2904 65972 -2632 66204
rect 294594 65972 294866 66204
rect -3384 65532 -3112 65764
rect 295074 65532 295346 65764
rect -2424 65092 -2152 65324
rect 294114 65092 294386 65324
rect -1944 64652 -1672 64884
rect 293634 64652 293906 64884
rect -1464 64212 -1192 64444
rect 293154 64212 293426 64444
rect -984 63772 -712 64004
rect 292674 63772 292946 64004
rect -4344 56852 -4072 57084
rect 296034 56852 296306 57084
rect -3864 56412 -3592 56644
rect 295554 56412 295826 56644
rect -2904 55972 -2632 56204
rect 294594 55972 294866 56204
rect -3384 55532 -3112 55764
rect 295074 55532 295346 55764
rect 294114 55092 294386 55324
rect -1944 54652 -1672 54884
rect 293634 54652 293906 54884
rect -1464 54212 -1192 54444
rect 293154 54212 293426 54444
rect -984 53772 -712 54004
rect 292674 53772 292946 54004
rect -4344 46852 -4072 47084
rect 296034 46852 296306 47084
rect -3864 46412 -3592 46644
rect 295554 46412 295826 46644
rect -2904 45972 -2632 46204
rect 294594 45972 294866 46204
rect -3384 45532 -3112 45764
rect 295074 45532 295346 45764
rect -2424 45092 -2152 45324
rect 294114 45092 294386 45324
rect -1944 44652 -1672 44884
rect 293634 44652 293906 44884
rect -1464 44212 -1192 44444
rect 293154 44212 293426 44444
rect -984 43772 -712 44004
rect 292674 43772 292946 44004
rect -4344 36852 -4072 37084
rect 296034 36852 296306 37084
rect -3864 36412 -3592 36644
rect 295554 36412 295826 36644
rect -2904 35972 -2632 36204
rect 294594 35972 294866 36204
rect 295074 35532 295346 35764
rect -2424 35092 -2152 35324
rect 294114 35092 294386 35324
rect -1944 34652 -1672 34884
rect 293634 34652 293906 34884
rect -1464 34212 -1192 34444
rect 293154 34212 293426 34444
rect -984 33772 -712 34004
rect 292674 33772 292946 34004
rect -4344 26852 -4072 27084
rect 296034 26852 296306 27084
rect -3864 26412 -3592 26644
rect 295554 26412 295826 26644
rect -2904 25972 -2632 26204
rect 294594 25972 294866 26204
rect -3384 25532 -3112 25764
rect 295074 25532 295346 25764
rect -2424 25092 -2152 25324
rect 294114 25092 294386 25324
rect -1944 24652 -1672 24884
rect 293634 24652 293906 24884
rect -1464 24212 -1192 24444
rect 293154 24212 293426 24444
rect -984 23772 -712 24004
rect 292674 23772 292946 24004
rect -4344 16852 -4072 17084
rect 296034 16852 296306 17084
rect -3864 16412 -3592 16644
rect 295554 16412 295826 16644
rect 294594 15972 294866 16204
rect -3384 15532 -3112 15764
rect 295074 15532 295346 15764
rect -2424 15092 -2152 15324
rect 294114 15092 294386 15324
rect -1944 14652 -1672 14884
rect 293634 14652 293906 14884
rect -1464 14212 -1192 14444
rect 293154 14212 293426 14444
rect -984 13772 -712 14004
rect 292674 13772 292946 14004
<< properties >>
string FIXED_BBOX 0 0 100 100
<< end >>
