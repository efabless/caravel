VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gpio_control_block
  CLASS BLOCK ;
  FOREIGN gpio_control_block ;
  ORIGIN 0.000 0.000 ;
  SIZE 170.000 BY 70.000 ;
  PIN gpio_defaults[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 8.200 170.000 8.800 ;
    END
  END gpio_defaults[0]
  PIN gpio_defaults[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 24.520 170.000 25.120 ;
    END
  END gpio_defaults[10]
  PIN gpio_defaults[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 26.560 170.000 27.160 ;
    END
  END gpio_defaults[11]
  PIN gpio_defaults[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 27.920 170.000 28.520 ;
    END
  END gpio_defaults[12]
  PIN gpio_defaults[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 10.240 170.000 10.840 ;
    END
  END gpio_defaults[1]
  PIN gpio_defaults[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 11.600 170.000 12.200 ;
    END
  END gpio_defaults[2]
  PIN gpio_defaults[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 13.640 170.000 14.240 ;
    END
  END gpio_defaults[3]
  PIN gpio_defaults[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 15.000 170.000 15.600 ;
    END
  END gpio_defaults[4]
  PIN gpio_defaults[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 16.360 170.000 16.960 ;
    END
  END gpio_defaults[5]
  PIN gpio_defaults[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 18.400 170.000 19.000 ;
    END
  END gpio_defaults[6]
  PIN gpio_defaults[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 19.760 170.000 20.360 ;
    END
  END gpio_defaults[7]
  PIN gpio_defaults[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 21.800 170.000 22.400 ;
    END
  END gpio_defaults[8]
  PIN gpio_defaults[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 23.160 170.000 23.760 ;
    END
  END gpio_defaults[9]
  PIN mgmt_gpio_in
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 3.440 170.000 4.040 ;
    END
  END mgmt_gpio_in
  PIN mgmt_gpio_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 5.480 170.000 6.080 ;
    END
  END mgmt_gpio_oeb
  PIN mgmt_gpio_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 6.840 170.000 7.440 ;
    END
  END mgmt_gpio_out
  PIN one
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 2.080 170.000 2.680 ;
    END
  END one
  PIN pad_gpio_ana_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 29.960 170.000 30.560 ;
    END
  END pad_gpio_ana_en
  PIN pad_gpio_ana_pol
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 31.320 170.000 31.920 ;
    END
  END pad_gpio_ana_pol
  PIN pad_gpio_ana_sel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 32.680 170.000 33.280 ;
    END
  END pad_gpio_ana_sel
  PIN pad_gpio_dm[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 34.720 170.000 35.320 ;
    END
  END pad_gpio_dm[0]
  PIN pad_gpio_dm[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 36.080 170.000 36.680 ;
    END
  END pad_gpio_dm[1]
  PIN pad_gpio_dm[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 38.120 170.000 38.720 ;
    END
  END pad_gpio_dm[2]
  PIN pad_gpio_holdover
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 39.480 170.000 40.080 ;
    END
  END pad_gpio_holdover
  PIN pad_gpio_ib_mode_sel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 40.840 170.000 41.440 ;
    END
  END pad_gpio_ib_mode_sel
  PIN pad_gpio_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 42.880 170.000 43.480 ;
    END
  END pad_gpio_in
  PIN pad_gpio_inenb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 44.240 170.000 44.840 ;
    END
  END pad_gpio_inenb
  PIN pad_gpio_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 46.280 170.000 46.880 ;
    END
  END pad_gpio_out
  PIN pad_gpio_outenb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 47.640 170.000 48.240 ;
    END
  END pad_gpio_outenb
  PIN pad_gpio_slow_sel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 49.000 170.000 49.600 ;
    END
  END pad_gpio_slow_sel
  PIN pad_gpio_vtrip_sel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 51.040 170.000 51.640 ;
    END
  END pad_gpio_vtrip_sel
  PIN resetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 52.400 170.000 53.000 ;
    END
  END resetn
  PIN resetn_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 54.440 170.000 55.040 ;
    END
  END resetn_out
  PIN serial_clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 55.800 170.000 56.400 ;
    END
  END serial_clock
  PIN serial_clock_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 57.160 170.000 57.760 ;
    END
  END serial_clock_out
  PIN serial_data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 59.200 170.000 59.800 ;
    END
  END serial_data_in
  PIN serial_data_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 60.560 170.000 61.160 ;
    END
  END serial_data_out
  PIN serial_load
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 62.600 170.000 63.200 ;
    END
  END serial_load
  PIN serial_load_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 63.960 170.000 64.560 ;
    END
  END serial_load_out
  PIN user_gpio_in
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 65.320 170.000 65.920 ;
    END
  END user_gpio_in
  PIN user_gpio_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 67.360 170.000 67.960 ;
    END
  END user_gpio_oeb
  PIN user_gpio_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 68.720 170.000 69.320 ;
    END
  END user_gpio_out
  PIN vccd
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 1.800 8.080 52.020 9.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -1.500 12.080 55.320 13.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -1.500 27.580 55.320 29.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -1.500 43.080 55.320 44.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.800 58.320 52.020 59.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.800 8.080 3.400 59.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.420 8.080 52.020 59.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 12.800 4.780 14.400 63.220 ;
    END
    PORT
      LAYER met4 ;
        RECT 28.300 4.780 29.900 63.220 ;
    END
    PORT
      LAYER met4 ;
        RECT 43.800 4.780 45.400 63.220 ;
    END
  END vccd
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -4.800 1.480 58.620 3.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -8.100 16.580 61.920 18.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -8.100 32.080 61.920 33.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -8.100 47.580 61.920 49.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.800 64.920 58.620 66.520 ;
    END
    PORT
      LAYER met4 ;
        RECT -4.800 1.480 -3.200 66.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 57.020 1.480 58.620 66.520 ;
    END
  END vccd1
  PIN vssd
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -1.500 4.780 55.320 6.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -1.500 19.830 55.320 21.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -1.500 35.330 55.320 36.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -1.500 50.830 55.320 52.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -1.500 61.620 55.320 63.220 ;
    END
    PORT
      LAYER met4 ;
        RECT -1.500 4.780 0.100 63.220 ;
    END
    PORT
      LAYER met4 ;
        RECT 20.550 4.780 22.150 63.220 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.050 4.780 37.650 63.220 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.720 4.780 55.320 63.220 ;
    END
  END vssd
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -8.100 -1.820 61.920 -0.220 ;
    END
    PORT
      LAYER met5 ;
        RECT -8.100 24.330 61.920 25.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -8.100 39.830 61.920 41.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -8.100 68.220 61.920 69.820 ;
    END
    PORT
      LAYER met4 ;
        RECT -8.100 -1.820 -6.500 69.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.320 -1.820 61.920 69.820 ;
    END
  END vssd1
  PIN zero
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 0.720 170.000 1.320 ;
    END
  END zero
  OBS
      LAYER li1 ;
        RECT 4.600 10.795 49.535 57.205 ;
      LAYER met1 ;
        RECT 4.600 9.900 114.010 59.800 ;
      LAYER met2 ;
        RECT 5.150 0.835 113.990 69.205 ;
      LAYER met3 ;
        RECT 5.125 66.960 69.600 69.185 ;
        RECT 5.125 66.320 70.000 66.960 ;
        RECT 5.125 62.200 69.600 66.320 ;
        RECT 5.125 61.560 70.000 62.200 ;
        RECT 5.125 58.800 69.600 61.560 ;
        RECT 5.125 58.160 70.000 58.800 ;
        RECT 5.125 54.040 69.600 58.160 ;
        RECT 5.125 53.400 70.000 54.040 ;
        RECT 5.125 50.640 69.600 53.400 ;
        RECT 5.125 50.000 70.000 50.640 ;
        RECT 5.125 45.880 69.600 50.000 ;
        RECT 5.125 45.240 70.000 45.880 ;
        RECT 5.125 42.480 69.600 45.240 ;
        RECT 5.125 41.840 70.000 42.480 ;
        RECT 5.125 37.720 69.600 41.840 ;
        RECT 5.125 37.080 70.000 37.720 ;
        RECT 5.125 34.320 69.600 37.080 ;
        RECT 5.125 33.680 70.000 34.320 ;
        RECT 5.125 29.560 69.600 33.680 ;
        RECT 5.125 28.920 70.000 29.560 ;
        RECT 5.125 26.160 69.600 28.920 ;
        RECT 5.125 25.520 70.000 26.160 ;
        RECT 5.125 21.400 69.600 25.520 ;
        RECT 5.125 20.760 70.000 21.400 ;
        RECT 5.125 18.000 69.600 20.760 ;
        RECT 5.125 17.360 70.000 18.000 ;
        RECT 5.125 13.240 69.600 17.360 ;
        RECT 5.125 12.600 70.000 13.240 ;
        RECT 5.125 9.840 69.600 12.600 ;
        RECT 5.125 9.200 70.000 9.840 ;
        RECT 5.125 5.080 69.600 9.200 ;
        RECT 5.125 4.440 70.000 5.080 ;
        RECT 5.125 0.855 69.600 4.440 ;
      LAYER met4 ;
        RECT 6.280 13.160 11.380 27.240 ;
  END
END gpio_control_block
END LIBRARY

