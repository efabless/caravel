magic
tech sky130A
magscale 1 2
timestamp 1665967863
<< locali >>
rect 676332 721460 676338 721678
rect 41261 602778 41267 602996
rect 41261 601582 41267 601800
rect 41261 600386 41267 600604
rect 41261 599190 41267 599408
rect 41261 597994 41267 598212
rect 676332 447436 676338 447654
rect 676332 446240 676338 446458
rect 676332 445044 676338 445262
rect 676332 443848 676338 444066
rect 676332 442652 676338 442870
rect 676332 441456 676338 441674
rect 676332 440260 676338 440478
rect 41283 345197 41289 345415
rect 41283 344001 41289 344219
rect 41283 342805 41289 343023
rect 41283 341609 41289 341827
rect 41283 340413 41289 340631
rect 41283 339217 41289 339435
rect 41283 338021 41289 338239
rect 41283 336825 41289 337043
rect 41283 335629 41289 335847
rect 134848 43204 135066 43210
rect 136044 43204 136262 43210
rect 137240 43204 137458 43210
rect 138436 43204 138654 43210
rect 139632 43204 139850 43210
rect 140828 43204 141046 43210
rect 142024 43204 142242 43210
rect 143220 43204 143438 43210
rect 144416 43204 144634 43210
rect 152788 43204 153006 43210
rect 153984 43204 154202 43210
rect 155180 43204 155398 43210
rect 156376 43204 156594 43210
rect 157572 43204 157790 43210
rect 158768 43204 158986 43210
rect 430248 43204 430466 43210
rect 431444 43204 431662 43210
rect 432640 43204 432858 43210
rect 433836 43204 434054 43210
rect 435032 43204 435250 43210
rect 436228 43204 436446 43210
rect 437424 43204 437642 43210
rect 438620 43204 438838 43210
rect 439816 43204 440034 43210
rect 448188 43204 448406 43210
rect 449384 43204 449602 43210
rect 450580 43204 450798 43210
rect 451776 43204 451994 43210
rect 452972 43204 453190 43210
rect 454168 43204 454386 43210
<< viali >>
rect 676338 721460 676372 721678
rect 676882 721362 677052 721396
rect 676270 720716 676440 720750
rect 676950 720534 676984 720752
rect 41227 602778 41261 602996
rect 40547 602680 40717 602714
rect 40615 601852 40649 602070
rect 41159 602034 41329 602068
rect 41227 601582 41261 601800
rect 40547 601484 40717 601518
rect 40615 600656 40649 600874
rect 41159 600838 41329 600872
rect 41227 600386 41261 600604
rect 40547 600288 40717 600322
rect 40615 599460 40649 599678
rect 41159 599642 41329 599676
rect 41227 599190 41261 599408
rect 40547 599092 40717 599126
rect 40615 598264 40649 598482
rect 41159 598446 41329 598480
rect 41227 597994 41261 598212
rect 40547 597896 40717 597930
rect 40615 597068 40649 597286
rect 41159 597250 41329 597284
rect 676338 447436 676372 447654
rect 676882 447338 677052 447372
rect 676270 446692 676440 446726
rect 676950 446510 676984 446728
rect 676338 446240 676372 446458
rect 676882 446142 677052 446176
rect 676270 445496 676440 445530
rect 676950 445314 676984 445532
rect 676338 445044 676372 445262
rect 676882 444946 677052 444980
rect 676270 444300 676440 444334
rect 676950 444118 676984 444336
rect 676338 443848 676372 444066
rect 676882 443750 677052 443784
rect 676270 443104 676440 443138
rect 676950 442922 676984 443140
rect 676338 442652 676372 442870
rect 676882 442554 677052 442588
rect 676270 441908 676440 441942
rect 676950 441726 676984 441944
rect 676338 441456 676372 441674
rect 676882 441358 677052 441392
rect 676270 440712 676440 440746
rect 676950 440530 676984 440748
rect 676338 440260 676372 440478
rect 676882 440162 677052 440196
rect 676270 439516 676440 439550
rect 676950 439334 676984 439552
rect 41249 345197 41283 345415
rect 40569 345099 40739 345133
rect 40637 344271 40671 344489
rect 41181 344453 41351 344487
rect 41249 344001 41283 344219
rect 40569 343903 40739 343937
rect 40637 343075 40671 343293
rect 41181 343257 41351 343291
rect 41249 342805 41283 343023
rect 40569 342707 40739 342741
rect 40637 341879 40671 342097
rect 41181 342061 41351 342095
rect 41249 341609 41283 341827
rect 40569 341511 40739 341545
rect 40637 340683 40671 340901
rect 41181 340865 41351 340899
rect 41249 340413 41283 340631
rect 40569 340315 40739 340349
rect 40637 339487 40671 339705
rect 41181 339669 41351 339703
rect 41249 339217 41283 339435
rect 40569 339119 40739 339153
rect 40637 338291 40671 338509
rect 41181 338473 41351 338507
rect 41249 338021 41283 338239
rect 40569 337923 40739 337957
rect 40637 337095 40671 337313
rect 41181 337277 41351 337311
rect 41249 336825 41283 337043
rect 40569 336727 40739 336761
rect 40637 335899 40671 336117
rect 41181 336081 41351 336115
rect 41249 335629 41283 335847
rect 40569 335531 40739 335565
rect 40637 334703 40671 334921
rect 41181 334885 41351 334919
rect 134104 43102 134138 43272
rect 134848 43170 135066 43204
rect 135300 43102 135334 43272
rect 136044 43170 136262 43204
rect 136496 43102 136530 43272
rect 137240 43170 137458 43204
rect 137692 43102 137726 43272
rect 138436 43170 138654 43204
rect 138888 43102 138922 43272
rect 139632 43170 139850 43204
rect 140084 43102 140118 43272
rect 140828 43170 141046 43204
rect 141280 43102 141314 43272
rect 142024 43170 142242 43204
rect 142476 43102 142510 43272
rect 143220 43170 143438 43204
rect 143672 43102 143706 43272
rect 144416 43170 144634 43204
rect 152044 43102 152078 43272
rect 152788 43170 153006 43204
rect 153240 43102 153274 43272
rect 153984 43170 154202 43204
rect 154436 43102 154470 43272
rect 155180 43170 155398 43204
rect 155632 43102 155666 43272
rect 156376 43170 156594 43204
rect 156828 43102 156862 43272
rect 157572 43170 157790 43204
rect 158024 43102 158058 43272
rect 158768 43170 158986 43204
rect 429504 43102 429538 43272
rect 430248 43170 430466 43204
rect 430700 43102 430734 43272
rect 431444 43170 431662 43204
rect 431896 43102 431930 43272
rect 432640 43170 432858 43204
rect 433092 43102 433126 43272
rect 433836 43170 434054 43204
rect 434288 43102 434322 43272
rect 435032 43170 435250 43204
rect 435484 43102 435518 43272
rect 436228 43170 436446 43204
rect 436680 43102 436714 43272
rect 437424 43170 437642 43204
rect 437876 43102 437910 43272
rect 438620 43170 438838 43204
rect 439072 43102 439106 43272
rect 439816 43170 440034 43204
rect 447444 43102 447478 43272
rect 448188 43170 448406 43204
rect 448640 43102 448674 43272
rect 449384 43170 449602 43204
rect 449836 43102 449870 43272
rect 450580 43170 450798 43204
rect 451032 43102 451066 43272
rect 451776 43170 451994 43204
rect 452228 43102 452262 43272
rect 452972 43170 453190 43204
rect 453424 43102 453458 43272
rect 454168 43170 454386 43204
rect 135118 42558 135336 42592
rect 135946 42490 135980 42660
rect 136314 42558 136532 42592
rect 137142 42490 137176 42660
rect 137510 42558 137728 42592
rect 138338 42490 138372 42660
rect 138706 42558 138924 42592
rect 139534 42490 139568 42660
rect 139902 42558 140120 42592
rect 140730 42490 140764 42660
rect 141098 42558 141316 42592
rect 141926 42490 141960 42660
rect 142294 42558 142512 42592
rect 143122 42490 143156 42660
rect 143490 42558 143708 42592
rect 144318 42490 144352 42660
rect 144686 42558 144904 42592
rect 145514 42490 145548 42660
rect 153058 42558 153276 42592
rect 153886 42490 153920 42660
rect 154254 42558 154472 42592
rect 155082 42490 155116 42660
rect 155450 42558 155668 42592
rect 156278 42490 156312 42660
rect 156646 42558 156864 42592
rect 157474 42490 157508 42660
rect 158024 42490 158058 42660
rect 158668 42558 158886 42592
rect 430518 42558 430736 42592
rect 431346 42490 431380 42660
rect 431714 42558 431932 42592
rect 432542 42490 432576 42660
rect 432910 42558 433128 42592
rect 433738 42490 433772 42660
rect 434106 42558 434324 42592
rect 434934 42490 434968 42660
rect 435302 42558 435520 42592
rect 436130 42490 436164 42660
rect 436498 42558 436716 42592
rect 437326 42490 437360 42660
rect 437694 42558 437912 42592
rect 438522 42490 438556 42660
rect 438890 42558 439108 42592
rect 439718 42490 439752 42660
rect 440086 42558 440304 42592
rect 440914 42490 440948 42660
rect 448458 42558 448676 42592
rect 449286 42490 449320 42660
rect 449654 42558 449872 42592
rect 450482 42490 450516 42660
rect 450850 42558 451068 42592
rect 451678 42490 451712 42660
rect 452046 42558 452264 42592
rect 452874 42490 452908 42660
rect 453424 42490 453458 42660
rect 454068 42558 454286 42592
<< metal1 >>
rect 674044 727707 674072 728121
rect 674044 727679 674128 727707
rect 674100 721423 674128 727679
rect 674156 721617 674184 728321
rect 676069 724853 676165 724882
rect 676069 724496 676093 724853
rect 676153 724496 676165 724853
rect 675525 723657 675621 723694
rect 675525 723300 675546 723657
rect 675606 723300 675621 723657
rect 675525 721688 675621 723300
rect 676069 721680 676165 724496
rect 677157 724853 677253 724894
rect 677157 724496 677175 724853
rect 677235 724496 677253 724853
rect 676613 723657 676709 723700
rect 676613 723300 676634 723657
rect 676694 723300 676709 723657
rect 676328 721678 676380 721690
rect 676613 721682 676709 723300
rect 677157 721682 677253 724496
rect 674156 721611 674208 721617
rect 674156 721553 674208 721559
rect 676328 721448 676380 721460
rect 674100 721417 674152 721423
rect 674100 721359 674152 721365
rect 676870 721352 676882 721404
rect 677052 721352 677064 721404
rect 674160 720768 674212 720774
rect 674160 720710 674212 720716
rect 674128 720650 674156 720655
rect 674104 720644 674156 720650
rect 674104 720586 674156 720592
rect 40346 604967 40442 604988
rect 40346 604610 40371 604967
rect 40431 604610 40442 604967
rect 40346 603012 40442 604610
rect 41434 604967 41530 604988
rect 41434 604610 41453 604967
rect 41513 604610 41530 604967
rect 40890 603771 40986 603804
rect 40890 603414 40912 603771
rect 40972 603414 40986 603771
rect 40890 603004 40986 603414
rect 41434 603012 41530 604610
rect 41978 603771 42074 603806
rect 41978 603414 42000 603771
rect 42060 603414 42074 603771
rect 41219 602996 41271 603008
rect 41978 603006 42074 603414
rect 43551 602935 43579 612568
rect 43663 611847 43691 612368
rect 43527 602929 43579 602935
rect 43527 602871 43579 602877
rect 43607 611819 43691 611847
rect 41219 602766 41271 602778
rect 43607 602741 43635 611819
rect 43583 602735 43635 602741
rect 40535 602670 40547 602722
rect 40717 602670 40729 602722
rect 43583 602677 43635 602683
rect 43523 602086 43575 602092
rect 40607 602070 40659 602082
rect 41147 602024 41159 602076
rect 41329 602024 41341 602076
rect 43523 602028 43575 602034
rect 40607 601840 40659 601852
rect 41219 601800 41271 601812
rect 41219 601570 41271 601582
rect 40535 601474 40547 601526
rect 40717 601474 40729 601526
rect 40607 600874 40659 600886
rect 41147 600828 41159 600880
rect 41329 600828 41341 600880
rect 40607 600644 40659 600656
rect 41219 600604 41271 600616
rect 41219 600374 41271 600386
rect 40535 600278 40547 600330
rect 40717 600278 40729 600330
rect 40607 599678 40659 599690
rect 41147 599632 41159 599684
rect 41329 599632 41341 599684
rect 40607 599448 40659 599460
rect 41219 599408 41271 599420
rect 41219 599178 41271 599190
rect 40535 599082 40547 599134
rect 40717 599082 40729 599134
rect 40607 598482 40659 598494
rect 41147 598436 41159 598488
rect 41329 598436 41341 598488
rect 40607 598252 40659 598264
rect 41219 598212 41271 598224
rect 41219 597982 41271 597994
rect 40535 597886 40547 597938
rect 40717 597886 40729 597938
rect 40607 597286 40659 597298
rect 41147 597240 41159 597292
rect 41329 597240 41341 597292
rect 40607 597056 40659 597068
rect 40368 347316 40464 347348
rect 40368 346959 40390 347316
rect 40450 346959 40464 347316
rect 40368 345430 40464 346959
rect 41456 347316 41552 347340
rect 41456 346959 41472 347316
rect 41532 346959 41552 347316
rect 40912 346120 41008 346158
rect 40912 345763 40931 346120
rect 40991 345763 41008 346120
rect 40912 345428 41008 345763
rect 41241 345415 41293 345427
rect 41456 345422 41552 346959
rect 42000 346120 42096 346160
rect 42000 345763 42019 346120
rect 42079 345763 42096 346120
rect 42000 345430 42096 345763
rect 43523 345354 43551 602028
rect 43499 345348 43551 345354
rect 43499 345290 43551 345296
rect 43579 601962 43631 601968
rect 43579 601904 43631 601910
rect 41241 345185 41293 345197
rect 43579 345160 43607 601904
rect 43775 601739 43803 612195
rect 43887 611474 43915 611995
rect 43751 601733 43803 601739
rect 43751 601675 43803 601681
rect 43831 611446 43915 611474
rect 43831 601545 43859 611446
rect 43807 601539 43859 601545
rect 43807 601481 43859 601487
rect 43555 345154 43607 345160
rect 40557 345089 40569 345141
rect 40739 345089 40751 345141
rect 43555 345096 43607 345102
rect 43747 600890 43799 600896
rect 43747 600832 43799 600838
rect 43495 344505 43547 344511
rect 40629 344489 40681 344501
rect 41169 344443 41181 344495
rect 41351 344443 41363 344495
rect 43495 344447 43547 344453
rect 40629 344259 40681 344271
rect 41241 344219 41293 344231
rect 41241 343989 41293 344001
rect 40557 343893 40569 343945
rect 40739 343893 40751 343945
rect 40629 343293 40681 343305
rect 41169 343247 41181 343299
rect 41351 343247 41363 343299
rect 40629 343133 40637 343161
rect 40671 343133 40681 343161
rect 40629 343063 40681 343075
rect 41241 343023 41293 343035
rect 41241 342793 41293 342805
rect 40557 342697 40569 342749
rect 40739 342697 40751 342749
rect 40629 342097 40681 342109
rect 41169 342051 41181 342103
rect 41351 342051 41363 342103
rect 40629 341867 40681 341879
rect 41241 341827 41293 341839
rect 41241 341597 41293 341609
rect 40557 341501 40569 341553
rect 40739 341501 40751 341553
rect 40629 340901 40681 340913
rect 41169 340855 41181 340907
rect 41351 340855 41363 340907
rect 40629 340671 40681 340683
rect 41241 340631 41293 340643
rect 41241 340401 41293 340413
rect 40557 340305 40569 340357
rect 40739 340305 40751 340357
rect 40629 339705 40681 339717
rect 41169 339659 41181 339711
rect 41351 339659 41363 339711
rect 40629 339475 40681 339487
rect 41241 339435 41293 339447
rect 41241 339205 41293 339217
rect 40557 339109 40569 339161
rect 40739 339109 40751 339161
rect 40629 338509 40681 338521
rect 41169 338463 41181 338515
rect 41351 338463 41363 338515
rect 40629 338279 40681 338291
rect 41241 338239 41293 338251
rect 41241 338009 41293 338021
rect 40557 337913 40569 337965
rect 40739 337913 40751 337965
rect 40629 337313 40681 337325
rect 41169 337267 41181 337319
rect 41351 337267 41363 337319
rect 40629 337083 40681 337095
rect 41241 337043 41293 337055
rect 41241 336813 41293 336825
rect 40557 336717 40569 336769
rect 40739 336717 40751 336769
rect 40629 336117 40681 336129
rect 41169 336071 41181 336123
rect 41351 336071 41363 336123
rect 40629 335887 40681 335899
rect 41241 335847 41293 335859
rect 41241 335617 41293 335629
rect 40557 335521 40569 335573
rect 40739 335521 40751 335573
rect 40629 334921 40681 334933
rect 41169 334875 41181 334927
rect 41351 334875 41363 334927
rect 40629 334691 40681 334703
rect 43495 46196 43523 344447
rect 43551 344381 43603 344387
rect 43551 344323 43603 344329
rect 43551 46252 43579 344323
rect 43747 344158 43775 600832
rect 43723 344152 43775 344158
rect 43723 344094 43775 344100
rect 43803 600766 43855 600772
rect 43803 600708 43855 600714
rect 43803 343964 43831 600708
rect 43999 600543 44027 611795
rect 44111 611031 44139 611595
rect 43975 600537 44027 600543
rect 43975 600479 44027 600485
rect 44055 611003 44139 611031
rect 44055 600349 44083 611003
rect 44031 600343 44083 600349
rect 44031 600285 44083 600291
rect 43779 343958 43831 343964
rect 43779 343900 43831 343906
rect 43971 599694 44023 599700
rect 43971 599636 44023 599642
rect 43719 343309 43771 343315
rect 43719 343251 43771 343257
rect 43719 46364 43747 343251
rect 43775 343185 43827 343191
rect 43775 343127 43827 343133
rect 43775 46420 43803 343127
rect 43971 342962 43999 599636
rect 43947 342956 43999 342962
rect 43947 342898 43999 342904
rect 44027 599570 44079 599576
rect 44027 599512 44079 599518
rect 44027 342768 44055 599512
rect 44223 599347 44251 611356
rect 44335 610635 44363 611156
rect 44199 599341 44251 599347
rect 44199 599283 44251 599289
rect 44279 610607 44363 610635
rect 44279 599153 44307 610607
rect 44255 599147 44307 599153
rect 44255 599089 44307 599095
rect 44003 342762 44055 342768
rect 44003 342704 44055 342710
rect 44195 598498 44247 598504
rect 44195 598440 44247 598446
rect 43943 342113 43995 342119
rect 43943 342055 43995 342061
rect 43943 46532 43971 342055
rect 43999 341989 44051 341995
rect 43999 341931 44051 341937
rect 43999 46588 44027 341931
rect 44195 341766 44223 598440
rect 44171 341760 44223 341766
rect 44171 341702 44223 341708
rect 44251 598374 44303 598380
rect 44251 598316 44303 598322
rect 44251 341572 44279 598316
rect 44447 598151 44475 610956
rect 44559 610222 44587 610756
rect 44423 598145 44475 598151
rect 44423 598087 44475 598093
rect 44503 610194 44587 610222
rect 44503 597957 44531 610194
rect 44479 597951 44531 597957
rect 44479 597893 44531 597899
rect 44227 341566 44279 341572
rect 44227 341508 44279 341514
rect 44419 597302 44471 597308
rect 44419 597244 44471 597250
rect 44167 340917 44219 340923
rect 44167 340859 44219 340865
rect 44167 46700 44195 340859
rect 44223 340793 44275 340799
rect 44223 340735 44275 340741
rect 44223 46756 44251 340735
rect 44419 340570 44447 597244
rect 44395 340564 44447 340570
rect 44395 340506 44447 340512
rect 44475 597178 44527 597184
rect 44475 597120 44527 597126
rect 44475 340376 44503 597120
rect 672728 453527 672756 454055
rect 672728 453499 672812 453527
rect 672784 440223 672812 453499
rect 672840 440417 672868 454255
rect 672952 453932 672980 454455
rect 672952 453904 673036 453932
rect 673008 441419 673036 453904
rect 673064 441613 673092 454655
rect 673176 454333 673204 454855
rect 673176 454305 673260 454333
rect 673232 442615 673260 454305
rect 673288 442809 673316 455055
rect 673400 454779 673428 455255
rect 673400 454751 673484 454779
rect 673456 443811 673484 454751
rect 673512 444005 673540 455455
rect 673624 455131 673652 455655
rect 673624 455103 673708 455131
rect 673680 445007 673708 455103
rect 673736 445201 673764 455855
rect 673848 455533 673876 456055
rect 673848 455505 673932 455533
rect 673904 446203 673932 455505
rect 673960 446397 673988 456255
rect 674128 447399 674156 720586
rect 674184 447593 674212 720710
rect 676258 720706 676270 720758
rect 676440 720706 676452 720758
rect 676940 720752 676992 720764
rect 676940 720522 676992 720534
rect 676069 448452 676165 448478
rect 676069 448095 676085 448452
rect 676145 448095 676165 448452
rect 676069 447672 676165 448095
rect 677157 448452 677253 448476
rect 677157 448095 677167 448452
rect 677227 448095 677253 448452
rect 677157 447670 677253 448095
rect 676328 447654 676380 447666
rect 674184 447587 674236 447593
rect 674184 447529 674236 447535
rect 676328 447424 676380 447436
rect 674128 447393 674180 447399
rect 674128 447335 674180 447341
rect 676870 447328 676882 447380
rect 677052 447328 677064 447380
rect 674188 446744 674240 446750
rect 674188 446686 674240 446692
rect 674132 446620 674184 446626
rect 674132 446562 674184 446568
rect 673960 446391 674012 446397
rect 673960 446333 674012 446339
rect 673904 446197 673956 446203
rect 673904 446139 673956 446145
rect 673964 445548 674016 445554
rect 673964 445490 674016 445496
rect 673908 445424 673960 445430
rect 673908 445366 673960 445372
rect 673736 445195 673788 445201
rect 673736 445137 673788 445143
rect 673680 445001 673732 445007
rect 673680 444943 673732 444949
rect 673740 444352 673792 444358
rect 673740 444294 673792 444300
rect 673684 444228 673736 444234
rect 673684 444170 673736 444176
rect 673512 443999 673564 444005
rect 673512 443941 673564 443947
rect 673456 443805 673508 443811
rect 673456 443747 673508 443753
rect 673516 443156 673568 443162
rect 673516 443098 673568 443104
rect 673460 443032 673512 443038
rect 673460 442974 673512 442980
rect 673288 442803 673340 442809
rect 673288 442745 673340 442751
rect 673232 442609 673284 442615
rect 673232 442551 673284 442557
rect 673292 441960 673344 441966
rect 673292 441902 673344 441908
rect 673236 441836 673288 441842
rect 673236 441778 673288 441784
rect 673064 441607 673116 441613
rect 673064 441549 673116 441555
rect 673008 441413 673060 441419
rect 673008 441355 673060 441361
rect 673068 440764 673120 440770
rect 673068 440706 673120 440712
rect 673012 440640 673064 440646
rect 673012 440582 673064 440588
rect 672840 440411 672892 440417
rect 672840 440353 672892 440359
rect 672784 440217 672836 440223
rect 672784 440159 672836 440165
rect 672844 439568 672896 439574
rect 672844 439510 672896 439516
rect 672788 439444 672840 439450
rect 672788 439386 672840 439392
rect 44451 340370 44503 340376
rect 44451 340312 44503 340318
rect 44391 339721 44443 339727
rect 44391 339663 44443 339669
rect 44391 46868 44419 339663
rect 44447 339597 44499 339603
rect 44447 339539 44499 339545
rect 44447 46924 44475 339539
rect 44643 339374 44671 354730
rect 44755 353903 44783 354530
rect 44619 339368 44671 339374
rect 44619 339310 44671 339316
rect 44699 353875 44783 353903
rect 44699 339180 44727 353875
rect 44675 339174 44727 339180
rect 44675 339116 44727 339122
rect 44615 338525 44667 338531
rect 44615 338467 44667 338473
rect 44615 47036 44643 338467
rect 44671 338401 44723 338407
rect 44671 338343 44723 338349
rect 44671 47092 44699 338343
rect 44867 338178 44895 354330
rect 44979 353506 45007 354130
rect 44843 338172 44895 338178
rect 44843 338114 44895 338120
rect 44923 353478 45007 353506
rect 44923 337984 44951 353478
rect 44899 337978 44951 337984
rect 44899 337920 44951 337926
rect 44839 337329 44891 337335
rect 44839 337271 44891 337277
rect 44839 47204 44867 337271
rect 44895 337205 44947 337211
rect 44895 337147 44947 337153
rect 44895 47260 44923 337147
rect 45091 336958 45119 353930
rect 45203 353120 45231 353730
rect 45067 336952 45119 336958
rect 45067 336894 45119 336900
rect 45147 353092 45231 353120
rect 45147 336788 45175 353092
rect 45123 336782 45175 336788
rect 45123 336724 45175 336730
rect 45063 336133 45115 336139
rect 45063 336075 45115 336081
rect 45063 47372 45091 336075
rect 45119 336009 45171 336015
rect 45119 335951 45171 335957
rect 45119 47428 45147 335951
rect 45315 335786 45343 353530
rect 45427 352705 45455 353330
rect 45291 335780 45343 335786
rect 45291 335722 45343 335728
rect 45371 352677 45455 352705
rect 45371 335592 45399 352677
rect 45347 335586 45399 335592
rect 45347 335528 45399 335534
rect 45287 334937 45339 334943
rect 45287 334879 45339 334885
rect 45287 47540 45315 334879
rect 45343 334813 45395 334819
rect 45343 334755 45395 334761
rect 45343 47596 45371 334755
rect 672812 237645 672840 439386
rect 672756 237617 672840 237645
rect 672756 237050 672784 237617
rect 672868 236850 672896 439510
rect 673036 237300 673064 440582
rect 672980 237272 673064 237300
rect 672980 236650 673008 237272
rect 673092 236450 673120 440706
rect 673260 236897 673288 441778
rect 673204 236869 673288 236897
rect 673204 236250 673232 236869
rect 673316 236050 673344 441902
rect 673484 236488 673512 442974
rect 673428 236460 673512 236488
rect 673428 235850 673456 236460
rect 673540 235650 673568 443098
rect 673708 236094 673736 444170
rect 673652 236066 673736 236094
rect 673652 235450 673680 236066
rect 673764 235250 673792 444294
rect 673932 235700 673960 445366
rect 673876 235672 673960 235700
rect 673876 235050 673904 235672
rect 673988 234850 674016 445490
rect 674156 235298 674184 446562
rect 674100 235270 674184 235298
rect 674100 234650 674128 235270
rect 674212 234450 674240 446686
rect 676258 446682 676270 446734
rect 676440 446682 676452 446734
rect 676940 446728 676992 446740
rect 676940 446498 676992 446510
rect 676328 446458 676380 446470
rect 676328 446228 676380 446240
rect 676870 446132 676882 446184
rect 677052 446132 677064 446184
rect 676258 445486 676270 445538
rect 676440 445486 676452 445538
rect 676940 445532 676992 445544
rect 676940 445302 676992 445314
rect 676328 445262 676380 445274
rect 676328 445032 676380 445044
rect 676870 444936 676882 444988
rect 677052 444936 677064 444988
rect 676258 444290 676270 444342
rect 676440 444290 676452 444342
rect 676940 444336 676992 444348
rect 676940 444106 676992 444118
rect 676328 444066 676380 444078
rect 676328 443836 676380 443848
rect 676870 443740 676882 443792
rect 677052 443740 677064 443792
rect 676258 443094 676270 443146
rect 676440 443094 676452 443146
rect 676940 443140 676992 443152
rect 676940 442910 676992 442922
rect 676328 442870 676380 442882
rect 676328 442640 676380 442652
rect 676870 442544 676882 442596
rect 677052 442544 677064 442596
rect 676258 441898 676270 441950
rect 676440 441898 676452 441950
rect 676940 441944 676992 441956
rect 676940 441714 676992 441726
rect 676328 441674 676380 441686
rect 676328 441444 676380 441456
rect 676870 441348 676882 441400
rect 677052 441348 677064 441400
rect 676258 440702 676270 440754
rect 676440 440702 676452 440754
rect 676940 440748 676992 440760
rect 676940 440518 676992 440530
rect 676328 440478 676380 440490
rect 676328 440248 676380 440260
rect 676870 440152 676882 440204
rect 677052 440152 677064 440204
rect 676258 439506 676270 439558
rect 676440 439506 676452 439558
rect 676940 439552 676992 439564
rect 676940 439322 676992 439334
rect 674240 228608 674268 229288
rect 674240 228580 674324 228608
rect 429498 47624 429504 47648
rect 134098 47596 134104 47620
rect 45343 47568 134104 47596
rect 134156 47568 134162 47620
rect 134941 47572 134947 47624
rect 134999 47596 141269 47624
rect 134999 47572 135005 47596
rect 135170 47540 135176 47564
rect 45287 47512 135176 47540
rect 135228 47512 135234 47564
rect 135943 47516 135949 47568
rect 136001 47540 141213 47568
rect 136001 47516 136007 47540
rect 135294 47428 135300 47452
rect 45119 47400 135300 47428
rect 135352 47400 135358 47452
rect 136137 47404 136143 47456
rect 136195 47428 141101 47456
rect 136195 47404 136201 47428
rect 136366 47372 136372 47396
rect 45063 47344 136372 47372
rect 136424 47344 136430 47396
rect 137139 47348 137145 47400
rect 137197 47372 141045 47400
rect 137197 47348 137203 47372
rect 136490 47260 136496 47284
rect 44895 47232 136496 47260
rect 136548 47232 136554 47284
rect 137333 47236 137339 47288
rect 137391 47260 140933 47288
rect 137391 47236 137397 47260
rect 137562 47204 137568 47228
rect 44839 47176 137568 47204
rect 137620 47176 137626 47228
rect 138335 47180 138341 47232
rect 138393 47204 140877 47232
rect 138393 47180 138399 47204
rect 137686 47092 137692 47116
rect 44671 47064 137692 47092
rect 137744 47064 137750 47116
rect 138529 47068 138535 47120
rect 138587 47092 140765 47120
rect 138587 47068 138593 47092
rect 138758 47036 138764 47060
rect 44615 47008 138764 47036
rect 138816 47008 138822 47060
rect 139531 47012 139537 47064
rect 139589 47036 140709 47064
rect 139589 47012 139595 47036
rect 138882 46924 138888 46948
rect 44447 46896 138888 46924
rect 138940 46896 138946 46948
rect 139725 46900 139731 46952
rect 139783 46924 140651 46952
rect 139783 46900 139789 46924
rect 139954 46868 139960 46892
rect 44391 46840 139960 46868
rect 140012 46840 140018 46892
rect 140078 46756 140084 46780
rect 44223 46728 140084 46756
rect 140136 46728 140142 46780
rect 44167 46672 140585 46700
rect 43999 46560 140526 46588
rect 43943 46504 140462 46532
rect 43775 46392 140403 46420
rect 43719 46336 140347 46364
rect 43551 46224 140287 46252
rect 43495 46168 140231 46196
rect 140203 46084 140231 46168
rect 140259 46140 140287 46224
rect 140319 46196 140347 46336
rect 140375 46252 140403 46392
rect 140434 46308 140462 46504
rect 140498 46364 140526 46560
rect 140557 46420 140585 46672
rect 140623 46616 140651 46924
rect 140681 46672 140709 47036
rect 140737 46728 140765 47092
rect 140849 46784 140877 47204
rect 140905 46840 140933 47260
rect 141017 46896 141045 47372
rect 141073 46952 141101 47428
rect 141185 47008 141213 47540
rect 141241 47064 141269 47596
rect 155603 47596 429504 47624
rect 429556 47596 429562 47648
rect 430341 47600 430347 47652
rect 430399 47624 487832 47652
rect 430399 47600 430405 47624
rect 155603 47064 155631 47596
rect 430570 47568 430576 47592
rect 141241 47036 155631 47064
rect 155659 47540 430576 47568
rect 430628 47540 430634 47592
rect 431343 47544 431349 47596
rect 431401 47568 487776 47596
rect 431401 47544 431407 47568
rect 155659 47008 155687 47540
rect 430694 47456 430700 47480
rect 141185 46980 155687 47008
rect 155771 47428 430700 47456
rect 430752 47428 430758 47480
rect 431537 47432 431543 47484
rect 431595 47456 487608 47484
rect 431595 47432 431601 47456
rect 155771 46952 155799 47428
rect 431766 47400 431772 47424
rect 141073 46924 155799 46952
rect 155827 47372 431772 47400
rect 431824 47372 431830 47424
rect 432539 47376 432545 47428
rect 432597 47400 487552 47428
rect 432597 47376 432603 47400
rect 155827 46896 155855 47372
rect 431890 47288 431896 47312
rect 141017 46868 155855 46896
rect 155939 47260 431896 47288
rect 431948 47260 431954 47312
rect 432733 47264 432739 47316
rect 432791 47288 487384 47316
rect 432791 47264 432797 47288
rect 155939 46840 155967 47260
rect 432962 47232 432968 47256
rect 140905 46812 155967 46840
rect 155995 47204 432968 47232
rect 433020 47204 433026 47256
rect 433735 47208 433741 47260
rect 433793 47232 487328 47260
rect 433793 47208 433799 47232
rect 155995 46784 156023 47204
rect 433086 47120 433092 47144
rect 140849 46756 156023 46784
rect 156107 47092 433092 47120
rect 433144 47092 433150 47144
rect 433929 47096 433935 47148
rect 433987 47120 487160 47148
rect 433987 47096 433993 47120
rect 156107 46728 156135 47092
rect 434158 47064 434164 47088
rect 140737 46700 156135 46728
rect 156163 47036 434164 47064
rect 434216 47036 434222 47088
rect 434931 47040 434937 47092
rect 434989 47064 487104 47092
rect 434989 47040 434995 47064
rect 156163 46672 156191 47036
rect 434282 46952 434288 46976
rect 140681 46644 156191 46672
rect 156275 46924 434288 46952
rect 434340 46924 434346 46976
rect 435125 46928 435131 46980
rect 435183 46952 486936 46980
rect 435183 46928 435189 46952
rect 156275 46616 156303 46924
rect 435354 46896 435360 46920
rect 140623 46588 156303 46616
rect 156331 46868 435360 46896
rect 435412 46868 435418 46920
rect 436127 46872 436133 46924
rect 436185 46896 486880 46924
rect 436185 46872 436191 46896
rect 156331 46560 156359 46868
rect 435478 46784 435484 46808
rect 140727 46508 140733 46560
rect 140785 46532 156359 46560
rect 156443 46756 435484 46784
rect 435536 46756 435542 46808
rect 436297 46760 436303 46812
rect 436355 46784 486712 46812
rect 436355 46760 436361 46784
rect 140785 46508 140791 46532
rect 156443 46504 156471 46756
rect 436550 46728 436556 46752
rect 140897 46452 140903 46504
rect 140955 46476 156471 46504
rect 156499 46700 436556 46728
rect 436608 46700 436614 46752
rect 437323 46704 437329 46756
rect 437381 46728 486656 46756
rect 437381 46704 437387 46728
rect 140955 46452 140961 46476
rect 156499 46448 156527 46700
rect 436674 46616 436680 46640
rect 141150 46420 141156 46444
rect 140557 46392 141156 46420
rect 141208 46392 141214 46444
rect 141923 46396 141929 46448
rect 141981 46420 156527 46448
rect 156611 46588 436680 46616
rect 436732 46588 436738 46640
rect 437517 46592 437523 46644
rect 437575 46616 486488 46644
rect 437575 46592 437581 46616
rect 141981 46396 141987 46420
rect 156611 46392 156639 46588
rect 437746 46560 437752 46584
rect 141274 46364 141280 46388
rect 140498 46336 141280 46364
rect 141332 46336 141338 46388
rect 142117 46340 142123 46392
rect 142175 46364 156639 46392
rect 156667 46532 437752 46560
rect 437804 46532 437810 46584
rect 438519 46536 438525 46588
rect 438577 46560 486432 46588
rect 438577 46536 438583 46560
rect 142175 46340 142181 46364
rect 156667 46336 156695 46532
rect 437870 46448 437876 46472
rect 142346 46308 142352 46332
rect 140434 46280 142352 46308
rect 142404 46280 142410 46332
rect 143119 46284 143125 46336
rect 143177 46308 156695 46336
rect 156779 46420 437876 46448
rect 437928 46420 437934 46472
rect 438689 46424 438695 46476
rect 438747 46448 486264 46476
rect 438747 46424 438753 46448
rect 143177 46284 143183 46308
rect 156779 46280 156807 46420
rect 438942 46392 438948 46416
rect 142470 46252 142476 46276
rect 140375 46224 142476 46252
rect 142528 46224 142534 46276
rect 143289 46228 143295 46280
rect 143347 46252 156807 46280
rect 156835 46364 438948 46392
rect 439000 46364 439006 46416
rect 439715 46368 439721 46420
rect 439773 46392 486208 46420
rect 439773 46368 439779 46392
rect 143347 46228 143353 46252
rect 156835 46224 156863 46364
rect 439066 46280 439072 46304
rect 143542 46196 143548 46220
rect 140319 46168 143548 46196
rect 143600 46168 143606 46220
rect 144315 46172 144321 46224
rect 144373 46196 156863 46224
rect 156947 46252 439072 46280
rect 439124 46252 439130 46304
rect 439909 46256 439915 46308
rect 439967 46280 486040 46308
rect 439967 46256 439973 46280
rect 144373 46172 144379 46196
rect 156947 46168 156975 46252
rect 440138 46224 440144 46248
rect 143666 46140 143672 46164
rect 140259 46112 143672 46140
rect 143724 46112 143730 46164
rect 144509 46116 144515 46168
rect 144567 46140 156975 46168
rect 157003 46196 440144 46224
rect 440196 46196 440202 46248
rect 440911 46200 440917 46252
rect 440969 46224 485984 46252
rect 440969 46200 440975 46224
rect 144567 46116 144573 46140
rect 157003 46112 157031 46196
rect 144738 46084 144744 46108
rect 140203 46056 144744 46084
rect 144796 46056 144802 46108
rect 145511 46060 145517 46112
rect 145569 46084 157031 46112
rect 145569 46060 145575 46084
rect 447438 45104 447444 45128
rect 131151 45076 131920 45104
rect 152038 45076 152044 45100
rect 131892 45048 152044 45076
rect 152096 45048 152102 45100
rect 152881 45052 152887 45104
rect 152939 45076 447444 45104
rect 447496 45076 447502 45128
rect 448281 45080 448287 45132
rect 448339 45104 484472 45132
rect 448339 45080 448345 45104
rect 152939 45052 152945 45076
rect 448510 45048 448516 45072
rect 153110 45020 153116 45044
rect 131323 44992 153116 45020
rect 153168 44992 153174 45044
rect 153883 44996 153889 45048
rect 153941 45020 448516 45048
rect 448568 45020 448574 45072
rect 449283 45024 449289 45076
rect 449341 45048 484416 45076
rect 449341 45024 449347 45048
rect 153941 44996 153947 45020
rect 448634 44936 448640 44960
rect 131551 44908 132328 44936
rect 153234 44908 153240 44932
rect 132300 44880 153240 44908
rect 153292 44880 153298 44932
rect 154077 44884 154083 44936
rect 154135 44908 448640 44936
rect 448692 44908 448698 44960
rect 449477 44912 449483 44964
rect 449535 44936 484248 44964
rect 449535 44912 449541 44936
rect 154135 44884 154141 44908
rect 449706 44880 449712 44904
rect 154306 44852 154312 44876
rect 131723 44824 154312 44852
rect 154364 44824 154370 44876
rect 155079 44828 155085 44880
rect 155137 44852 449712 44880
rect 449764 44852 449770 44904
rect 450479 44856 450485 44908
rect 450537 44880 484192 44908
rect 450537 44856 450543 44880
rect 155137 44828 155143 44852
rect 449830 44768 449836 44792
rect 131951 44740 132727 44768
rect 154430 44740 154436 44764
rect 132699 44712 154436 44740
rect 154488 44712 154494 44764
rect 155249 44716 155255 44768
rect 155307 44740 449836 44768
rect 449888 44740 449894 44792
rect 450649 44744 450655 44796
rect 450707 44768 484024 44796
rect 450707 44744 450713 44768
rect 155307 44716 155313 44740
rect 450902 44712 450908 44736
rect 155502 44684 155508 44708
rect 132123 44656 155508 44684
rect 155560 44656 155566 44708
rect 156275 44660 156281 44712
rect 156333 44684 450908 44712
rect 450960 44684 450966 44736
rect 451675 44688 451681 44740
rect 451733 44712 483968 44740
rect 451733 44688 451739 44712
rect 156333 44660 156339 44684
rect 451026 44600 451032 44624
rect 132351 44572 133117 44600
rect 155626 44572 155632 44596
rect 133089 44544 155632 44572
rect 155684 44544 155690 44596
rect 156469 44548 156475 44600
rect 156527 44572 451032 44600
rect 451084 44572 451090 44624
rect 451869 44576 451875 44628
rect 451927 44600 483800 44628
rect 451927 44576 451933 44600
rect 156527 44548 156533 44572
rect 452098 44544 452104 44568
rect 156698 44516 156704 44540
rect 132523 44488 156704 44516
rect 156756 44488 156762 44540
rect 157471 44492 157477 44544
rect 157529 44516 452104 44544
rect 452156 44516 452162 44568
rect 452871 44520 452877 44572
rect 452929 44544 483744 44572
rect 452929 44520 452935 44544
rect 157529 44492 157535 44516
rect 452222 44432 452228 44456
rect 156822 44404 156828 44428
rect 132723 44376 156828 44404
rect 156880 44376 156886 44428
rect 157641 44380 157647 44432
rect 157699 44404 452228 44432
rect 452280 44404 452286 44456
rect 453041 44408 453047 44460
rect 453099 44432 483576 44460
rect 453099 44408 453105 44432
rect 157699 44380 157705 44404
rect 453294 44320 453300 44344
rect 157894 44292 157900 44316
rect 132923 44264 157900 44292
rect 157952 44264 157958 44316
rect 158667 44268 158673 44320
rect 158725 44292 453300 44320
rect 453352 44292 453358 44344
rect 454067 44296 454073 44348
rect 454125 44320 483408 44348
rect 454125 44296 454131 44320
rect 158725 44268 158731 44292
rect 453418 44208 453424 44232
rect 158018 44180 158024 44204
rect 133123 44152 158024 44180
rect 158076 44152 158082 44204
rect 158861 44156 158867 44208
rect 158919 44180 453424 44208
rect 453476 44180 453482 44232
rect 454261 44184 454267 44236
rect 454319 44208 483240 44236
rect 454319 44184 454325 44208
rect 158919 44156 158925 44180
rect 145832 44004 151750 44017
rect 145832 43944 146199 44004
rect 146556 43944 151750 44004
rect 145832 43921 151750 43944
rect 441228 43921 447154 44017
rect 145840 43457 151748 43473
rect 145840 43397 147395 43457
rect 147752 43397 151748 43457
rect 145840 43377 151748 43397
rect 441228 43450 447154 43473
rect 441228 43390 441626 43450
rect 441983 43390 447154 43450
rect 441228 43377 447154 43390
rect 134094 43272 134146 43284
rect 135290 43272 135342 43284
rect 134836 43162 134848 43214
rect 135066 43162 135078 43214
rect 134094 43090 134146 43102
rect 136486 43272 136538 43284
rect 136032 43162 136044 43214
rect 136262 43162 136274 43214
rect 135290 43090 135342 43102
rect 137682 43272 137734 43284
rect 137228 43162 137240 43214
rect 137458 43162 137470 43214
rect 136486 43090 136538 43102
rect 138878 43272 138930 43284
rect 138424 43162 138436 43214
rect 138654 43162 138666 43214
rect 137682 43090 137734 43102
rect 140074 43272 140126 43284
rect 139620 43162 139632 43214
rect 139850 43162 139862 43214
rect 138878 43090 138930 43102
rect 141270 43272 141322 43284
rect 140816 43162 140828 43214
rect 141046 43162 141058 43214
rect 140074 43090 140126 43102
rect 142466 43272 142518 43284
rect 142012 43162 142024 43214
rect 142242 43162 142254 43214
rect 141270 43090 141322 43102
rect 143662 43272 143714 43284
rect 143208 43162 143220 43214
rect 143438 43162 143450 43214
rect 142466 43090 142518 43102
rect 152034 43272 152086 43284
rect 144404 43162 144416 43214
rect 144634 43162 144646 43214
rect 143662 43090 143714 43102
rect 153230 43272 153282 43284
rect 152776 43162 152788 43214
rect 153006 43162 153018 43214
rect 152034 43090 152086 43102
rect 154426 43272 154478 43284
rect 153972 43162 153984 43214
rect 154202 43162 154214 43214
rect 153230 43090 153282 43102
rect 155622 43272 155674 43284
rect 155168 43162 155180 43214
rect 155398 43162 155410 43214
rect 154426 43090 154478 43102
rect 156818 43272 156870 43284
rect 156364 43162 156376 43214
rect 156594 43162 156606 43214
rect 155622 43090 155674 43102
rect 158014 43272 158066 43284
rect 157560 43162 157572 43214
rect 157790 43162 157802 43214
rect 156818 43090 156870 43102
rect 429494 43272 429546 43284
rect 158756 43162 158768 43214
rect 158986 43162 158998 43214
rect 158014 43090 158066 43102
rect 430690 43272 430742 43284
rect 430236 43162 430248 43214
rect 430466 43162 430478 43214
rect 429494 43090 429546 43102
rect 431886 43272 431938 43284
rect 431432 43162 431444 43214
rect 431662 43162 431674 43214
rect 430690 43090 430742 43102
rect 433082 43272 433134 43284
rect 432628 43162 432640 43214
rect 432858 43162 432870 43214
rect 431886 43090 431938 43102
rect 434278 43272 434330 43284
rect 433824 43162 433836 43214
rect 434054 43162 434066 43214
rect 433082 43090 433134 43102
rect 435474 43272 435526 43284
rect 435020 43162 435032 43214
rect 435250 43162 435262 43214
rect 434278 43090 434330 43102
rect 436670 43272 436722 43284
rect 436216 43162 436228 43214
rect 436446 43162 436458 43214
rect 435474 43090 435526 43102
rect 437866 43272 437918 43284
rect 437412 43162 437424 43214
rect 437642 43162 437654 43214
rect 436670 43090 436722 43102
rect 439062 43272 439114 43284
rect 438608 43162 438620 43214
rect 438838 43162 438850 43214
rect 437866 43090 437918 43102
rect 447434 43272 447486 43284
rect 439804 43162 439816 43214
rect 440034 43162 440046 43214
rect 439062 43090 439114 43102
rect 448630 43272 448682 43284
rect 448176 43162 448188 43214
rect 448406 43162 448418 43214
rect 447434 43090 447486 43102
rect 449826 43272 449878 43284
rect 449372 43162 449384 43214
rect 449602 43162 449614 43214
rect 448630 43090 448682 43102
rect 451022 43272 451074 43284
rect 450568 43162 450580 43214
rect 450798 43162 450810 43214
rect 449826 43090 449878 43102
rect 452218 43272 452270 43284
rect 451764 43162 451776 43214
rect 451994 43162 452006 43214
rect 451022 43090 451074 43102
rect 453414 43272 453466 43284
rect 452960 43162 452972 43214
rect 453190 43162 453202 43214
rect 452218 43090 452270 43102
rect 454156 43162 454168 43214
rect 454386 43162 454398 43214
rect 453414 43090 453466 43102
rect 145840 42916 151748 42929
rect 145840 42856 146199 42916
rect 146556 42856 151748 42916
rect 145840 42833 151748 42856
rect 441228 42833 447154 42929
rect 135936 42660 135988 42672
rect 135106 42550 135118 42602
rect 135336 42550 135348 42602
rect 137132 42660 137184 42672
rect 136302 42550 136314 42602
rect 136532 42550 136544 42602
rect 135936 42478 135988 42490
rect 138328 42660 138380 42672
rect 137498 42550 137510 42602
rect 137728 42550 137740 42602
rect 137132 42478 137184 42490
rect 139524 42660 139576 42672
rect 138694 42550 138706 42602
rect 138924 42550 138936 42602
rect 138328 42478 138380 42490
rect 140720 42660 140772 42672
rect 139890 42550 139902 42602
rect 140120 42550 140132 42602
rect 139524 42478 139576 42490
rect 141916 42660 141968 42672
rect 141086 42550 141098 42602
rect 141316 42550 141328 42602
rect 140720 42478 140772 42490
rect 143112 42660 143164 42672
rect 142282 42550 142294 42602
rect 142512 42550 142524 42602
rect 141916 42478 141968 42490
rect 144308 42660 144360 42672
rect 143478 42550 143490 42602
rect 143708 42550 143720 42602
rect 143112 42478 143164 42490
rect 145504 42660 145556 42672
rect 144674 42550 144686 42602
rect 144904 42550 144916 42602
rect 144308 42478 144360 42490
rect 153876 42660 153928 42672
rect 153046 42550 153058 42602
rect 153276 42550 153288 42602
rect 145504 42478 145556 42490
rect 155072 42660 155124 42672
rect 154242 42550 154254 42602
rect 154472 42550 154484 42602
rect 153876 42478 153928 42490
rect 156268 42660 156320 42672
rect 155438 42550 155450 42602
rect 155668 42550 155680 42602
rect 155072 42478 155124 42490
rect 157464 42660 157516 42672
rect 156634 42550 156646 42602
rect 156864 42550 156876 42602
rect 156268 42478 156320 42490
rect 157464 42478 157516 42490
rect 158016 42660 158068 42672
rect 431336 42660 431388 42672
rect 158656 42550 158668 42602
rect 158886 42550 158898 42602
rect 430506 42550 430518 42602
rect 430736 42550 430748 42602
rect 158016 42478 158068 42490
rect 432532 42660 432584 42672
rect 431702 42550 431714 42602
rect 431932 42550 431944 42602
rect 431336 42478 431388 42490
rect 433728 42660 433780 42672
rect 432898 42550 432910 42602
rect 433128 42550 433140 42602
rect 432532 42478 432584 42490
rect 434924 42660 434976 42672
rect 434094 42550 434106 42602
rect 434324 42550 434336 42602
rect 433728 42478 433780 42490
rect 436120 42660 436172 42672
rect 435290 42550 435302 42602
rect 435520 42550 435532 42602
rect 434924 42478 434976 42490
rect 437316 42660 437368 42672
rect 436486 42550 436498 42602
rect 436716 42550 436728 42602
rect 436120 42478 436172 42490
rect 438512 42660 438564 42672
rect 437682 42550 437694 42602
rect 437912 42550 437924 42602
rect 437316 42478 437368 42490
rect 439708 42660 439760 42672
rect 438878 42550 438890 42602
rect 439108 42550 439120 42602
rect 438512 42478 438564 42490
rect 440904 42660 440956 42672
rect 440074 42550 440086 42602
rect 440304 42550 440316 42602
rect 439708 42478 439760 42490
rect 449276 42660 449328 42672
rect 448446 42550 448458 42602
rect 448676 42550 448688 42602
rect 440904 42478 440956 42490
rect 450472 42660 450524 42672
rect 449642 42550 449654 42602
rect 449872 42550 449884 42602
rect 449276 42478 449328 42490
rect 451668 42660 451720 42672
rect 450838 42550 450850 42602
rect 451068 42550 451080 42602
rect 450472 42478 450524 42490
rect 452864 42660 452916 42672
rect 452034 42550 452046 42602
rect 452264 42550 452276 42602
rect 451668 42478 451720 42490
rect 452864 42478 452916 42490
rect 453416 42660 453468 42672
rect 454056 42550 454068 42602
rect 454286 42550 454298 42602
rect 453416 42478 453468 42490
rect 145840 42375 151748 42385
rect 145840 42315 147395 42375
rect 147752 42315 151748 42375
rect 145840 42289 151748 42315
rect 441228 42368 447154 42385
rect 441228 42308 441626 42368
rect 441983 42308 447154 42368
rect 483212 42356 483240 44208
rect 483380 42412 483408 44320
rect 483548 42468 483576 44432
rect 483716 42524 483744 44544
rect 483772 42580 483800 44600
rect 483939 42636 483967 44712
rect 483996 42692 484024 44768
rect 484164 42748 484192 44880
rect 484220 42804 484248 44936
rect 484388 42860 484416 45048
rect 484444 42916 484472 45104
rect 485956 43644 485984 46224
rect 486012 43700 486040 46280
rect 486180 43756 486208 46392
rect 486236 43812 486264 46448
rect 486404 43868 486432 46560
rect 486460 43924 486488 46616
rect 486628 43980 486656 46728
rect 486684 44036 486712 46784
rect 486852 44092 486880 46896
rect 486908 44148 486936 46952
rect 487076 44204 487104 47064
rect 487132 44260 487160 47120
rect 487300 44316 487328 47232
rect 487356 44372 487384 47288
rect 487524 44428 487552 47400
rect 487580 44484 487608 47456
rect 487748 44540 487776 47568
rect 487804 44596 487832 47624
rect 670936 45852 670964 223350
rect 671048 222856 671076 223546
rect 502852 45824 670964 45852
rect 670992 222828 671076 222856
rect 502852 44596 502880 45824
rect 670992 45796 671020 222828
rect 487804 44568 502880 44596
rect 502908 45768 671020 45796
rect 502908 44540 502936 45768
rect 671160 45684 671188 223740
rect 671272 223241 671300 223938
rect 487748 44512 502936 44540
rect 503076 45656 671188 45684
rect 671216 223213 671300 223241
rect 503076 44484 503104 45656
rect 671216 45628 671244 223213
rect 487580 44456 503104 44484
rect 503132 45600 671244 45628
rect 503132 44428 503160 45600
rect 671384 45516 671412 224138
rect 671496 223642 671524 224348
rect 487524 44400 503160 44428
rect 503300 45488 671412 45516
rect 671440 223614 671524 223642
rect 503300 44372 503328 45488
rect 671440 45460 671468 223614
rect 487356 44344 503328 44372
rect 503356 45432 671468 45460
rect 503356 44316 503384 45432
rect 671608 45348 671636 224542
rect 671720 224066 671748 224744
rect 487300 44288 503384 44316
rect 503524 45320 671636 45348
rect 671664 224038 671748 224066
rect 503524 44260 503552 45320
rect 671664 45292 671692 224038
rect 487132 44232 503552 44260
rect 503580 45264 671692 45292
rect 503580 44204 503608 45264
rect 671832 45180 671860 224936
rect 671944 224443 671972 225140
rect 487076 44176 503608 44204
rect 503748 45152 671860 45180
rect 671888 224415 671972 224443
rect 503748 44148 503776 45152
rect 671888 45124 671916 224415
rect 486908 44120 503776 44148
rect 503804 45096 671916 45124
rect 503804 44092 503832 45096
rect 672056 45012 672084 225340
rect 672168 224833 672196 225536
rect 486852 44064 503832 44092
rect 503972 44984 672084 45012
rect 672112 224805 672196 224833
rect 503972 44036 504000 44984
rect 672112 44956 672140 224805
rect 486684 44008 504000 44036
rect 504028 44928 672140 44956
rect 504028 43980 504056 44928
rect 672280 44844 672308 225738
rect 672392 225255 672420 225942
rect 486628 43952 504056 43980
rect 504196 44816 672308 44844
rect 672336 225227 672420 225255
rect 504196 43924 504224 44816
rect 672336 44788 672364 225227
rect 486460 43896 504224 43924
rect 504252 44760 672364 44788
rect 504252 43868 504280 44760
rect 672504 44676 672532 226138
rect 672616 225654 672644 226336
rect 486404 43840 504280 43868
rect 504420 44648 672532 44676
rect 672560 225626 672644 225654
rect 504420 43812 504448 44648
rect 672560 44620 672588 225626
rect 486236 43784 504448 43812
rect 504476 44592 672588 44620
rect 504476 43756 504504 44592
rect 672728 44508 672756 226538
rect 672840 226029 672868 226736
rect 486180 43728 504504 43756
rect 504644 44480 672756 44508
rect 672784 226001 672868 226029
rect 504644 43700 504672 44480
rect 672784 44452 672812 226001
rect 486012 43672 504672 43700
rect 504700 44424 672812 44452
rect 504700 43644 504728 44424
rect 485956 43616 504728 43644
rect 674296 43332 674324 228580
rect 506212 43304 674324 43332
rect 506212 42916 506240 43304
rect 674352 43276 674380 229488
rect 674464 229001 674492 229690
rect 674464 228973 674548 229001
rect 484444 42888 506240 42916
rect 506268 43248 674380 43276
rect 506268 42860 506296 43248
rect 674520 43164 674548 228973
rect 484388 42832 506296 42860
rect 506436 43136 674548 43164
rect 506436 42804 506464 43136
rect 674576 43108 674604 229888
rect 674688 229397 674716 230088
rect 674688 229369 674772 229397
rect 484220 42776 506464 42804
rect 506492 43080 674604 43108
rect 506492 42748 506520 43080
rect 674744 42996 674772 229369
rect 484164 42720 506520 42748
rect 506660 42968 674772 42996
rect 506660 42692 506688 42968
rect 674800 42940 674828 230290
rect 674912 229796 674940 230490
rect 674912 229768 674996 229796
rect 483996 42664 506688 42692
rect 506716 42912 674828 42940
rect 506716 42636 506744 42912
rect 674968 42828 674996 229768
rect 483939 42608 506744 42636
rect 506884 42800 674996 42828
rect 506884 42580 506912 42800
rect 675024 42772 675052 230690
rect 483772 42552 506912 42580
rect 506940 42744 675052 42772
rect 506940 42524 506968 42744
rect 675192 42660 675220 230888
rect 483716 42496 506968 42524
rect 507108 42632 675220 42660
rect 507108 42468 507136 42632
rect 675360 42548 675388 231090
rect 483548 42440 507136 42468
rect 507276 42520 675388 42548
rect 507276 42412 507304 42520
rect 675528 42449 675556 231290
rect 483380 42384 507304 42412
rect 507444 42421 675556 42449
rect 507444 42356 507472 42421
rect 483212 42328 507472 42356
rect 441228 42289 447154 42308
<< via1 >>
rect 676093 724496 676153 724853
rect 675546 723300 675606 723657
rect 677175 724496 677235 724853
rect 676634 723300 676694 723657
rect 674156 721559 674208 721611
rect 676328 721460 676338 721678
rect 676338 721460 676372 721678
rect 676372 721460 676380 721678
rect 674100 721365 674152 721417
rect 676882 721396 677052 721404
rect 676882 721362 677052 721396
rect 676882 721352 677052 721362
rect 674160 720716 674212 720768
rect 674104 720592 674156 720644
rect 40371 604610 40431 604967
rect 41453 604610 41513 604967
rect 40912 603414 40972 603771
rect 42000 603414 42060 603771
rect 41219 602778 41227 602996
rect 41227 602778 41261 602996
rect 41261 602778 41271 602996
rect 43527 602877 43579 602929
rect 40547 602714 40717 602722
rect 40547 602680 40717 602714
rect 40547 602670 40717 602680
rect 43583 602683 43635 602735
rect 40607 601852 40615 602070
rect 40615 601852 40649 602070
rect 40649 601852 40659 602070
rect 41159 602068 41329 602076
rect 41159 602034 41329 602068
rect 41159 602024 41329 602034
rect 43523 602034 43575 602086
rect 41219 601582 41227 601800
rect 41227 601582 41261 601800
rect 41261 601582 41271 601800
rect 40547 601518 40717 601526
rect 40547 601484 40717 601518
rect 40547 601474 40717 601484
rect 40607 600656 40615 600874
rect 40615 600656 40649 600874
rect 40649 600656 40659 600874
rect 41159 600872 41329 600880
rect 41159 600838 41329 600872
rect 41159 600828 41329 600838
rect 41219 600386 41227 600604
rect 41227 600386 41261 600604
rect 41261 600386 41271 600604
rect 40547 600322 40717 600330
rect 40547 600288 40717 600322
rect 40547 600278 40717 600288
rect 40607 599460 40615 599678
rect 40615 599460 40649 599678
rect 40649 599460 40659 599678
rect 41159 599676 41329 599684
rect 41159 599642 41329 599676
rect 41159 599632 41329 599642
rect 41219 599190 41227 599408
rect 41227 599190 41261 599408
rect 41261 599190 41271 599408
rect 40547 599126 40717 599134
rect 40547 599092 40717 599126
rect 40547 599082 40717 599092
rect 40607 598264 40615 598482
rect 40615 598264 40649 598482
rect 40649 598264 40659 598482
rect 41159 598480 41329 598488
rect 41159 598446 41329 598480
rect 41159 598436 41329 598446
rect 41219 597994 41227 598212
rect 41227 597994 41261 598212
rect 41261 597994 41271 598212
rect 40547 597930 40717 597938
rect 40547 597896 40717 597930
rect 40547 597886 40717 597896
rect 40607 597068 40615 597286
rect 40615 597068 40649 597286
rect 40649 597068 40659 597286
rect 41159 597284 41329 597292
rect 41159 597250 41329 597284
rect 41159 597240 41329 597250
rect 40390 346959 40450 347316
rect 41472 346959 41532 347316
rect 40931 345763 40991 346120
rect 42019 345763 42079 346120
rect 41241 345197 41249 345415
rect 41249 345197 41283 345415
rect 41283 345197 41293 345415
rect 43499 345296 43551 345348
rect 43579 601910 43631 601962
rect 43751 601681 43803 601733
rect 43807 601487 43859 601539
rect 40569 345133 40739 345141
rect 40569 345099 40739 345133
rect 40569 345089 40739 345099
rect 43555 345102 43607 345154
rect 43747 600838 43799 600890
rect 40629 344271 40637 344489
rect 40637 344271 40671 344489
rect 40671 344271 40681 344489
rect 41181 344487 41351 344495
rect 41181 344453 41351 344487
rect 41181 344443 41351 344453
rect 43495 344453 43547 344505
rect 41241 344001 41249 344219
rect 41249 344001 41283 344219
rect 41283 344001 41293 344219
rect 40569 343937 40739 343945
rect 40569 343903 40739 343937
rect 40569 343893 40739 343903
rect 40629 343161 40637 343293
rect 40637 343161 40671 343293
rect 40671 343161 40681 343293
rect 41181 343291 41351 343299
rect 41181 343257 41351 343291
rect 41181 343247 41351 343257
rect 40629 343075 40637 343133
rect 40637 343075 40671 343133
rect 40671 343075 40681 343133
rect 41241 342805 41249 343023
rect 41249 342805 41283 343023
rect 41283 342805 41293 343023
rect 40569 342741 40739 342749
rect 40569 342707 40739 342741
rect 40569 342697 40739 342707
rect 40629 341879 40637 342097
rect 40637 341879 40671 342097
rect 40671 341879 40681 342097
rect 41181 342095 41351 342103
rect 41181 342061 41351 342095
rect 41181 342051 41351 342061
rect 41241 341609 41249 341827
rect 41249 341609 41283 341827
rect 41283 341609 41293 341827
rect 40569 341545 40739 341553
rect 40569 341511 40739 341545
rect 40569 341501 40739 341511
rect 40629 340683 40637 340901
rect 40637 340683 40671 340901
rect 40671 340683 40681 340901
rect 41181 340899 41351 340907
rect 41181 340865 41351 340899
rect 41181 340855 41351 340865
rect 41241 340413 41249 340631
rect 41249 340413 41283 340631
rect 41283 340413 41293 340631
rect 40569 340349 40739 340357
rect 40569 340315 40739 340349
rect 40569 340305 40739 340315
rect 40629 339487 40637 339705
rect 40637 339487 40671 339705
rect 40671 339487 40681 339705
rect 41181 339703 41351 339711
rect 41181 339669 41351 339703
rect 41181 339659 41351 339669
rect 41241 339217 41249 339435
rect 41249 339217 41283 339435
rect 41283 339217 41293 339435
rect 40569 339153 40739 339161
rect 40569 339119 40739 339153
rect 40569 339109 40739 339119
rect 40629 338291 40637 338509
rect 40637 338291 40671 338509
rect 40671 338291 40681 338509
rect 41181 338507 41351 338515
rect 41181 338473 41351 338507
rect 41181 338463 41351 338473
rect 41241 338021 41249 338239
rect 41249 338021 41283 338239
rect 41283 338021 41293 338239
rect 40569 337957 40739 337965
rect 40569 337923 40739 337957
rect 40569 337913 40739 337923
rect 40629 337095 40637 337313
rect 40637 337095 40671 337313
rect 40671 337095 40681 337313
rect 41181 337311 41351 337319
rect 41181 337277 41351 337311
rect 41181 337267 41351 337277
rect 41241 336825 41249 337043
rect 41249 336825 41283 337043
rect 41283 336825 41293 337043
rect 40569 336761 40739 336769
rect 40569 336727 40739 336761
rect 40569 336717 40739 336727
rect 40629 335899 40637 336117
rect 40637 335899 40671 336117
rect 40671 335899 40681 336117
rect 41181 336115 41351 336123
rect 41181 336081 41351 336115
rect 41181 336071 41351 336081
rect 41241 335629 41249 335847
rect 41249 335629 41283 335847
rect 41283 335629 41293 335847
rect 40569 335565 40739 335573
rect 40569 335531 40739 335565
rect 40569 335521 40739 335531
rect 40629 334703 40637 334921
rect 40637 334703 40671 334921
rect 40671 334703 40681 334921
rect 41181 334919 41351 334927
rect 41181 334885 41351 334919
rect 41181 334875 41351 334885
rect 43551 344329 43603 344381
rect 43723 344100 43775 344152
rect 43803 600714 43855 600766
rect 43975 600485 44027 600537
rect 44031 600291 44083 600343
rect 43779 343906 43831 343958
rect 43971 599642 44023 599694
rect 43719 343257 43771 343309
rect 43775 343133 43827 343185
rect 43947 342904 43999 342956
rect 44027 599518 44079 599570
rect 44199 599289 44251 599341
rect 44255 599095 44307 599147
rect 44003 342710 44055 342762
rect 44195 598446 44247 598498
rect 43943 342061 43995 342113
rect 43999 341937 44051 341989
rect 44171 341708 44223 341760
rect 44251 598322 44303 598374
rect 44423 598093 44475 598145
rect 44479 597899 44531 597951
rect 44227 341514 44279 341566
rect 44419 597250 44471 597302
rect 44167 340865 44219 340917
rect 44223 340741 44275 340793
rect 44395 340512 44447 340564
rect 44475 597126 44527 597178
rect 676270 720750 676440 720758
rect 676270 720716 676440 720750
rect 676270 720706 676440 720716
rect 676940 720534 676950 720752
rect 676950 720534 676984 720752
rect 676984 720534 676992 720752
rect 676085 448095 676145 448452
rect 677167 448095 677227 448452
rect 674184 447535 674236 447587
rect 676328 447436 676338 447654
rect 676338 447436 676372 447654
rect 676372 447436 676380 447654
rect 674128 447341 674180 447393
rect 676882 447372 677052 447380
rect 676882 447338 677052 447372
rect 676882 447328 677052 447338
rect 675538 446899 675598 447256
rect 676626 446899 676686 447256
rect 674188 446692 674240 446744
rect 674132 446568 674184 446620
rect 673960 446339 674012 446391
rect 673904 446145 673956 446197
rect 673964 445496 674016 445548
rect 673908 445372 673960 445424
rect 673736 445143 673788 445195
rect 673680 444949 673732 445001
rect 673740 444300 673792 444352
rect 673684 444176 673736 444228
rect 673512 443947 673564 443999
rect 673456 443753 673508 443805
rect 673516 443104 673568 443156
rect 673460 442980 673512 443032
rect 673288 442751 673340 442803
rect 673232 442557 673284 442609
rect 673292 441908 673344 441960
rect 673236 441784 673288 441836
rect 673064 441555 673116 441607
rect 673008 441361 673060 441413
rect 673068 440712 673120 440764
rect 673012 440588 673064 440640
rect 672840 440359 672892 440411
rect 672784 440165 672836 440217
rect 672844 439516 672896 439568
rect 672788 439392 672840 439444
rect 44451 340318 44503 340370
rect 44391 339669 44443 339721
rect 44447 339545 44499 339597
rect 44619 339316 44671 339368
rect 44675 339122 44727 339174
rect 44615 338473 44667 338525
rect 44671 338349 44723 338401
rect 44843 338120 44895 338172
rect 44899 337926 44951 337978
rect 44839 337277 44891 337329
rect 44895 337153 44947 337205
rect 45067 336900 45119 336952
rect 45123 336730 45175 336782
rect 45063 336081 45115 336133
rect 45119 335957 45171 336009
rect 45291 335728 45343 335780
rect 45347 335534 45399 335586
rect 45287 334885 45339 334937
rect 45343 334761 45395 334813
rect 676270 446726 676440 446734
rect 676270 446692 676440 446726
rect 676270 446682 676440 446692
rect 676940 446510 676950 446728
rect 676950 446510 676984 446728
rect 676984 446510 676992 446728
rect 676328 446240 676338 446458
rect 676338 446240 676372 446458
rect 676372 446240 676380 446458
rect 676882 446176 677052 446184
rect 676882 446142 677052 446176
rect 676882 446132 677052 446142
rect 676270 445530 676440 445538
rect 676270 445496 676440 445530
rect 676270 445486 676440 445496
rect 676940 445314 676950 445532
rect 676950 445314 676984 445532
rect 676984 445314 676992 445532
rect 676328 445044 676338 445262
rect 676338 445044 676372 445262
rect 676372 445044 676380 445262
rect 676882 444980 677052 444988
rect 676882 444946 677052 444980
rect 676882 444936 677052 444946
rect 676270 444334 676440 444342
rect 676270 444300 676440 444334
rect 676270 444290 676440 444300
rect 676940 444118 676950 444336
rect 676950 444118 676984 444336
rect 676984 444118 676992 444336
rect 676328 443848 676338 444066
rect 676338 443848 676372 444066
rect 676372 443848 676380 444066
rect 676882 443784 677052 443792
rect 676882 443750 677052 443784
rect 676882 443740 677052 443750
rect 676270 443138 676440 443146
rect 676270 443104 676440 443138
rect 676270 443094 676440 443104
rect 676940 442922 676950 443140
rect 676950 442922 676984 443140
rect 676984 442922 676992 443140
rect 676328 442652 676338 442870
rect 676338 442652 676372 442870
rect 676372 442652 676380 442870
rect 676882 442588 677052 442596
rect 676882 442554 677052 442588
rect 676882 442544 677052 442554
rect 676270 441942 676440 441950
rect 676270 441908 676440 441942
rect 676270 441898 676440 441908
rect 676940 441726 676950 441944
rect 676950 441726 676984 441944
rect 676984 441726 676992 441944
rect 676328 441456 676338 441674
rect 676338 441456 676372 441674
rect 676372 441456 676380 441674
rect 676882 441392 677052 441400
rect 676882 441358 677052 441392
rect 676882 441348 677052 441358
rect 676270 440746 676440 440754
rect 676270 440712 676440 440746
rect 676270 440702 676440 440712
rect 676940 440530 676950 440748
rect 676950 440530 676984 440748
rect 676984 440530 676992 440748
rect 676328 440260 676338 440478
rect 676338 440260 676372 440478
rect 676372 440260 676380 440478
rect 676882 440196 677052 440204
rect 676882 440162 677052 440196
rect 676882 440152 677052 440162
rect 676270 439550 676440 439558
rect 676270 439516 676440 439550
rect 676270 439506 676440 439516
rect 676940 439334 676950 439552
rect 676950 439334 676984 439552
rect 676984 439334 676992 439552
rect 134104 47568 134156 47620
rect 134947 47572 134999 47624
rect 135176 47512 135228 47564
rect 135949 47516 136001 47568
rect 135300 47400 135352 47452
rect 136143 47404 136195 47456
rect 136372 47344 136424 47396
rect 137145 47348 137197 47400
rect 136496 47232 136548 47284
rect 137339 47236 137391 47288
rect 137568 47176 137620 47228
rect 138341 47180 138393 47232
rect 137692 47064 137744 47116
rect 138535 47068 138587 47120
rect 138764 47008 138816 47060
rect 139537 47012 139589 47064
rect 138888 46896 138940 46948
rect 139731 46900 139783 46952
rect 139960 46840 140012 46892
rect 140084 46728 140136 46780
rect 429504 47596 429556 47648
rect 430347 47600 430399 47652
rect 430576 47540 430628 47592
rect 431349 47544 431401 47596
rect 430700 47428 430752 47480
rect 431543 47432 431595 47484
rect 431772 47372 431824 47424
rect 432545 47376 432597 47428
rect 431896 47260 431948 47312
rect 432739 47264 432791 47316
rect 432968 47204 433020 47256
rect 433741 47208 433793 47260
rect 433092 47092 433144 47144
rect 433935 47096 433987 47148
rect 434164 47036 434216 47088
rect 434937 47040 434989 47092
rect 434288 46924 434340 46976
rect 435131 46928 435183 46980
rect 435360 46868 435412 46920
rect 436133 46872 436185 46924
rect 140733 46508 140785 46560
rect 435484 46756 435536 46808
rect 436303 46760 436355 46812
rect 140903 46452 140955 46504
rect 436556 46700 436608 46752
rect 437329 46704 437381 46756
rect 141156 46392 141208 46444
rect 141929 46396 141981 46448
rect 436680 46588 436732 46640
rect 437523 46592 437575 46644
rect 141280 46336 141332 46388
rect 142123 46340 142175 46392
rect 437752 46532 437804 46584
rect 438525 46536 438577 46588
rect 142352 46280 142404 46332
rect 143125 46284 143177 46336
rect 437876 46420 437928 46472
rect 438695 46424 438747 46476
rect 142476 46224 142528 46276
rect 143295 46228 143347 46280
rect 438948 46364 439000 46416
rect 439721 46368 439773 46420
rect 143548 46168 143600 46220
rect 144321 46172 144373 46224
rect 439072 46252 439124 46304
rect 439915 46256 439967 46308
rect 143672 46112 143724 46164
rect 144515 46116 144567 46168
rect 440144 46196 440196 46248
rect 440917 46200 440969 46252
rect 144744 46056 144796 46108
rect 145517 46060 145569 46112
rect 152044 45048 152096 45100
rect 152887 45052 152939 45104
rect 447444 45076 447496 45128
rect 448287 45080 448339 45132
rect 153116 44992 153168 45044
rect 153889 44996 153941 45048
rect 448516 45020 448568 45072
rect 449289 45024 449341 45076
rect 153240 44880 153292 44932
rect 154083 44884 154135 44936
rect 448640 44908 448692 44960
rect 449483 44912 449535 44964
rect 154312 44824 154364 44876
rect 155085 44828 155137 44880
rect 449712 44852 449764 44904
rect 450485 44856 450537 44908
rect 154436 44712 154488 44764
rect 155255 44716 155307 44768
rect 449836 44740 449888 44792
rect 450655 44744 450707 44796
rect 155508 44656 155560 44708
rect 156281 44660 156333 44712
rect 450908 44684 450960 44736
rect 451681 44688 451733 44740
rect 155632 44544 155684 44596
rect 156475 44548 156527 44600
rect 451032 44572 451084 44624
rect 451875 44576 451927 44628
rect 156704 44488 156756 44540
rect 157477 44492 157529 44544
rect 452104 44516 452156 44568
rect 452877 44520 452929 44572
rect 156828 44376 156880 44428
rect 157647 44380 157699 44432
rect 452228 44404 452280 44456
rect 453047 44408 453099 44460
rect 157900 44264 157952 44316
rect 158673 44268 158725 44320
rect 453300 44292 453352 44344
rect 454073 44296 454125 44348
rect 158024 44152 158076 44204
rect 158867 44156 158919 44208
rect 453424 44180 453476 44232
rect 454267 44184 454319 44236
rect 146199 43944 146556 44004
rect 440430 43937 440787 43997
rect 147395 43397 147752 43457
rect 441626 43390 441983 43450
rect 134094 43102 134104 43272
rect 134104 43102 134138 43272
rect 134138 43102 134146 43272
rect 134848 43204 135066 43214
rect 134848 43170 135066 43204
rect 134848 43162 135066 43170
rect 135290 43102 135300 43272
rect 135300 43102 135334 43272
rect 135334 43102 135342 43272
rect 136044 43204 136262 43214
rect 136044 43170 136262 43204
rect 136044 43162 136262 43170
rect 136486 43102 136496 43272
rect 136496 43102 136530 43272
rect 136530 43102 136538 43272
rect 137240 43204 137458 43214
rect 137240 43170 137458 43204
rect 137240 43162 137458 43170
rect 137682 43102 137692 43272
rect 137692 43102 137726 43272
rect 137726 43102 137734 43272
rect 138436 43204 138654 43214
rect 138436 43170 138654 43204
rect 138436 43162 138654 43170
rect 138878 43102 138888 43272
rect 138888 43102 138922 43272
rect 138922 43102 138930 43272
rect 139632 43204 139850 43214
rect 139632 43170 139850 43204
rect 139632 43162 139850 43170
rect 140074 43102 140084 43272
rect 140084 43102 140118 43272
rect 140118 43102 140126 43272
rect 140828 43204 141046 43214
rect 140828 43170 141046 43204
rect 140828 43162 141046 43170
rect 141270 43102 141280 43272
rect 141280 43102 141314 43272
rect 141314 43102 141322 43272
rect 142024 43204 142242 43214
rect 142024 43170 142242 43204
rect 142024 43162 142242 43170
rect 142466 43102 142476 43272
rect 142476 43102 142510 43272
rect 142510 43102 142518 43272
rect 143220 43204 143438 43214
rect 143220 43170 143438 43204
rect 143220 43162 143438 43170
rect 143662 43102 143672 43272
rect 143672 43102 143706 43272
rect 143706 43102 143714 43272
rect 144416 43204 144634 43214
rect 144416 43170 144634 43204
rect 144416 43162 144634 43170
rect 152034 43102 152044 43272
rect 152044 43102 152078 43272
rect 152078 43102 152086 43272
rect 152788 43204 153006 43214
rect 152788 43170 153006 43204
rect 152788 43162 153006 43170
rect 153230 43102 153240 43272
rect 153240 43102 153274 43272
rect 153274 43102 153282 43272
rect 153984 43204 154202 43214
rect 153984 43170 154202 43204
rect 153984 43162 154202 43170
rect 154426 43102 154436 43272
rect 154436 43102 154470 43272
rect 154470 43102 154478 43272
rect 155180 43204 155398 43214
rect 155180 43170 155398 43204
rect 155180 43162 155398 43170
rect 155622 43102 155632 43272
rect 155632 43102 155666 43272
rect 155666 43102 155674 43272
rect 156376 43204 156594 43214
rect 156376 43170 156594 43204
rect 156376 43162 156594 43170
rect 156818 43102 156828 43272
rect 156828 43102 156862 43272
rect 156862 43102 156870 43272
rect 157572 43204 157790 43214
rect 157572 43170 157790 43204
rect 157572 43162 157790 43170
rect 158014 43102 158024 43272
rect 158024 43102 158058 43272
rect 158058 43102 158066 43272
rect 158768 43204 158986 43214
rect 158768 43170 158986 43204
rect 158768 43162 158986 43170
rect 429494 43102 429504 43272
rect 429504 43102 429538 43272
rect 429538 43102 429546 43272
rect 430248 43204 430466 43214
rect 430248 43170 430466 43204
rect 430248 43162 430466 43170
rect 430690 43102 430700 43272
rect 430700 43102 430734 43272
rect 430734 43102 430742 43272
rect 431444 43204 431662 43214
rect 431444 43170 431662 43204
rect 431444 43162 431662 43170
rect 431886 43102 431896 43272
rect 431896 43102 431930 43272
rect 431930 43102 431938 43272
rect 432640 43204 432858 43214
rect 432640 43170 432858 43204
rect 432640 43162 432858 43170
rect 433082 43102 433092 43272
rect 433092 43102 433126 43272
rect 433126 43102 433134 43272
rect 433836 43204 434054 43214
rect 433836 43170 434054 43204
rect 433836 43162 434054 43170
rect 434278 43102 434288 43272
rect 434288 43102 434322 43272
rect 434322 43102 434330 43272
rect 435032 43204 435250 43214
rect 435032 43170 435250 43204
rect 435032 43162 435250 43170
rect 435474 43102 435484 43272
rect 435484 43102 435518 43272
rect 435518 43102 435526 43272
rect 436228 43204 436446 43214
rect 436228 43170 436446 43204
rect 436228 43162 436446 43170
rect 436670 43102 436680 43272
rect 436680 43102 436714 43272
rect 436714 43102 436722 43272
rect 437424 43204 437642 43214
rect 437424 43170 437642 43204
rect 437424 43162 437642 43170
rect 437866 43102 437876 43272
rect 437876 43102 437910 43272
rect 437910 43102 437918 43272
rect 438620 43204 438838 43214
rect 438620 43170 438838 43204
rect 438620 43162 438838 43170
rect 439062 43102 439072 43272
rect 439072 43102 439106 43272
rect 439106 43102 439114 43272
rect 439816 43204 440034 43214
rect 439816 43170 440034 43204
rect 439816 43162 440034 43170
rect 447434 43102 447444 43272
rect 447444 43102 447478 43272
rect 447478 43102 447486 43272
rect 448188 43204 448406 43214
rect 448188 43170 448406 43204
rect 448188 43162 448406 43170
rect 448630 43102 448640 43272
rect 448640 43102 448674 43272
rect 448674 43102 448682 43272
rect 449384 43204 449602 43214
rect 449384 43170 449602 43204
rect 449384 43162 449602 43170
rect 449826 43102 449836 43272
rect 449836 43102 449870 43272
rect 449870 43102 449878 43272
rect 450580 43204 450798 43214
rect 450580 43170 450798 43204
rect 450580 43162 450798 43170
rect 451022 43102 451032 43272
rect 451032 43102 451066 43272
rect 451066 43102 451074 43272
rect 451776 43204 451994 43214
rect 451776 43170 451994 43204
rect 451776 43162 451994 43170
rect 452218 43102 452228 43272
rect 452228 43102 452262 43272
rect 452262 43102 452270 43272
rect 452972 43204 453190 43214
rect 452972 43170 453190 43204
rect 452972 43162 453190 43170
rect 453414 43102 453424 43272
rect 453424 43102 453458 43272
rect 453458 43102 453466 43272
rect 454168 43204 454386 43214
rect 454168 43170 454386 43204
rect 454168 43162 454386 43170
rect 146199 42856 146556 42916
rect 440430 42849 440787 42909
rect 135118 42592 135336 42602
rect 135118 42558 135336 42592
rect 135118 42550 135336 42558
rect 135936 42490 135946 42660
rect 135946 42490 135980 42660
rect 135980 42490 135988 42660
rect 136314 42592 136532 42602
rect 136314 42558 136532 42592
rect 136314 42550 136532 42558
rect 137132 42490 137142 42660
rect 137142 42490 137176 42660
rect 137176 42490 137184 42660
rect 137510 42592 137728 42602
rect 137510 42558 137728 42592
rect 137510 42550 137728 42558
rect 138328 42490 138338 42660
rect 138338 42490 138372 42660
rect 138372 42490 138380 42660
rect 138706 42592 138924 42602
rect 138706 42558 138924 42592
rect 138706 42550 138924 42558
rect 139524 42490 139534 42660
rect 139534 42490 139568 42660
rect 139568 42490 139576 42660
rect 139902 42592 140120 42602
rect 139902 42558 140120 42592
rect 139902 42550 140120 42558
rect 140720 42490 140730 42660
rect 140730 42490 140764 42660
rect 140764 42490 140772 42660
rect 141098 42592 141316 42602
rect 141098 42558 141316 42592
rect 141098 42550 141316 42558
rect 141916 42490 141926 42660
rect 141926 42490 141960 42660
rect 141960 42490 141968 42660
rect 142294 42592 142512 42602
rect 142294 42558 142512 42592
rect 142294 42550 142512 42558
rect 143112 42490 143122 42660
rect 143122 42490 143156 42660
rect 143156 42490 143164 42660
rect 143490 42592 143708 42602
rect 143490 42558 143708 42592
rect 143490 42550 143708 42558
rect 144308 42490 144318 42660
rect 144318 42490 144352 42660
rect 144352 42490 144360 42660
rect 144686 42592 144904 42602
rect 144686 42558 144904 42592
rect 144686 42550 144904 42558
rect 145504 42490 145514 42660
rect 145514 42490 145548 42660
rect 145548 42490 145556 42660
rect 153058 42592 153276 42602
rect 153058 42558 153276 42592
rect 153058 42550 153276 42558
rect 153876 42490 153886 42660
rect 153886 42490 153920 42660
rect 153920 42490 153928 42660
rect 154254 42592 154472 42602
rect 154254 42558 154472 42592
rect 154254 42550 154472 42558
rect 155072 42490 155082 42660
rect 155082 42490 155116 42660
rect 155116 42490 155124 42660
rect 155450 42592 155668 42602
rect 155450 42558 155668 42592
rect 155450 42550 155668 42558
rect 156268 42490 156278 42660
rect 156278 42490 156312 42660
rect 156312 42490 156320 42660
rect 156646 42592 156864 42602
rect 156646 42558 156864 42592
rect 156646 42550 156864 42558
rect 157464 42490 157474 42660
rect 157474 42490 157508 42660
rect 157508 42490 157516 42660
rect 158016 42490 158024 42660
rect 158024 42490 158058 42660
rect 158058 42490 158068 42660
rect 158668 42592 158886 42602
rect 158668 42558 158886 42592
rect 158668 42550 158886 42558
rect 430518 42592 430736 42602
rect 430518 42558 430736 42592
rect 430518 42550 430736 42558
rect 431336 42490 431346 42660
rect 431346 42490 431380 42660
rect 431380 42490 431388 42660
rect 431714 42592 431932 42602
rect 431714 42558 431932 42592
rect 431714 42550 431932 42558
rect 432532 42490 432542 42660
rect 432542 42490 432576 42660
rect 432576 42490 432584 42660
rect 432910 42592 433128 42602
rect 432910 42558 433128 42592
rect 432910 42550 433128 42558
rect 433728 42490 433738 42660
rect 433738 42490 433772 42660
rect 433772 42490 433780 42660
rect 434106 42592 434324 42602
rect 434106 42558 434324 42592
rect 434106 42550 434324 42558
rect 434924 42490 434934 42660
rect 434934 42490 434968 42660
rect 434968 42490 434976 42660
rect 435302 42592 435520 42602
rect 435302 42558 435520 42592
rect 435302 42550 435520 42558
rect 436120 42490 436130 42660
rect 436130 42490 436164 42660
rect 436164 42490 436172 42660
rect 436498 42592 436716 42602
rect 436498 42558 436716 42592
rect 436498 42550 436716 42558
rect 437316 42490 437326 42660
rect 437326 42490 437360 42660
rect 437360 42490 437368 42660
rect 437694 42592 437912 42602
rect 437694 42558 437912 42592
rect 437694 42550 437912 42558
rect 438512 42490 438522 42660
rect 438522 42490 438556 42660
rect 438556 42490 438564 42660
rect 438890 42592 439108 42602
rect 438890 42558 439108 42592
rect 438890 42550 439108 42558
rect 439708 42490 439718 42660
rect 439718 42490 439752 42660
rect 439752 42490 439760 42660
rect 440086 42592 440304 42602
rect 440086 42558 440304 42592
rect 440086 42550 440304 42558
rect 440904 42490 440914 42660
rect 440914 42490 440948 42660
rect 440948 42490 440956 42660
rect 448458 42592 448676 42602
rect 448458 42558 448676 42592
rect 448458 42550 448676 42558
rect 449276 42490 449286 42660
rect 449286 42490 449320 42660
rect 449320 42490 449328 42660
rect 449654 42592 449872 42602
rect 449654 42558 449872 42592
rect 449654 42550 449872 42558
rect 450472 42490 450482 42660
rect 450482 42490 450516 42660
rect 450516 42490 450524 42660
rect 450850 42592 451068 42602
rect 450850 42558 451068 42592
rect 450850 42550 451068 42558
rect 451668 42490 451678 42660
rect 451678 42490 451712 42660
rect 451712 42490 451720 42660
rect 452046 42592 452264 42602
rect 452046 42558 452264 42592
rect 452046 42550 452264 42558
rect 452864 42490 452874 42660
rect 452874 42490 452908 42660
rect 452908 42490 452916 42660
rect 453416 42490 453424 42660
rect 453424 42490 453458 42660
rect 453458 42490 453468 42660
rect 454068 42592 454286 42602
rect 454068 42558 454286 42592
rect 454068 42550 454286 42558
rect 147395 42315 147752 42375
rect 441626 42308 441983 42368
<< metal2 >>
rect 676081 724853 676167 724861
rect 676081 724496 676093 724853
rect 676153 724496 676167 724853
rect 676081 724488 676167 724496
rect 677166 724853 677252 724861
rect 677166 724496 677175 724853
rect 677235 724496 677252 724853
rect 677166 724488 677252 724496
rect 675532 723657 675618 723665
rect 675532 723300 675546 723657
rect 675606 723300 675618 723657
rect 675532 723292 675618 723300
rect 676620 723657 676706 723665
rect 676620 723300 676634 723657
rect 676694 723300 676706 723657
rect 676620 723292 676706 723300
rect 674150 721587 674156 721611
rect 674066 721559 674156 721587
rect 674208 721587 674214 721611
rect 676322 721587 676328 721678
rect 674208 721559 676328 721587
rect 676322 721460 676328 721559
rect 676380 721460 676386 721678
rect 674094 721393 674100 721417
rect 674066 721365 674100 721393
rect 674152 721393 674158 721417
rect 676882 721404 677052 721410
rect 674152 721365 676882 721393
rect 676882 721346 677052 721352
rect 674154 720744 674160 720768
rect 674066 720716 674160 720744
rect 674212 720744 674218 720768
rect 676270 720758 676440 720764
rect 674212 720716 676270 720744
rect 676270 720700 676440 720706
rect 674098 720620 674104 720644
rect 674066 720592 674104 720620
rect 674156 720620 674162 720644
rect 676934 720620 676940 720752
rect 674156 720592 676940 720620
rect 676934 720534 676940 720592
rect 676992 720534 676998 720752
rect 40354 604967 40440 604975
rect 40354 604610 40371 604967
rect 40431 604610 40440 604967
rect 40354 604602 40440 604610
rect 41439 604967 41525 604975
rect 41439 604610 41453 604967
rect 41513 604610 41525 604967
rect 41439 604602 41525 604610
rect 40900 603771 40986 603779
rect 40900 603414 40912 603771
rect 40972 603414 40986 603771
rect 40900 603406 40986 603414
rect 41988 603771 42074 603779
rect 41988 603414 42000 603771
rect 42060 603414 42074 603771
rect 41988 603406 42074 603414
rect 41213 602778 41219 602996
rect 41271 602905 41277 602996
rect 43521 602905 43527 602929
rect 41271 602877 43527 602905
rect 43579 602905 43585 602929
rect 43579 602877 44320 602905
rect 41271 602778 41277 602877
rect 40547 602722 40717 602728
rect 43577 602711 43583 602735
rect 40717 602683 43583 602711
rect 43635 602711 43641 602735
rect 43635 602683 44320 602711
rect 40547 602664 40717 602670
rect 41159 602076 41329 602082
rect 40601 601852 40607 602070
rect 40659 601938 40665 602070
rect 43517 602062 43523 602086
rect 41329 602034 43523 602062
rect 43575 602062 43581 602086
rect 43575 602034 44320 602062
rect 41159 602018 41329 602024
rect 43573 601938 43579 601962
rect 40659 601910 43579 601938
rect 43631 601938 43637 601962
rect 43631 601910 44320 601938
rect 40659 601852 40665 601910
rect 41213 601582 41219 601800
rect 41271 601709 41277 601800
rect 43745 601709 43751 601733
rect 41271 601681 43751 601709
rect 43803 601709 43809 601733
rect 43803 601681 44320 601709
rect 41271 601582 41277 601681
rect 40547 601526 40717 601532
rect 43801 601515 43807 601539
rect 40717 601487 43807 601515
rect 43859 601515 43865 601539
rect 43859 601487 44320 601515
rect 40547 601468 40717 601474
rect 41159 600880 41329 600886
rect 40601 600656 40607 600874
rect 40659 600742 40665 600874
rect 43741 600866 43747 600890
rect 41329 600838 43747 600866
rect 43799 600866 43805 600890
rect 43799 600838 44320 600866
rect 41159 600822 41329 600828
rect 43797 600742 43803 600766
rect 40659 600714 43803 600742
rect 43855 600742 43861 600766
rect 43855 600714 44320 600742
rect 40659 600656 40665 600714
rect 41213 600386 41219 600604
rect 41271 600513 41277 600604
rect 43969 600513 43975 600537
rect 41271 600485 43975 600513
rect 44027 600513 44033 600537
rect 44027 600485 44320 600513
rect 41271 600386 41277 600485
rect 40547 600330 40717 600336
rect 44025 600319 44031 600343
rect 40717 600291 44031 600319
rect 44083 600319 44089 600343
rect 44083 600291 44320 600319
rect 40547 600272 40717 600278
rect 41159 599684 41329 599690
rect 40601 599460 40607 599678
rect 40659 599546 40665 599678
rect 43965 599670 43971 599694
rect 41329 599642 43971 599670
rect 44023 599670 44029 599694
rect 44023 599642 44320 599670
rect 41159 599626 41329 599632
rect 44021 599546 44027 599570
rect 40659 599518 44027 599546
rect 44079 599546 44085 599570
rect 44079 599518 44320 599546
rect 40659 599460 40665 599518
rect 41213 599190 41219 599408
rect 41271 599317 41277 599408
rect 44193 599317 44199 599341
rect 41271 599289 44199 599317
rect 44251 599317 44257 599341
rect 44251 599289 44321 599317
rect 41271 599190 41277 599289
rect 40547 599134 40717 599140
rect 44249 599123 44255 599147
rect 40717 599095 44255 599123
rect 44307 599123 44313 599147
rect 44307 599095 44321 599123
rect 40547 599076 40717 599082
rect 41159 598488 41329 598494
rect 40601 598264 40607 598482
rect 40659 598350 40665 598482
rect 44189 598474 44195 598498
rect 41329 598446 44195 598474
rect 44247 598474 44253 598498
rect 44247 598446 44335 598474
rect 41159 598430 41329 598436
rect 44245 598350 44251 598374
rect 40659 598322 44251 598350
rect 44303 598350 44309 598374
rect 44303 598322 44335 598350
rect 40659 598264 40665 598322
rect 41213 597994 41219 598212
rect 41271 598121 41277 598212
rect 44417 598121 44423 598145
rect 41271 598093 44423 598121
rect 44475 598121 44481 598145
rect 44475 598093 44544 598121
rect 41271 597994 41277 598093
rect 40547 597938 40717 597944
rect 44473 597927 44479 597951
rect 40717 597899 44479 597927
rect 44531 597927 44537 597951
rect 44531 597899 44544 597927
rect 40547 597880 40717 597886
rect 41159 597292 41329 597298
rect 40601 597068 40607 597286
rect 40659 597154 40665 597286
rect 44413 597278 44419 597302
rect 41329 597250 44419 597278
rect 44471 597278 44477 597302
rect 44471 597250 44544 597278
rect 41159 597234 41329 597240
rect 44469 597154 44475 597178
rect 40659 597126 44475 597154
rect 44527 597154 44533 597178
rect 44527 597126 44544 597154
rect 40659 597068 40665 597126
rect 676073 448452 676159 448460
rect 676073 448095 676085 448452
rect 676145 448095 676159 448452
rect 676073 448087 676159 448095
rect 677158 448452 677244 448460
rect 677158 448095 677167 448452
rect 677227 448095 677244 448452
rect 677158 448087 677244 448095
rect 674178 447563 674184 447587
rect 673198 447535 674184 447563
rect 674236 447563 674242 447587
rect 676322 447563 676328 447654
rect 674236 447535 676328 447563
rect 676322 447436 676328 447535
rect 676380 447436 676386 447654
rect 674122 447369 674128 447393
rect 673198 447341 674128 447369
rect 674180 447369 674186 447393
rect 676882 447380 677052 447386
rect 674180 447341 676882 447369
rect 676882 447322 677052 447328
rect 675524 447256 675610 447264
rect 675524 446899 675538 447256
rect 675598 446899 675610 447256
rect 675524 446891 675610 446899
rect 676612 447256 676698 447264
rect 676612 446899 676626 447256
rect 676686 446899 676698 447256
rect 676612 446891 676698 446899
rect 674182 446720 674188 446744
rect 673198 446692 674188 446720
rect 674240 446720 674246 446744
rect 676270 446734 676440 446740
rect 674240 446692 676270 446720
rect 676270 446676 676440 446682
rect 674126 446596 674132 446620
rect 673198 446568 674132 446596
rect 674184 446596 674190 446620
rect 676934 446596 676940 446728
rect 674184 446568 676940 446596
rect 676934 446510 676940 446568
rect 676992 446510 676998 446728
rect 673954 446367 673960 446391
rect 673198 446339 673960 446367
rect 674012 446367 674018 446391
rect 676322 446367 676328 446458
rect 674012 446339 676328 446367
rect 676322 446240 676328 446339
rect 676380 446240 676386 446458
rect 673898 446173 673904 446197
rect 673198 446145 673904 446173
rect 673956 446173 673962 446197
rect 676882 446184 677052 446190
rect 673956 446145 676882 446173
rect 676882 446126 677052 446132
rect 673958 445524 673964 445548
rect 673198 445496 673964 445524
rect 674016 445524 674022 445548
rect 676270 445538 676440 445544
rect 674016 445496 676270 445524
rect 676270 445480 676440 445486
rect 673902 445400 673908 445424
rect 673198 445372 673908 445400
rect 673960 445400 673966 445424
rect 676934 445400 676940 445532
rect 673960 445372 676940 445400
rect 676934 445314 676940 445372
rect 676992 445314 676998 445532
rect 673730 445171 673736 445195
rect 673198 445143 673736 445171
rect 673788 445171 673794 445195
rect 676322 445171 676328 445262
rect 673788 445143 676328 445171
rect 676322 445044 676328 445143
rect 676380 445044 676386 445262
rect 673674 444977 673680 445001
rect 673198 444949 673680 444977
rect 673732 444977 673738 445001
rect 676882 444988 677052 444994
rect 673732 444949 676882 444977
rect 676882 444930 677052 444936
rect 673734 444328 673740 444352
rect 673198 444300 673740 444328
rect 673792 444328 673798 444352
rect 676270 444342 676440 444348
rect 673792 444300 676270 444328
rect 676270 444284 676440 444290
rect 673678 444204 673684 444228
rect 673198 444176 673684 444204
rect 673736 444204 673742 444228
rect 676934 444204 676940 444336
rect 673736 444176 676940 444204
rect 676934 444118 676940 444176
rect 676992 444118 676998 444336
rect 673506 443975 673512 443999
rect 673198 443947 673512 443975
rect 673564 443975 673570 443999
rect 676322 443975 676328 444066
rect 673564 443947 676328 443975
rect 676322 443848 676328 443947
rect 676380 443848 676386 444066
rect 673450 443781 673456 443805
rect 673198 443753 673456 443781
rect 673508 443781 673514 443805
rect 676882 443792 677052 443798
rect 673508 443753 676882 443781
rect 676882 443734 677052 443740
rect 673510 443132 673516 443156
rect 673198 443104 673516 443132
rect 673568 443132 673574 443156
rect 676270 443146 676440 443152
rect 673568 443104 676270 443132
rect 676270 443088 676440 443094
rect 673454 443008 673460 443032
rect 673198 442980 673460 443008
rect 673512 443008 673518 443032
rect 676934 443008 676940 443140
rect 673512 442980 676940 443008
rect 676934 442922 676940 442980
rect 676992 442922 676998 443140
rect 673282 442779 673288 442803
rect 673198 442751 673288 442779
rect 673340 442779 673346 442803
rect 676322 442779 676328 442870
rect 673340 442751 676328 442779
rect 676322 442652 676328 442751
rect 676380 442652 676386 442870
rect 673226 442585 673232 442609
rect 673198 442557 673232 442585
rect 673284 442585 673290 442609
rect 676882 442596 677052 442602
rect 673284 442557 676882 442585
rect 676882 442538 677052 442544
rect 673286 441936 673292 441960
rect 673198 441908 673292 441936
rect 673344 441936 673350 441960
rect 676270 441950 676440 441956
rect 673344 441908 676270 441936
rect 676270 441892 676440 441898
rect 673230 441812 673236 441836
rect 673198 441784 673236 441812
rect 673288 441812 673294 441836
rect 676934 441812 676940 441944
rect 673288 441784 676940 441812
rect 676934 441726 676940 441784
rect 676992 441726 676998 441944
rect 673058 441583 673064 441607
rect 672973 441555 673064 441583
rect 673116 441583 673122 441607
rect 676322 441583 676328 441674
rect 673116 441555 676328 441583
rect 676322 441456 676328 441555
rect 676380 441456 676386 441674
rect 673002 441389 673008 441413
rect 672973 441361 673008 441389
rect 673060 441389 673066 441413
rect 676882 441400 677052 441406
rect 673060 441361 676882 441389
rect 676882 441342 677052 441348
rect 673062 440740 673068 440764
rect 672980 440712 673068 440740
rect 673120 440740 673126 440764
rect 676270 440754 676440 440760
rect 673120 440712 676270 440740
rect 676270 440696 676440 440702
rect 673006 440616 673012 440640
rect 672980 440588 673012 440616
rect 673064 440616 673070 440640
rect 676934 440616 676940 440748
rect 673064 440588 676940 440616
rect 676934 440530 676940 440588
rect 676992 440530 676998 440748
rect 672834 440387 672840 440411
rect 672750 440359 672840 440387
rect 672892 440387 672898 440411
rect 676322 440387 676328 440478
rect 672892 440359 676328 440387
rect 676322 440260 676328 440359
rect 676380 440260 676386 440478
rect 672778 440193 672784 440217
rect 672750 440165 672784 440193
rect 672836 440193 672842 440217
rect 676882 440204 677052 440210
rect 672836 440165 676882 440193
rect 676882 440146 677052 440152
rect 672838 439544 672844 439568
rect 672750 439516 672844 439544
rect 672896 439544 672902 439568
rect 676270 439558 676440 439564
rect 672896 439516 676270 439544
rect 676270 439500 676440 439506
rect 672782 439420 672788 439444
rect 672750 439392 672788 439420
rect 672840 439420 672846 439444
rect 676934 439420 676940 439552
rect 672840 439392 676940 439420
rect 676934 439334 676940 439392
rect 676992 439334 676998 439552
rect 40373 347316 40459 347324
rect 40373 346959 40390 347316
rect 40450 346959 40459 347316
rect 40373 346951 40459 346959
rect 41458 347316 41544 347324
rect 41458 346959 41472 347316
rect 41532 346959 41544 347316
rect 41458 346951 41544 346959
rect 40919 346120 41005 346128
rect 40919 345763 40931 346120
rect 40991 345763 41005 346120
rect 40919 345755 41005 345763
rect 42007 346120 42093 346128
rect 42007 345763 42019 346120
rect 42079 345763 42093 346120
rect 42007 345755 42093 345763
rect 41235 345197 41241 345415
rect 41293 345324 41299 345415
rect 43493 345324 43499 345348
rect 41293 345296 43499 345324
rect 43551 345324 43557 345348
rect 43551 345296 44748 345324
rect 41293 345197 41299 345296
rect 40569 345141 40739 345147
rect 43549 345130 43555 345154
rect 40739 345102 43555 345130
rect 43607 345130 43613 345154
rect 43607 345102 44748 345130
rect 40569 345083 40739 345089
rect 41181 344495 41351 344501
rect 40623 344271 40629 344489
rect 40681 344357 40687 344489
rect 43489 344481 43495 344505
rect 41351 344453 43495 344481
rect 43547 344481 43553 344505
rect 43547 344453 44748 344481
rect 41181 344437 41351 344443
rect 43545 344357 43551 344381
rect 40681 344329 43551 344357
rect 43603 344357 43609 344381
rect 43603 344329 44748 344357
rect 40681 344271 40687 344329
rect 41235 344001 41241 344219
rect 41293 344128 41299 344219
rect 43717 344128 43723 344152
rect 41293 344100 43723 344128
rect 43775 344128 43781 344152
rect 43775 344100 44748 344128
rect 41293 344001 41299 344100
rect 40569 343945 40739 343951
rect 43773 343934 43779 343958
rect 40739 343906 43779 343934
rect 43831 343934 43837 343958
rect 43831 343906 44748 343934
rect 40569 343887 40739 343893
rect 41181 343299 41351 343305
rect 40623 343161 40629 343293
rect 40681 343161 40687 343293
rect 43713 343285 43719 343309
rect 41351 343257 43719 343285
rect 43771 343285 43777 343309
rect 43771 343257 44748 343285
rect 41181 343241 41351 343247
rect 43769 343161 43775 343185
rect 40569 343133 43775 343161
rect 43827 343161 43833 343185
rect 43827 343133 44748 343161
rect 40623 343075 40629 343133
rect 40681 343075 40687 343133
rect 41235 342805 41241 343023
rect 41293 342932 41299 343023
rect 43941 342932 43947 342956
rect 41293 342904 43947 342932
rect 43999 342932 44005 342956
rect 43999 342904 44748 342932
rect 41293 342805 41299 342904
rect 40569 342749 40739 342755
rect 43997 342738 44003 342762
rect 40739 342710 44003 342738
rect 44055 342738 44061 342762
rect 44055 342710 44748 342738
rect 40569 342691 40739 342697
rect 41181 342103 41351 342109
rect 40623 341879 40629 342097
rect 40681 341965 40687 342097
rect 43937 342089 43943 342113
rect 41351 342061 43943 342089
rect 43995 342089 44001 342113
rect 43995 342061 44748 342089
rect 41181 342045 41351 342051
rect 43993 341965 43999 341989
rect 40681 341937 43999 341965
rect 44051 341965 44057 341989
rect 44051 341937 44748 341965
rect 40681 341879 40687 341937
rect 41235 341609 41241 341827
rect 41293 341736 41299 341827
rect 44165 341736 44171 341760
rect 41293 341708 44171 341736
rect 44223 341736 44229 341760
rect 44223 341708 44748 341736
rect 41293 341609 41299 341708
rect 40569 341553 40739 341559
rect 44221 341542 44227 341566
rect 40739 341514 44227 341542
rect 44279 341542 44285 341566
rect 44279 341514 44748 341542
rect 40569 341495 40739 341501
rect 41181 340907 41351 340913
rect 40623 340683 40629 340901
rect 40681 340769 40687 340901
rect 44161 340893 44167 340917
rect 41351 340865 44167 340893
rect 44219 340893 44225 340917
rect 44219 340865 44748 340893
rect 41181 340849 41351 340855
rect 44217 340769 44223 340793
rect 40681 340741 44223 340769
rect 44275 340769 44281 340793
rect 44275 340741 44748 340769
rect 40681 340683 40687 340741
rect 41235 340413 41241 340631
rect 41293 340540 41299 340631
rect 44389 340540 44395 340564
rect 41293 340512 44395 340540
rect 44447 340540 44453 340564
rect 44447 340512 44748 340540
rect 41293 340413 41299 340512
rect 40569 340357 40739 340363
rect 44445 340346 44451 340370
rect 40739 340318 44451 340346
rect 44503 340346 44509 340370
rect 44503 340318 44748 340346
rect 40569 340299 40739 340305
rect 41181 339711 41351 339717
rect 40623 339487 40629 339705
rect 40681 339573 40687 339705
rect 44385 339697 44391 339721
rect 41351 339669 44391 339697
rect 44443 339697 44449 339721
rect 44443 339669 44748 339697
rect 41181 339653 41351 339659
rect 44441 339573 44447 339597
rect 40681 339545 44447 339573
rect 44499 339573 44505 339597
rect 44499 339545 44748 339573
rect 40681 339487 40687 339545
rect 41235 339217 41241 339435
rect 41293 339344 41299 339435
rect 44613 339344 44619 339368
rect 41293 339316 44619 339344
rect 44671 339344 44677 339368
rect 44671 339316 44768 339344
rect 41293 339217 41299 339316
rect 40569 339161 40739 339167
rect 44669 339150 44675 339174
rect 40739 339122 44675 339150
rect 44727 339150 44733 339174
rect 44727 339122 44768 339150
rect 40569 339103 40739 339109
rect 41181 338515 41351 338521
rect 40623 338291 40629 338509
rect 40681 338377 40687 338509
rect 44609 338501 44615 338525
rect 41351 338473 44615 338501
rect 44667 338501 44673 338525
rect 44667 338473 44749 338501
rect 41181 338457 41351 338463
rect 44665 338377 44671 338401
rect 40681 338349 44671 338377
rect 44723 338377 44729 338401
rect 44723 338349 44749 338377
rect 40681 338291 40687 338349
rect 41235 338021 41241 338239
rect 41293 338148 41299 338239
rect 44837 338148 44843 338172
rect 41293 338120 44843 338148
rect 44895 338148 44901 338172
rect 44895 338120 44982 338148
rect 41293 338021 41299 338120
rect 40569 337965 40739 337971
rect 44893 337954 44899 337978
rect 40739 337926 44899 337954
rect 44951 337954 44957 337978
rect 44951 337926 44982 337954
rect 40569 337907 40739 337913
rect 41181 337319 41351 337325
rect 40623 337095 40629 337313
rect 40681 337181 40687 337313
rect 44833 337305 44839 337329
rect 41351 337277 44839 337305
rect 44891 337305 44897 337329
rect 44891 337277 44961 337305
rect 41181 337261 41351 337267
rect 44889 337181 44895 337205
rect 40681 337153 44895 337181
rect 44947 337181 44953 337205
rect 44947 337153 44961 337181
rect 40681 337095 40687 337153
rect 41235 336825 41241 337043
rect 41293 336952 41299 337043
rect 41293 336924 45067 336952
rect 41293 336825 41299 336924
rect 45061 336900 45067 336924
rect 45119 336924 45195 336952
rect 45119 336900 45125 336924
rect 40569 336769 40739 336775
rect 45117 336758 45123 336782
rect 40739 336730 45123 336758
rect 45175 336758 45181 336782
rect 45175 336730 45195 336758
rect 40569 336711 40739 336717
rect 41181 336123 41351 336129
rect 40623 335899 40629 336117
rect 40681 335985 40687 336117
rect 45057 336109 45063 336133
rect 41351 336081 45063 336109
rect 45115 336109 45121 336133
rect 45115 336081 45206 336109
rect 41181 336065 41351 336071
rect 45113 335985 45119 336009
rect 40681 335957 45119 335985
rect 45171 335985 45177 336009
rect 45171 335957 45206 335985
rect 40681 335899 40687 335957
rect 41235 335629 41241 335847
rect 41293 335756 41299 335847
rect 45285 335756 45291 335780
rect 41293 335728 45291 335756
rect 45343 335756 45349 335780
rect 45343 335728 45420 335756
rect 41293 335629 41299 335728
rect 40569 335573 40739 335579
rect 45341 335562 45347 335586
rect 40739 335534 45347 335562
rect 45399 335562 45405 335586
rect 45399 335534 45420 335562
rect 40569 335515 40739 335521
rect 41181 334927 41351 334933
rect 40623 334703 40629 334921
rect 40681 334789 40687 334921
rect 45281 334913 45287 334937
rect 41351 334885 45287 334913
rect 45339 334913 45345 334937
rect 45339 334885 45420 334913
rect 41181 334869 41351 334875
rect 45337 334789 45343 334813
rect 40681 334761 45343 334789
rect 45395 334789 45401 334813
rect 45395 334761 45420 334789
rect 40681 334703 40687 334761
rect 429504 47654 429532 47673
rect 430347 47658 430375 47673
rect 429504 47648 429556 47654
rect 134104 47626 134132 47645
rect 134947 47630 134975 47645
rect 134104 47620 134156 47626
rect 134104 47562 134156 47568
rect 134947 47624 134999 47630
rect 429504 47590 429556 47596
rect 430347 47652 430399 47658
rect 430347 47594 430399 47600
rect 430576 47598 430604 47610
rect 431349 47602 431377 47617
rect 134947 47566 134999 47572
rect 135176 47570 135204 47580
rect 135949 47574 135977 47585
rect 134104 43272 134132 47562
rect 134088 43102 134094 43272
rect 134146 43102 134152 43272
rect 134947 43220 134975 47566
rect 135176 47564 135228 47570
rect 135176 47506 135228 47512
rect 135949 47568 136001 47574
rect 135949 47510 136001 47516
rect 134848 43214 135066 43220
rect 134848 43156 135066 43162
rect 135176 42608 135204 47506
rect 135300 47458 135328 47480
rect 135300 47452 135352 47458
rect 135300 47394 135352 47400
rect 135300 43272 135328 47394
rect 135284 43102 135290 43272
rect 135342 43102 135348 43272
rect 135949 42660 135977 47510
rect 136143 47462 136171 47480
rect 136143 47456 136195 47462
rect 136143 47398 136195 47404
rect 136372 47402 136400 47410
rect 137145 47406 137173 47417
rect 136143 43220 136171 47398
rect 136372 47396 136424 47402
rect 136372 47338 136424 47344
rect 137145 47400 137197 47406
rect 137145 47342 137197 47348
rect 136044 43214 136262 43220
rect 136044 43156 136262 43162
rect 135118 42602 135336 42608
rect 135118 42544 135336 42550
rect 135930 42490 135936 42660
rect 135988 42490 135994 42660
rect 136372 42608 136400 47338
rect 136496 47290 136524 47309
rect 136496 47284 136548 47290
rect 136496 47226 136548 47232
rect 136496 43272 136524 47226
rect 136480 43102 136486 43272
rect 136538 43102 136544 43272
rect 137145 42660 137173 47342
rect 137339 47294 137367 47304
rect 137339 47288 137391 47294
rect 137339 47230 137391 47236
rect 137568 47234 137596 47247
rect 138341 47238 138369 47252
rect 137339 43220 137367 47230
rect 137568 47228 137620 47234
rect 137568 47170 137620 47176
rect 138341 47232 138393 47238
rect 138341 47174 138393 47180
rect 137240 43214 137458 43220
rect 137240 43156 137458 43162
rect 136314 42602 136532 42608
rect 136314 42544 136532 42550
rect 137126 42490 137132 42660
rect 137184 42490 137190 42660
rect 137568 42608 137596 47170
rect 137692 47122 137720 47163
rect 137692 47116 137744 47122
rect 137692 47058 137744 47064
rect 137692 43272 137720 47058
rect 137676 43102 137682 43272
rect 137734 43102 137740 43272
rect 138341 42660 138369 47174
rect 138535 47126 138563 47139
rect 138535 47120 138587 47126
rect 138535 47062 138587 47068
rect 138764 47066 138792 47090
rect 139537 47070 139565 47094
rect 138535 43220 138563 47062
rect 138764 47060 138816 47066
rect 138764 47002 138816 47008
rect 139537 47064 139589 47070
rect 139537 47006 139589 47012
rect 138436 43214 138654 43220
rect 138436 43156 138654 43162
rect 137510 42602 137728 42608
rect 137510 42544 137728 42550
rect 138322 42490 138328 42660
rect 138380 42490 138386 42660
rect 138764 42608 138792 47002
rect 138888 46954 138916 46974
rect 138888 46948 138940 46954
rect 138888 46890 138940 46896
rect 138888 43272 138916 46890
rect 138872 43102 138878 43272
rect 138930 43102 138936 43272
rect 139537 42660 139565 47006
rect 139731 46958 139759 46981
rect 139731 46952 139783 46958
rect 139731 46894 139783 46900
rect 139960 46898 139988 46903
rect 139731 43220 139759 46894
rect 139960 46892 140012 46898
rect 139960 46834 140012 46840
rect 139632 43214 139850 43220
rect 139632 43156 139850 43162
rect 138706 42602 138924 42608
rect 138706 42544 138924 42550
rect 139518 42490 139524 42660
rect 139576 42490 139582 42660
rect 139960 42608 139988 46834
rect 140084 46786 140112 46812
rect 140084 46780 140136 46786
rect 140084 46722 140136 46728
rect 140084 43272 140112 46722
rect 140733 46566 140761 46578
rect 140733 46560 140785 46566
rect 140927 46510 140955 46536
rect 140733 46502 140785 46508
rect 140903 46504 140955 46510
rect 140068 43102 140074 43272
rect 140126 43102 140132 43272
rect 140733 42660 140761 46502
rect 140903 46446 140955 46452
rect 140927 43220 140955 46446
rect 141156 46450 141184 46463
rect 141929 46454 141957 46462
rect 141156 46444 141208 46450
rect 141929 46448 141981 46454
rect 141156 46386 141208 46392
rect 141280 46394 141308 46430
rect 141280 46388 141332 46394
rect 140828 43214 141046 43220
rect 140828 43156 141046 43162
rect 139902 42602 140120 42608
rect 139902 42544 140120 42550
rect 140714 42490 140720 42660
rect 140772 42490 140778 42660
rect 141156 42608 141184 46386
rect 141280 46330 141332 46336
rect 141929 46390 141981 46396
rect 142123 46398 142151 46438
rect 142123 46392 142175 46398
rect 141280 43272 141308 46330
rect 141264 43102 141270 43272
rect 141322 43102 141328 43272
rect 141929 42660 141957 46390
rect 142123 46334 142175 46340
rect 142352 46338 142380 46350
rect 143125 46342 143153 46356
rect 142123 43220 142151 46334
rect 142352 46332 142404 46338
rect 143125 46336 143177 46342
rect 142352 46274 142404 46280
rect 142476 46282 142504 46301
rect 143319 46286 143347 46305
rect 142476 46276 142528 46282
rect 142024 43214 142242 43220
rect 142024 43156 142242 43162
rect 141098 42602 141316 42608
rect 141098 42544 141316 42550
rect 141910 42490 141916 42660
rect 141968 42490 141974 42660
rect 142352 42608 142380 46274
rect 142476 46218 142528 46224
rect 143125 46278 143177 46284
rect 143295 46280 143347 46286
rect 142476 43272 142504 46218
rect 142460 43102 142466 43272
rect 142518 43102 142524 43272
rect 143125 42660 143153 46278
rect 143295 46222 143347 46228
rect 143319 43220 143347 46222
rect 143548 46226 143576 46469
rect 143548 46220 143600 46226
rect 143548 46162 143600 46168
rect 143672 46170 143700 46469
rect 144321 46230 144349 46469
rect 144321 46224 144373 46230
rect 143672 46164 143724 46170
rect 143220 43214 143438 43220
rect 143220 43156 143438 43162
rect 142294 42602 142512 42608
rect 142294 42544 142512 42550
rect 143106 42490 143112 42660
rect 143164 42490 143170 42660
rect 143548 42608 143576 46162
rect 143672 46106 143724 46112
rect 144321 46166 144373 46172
rect 144515 46174 144543 46469
rect 144515 46168 144567 46174
rect 143672 43272 143700 46106
rect 143656 43102 143662 43272
rect 143714 43102 143720 43272
rect 144321 42660 144349 46166
rect 144515 46110 144567 46116
rect 144744 46114 144772 46469
rect 145517 46118 145545 46469
rect 144515 43220 144543 46110
rect 144744 46108 144796 46114
rect 144744 46050 144796 46056
rect 145517 46112 145569 46118
rect 145517 46054 145569 46060
rect 144416 43214 144634 43220
rect 144416 43156 144634 43162
rect 143490 42602 143708 42608
rect 143490 42544 143708 42550
rect 144302 42490 144308 42660
rect 144360 42490 144366 42660
rect 144744 42608 144772 46050
rect 145517 42660 145545 46054
rect 152044 45106 152072 46469
rect 152887 45110 152915 46469
rect 152044 45100 152096 45106
rect 152044 45042 152096 45048
rect 152887 45104 152939 45110
rect 152887 45046 152939 45052
rect 153116 45050 153144 46469
rect 146191 44004 146564 44018
rect 146191 43944 146199 44004
rect 146556 43944 146564 44004
rect 146191 43932 146564 43944
rect 147387 43457 147760 43469
rect 147387 43397 147395 43457
rect 147752 43397 147760 43457
rect 147387 43383 147760 43397
rect 152044 43272 152072 45042
rect 152028 43102 152034 43272
rect 152086 43102 152092 43272
rect 152887 43220 152915 45046
rect 153116 45044 153168 45050
rect 153116 44986 153168 44992
rect 152788 43214 153006 43220
rect 152788 43156 153006 43162
rect 146191 42916 146564 42930
rect 146191 42856 146199 42916
rect 146556 42856 146564 42916
rect 146191 42844 146564 42856
rect 144686 42602 144904 42608
rect 144686 42544 144904 42550
rect 145498 42490 145504 42660
rect 145556 42490 145562 42660
rect 153116 42608 153144 44986
rect 153240 44938 153268 46469
rect 153889 45054 153917 46469
rect 153889 45048 153941 45054
rect 153889 44990 153941 44996
rect 153240 44932 153292 44938
rect 153240 44874 153292 44880
rect 153240 43272 153268 44874
rect 153224 43102 153230 43272
rect 153282 43102 153288 43272
rect 153889 42660 153917 44990
rect 154083 44942 154111 46469
rect 154083 44936 154135 44942
rect 154083 44878 154135 44884
rect 154312 44882 154340 46469
rect 154083 43220 154111 44878
rect 154312 44876 154364 44882
rect 154312 44818 154364 44824
rect 153984 43214 154202 43220
rect 153984 43156 154202 43162
rect 153058 42602 153276 42608
rect 153058 42544 153276 42550
rect 153870 42490 153876 42660
rect 153928 42490 153934 42660
rect 154312 42608 154340 44818
rect 154436 44770 154464 46469
rect 155085 44886 155113 46469
rect 155085 44880 155137 44886
rect 155085 44822 155137 44828
rect 154436 44764 154488 44770
rect 154436 44706 154488 44712
rect 154436 43272 154464 44706
rect 154420 43102 154426 43272
rect 154478 43102 154484 43272
rect 155085 42660 155113 44822
rect 155279 44774 155307 46469
rect 155255 44768 155307 44774
rect 155255 44710 155307 44716
rect 155279 43220 155307 44710
rect 155508 44714 155536 46469
rect 155508 44708 155560 44714
rect 155508 44650 155560 44656
rect 155180 43214 155398 43220
rect 155180 43156 155398 43162
rect 154254 42602 154472 42608
rect 154254 42544 154472 42550
rect 155066 42490 155072 42660
rect 155124 42490 155130 42660
rect 155508 42608 155536 44650
rect 155632 44602 155660 46469
rect 156281 44718 156309 46469
rect 156281 44712 156333 44718
rect 156281 44654 156333 44660
rect 155632 44596 155684 44602
rect 155632 44538 155684 44544
rect 155632 43272 155660 44538
rect 155616 43102 155622 43272
rect 155674 43102 155680 43272
rect 156281 42660 156309 44654
rect 156475 44606 156503 46469
rect 156475 44600 156527 44606
rect 156475 44542 156527 44548
rect 156704 44546 156732 46469
rect 156475 43220 156503 44542
rect 156704 44540 156756 44546
rect 156704 44482 156756 44488
rect 156376 43214 156594 43220
rect 156376 43156 156594 43162
rect 155450 42602 155668 42608
rect 155450 42544 155668 42550
rect 156262 42490 156268 42660
rect 156320 42490 156326 42660
rect 156704 42608 156732 44482
rect 156828 44434 156856 46469
rect 157477 44550 157505 46469
rect 157477 44544 157529 44550
rect 157477 44486 157529 44492
rect 156828 44428 156880 44434
rect 156828 44370 156880 44376
rect 156828 43272 156856 44370
rect 156812 43102 156818 43272
rect 156870 43102 156876 43272
rect 157477 42660 157505 44486
rect 157671 44438 157699 46469
rect 157647 44432 157699 44438
rect 157647 44374 157699 44380
rect 157671 43220 157699 44374
rect 157900 44322 157928 46469
rect 157900 44316 157952 44322
rect 157900 44258 157952 44264
rect 157572 43214 157790 43220
rect 157572 43156 157790 43162
rect 157900 42848 157928 44258
rect 158024 44210 158052 46469
rect 158673 44326 158701 46469
rect 158673 44320 158725 44326
rect 158673 44262 158725 44268
rect 158024 44204 158076 44210
rect 158024 44146 158076 44152
rect 158024 43272 158052 44146
rect 158008 43102 158014 43272
rect 158066 43102 158072 43272
rect 158673 42848 158701 44262
rect 158867 44214 158895 46469
rect 158867 44208 158919 44214
rect 158867 44150 158919 44156
rect 158867 43220 158895 44150
rect 429504 43272 429532 47590
rect 158768 43214 158986 43220
rect 158768 43156 158986 43162
rect 429488 43102 429494 43272
rect 429546 43102 429552 43272
rect 430347 43220 430375 47594
rect 430576 47592 430628 47598
rect 430576 47534 430628 47540
rect 431349 47596 431401 47602
rect 431349 47538 431401 47544
rect 430248 43214 430466 43220
rect 430248 43156 430466 43162
rect 157900 42820 158055 42848
rect 158673 42820 158828 42848
rect 158027 42660 158055 42820
rect 156646 42602 156864 42608
rect 156646 42544 156864 42550
rect 157458 42490 157464 42660
rect 157516 42490 157522 42660
rect 158010 42490 158016 42660
rect 158068 42490 158074 42660
rect 158800 42608 158828 42820
rect 430576 42608 430604 47534
rect 430700 47486 430728 47505
rect 430700 47480 430752 47486
rect 430700 47422 430752 47428
rect 430700 43272 430728 47422
rect 430684 43102 430690 43272
rect 430742 43102 430748 43272
rect 431349 42660 431377 47538
rect 431543 47490 431571 47515
rect 431543 47484 431595 47490
rect 431543 47426 431595 47432
rect 431772 47430 431800 47447
rect 432545 47434 432573 47445
rect 431543 43220 431571 47426
rect 431772 47424 431824 47430
rect 431772 47366 431824 47372
rect 432545 47428 432597 47434
rect 432545 47370 432597 47376
rect 431444 43214 431662 43220
rect 431444 43156 431662 43162
rect 158668 42602 158886 42608
rect 158668 42544 158886 42550
rect 430518 42602 430736 42608
rect 430518 42544 430736 42550
rect 431330 42490 431336 42660
rect 431388 42490 431394 42660
rect 431772 42608 431800 47366
rect 431896 47318 431924 47341
rect 431896 47312 431948 47318
rect 431896 47254 431948 47260
rect 431896 43272 431924 47254
rect 431880 43102 431886 43272
rect 431938 43102 431944 43272
rect 432545 42660 432573 47370
rect 432739 47322 432767 47344
rect 432739 47316 432791 47322
rect 432739 47258 432791 47264
rect 432968 47262 432996 47279
rect 433741 47266 433769 47280
rect 432739 43220 432767 47258
rect 432968 47256 433020 47262
rect 432968 47198 433020 47204
rect 433741 47260 433793 47266
rect 433741 47202 433793 47208
rect 432640 43214 432858 43220
rect 432640 43156 432858 43162
rect 431714 42602 431932 42608
rect 431714 42544 431932 42550
rect 432526 42490 432532 42660
rect 432584 42490 432590 42660
rect 432968 42608 432996 47198
rect 433092 47150 433120 47163
rect 433092 47144 433144 47150
rect 433092 47086 433144 47092
rect 433092 43272 433120 47086
rect 433076 43102 433082 43272
rect 433134 43102 433140 43272
rect 433741 42660 433769 47202
rect 433935 47154 433963 47186
rect 433935 47148 433987 47154
rect 433935 47090 433987 47096
rect 434164 47094 434192 47108
rect 434937 47098 434965 47106
rect 433935 43220 433963 47090
rect 434164 47088 434216 47094
rect 434164 47030 434216 47036
rect 434937 47092 434989 47098
rect 434937 47034 434989 47040
rect 433836 43214 434054 43220
rect 433836 43156 434054 43162
rect 432910 42602 433128 42608
rect 432910 42544 433128 42550
rect 433722 42490 433728 42660
rect 433780 42490 433786 42660
rect 434164 42608 434192 47030
rect 434288 46982 434316 46998
rect 434288 46976 434340 46982
rect 434288 46918 434340 46924
rect 434288 43272 434316 46918
rect 434272 43102 434278 43272
rect 434330 43102 434336 43272
rect 434937 42660 434965 47034
rect 435131 46986 435159 47002
rect 435131 46980 435183 46986
rect 435131 46922 435183 46928
rect 435360 46926 435388 46935
rect 436133 46930 436161 46941
rect 435131 43220 435159 46922
rect 435360 46920 435412 46926
rect 435360 46862 435412 46868
rect 436133 46924 436185 46930
rect 436133 46866 436185 46872
rect 435032 43214 435250 43220
rect 435032 43156 435250 43162
rect 434106 42602 434324 42608
rect 434106 42544 434324 42550
rect 434918 42490 434924 42660
rect 434976 42490 434982 42660
rect 435360 42608 435388 46862
rect 435484 46814 435512 46836
rect 435484 46808 435536 46814
rect 435484 46750 435536 46756
rect 435484 43272 435512 46750
rect 435468 43102 435474 43272
rect 435526 43102 435532 43272
rect 436133 42660 436161 46866
rect 436327 46818 436355 46840
rect 436303 46812 436355 46818
rect 436303 46754 436355 46760
rect 436327 43220 436355 46754
rect 436556 46758 436584 46769
rect 437329 46762 437357 46774
rect 436556 46752 436608 46758
rect 436556 46694 436608 46700
rect 437329 46756 437381 46762
rect 437329 46698 437381 46704
rect 436228 43214 436446 43220
rect 436228 43156 436446 43162
rect 435302 42602 435520 42608
rect 435302 42544 435520 42550
rect 436114 42490 436120 42660
rect 436172 42490 436178 42660
rect 436556 42608 436584 46694
rect 436680 46646 436708 46662
rect 436680 46640 436732 46646
rect 436680 46582 436732 46588
rect 436680 43272 436708 46582
rect 436664 43102 436670 43272
rect 436722 43102 436728 43272
rect 437329 42660 437357 46698
rect 437523 46650 437551 46673
rect 437523 46644 437575 46650
rect 437523 46586 437575 46592
rect 437752 46590 437780 46600
rect 438525 46594 438553 46602
rect 437523 43220 437551 46586
rect 437752 46584 437804 46590
rect 437752 46526 437804 46532
rect 438525 46588 438577 46594
rect 438525 46530 438577 46536
rect 437424 43214 437642 43220
rect 437424 43156 437642 43162
rect 436498 42602 436716 42608
rect 436498 42544 436716 42550
rect 437310 42490 437316 42660
rect 437368 42490 437374 42660
rect 437752 42608 437780 46526
rect 437876 46478 437904 46497
rect 437876 46472 437928 46478
rect 437876 46414 437928 46420
rect 437876 43272 437904 46414
rect 437860 43102 437866 43272
rect 437918 43102 437924 43272
rect 438525 42660 438553 46530
rect 438719 46482 438747 46497
rect 438695 46476 438747 46482
rect 438695 46418 438747 46424
rect 438719 43220 438747 46418
rect 438948 46422 438976 46497
rect 438948 46416 439000 46422
rect 438948 46358 439000 46364
rect 438620 43214 438838 43220
rect 438620 43156 438838 43162
rect 437694 42602 437912 42608
rect 437694 42544 437912 42550
rect 438506 42490 438512 42660
rect 438564 42490 438570 42660
rect 438948 42608 438976 46358
rect 439072 46310 439100 46497
rect 439721 46426 439749 46497
rect 439721 46420 439773 46426
rect 439721 46362 439773 46368
rect 439072 46304 439124 46310
rect 439072 46246 439124 46252
rect 439072 43272 439100 46246
rect 439056 43102 439062 43272
rect 439114 43102 439120 43272
rect 439721 42660 439749 46362
rect 439915 46314 439943 46497
rect 439915 46308 439967 46314
rect 439915 46250 439967 46256
rect 440144 46254 440172 46497
rect 440917 46258 440945 46497
rect 439915 43220 439943 46250
rect 440144 46248 440196 46254
rect 440144 46190 440196 46196
rect 440917 46252 440969 46258
rect 440917 46194 440969 46200
rect 439816 43214 440034 43220
rect 439816 43156 440034 43162
rect 438890 42602 439108 42608
rect 438890 42544 439108 42550
rect 439702 42490 439708 42660
rect 439760 42490 439766 42660
rect 440144 42608 440172 46190
rect 440422 43997 440795 44011
rect 440422 43937 440430 43997
rect 440787 43937 440795 43997
rect 440422 43925 440795 43937
rect 440422 42909 440795 42923
rect 440422 42849 440430 42909
rect 440787 42849 440795 42909
rect 440422 42837 440795 42849
rect 440917 42660 440945 46194
rect 447444 45134 447472 46497
rect 448287 45138 448315 46497
rect 447444 45128 447496 45134
rect 447444 45070 447496 45076
rect 448287 45132 448339 45138
rect 448287 45074 448339 45080
rect 448516 45078 448544 46497
rect 441618 43450 441991 43462
rect 441618 43390 441626 43450
rect 441983 43390 441991 43450
rect 441618 43376 441991 43390
rect 447444 43272 447472 45070
rect 447428 43102 447434 43272
rect 447486 43102 447492 43272
rect 448287 43220 448315 45074
rect 448516 45072 448568 45078
rect 448516 45014 448568 45020
rect 448188 43214 448406 43220
rect 448188 43156 448406 43162
rect 440086 42602 440304 42608
rect 440086 42544 440304 42550
rect 440898 42490 440904 42660
rect 440956 42490 440962 42660
rect 448516 42608 448544 45014
rect 448640 44966 448668 46497
rect 449289 45082 449317 46497
rect 449289 45076 449341 45082
rect 449289 45018 449341 45024
rect 448640 44960 448692 44966
rect 448640 44902 448692 44908
rect 448640 43272 448668 44902
rect 448624 43102 448630 43272
rect 448682 43102 448688 43272
rect 449289 42660 449317 45018
rect 449483 44970 449511 46497
rect 449483 44964 449535 44970
rect 449483 44906 449535 44912
rect 449712 44910 449740 46497
rect 449483 43220 449511 44906
rect 449712 44904 449764 44910
rect 449712 44846 449764 44852
rect 449384 43214 449602 43220
rect 449384 43156 449602 43162
rect 448458 42602 448676 42608
rect 448458 42544 448676 42550
rect 449270 42490 449276 42660
rect 449328 42490 449334 42660
rect 449712 42608 449740 44846
rect 449836 44798 449864 46497
rect 450485 44914 450513 46497
rect 450485 44908 450537 44914
rect 450485 44850 450537 44856
rect 449836 44792 449888 44798
rect 449836 44734 449888 44740
rect 449836 43272 449864 44734
rect 449820 43102 449826 43272
rect 449878 43102 449884 43272
rect 450485 42660 450513 44850
rect 450679 44802 450707 46497
rect 450655 44796 450707 44802
rect 450655 44738 450707 44744
rect 450679 43220 450707 44738
rect 450908 44742 450936 46497
rect 450908 44736 450960 44742
rect 450908 44678 450960 44684
rect 450580 43214 450798 43220
rect 450580 43156 450798 43162
rect 449654 42602 449872 42608
rect 449654 42544 449872 42550
rect 450466 42490 450472 42660
rect 450524 42490 450530 42660
rect 450908 42608 450936 44678
rect 451032 44630 451060 46497
rect 451681 44746 451709 46497
rect 451681 44740 451733 44746
rect 451681 44682 451733 44688
rect 451032 44624 451084 44630
rect 451032 44566 451084 44572
rect 451032 43272 451060 44566
rect 451016 43102 451022 43272
rect 451074 43102 451080 43272
rect 451681 42660 451709 44682
rect 451875 44634 451903 46497
rect 451875 44628 451927 44634
rect 451875 44570 451927 44576
rect 452104 44574 452132 46497
rect 451875 43220 451903 44570
rect 452104 44568 452156 44574
rect 452104 44510 452156 44516
rect 451776 43214 451994 43220
rect 451776 43156 451994 43162
rect 450850 42602 451068 42608
rect 450850 42544 451068 42550
rect 451662 42490 451668 42660
rect 451720 42490 451726 42660
rect 452104 42608 452132 44510
rect 452228 44462 452256 46497
rect 452877 44578 452905 46497
rect 452877 44572 452929 44578
rect 452877 44514 452929 44520
rect 452228 44456 452280 44462
rect 452228 44398 452280 44404
rect 452228 43272 452256 44398
rect 452212 43102 452218 43272
rect 452270 43102 452276 43272
rect 452877 42660 452905 44514
rect 453071 44466 453099 46497
rect 453047 44460 453099 44466
rect 453047 44402 453099 44408
rect 453071 43220 453099 44402
rect 453300 44350 453328 46497
rect 453300 44344 453352 44350
rect 453300 44286 453352 44292
rect 452972 43214 453190 43220
rect 452972 43156 453190 43162
rect 453300 42834 453328 44286
rect 453424 44238 453452 46497
rect 454073 44354 454101 46497
rect 454073 44348 454125 44354
rect 454073 44290 454125 44296
rect 453424 44232 453476 44238
rect 453424 44174 453476 44180
rect 453424 43272 453452 44174
rect 453408 43102 453414 43272
rect 453466 43102 453472 43272
rect 454073 42834 454101 44290
rect 454267 44242 454295 46497
rect 454267 44236 454319 44242
rect 454267 44178 454319 44184
rect 454267 43220 454295 44178
rect 454168 43214 454386 43220
rect 454168 43156 454386 43162
rect 453300 42806 453455 42834
rect 454073 42806 454228 42834
rect 453427 42660 453455 42806
rect 452046 42602 452264 42608
rect 452046 42544 452264 42550
rect 452858 42490 452864 42660
rect 452916 42490 452922 42660
rect 453410 42490 453416 42660
rect 453468 42490 453474 42660
rect 454200 42608 454228 42806
rect 454068 42602 454286 42608
rect 454068 42544 454286 42550
rect 147387 42375 147760 42384
rect 147387 42315 147395 42375
rect 147752 42315 147760 42375
rect 147387 42298 147760 42315
rect 441618 42368 441991 42377
rect 441618 42308 441626 42368
rect 441983 42308 441991 42368
rect 441618 42291 441991 42308
<< via2 >>
rect 676093 724496 676153 724853
rect 677175 724496 677235 724853
rect 675546 723300 675606 723657
rect 676634 723300 676694 723657
rect 40371 604610 40431 604967
rect 41453 604610 41513 604967
rect 40912 603414 40972 603771
rect 42000 603414 42060 603771
rect 676085 448095 676145 448452
rect 677167 448095 677227 448452
rect 675538 446899 675598 447256
rect 676626 446899 676686 447256
rect 40390 346959 40450 347316
rect 41472 346959 41532 347316
rect 40931 345763 40991 346120
rect 42019 345763 42079 346120
rect 146199 43944 146556 44004
rect 147395 43397 147752 43457
rect 146199 42856 146556 42916
rect 440430 43937 440787 43997
rect 440430 42849 440787 42909
rect 441626 43390 441983 43450
rect 147395 42315 147752 42375
rect 441626 42308 441983 42368
<< metal3 >>
rect 676078 724853 677583 724862
rect 676078 724496 676093 724853
rect 676153 724496 677175 724853
rect 677235 724496 677583 724853
rect 676078 724489 677583 724496
rect 675532 723657 677583 723664
rect 675532 723300 675546 723657
rect 675606 723300 676634 723657
rect 676694 723300 677583 723657
rect 675532 723294 677583 723300
rect 40023 604967 41528 604974
rect 40023 604610 40371 604967
rect 40431 604610 41453 604967
rect 41513 604610 41528 604967
rect 40023 604601 41528 604610
rect 40023 603771 42074 603777
rect 40023 603414 40912 603771
rect 40972 603414 42000 603771
rect 42060 603414 42074 603771
rect 40023 603407 42074 603414
rect 676070 448452 677575 448461
rect 676070 448095 676085 448452
rect 676145 448095 677167 448452
rect 677227 448095 677575 448452
rect 676070 448088 677575 448095
rect 675524 447256 677575 447263
rect 675524 446899 675538 447256
rect 675598 446899 676626 447256
rect 676686 446899 677575 447256
rect 675524 446893 677575 446899
rect 40042 347316 41547 347323
rect 40042 346959 40390 347316
rect 40450 346959 41472 347316
rect 41532 346959 41547 347316
rect 40042 346950 41547 346959
rect 40042 346120 42093 346126
rect 40042 345763 40931 346120
rect 40991 345763 42019 346120
rect 42079 345763 42093 346120
rect 40042 345756 42093 345763
rect 146193 44004 146563 44018
rect 146193 43944 146199 44004
rect 146556 43944 146563 44004
rect 146193 42916 146563 43944
rect 440424 43997 440794 44011
rect 440424 43937 440430 43997
rect 440787 43937 440794 43997
rect 146193 42856 146199 42916
rect 146556 42856 146563 42916
rect 146193 41967 146563 42856
rect 147388 43457 147761 43472
rect 147388 43397 147395 43457
rect 147752 43397 147761 43457
rect 147388 42375 147761 43397
rect 147388 42315 147395 42375
rect 147752 42315 147761 42375
rect 147388 41967 147761 42315
rect 440424 42909 440794 43937
rect 440424 42849 440430 42909
rect 440787 42849 440794 42909
rect 440424 41960 440794 42849
rect 441619 43450 441992 43465
rect 441619 43390 441626 43450
rect 441983 43390 441992 43450
rect 441619 42368 441992 43390
rect 441619 42308 441626 42368
rect 441983 42308 441992 42368
rect 441619 41960 441992 42308
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform 1 0 434076 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_1
timestamp 1663859327
transform 1 0 429292 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_2
timestamp 1663859327
transform 1 0 430488 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_3
timestamp 1663859327
transform 1 0 431684 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_4
timestamp 1663859327
transform 1 0 432880 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_5
timestamp 1663859327
transform 1 0 447232 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_6
timestamp 1663859327
transform 1 0 435272 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_7
timestamp 1663859327
transform 1 0 436468 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_8
timestamp 1663859327
transform 1 0 437664 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_9
timestamp 1663859327
transform 1 0 438860 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_10
timestamp 1663859327
transform 1 0 440056 0 -1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_11
timestamp 1663859327
transform 1 0 440056 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_12
timestamp 1663859327
transform 0 1 41504 -1 0 336973
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_13
timestamp 1663859327
transform 0 -1 676117 -1 0 721608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_14
timestamp 1663859327
transform 0 1 41504 -1 0 335777
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_15
timestamp 1663859327
transform 1 0 447232 0 1 42337
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_16
timestamp 1663859327
transform 1 0 448428 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_17
timestamp 1663859327
transform 1 0 450820 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_18
timestamp 1663859327
transform 1 0 449624 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_19
timestamp 1663859327
transform 1 0 452016 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_20
timestamp 1663859327
transform 1 0 453212 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_21
timestamp 1663859327
transform 1 0 133892 0 1 42337
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_22
timestamp 1663859327
transform 1 0 429292 0 1 42337
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_23
timestamp 1663859327
transform 1 0 135088 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_24
timestamp 1663859327
transform 1 0 133892 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_25
timestamp 1663859327
transform 1 0 137480 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_26
timestamp 1663859327
transform 1 0 136284 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_27
timestamp 1663859327
transform 1 0 138676 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_28
timestamp 1663859327
transform 1 0 141068 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_29
timestamp 1663859327
transform 1 0 139872 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_30
timestamp 1663859327
transform 1 0 142264 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_31
timestamp 1663859327
transform 1 0 144656 0 -1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_32
timestamp 1663859327
transform 1 0 143460 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_33
timestamp 1663859327
transform 1 0 144656 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_34
timestamp 1663859327
transform 1 0 151832 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_35
timestamp 1663859327
transform 0 1 41482 -1 0 600534
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_36
timestamp 1663859327
transform 0 1 41482 -1 0 602926
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_37
timestamp 1663859327
transform 0 1 41482 -1 0 601730
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_38
timestamp 1663859327
transform 1 0 154224 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_39
timestamp 1663859327
transform 1 0 151832 0 1 42337
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_40
timestamp 1663859327
transform 1 0 153028 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_41
timestamp 1663859327
transform 1 0 156616 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_42
timestamp 1663859327
transform 1 0 155420 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_43
timestamp 1663859327
transform 1 0 157812 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_44
timestamp 1663859327
transform 0 1 41504 -1 0 338169
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_45
timestamp 1663859327
transform 0 1 41504 -1 0 340561
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_46
timestamp 1663859327
transform 0 1 41504 -1 0 339365
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_47
timestamp 1663859327
transform 0 1 41504 -1 0 341757
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_48
timestamp 1663859327
transform 0 1 41504 -1 0 344149
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_49
timestamp 1663859327
transform 0 1 41504 -1 0 342953
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_50
timestamp 1663859327
transform 0 1 41504 -1 0 345345
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_51
timestamp 1663859327
transform 0 1 41482 -1 0 599338
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_52
timestamp 1663859327
transform 0 1 41482 -1 0 598142
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_53
timestamp 1663859327
transform 0 -1 676117 -1 0 446388
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_54
timestamp 1663859327
transform 0 -1 676117 -1 0 447584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_55
timestamp 1663859327
transform 0 -1 676117 -1 0 445192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_56
timestamp 1663859327
transform 0 -1 676117 -1 0 442800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_57
timestamp 1663859327
transform 0 -1 676117 -1 0 443996
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_58
timestamp 1663859327
transform 0 -1 676117 -1 0 440408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_59
timestamp 1663859327
transform 0 -1 676117 -1 0 441604
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform -1 0 134996 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_2
timestamp 1663859327
transform 1 0 153028 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_3
timestamp 1663859327
transform -1 0 154132 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_4
timestamp 1663859327
transform 1 0 155420 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_5
timestamp 1663859327
transform -1 0 156524 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_6
timestamp 1663859327
transform 1 0 156616 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_7
timestamp 1663859327
transform -1 0 157720 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_8
timestamp 1663859327
transform -1 0 158916 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_9
timestamp 1663859327
transform -1 0 158916 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_12
timestamp 1663859327
transform 0 -1 677205 1 0 439304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_13
timestamp 1663859327
transform 0 1 676117 -1 0 440408
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_24
timestamp 1663859327
transform 0 -1 677205 1 0 720504
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_25
timestamp 1663859327
transform 0 1 676117 -1 0 721608
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_34
timestamp 1663859327
transform 0 1 676117 -1 0 446388
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_35
timestamp 1663859327
transform 0 -1 677205 1 0 445284
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_36
timestamp 1663859327
transform 0 1 676117 -1 0 447584
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_37
timestamp 1663859327
transform 0 -1 677205 1 0 446480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_46
timestamp 1663859327
transform 0 1 676117 -1 0 441604
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_47
timestamp 1663859327
transform 0 -1 677205 1 0 440500
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_48
timestamp 1663859327
transform 0 -1 677205 1 0 441696
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_49
timestamp 1663859327
transform 0 1 676117 -1 0 442800
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_50
timestamp 1663859327
transform 0 -1 677205 1 0 442892
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_51
timestamp 1663859327
transform 0 1 676117 -1 0 443996
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_52
timestamp 1663859327
transform 0 -1 677205 1 0 444088
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_53
timestamp 1663859327
transform 0 1 676117 -1 0 445192
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_55
timestamp 1663859327
transform -1 0 152936 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_67
timestamp 1663859327
transform 1 0 144656 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_68
timestamp 1663859327
transform 1 0 143460 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_69
timestamp 1663859327
transform -1 0 144564 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_70
timestamp 1663859327
transform 1 0 142264 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_71
timestamp 1663859327
transform -1 0 143368 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_72
timestamp 1663859327
transform 1 0 141068 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_73
timestamp 1663859327
transform -1 0 142172 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_74
timestamp 1663859327
transform 1 0 139872 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_75
timestamp 1663859327
transform -1 0 140976 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_76
timestamp 1663859327
transform 1 0 138676 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_77
timestamp 1663859327
transform -1 0 139780 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_78
timestamp 1663859327
transform -1 0 138584 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_79
timestamp 1663859327
transform 1 0 137480 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_80
timestamp 1663859327
transform 1 0 136284 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_81
timestamp 1663859327
transform -1 0 137388 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_82
timestamp 1663859327
transform 1 0 135088 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_83
timestamp 1663859327
transform -1 0 136192 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_84
timestamp 1663859327
transform -1 0 155328 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_85
timestamp 1663859327
transform 1 0 154224 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_86
timestamp 1663859327
transform -1 0 430396 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_88
timestamp 1663859327
transform -1 0 431592 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_89
timestamp 1663859327
transform 1 0 430488 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_90
timestamp 1663859327
transform 1 0 431684 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_91
timestamp 1663859327
transform -1 0 432788 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_92
timestamp 1663859327
transform -1 0 433984 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_93
timestamp 1663859327
transform 1 0 432880 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_94
timestamp 1663859327
transform -1 0 435180 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_95
timestamp 1663859327
transform 1 0 434076 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_96
timestamp 1663859327
transform 1 0 435272 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_97
timestamp 1663859327
transform 1 0 436468 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_98
timestamp 1663859327
transform -1 0 436376 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_99
timestamp 1663859327
transform -1 0 437572 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_100
timestamp 1663859327
transform 1 0 437664 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_101
timestamp 1663859327
transform 1 0 438860 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_102
timestamp 1663859327
transform 1 0 440056 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_103
timestamp 1663859327
transform -1 0 438768 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_104
timestamp 1663859327
transform -1 0 439964 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_117
timestamp 1663859327
transform -1 0 448336 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_118
timestamp 1663859327
transform -1 0 449532 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_119
timestamp 1663859327
transform 1 0 448428 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_120
timestamp 1663859327
transform -1 0 450728 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_121
timestamp 1663859327
transform 1 0 449624 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_122
timestamp 1663859327
transform 1 0 450820 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_123
timestamp 1663859327
transform -1 0 451924 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_124
timestamp 1663859327
transform 1 0 452016 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_125
timestamp 1663859327
transform -1 0 454316 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_126
timestamp 1663859327
transform -1 0 453120 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_127
timestamp 1663859327
transform -1 0 454316 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_128
timestamp 1663859327
transform 0 -1 41504 -1 0 335777
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_129
timestamp 1663859327
transform 0 1 40416 1 0 334673
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_130
timestamp 1663859327
transform 0 -1 41504 -1 0 336973
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_131
timestamp 1663859327
transform 0 1 40416 1 0 335869
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_132
timestamp 1663859327
transform 0 -1 41504 -1 0 338169
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_133
timestamp 1663859327
transform 0 1 40416 1 0 337065
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_134
timestamp 1663859327
transform 0 -1 41504 -1 0 341757
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_135
timestamp 1663859327
transform 0 1 40416 1 0 340653
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_136
timestamp 1663859327
transform 0 -1 41504 -1 0 340561
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_137
timestamp 1663859327
transform 0 1 40416 1 0 339457
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_138
timestamp 1663859327
transform 0 1 40416 1 0 338261
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_139
timestamp 1663859327
transform 0 -1 41504 -1 0 339365
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_140
timestamp 1663859327
transform 0 1 40416 1 0 343045
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_141
timestamp 1663859327
transform 0 -1 41504 -1 0 344149
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_142
timestamp 1663859327
transform 0 1 40416 1 0 341849
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_143
timestamp 1663859327
transform 0 -1 41504 -1 0 342953
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_148
timestamp 1663859327
transform 0 1 40416 1 0 344241
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_149
timestamp 1663859327
transform 0 -1 41504 -1 0 345345
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_170
timestamp 1663859327
transform 0 1 40394 1 0 601822
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_171
timestamp 1663859327
transform 0 -1 41482 -1 0 602926
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_172
timestamp 1663859327
transform 0 -1 41482 -1 0 601730
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_173
timestamp 1663859327
transform 0 1 40394 1 0 600626
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_174
timestamp 1663859327
transform 0 1 40394 1 0 599430
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_175
timestamp 1663859327
transform 0 -1 41482 -1 0 600534
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_176
timestamp 1663859327
transform 0 1 40394 1 0 598234
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_177
timestamp 1663859327
transform 0 -1 41482 -1 0 599338
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_178
timestamp 1663859327
transform 0 1 40394 1 0 597038
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_179
timestamp 1663859327
transform 0 -1 41482 -1 0 598142
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform 0 -1 677205 -1 0 721700
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1663859327
transform -1 0 434076 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1663859327
transform -1 0 133892 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1663859327
transform -1 0 155420 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1663859327
transform -1 0 155420 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1663859327
transform -1 0 153028 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1663859327
transform -1 0 153028 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1663859327
transform -1 0 156616 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1663859327
transform -1 0 156616 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_10
timestamp 1663859327
transform -1 0 157812 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_11
timestamp 1663859327
transform -1 0 157812 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_12
timestamp 1663859327
transform -1 0 159008 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_13
timestamp 1663859327
transform -1 0 159008 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_16
timestamp 1663859327
transform 0 1 676117 -1 0 447676
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_17
timestamp 1663859327
transform 0 -1 677205 -1 0 447676
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_28
timestamp 1663859327
transform 0 1 676117 -1 0 720504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_29
timestamp 1663859327
transform 0 1 676117 -1 0 721700
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_38
timestamp 1663859327
transform 0 1 676117 -1 0 446480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_39
timestamp 1663859327
transform 0 -1 677205 -1 0 446480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_52
timestamp 1663859327
transform 0 -1 676117 -1 0 440500
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_53
timestamp 1663859327
transform 0 1 676117 -1 0 439304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_54
timestamp 1663859327
transform 0 -1 677205 -1 0 440500
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_55
timestamp 1663859327
transform 0 1 676117 -1 0 440500
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_56
timestamp 1663859327
transform 0 -1 677205 -1 0 441696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_57
timestamp 1663859327
transform 0 1 676117 -1 0 441696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_58
timestamp 1663859327
transform 0 -1 677205 -1 0 442892
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_59
timestamp 1663859327
transform 0 1 676117 -1 0 442892
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_60
timestamp 1663859327
transform 0 -1 677205 -1 0 444088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_61
timestamp 1663859327
transform 0 1 676117 -1 0 444088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_62
timestamp 1663859327
transform 0 -1 677205 -1 0 445284
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_63
timestamp 1663859327
transform 0 1 676117 -1 0 445284
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_64
timestamp 1663859327
transform -1 0 151832 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_65
timestamp 1663859327
transform -1 0 151832 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_74
timestamp 1663859327
transform -1 0 145852 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_75
timestamp 1663859327
transform -1 0 145852 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_76
timestamp 1663859327
transform -1 0 144656 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_77
timestamp 1663859327
transform -1 0 144656 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_78
timestamp 1663859327
transform -1 0 143460 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_79
timestamp 1663859327
transform -1 0 143460 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_80
timestamp 1663859327
transform -1 0 142264 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_81
timestamp 1663859327
transform -1 0 142264 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_82
timestamp 1663859327
transform -1 0 141068 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_83
timestamp 1663859327
transform -1 0 141068 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_84
timestamp 1663859327
transform -1 0 139872 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_85
timestamp 1663859327
transform -1 0 139872 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_86
timestamp 1663859327
transform -1 0 138676 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_87
timestamp 1663859327
transform -1 0 138676 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_88
timestamp 1663859327
transform -1 0 137480 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_89
timestamp 1663859327
transform -1 0 137480 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_90
timestamp 1663859327
transform -1 0 136284 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_91
timestamp 1663859327
transform -1 0 136284 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_92
timestamp 1663859327
transform -1 0 135088 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_93
timestamp 1663859327
transform -1 0 135088 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_94
timestamp 1663859327
transform -1 0 154224 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_95
timestamp 1663859327
transform -1 0 154224 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_96
timestamp 1663859327
transform -1 0 429292 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_97
timestamp 1663859327
transform -1 0 429292 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_98
timestamp 1663859327
transform -1 0 430488 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_99
timestamp 1663859327
transform -1 0 430488 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_100
timestamp 1663859327
transform -1 0 431684 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_101
timestamp 1663859327
transform -1 0 431684 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_102
timestamp 1663859327
transform -1 0 434076 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_103
timestamp 1663859327
transform -1 0 434076 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_104
timestamp 1663859327
transform -1 0 432880 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_105
timestamp 1663859327
transform -1 0 432880 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_106
timestamp 1663859327
transform -1 0 435272 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_107
timestamp 1663859327
transform -1 0 436468 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_108
timestamp 1663859327
transform -1 0 437664 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_109
timestamp 1663859327
transform -1 0 435272 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_110
timestamp 1663859327
transform -1 0 436468 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_111
timestamp 1663859327
transform -1 0 437664 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_112
timestamp 1663859327
transform -1 0 438860 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_113
timestamp 1663859327
transform -1 0 440056 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_114
timestamp 1663859327
transform -1 0 438860 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_115
timestamp 1663859327
transform -1 0 440056 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_116
timestamp 1663859327
transform -1 0 441252 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_117
timestamp 1663859327
transform -1 0 441252 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_126
timestamp 1663859327
transform -1 0 447232 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_127
timestamp 1663859327
transform -1 0 447232 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_128
timestamp 1663859327
transform -1 0 448428 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_129
timestamp 1663859327
transform -1 0 448428 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_130
timestamp 1663859327
transform -1 0 449624 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_131
timestamp 1663859327
transform -1 0 449624 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_132
timestamp 1663859327
transform -1 0 450820 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_133
timestamp 1663859327
transform -1 0 450820 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_134
timestamp 1663859327
transform -1 0 452016 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_135
timestamp 1663859327
transform -1 0 453212 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_136
timestamp 1663859327
transform -1 0 454408 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_137
timestamp 1663859327
transform -1 0 452016 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_138
timestamp 1663859327
transform -1 0 453212 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_139
timestamp 1663859327
transform -1 0 454408 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_140
timestamp 1663859327
transform 0 -1 41504 -1 0 334673
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_141
timestamp 1663859327
transform 0 1 41504 -1 0 334673
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_142
timestamp 1663859327
transform 0 -1 41504 -1 0 335869
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_143
timestamp 1663859327
transform 0 1 40416 -1 0 335869
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_144
timestamp 1663859327
transform 0 -1 41504 -1 0 337065
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_145
timestamp 1663859327
transform 0 1 40416 -1 0 337065
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_146
timestamp 1663859327
transform 0 1 40416 -1 0 340653
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_147
timestamp 1663859327
transform 0 -1 41504 -1 0 340653
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_148
timestamp 1663859327
transform 0 1 40416 -1 0 339457
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_149
timestamp 1663859327
transform 0 -1 41504 -1 0 339457
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_150
timestamp 1663859327
transform 0 1 40416 -1 0 338261
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_151
timestamp 1663859327
transform 0 -1 41504 -1 0 338261
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_152
timestamp 1663859327
transform 0 -1 41504 -1 0 343045
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_153
timestamp 1663859327
transform 0 1 40416 -1 0 343045
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_154
timestamp 1663859327
transform 0 -1 41504 -1 0 341849
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_155
timestamp 1663859327
transform 0 1 40416 -1 0 341849
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_158
timestamp 1663859327
transform 0 -1 41504 -1 0 345437
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_159
timestamp 1663859327
transform 0 1 40416 -1 0 345437
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_160
timestamp 1663859327
transform 0 -1 41504 -1 0 344241
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_161
timestamp 1663859327
transform 0 1 40416 -1 0 344241
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_184
timestamp 1663859327
transform 0 1 40394 -1 0 603018
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_185
timestamp 1663859327
transform 0 -1 41482 -1 0 603018
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_186
timestamp 1663859327
transform 0 -1 41482 -1 0 601822
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_187
timestamp 1663859327
transform 0 1 40394 -1 0 601822
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_188
timestamp 1663859327
transform 0 1 40394 -1 0 600626
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_189
timestamp 1663859327
transform 0 -1 41482 -1 0 600626
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_190
timestamp 1663859327
transform 0 1 40394 -1 0 598234
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_191
timestamp 1663859327
transform 0 1 40394 -1 0 599430
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_192
timestamp 1663859327
transform 0 -1 41482 -1 0 598234
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_193
timestamp 1663859327
transform 0 -1 41482 -1 0 599430
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_194
timestamp 1663859327
transform 0 1 40394 -1 0 597038
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_195
timestamp 1663859327
transform 0 -1 41482 -1 0 597038
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_218
timestamp 1663859327
transform -1 0 430488 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_219
timestamp 1663859327
transform -1 0 431684 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_220
timestamp 1663859327
transform -1 0 432880 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_221
timestamp 1663859327
transform -1 0 441252 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_222
timestamp 1663859327
transform -1 0 435272 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_223
timestamp 1663859327
transform -1 0 436468 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_224
timestamp 1663859327
transform -1 0 437664 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_225
timestamp 1663859327
transform -1 0 438860 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_226
timestamp 1663859327
transform -1 0 440056 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_231
timestamp 1663859327
transform -1 0 447232 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_232
timestamp 1663859327
transform -1 0 448428 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_233
timestamp 1663859327
transform -1 0 450820 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_234
timestamp 1663859327
transform -1 0 449624 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_235
timestamp 1663859327
transform -1 0 453212 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_236
timestamp 1663859327
transform -1 0 452016 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_237
timestamp 1663859327
transform -1 0 454408 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_238
timestamp 1663859327
transform -1 0 133892 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_239
timestamp 1663859327
transform -1 0 429292 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_240
timestamp 1663859327
transform -1 0 135088 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_241
timestamp 1663859327
transform -1 0 133892 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_242
timestamp 1663859327
transform -1 0 136284 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_243
timestamp 1663859327
transform -1 0 137480 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_244
timestamp 1663859327
transform -1 0 138676 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_245
timestamp 1663859327
transform -1 0 141068 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_246
timestamp 1663859327
transform -1 0 139872 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_247
timestamp 1663859327
transform -1 0 142264 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_248
timestamp 1663859327
transform -1 0 144656 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_249
timestamp 1663859327
transform -1 0 143460 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_250
timestamp 1663859327
transform -1 0 145852 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_255
timestamp 1663859327
transform -1 0 154224 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_256
timestamp 1663859327
transform -1 0 151832 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_257
timestamp 1663859327
transform -1 0 153028 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_258
timestamp 1663859327
transform -1 0 156616 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_259
timestamp 1663859327
transform -1 0 155420 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_260
timestamp 1663859327
transform -1 0 157812 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_261
timestamp 1663859327
transform 0 -1 677205 -1 0 439304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_262
timestamp 1663859327
transform 0 -1 676117 -1 0 439304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_263
timestamp 1663859327
transform 0 -1 676117 -1 0 442892
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_264
timestamp 1663859327
transform 0 -1 676117 -1 0 441696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_265
timestamp 1663859327
transform 0 -1 676117 -1 0 444088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_266
timestamp 1663859327
transform 0 -1 676117 -1 0 446480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_267
timestamp 1663859327
transform 0 -1 676117 -1 0 445284
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_269
timestamp 1663859327
transform 0 -1 676117 -1 0 447676
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_272
timestamp 1663859327
transform 0 -1 677205 -1 0 720504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_274
timestamp 1663859327
transform 0 -1 676117 -1 0 720504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_275
timestamp 1663859327
transform 0 -1 676117 -1 0 721700
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_297
timestamp 1663859327
transform 0 1 41482 -1 0 597038
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_298
timestamp 1663859327
transform 0 1 41482 -1 0 599430
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_299
timestamp 1663859327
transform 0 1 41482 -1 0 598234
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_300
timestamp 1663859327
transform 0 1 41482 -1 0 600626
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_301
timestamp 1663859327
transform 0 1 41482 -1 0 603018
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_302
timestamp 1663859327
transform 0 1 41482 -1 0 601822
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_309
timestamp 1663859327
transform 0 1 40416 -1 0 334673
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_310
timestamp 1663859327
transform 0 1 41504 -1 0 335869
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_311
timestamp 1663859327
transform 0 1 41504 -1 0 338261
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_312
timestamp 1663859327
transform 0 1 41504 -1 0 337065
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_313
timestamp 1663859327
transform 0 1 41504 -1 0 339457
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_314
timestamp 1663859327
transform 0 1 41504 -1 0 340653
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_315
timestamp 1663859327
transform 0 1 41504 -1 0 343045
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_316
timestamp 1663859327
transform 0 1 41504 -1 0 341849
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_317
timestamp 1663859327
transform 0 1 41504 -1 0 344241
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_318
timestamp 1663859327
transform 0 1 41504 -1 0 345437
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_326
timestamp 1663859327
transform -1 0 159008 0 1 43425
box -38 -48 130 592
<< labels >>
flabel metal3 677462 446931 677552 447228 0 FreeSans 400 90 0 0 vccd
port 136 nsew power input
flabel metal3 677464 448130 677554 448427 0 FreeSans 400 90 0 0 vssd
port 135 nsew ground input
flabel metal3 677461 723330 677551 723627 0 FreeSans 400 90 0 0 vccd
port 136 nsew power input
flabel metal3 677470 724527 677560 724824 0 FreeSans 400 90 0 0 vssd
port 135 nsew ground input
flabel metal1 673736 455568 673764 455855 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[4]
port 14 nsew signal input
flabel metal1 674156 728034 674184 728321 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[6]
port 10 nsew signal input
flabel metal1 673960 455968 673988 456255 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[5]
port 13 nsew signal input
flabel metal1 672840 453968 672868 454255 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[0]
port 18 nsew signal input
flabel metal1 673064 454368 673092 454655 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[1]
port 17 nsew signal input
flabel metal1 673288 454768 673316 455055 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[2]
port 16 nsew signal input
flabel metal1 673512 455168 673540 455455 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[3]
port 15 nsew signal input
flabel metal3 147432 41997 147738 42091 0 FreeSans 400 0 0 0 vssd
port 135 nsew ground input
flabel metal3 146226 41997 146532 42091 0 FreeSans 400 0 0 0 vccd
port 136 nsew power input
flabel metal3 441644 41978 441950 42072 0 FreeSans 400 0 0 0 vssd
port 135 nsew ground input
flabel metal3 440451 41984 440757 42078 0 FreeSans 400 0 0 0 vccd
port 136 nsew power input
flabel metal1 133123 44152 133374 44180 0 FreeSans 288 0 0 0 mgmt_io_oeb_buf[2]
port 93 nsew signal output
flabel metal1 131323 44992 131574 45020 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[16]
port 90 nsew signal input
flabel metal1 131723 44824 131974 44852 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[17]
port 89 nsew signal input
flabel metal1 132123 44656 132374 44684 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[18]
port 88 nsew signal input
flabel metal1 132523 44488 132774 44516 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[19]
port 87 nsew signal input
flabel metal1 132723 44376 132974 44404 0 FreeSans 288 0 0 0 mgmt_io_oeb_buf[0]
port 91 nsew signal output
flabel metal1 132923 44264 133174 44292 0 FreeSans 288 0 0 0 mgmt_io_oeb_buf[1]
port 92 nsew signal output
flabel metal3 40074 346985 40164 347282 0 FreeSans 400 90 0 0 vssd
port 135 nsew ground input
flabel metal3 40076 345792 40166 346089 0 FreeSans 400 90 0 0 vccd
port 136 nsew power input
flabel metal3 40053 604641 40143 604938 0 FreeSans 400 90 0 0 vssd
port 135 nsew ground input
flabel metal3 40053 603440 40143 603737 0 FreeSans 400 90 0 0 vccd
port 136 nsew power input
flabel metal1 45315 353236 45343 353530 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[15]
port 78 nsew signal input
flabel metal1 45091 353636 45119 353930 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[14]
port 79 nsew signal input
flabel metal1 44867 354036 44895 354330 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[13]
port 80 nsew signal input
flabel metal1 44643 354436 44671 354730 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[12]
port 81 nsew signal input
flabel metal1 673764 235250 673792 235537 0 FreeSans 288 90 0 0 mgmt_io_in_buf[4]
port 44 nsew signal output
flabel metal1 674212 234450 674240 234737 0 FreeSans 288 90 0 0 mgmt_io_in_buf[6]
port 42 nsew signal output
flabel metal1 673988 234850 674016 235137 0 FreeSans 288 90 0 0 mgmt_io_in_buf[5]
port 43 nsew signal output
flabel metal1 672868 236850 672896 237137 0 FreeSans 288 90 0 0 mgmt_io_in_buf[0]
port 48 nsew signal output
flabel metal1 673092 236450 673120 236737 0 FreeSans 288 90 0 0 mgmt_io_in_buf[1]
port 47 nsew signal output
flabel metal1 673316 236050 673344 236337 0 FreeSans 288 90 0 0 mgmt_io_in_buf[2]
port 46 nsew signal output
flabel metal1 673540 235650 673568 235937 0 FreeSans 288 90 0 0 mgmt_io_in_buf[3]
port 45 nsew signal output
flabel metal1 674352 229250 674380 229487 0 FreeSans 288 90 0 0 mgmt_io_in_buf[16]
port 100 nsew signal output
flabel metal1 674576 229650 674604 229887 0 FreeSans 288 90 0 0 mgmt_io_in_buf[17]
port 99 nsew signal output
flabel metal1 674800 230050 674828 230287 0 FreeSans 288 90 0 0 mgmt_io_in_buf[18]
port 98 nsew signal output
flabel metal1 675024 230450 675052 230687 0 FreeSans 288 90 0 0 mgmt_io_in_buf[19]
port 97 nsew signal output
flabel metal1 670936 223050 670964 223333 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[15]
port 105 nsew signal input
flabel metal1 671160 223450 671188 223733 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[14]
port 106 nsew signal input
flabel metal1 671384 223850 671412 224133 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[13]
port 107 nsew signal input
flabel metal1 671608 224250 671636 224533 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[12]
port 108 nsew signal input
flabel metal1 671832 224650 671860 224933 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[11]
port 109 nsew signal input
flabel metal1 672056 225050 672084 225333 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[10]
port 110 nsew signal input
flabel metal1 672280 225450 672308 225733 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[9]
port 111 nsew signal input
flabel metal1 672504 225850 672532 226133 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[8]
port 112 nsew signal input
flabel metal1 672728 226250 672756 226533 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[7]
port 113 nsew signal input
flabel metal1 675192 230650 675220 230887 0 FreeSans 288 90 0 0 mgmt_io_oeb_unbuf[0]
port 96 nsew signal input
flabel metal1 675528 231050 675556 231287 0 FreeSans 288 90 0 0 mgmt_io_oeb_unbuf[2]
port 94 nsew signal input
flabel metal1 675360 230850 675388 231087 0 FreeSans 288 90 0 0 mgmt_io_oeb_unbuf[1]
port 95 nsew signal input
flabel metal1 671048 223250 671076 223533 0 FreeSans 288 90 0 0 mgmt_io_in_buf[15]
port 134 nsew signal output
flabel metal1 671272 223650 671300 223933 0 FreeSans 288 90 0 0 mgmt_io_in_buf[14]
port 133 nsew signal output
flabel metal1 671496 224050 671524 224333 0 FreeSans 288 90 0 0 mgmt_io_in_buf[13]
port 132 nsew signal output
flabel metal1 671720 224450 671748 224733 0 FreeSans 288 90 0 0 mgmt_io_in_buf[12]
port 131 nsew signal output
flabel metal1 671944 224850 671972 225133 0 FreeSans 288 90 0 0 mgmt_io_in_buf[11]
port 130 nsew signal output
flabel metal1 672168 225250 672196 225533 0 FreeSans 288 90 0 0 mgmt_io_in_buf[10]
port 129 nsew signal output
flabel metal1 672392 225650 672420 225933 0 FreeSans 288 90 0 0 mgmt_io_in_buf[9]
port 128 nsew signal output
flabel metal1 672616 226050 672644 226333 0 FreeSans 288 90 0 0 mgmt_io_in_buf[8]
port 127 nsew signal output
flabel metal1 672840 226450 672868 226733 0 FreeSans 288 90 0 0 mgmt_io_in_buf[7]
port 126 nsew signal output
flabel metal1 674688 229850 674716 230087 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[18]
port 103 nsew signal input
flabel metal1 674464 229450 674492 229687 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[17]
port 102 nsew signal input
flabel metal1 674240 229050 674268 229287 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[16]
port 101 nsew signal input
flabel metal1 674912 230250 674940 230487 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[19]
port 104 nsew signal input
flabel metal1 672756 237050 672784 237337 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[0]
port 25 nsew signal input
flabel metal1 672980 236650 673008 236937 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[1]
port 26 nsew signal input
flabel metal1 673204 236250 673232 236537 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[2]
port 27 nsew signal input
flabel metal1 673428 235850 673456 236137 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[3]
port 28 nsew signal input
flabel metal1 673652 235450 673680 235737 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[4]
port 29 nsew signal input
flabel metal1 673876 235050 673904 235337 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[5]
port 30 nsew signal input
flabel metal1 674100 234650 674128 234937 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[6]
port 31 nsew signal input
flabel metal1 672728 453768 672756 454055 0 FreeSans 288 90 0 0 mgmt_io_out_buf[0]
port 19 nsew signal output
flabel metal1 672952 454168 672980 454455 0 FreeSans 288 90 0 0 mgmt_io_out_buf[1]
port 20 nsew signal output
flabel metal1 673176 454568 673204 454855 0 FreeSans 288 90 0 0 mgmt_io_out_buf[2]
port 21 nsew signal output
flabel metal1 673400 454968 673428 455255 0 FreeSans 288 90 0 0 mgmt_io_out_buf[3]
port 22 nsew signal output
flabel metal1 673624 455368 673652 455655 0 FreeSans 288 90 0 0 mgmt_io_out_buf[4]
port 23 nsew signal output
flabel metal1 673848 455768 673876 456055 0 FreeSans 288 90 0 0 mgmt_io_out_buf[5]
port 24 nsew signal output
flabel metal1 674044 727834 674072 728121 0 FreeSans 288 90 0 0 mgmt_io_out_buf[6]
port 12 nsew signal output
flabel metal1 44755 354236 44783 354530 0 FreeSans 288 90 0 0 mgmt_io_out_buf[12]
port 74 nsew signal output
flabel metal1 44979 353836 45007 354130 0 FreeSans 288 90 0 0 mgmt_io_out_buf[13]
port 75 nsew signal output
flabel metal1 45203 353436 45231 353730 0 FreeSans 288 90 0 0 mgmt_io_out_buf[14]
port 76 nsew signal output
flabel metal1 45427 353036 45455 353330 0 FreeSans 288 90 0 0 mgmt_io_out_buf[15]
port 77 nsew signal output
flabel metal1 131151 45076 131402 45104 0 FreeSans 288 0 0 0 mgmt_io_out_buf[16]
port 83 nsew signal output
flabel metal1 131551 44908 131802 44936 0 FreeSans 288 0 0 0 mgmt_io_out_buf[17]
port 84 nsew signal output
flabel metal1 131951 44740 132202 44768 0 FreeSans 288 0 0 0 mgmt_io_out_buf[18]
port 85 nsew signal output
flabel metal1 132351 44572 132602 44600 0 FreeSans 288 0 0 0 mgmt_io_out_buf[19]
port 86 nsew signal output
flabel metal1 44559 610495 44587 610756 0 FreeSans 288 90 0 0 mgmt_io_out_buf[11]
port 67 nsew signal output
flabel metal1 44335 610895 44363 611156 0 FreeSans 288 90 0 0 mgmt_io_out_buf[10]
port 66 nsew signal output
flabel metal1 44223 611095 44251 611356 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[10]
port 69 nsew signal input
flabel metal1 44447 610695 44475 610956 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[11]
port 68 nsew signal input
flabel metal1 44111 611334 44139 611595 0 FreeSans 288 90 0 0 mgmt_io_out_buf[9]
port 137 nsew
flabel metal1 43999 611534 44027 611795 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[9]
port 138 nsew
flabel metal1 43887 611734 43915 611995 0 FreeSans 288 90 0 0 mgmt_io_out_buf[8]
port 140 nsew
flabel metal1 43775 611934 43803 612195 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[8]
port 141 nsew
flabel metal1 43663 612107 43691 612368 0 FreeSans 288 90 0 0 mgmt_io_out_buf[7]
port 142 nsew
flabel metal1 43551 612307 43579 612568 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[7]
port 143 nsew
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
