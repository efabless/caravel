VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mgmt_protect_hv
  CLASS BLOCK ;
  FOREIGN mgmt_protect_hv ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 20.000 ;
  PIN vccd
    PORT
      LAYER met3 ;
        RECT 4.800 15.365 149.760 15.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.800 4.565 149.760 5.065 ;
    END
    PORT
      LAYER met2 ;
        RECT 94.650 3.815 94.950 16.535 ;
    END
  END vccd
  PIN vssd
    PORT
      LAYER met3 ;
        RECT 4.800 9.965 149.760 10.465 ;
    END
    PORT
      LAYER met2 ;
        RECT 134.650 3.815 134.950 16.535 ;
    END
    PORT
      LAYER met2 ;
        RECT 54.650 3.815 54.950 16.535 ;
    END
  END vssd
  PIN vdda1
    PORT
      LAYER met3 ;
        RECT 4.800 6.820 149.760 7.320 ;
    END
    PORT
      LAYER met2 ;
        RECT 96.650 4.070 96.950 16.280 ;
    END
  END vdda1
  PIN vssa1
    PORT
      LAYER met3 ;
        RECT 4.800 12.220 149.760 12.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 136.650 4.070 136.950 16.280 ;
    END
    PORT
      LAYER met2 ;
        RECT 56.650 4.070 56.950 16.280 ;
    END
  END vssa1
  PIN vdda2
    PORT
      LAYER met3 ;
        RECT 4.800 8.820 149.760 9.320 ;
    END
    PORT
      LAYER met2 ;
        RECT 98.650 4.070 98.950 16.280 ;
    END
  END vdda2
  PIN vssa2
    PORT
      LAYER met3 ;
        RECT 4.800 14.220 149.760 14.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 138.650 4.070 138.950 16.280 ;
    END
    PORT
      LAYER met2 ;
        RECT 58.650 4.070 58.950 16.280 ;
    END
  END vssa2
  PIN mprj2_vdd_logic1
    PORT
      LAYER met3 ;
        RECT 0.000 4.510 4.000 5.110 ;
    END
  END mprj2_vdd_logic1
  PIN mprj_vdd_logic1
    PORT
      LAYER met3 ;
        RECT 0.000 14.130 4.000 14.730 ;
    END
  END mprj_vdd_logic1
  OBS
      LAYER nwell ;
        RECT 147.640 10.025 150.090 14.395 ;
      LAYER li1 ;
        RECT 31.680 8.055 149.760 16.365 ;
      LAYER met1 ;
        RECT 3.920 3.815 149.760 16.535 ;
      LAYER met2 ;
        RECT 3.940 4.625 54.370 14.855 ;
        RECT 55.230 4.625 56.370 14.855 ;
        RECT 57.230 4.625 58.370 14.855 ;
        RECT 59.230 4.625 94.370 14.855 ;
        RECT 95.230 4.625 96.370 14.855 ;
        RECT 97.230 4.625 98.370 14.855 ;
        RECT 99.230 4.625 134.370 14.855 ;
        RECT 135.230 4.625 136.370 14.855 ;
        RECT 137.230 4.625 138.370 14.855 ;
        RECT 139.230 4.625 146.560 14.855 ;
      LAYER met3 ;
        RECT 4.400 13.730 146.585 13.820 ;
        RECT 4.000 13.120 146.585 13.730 ;
        RECT 4.000 11.820 4.400 13.120 ;
        RECT 4.000 10.865 146.585 11.820 ;
        RECT 4.000 8.420 4.400 10.865 ;
        RECT 4.000 7.720 146.585 8.420 ;
        RECT 4.000 6.420 4.400 7.720 ;
        RECT 4.000 5.510 146.585 6.420 ;
        RECT 4.400 5.465 146.585 5.510 ;
  END
END mgmt_protect_hv
END LIBRARY

