magic
tech sky130A
timestamp 1598786981
<< metal5 >>
rect 0 3240 1620 3780
rect 0 540 540 3240
rect 1080 540 1620 3240
rect 0 0 1620 540
<< properties >>
string FIXED_BBOX 0 -1080 2160 3780
<< end >>
