VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mgmt_protect
  CLASS BLOCK ;
  FOREIGN mgmt_protect ;
  ORIGIN 0.000 0.000 ;
  SIZE 1900.000 BY 160.000 ;
  PIN caravel_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 6.160 1902.000 6.760 ;
    END
  END caravel_clk
  PIN caravel_clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 18.400 1902.000 19.000 ;
    END
  END caravel_clk2
  PIN caravel_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 30.640 1902.000 31.240 ;
    END
  END caravel_rstn
  PIN la_data_in_core[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 156.000 432.770 162.000 ;
    END
  END la_data_in_core[0]
  PIN la_data_in_core[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.490 156.000 1536.770 162.000 ;
    END
  END la_data_in_core[100]
  PIN la_data_in_core[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1547.530 156.000 1547.810 162.000 ;
    END
  END la_data_in_core[101]
  PIN la_data_in_core[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1558.570 156.000 1558.850 162.000 ;
    END
  END la_data_in_core[102]
  PIN la_data_in_core[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1569.610 156.000 1569.890 162.000 ;
    END
  END la_data_in_core[103]
  PIN la_data_in_core[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.650 156.000 1580.930 162.000 ;
    END
  END la_data_in_core[104]
  PIN la_data_in_core[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1591.690 156.000 1591.970 162.000 ;
    END
  END la_data_in_core[105]
  PIN la_data_in_core[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1602.730 156.000 1603.010 162.000 ;
    END
  END la_data_in_core[106]
  PIN la_data_in_core[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1613.770 156.000 1614.050 162.000 ;
    END
  END la_data_in_core[107]
  PIN la_data_in_core[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1624.810 156.000 1625.090 162.000 ;
    END
  END la_data_in_core[108]
  PIN la_data_in_core[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1635.850 156.000 1636.130 162.000 ;
    END
  END la_data_in_core[109]
  PIN la_data_in_core[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 156.000 543.170 162.000 ;
    END
  END la_data_in_core[10]
  PIN la_data_in_core[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1646.890 156.000 1647.170 162.000 ;
    END
  END la_data_in_core[110]
  PIN la_data_in_core[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.930 156.000 1658.210 162.000 ;
    END
  END la_data_in_core[111]
  PIN la_data_in_core[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.970 156.000 1669.250 162.000 ;
    END
  END la_data_in_core[112]
  PIN la_data_in_core[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1680.010 156.000 1680.290 162.000 ;
    END
  END la_data_in_core[113]
  PIN la_data_in_core[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.050 156.000 1691.330 162.000 ;
    END
  END la_data_in_core[114]
  PIN la_data_in_core[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1702.090 156.000 1702.370 162.000 ;
    END
  END la_data_in_core[115]
  PIN la_data_in_core[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1713.130 156.000 1713.410 162.000 ;
    END
  END la_data_in_core[116]
  PIN la_data_in_core[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1724.170 156.000 1724.450 162.000 ;
    END
  END la_data_in_core[117]
  PIN la_data_in_core[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1735.210 156.000 1735.490 162.000 ;
    END
  END la_data_in_core[118]
  PIN la_data_in_core[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.250 156.000 1746.530 162.000 ;
    END
  END la_data_in_core[119]
  PIN la_data_in_core[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 156.000 554.210 162.000 ;
    END
  END la_data_in_core[11]
  PIN la_data_in_core[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1757.290 156.000 1757.570 162.000 ;
    END
  END la_data_in_core[120]
  PIN la_data_in_core[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1768.330 156.000 1768.610 162.000 ;
    END
  END la_data_in_core[121]
  PIN la_data_in_core[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1779.370 156.000 1779.650 162.000 ;
    END
  END la_data_in_core[122]
  PIN la_data_in_core[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1790.410 156.000 1790.690 162.000 ;
    END
  END la_data_in_core[123]
  PIN la_data_in_core[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1801.450 156.000 1801.730 162.000 ;
    END
  END la_data_in_core[124]
  PIN la_data_in_core[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1812.490 156.000 1812.770 162.000 ;
    END
  END la_data_in_core[125]
  PIN la_data_in_core[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1823.530 156.000 1823.810 162.000 ;
    END
  END la_data_in_core[126]
  PIN la_data_in_core[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.570 156.000 1834.850 162.000 ;
    END
  END la_data_in_core[127]
  PIN la_data_in_core[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 156.000 565.250 162.000 ;
    END
  END la_data_in_core[12]
  PIN la_data_in_core[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 156.000 576.290 162.000 ;
    END
  END la_data_in_core[13]
  PIN la_data_in_core[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 156.000 587.330 162.000 ;
    END
  END la_data_in_core[14]
  PIN la_data_in_core[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 156.000 598.370 162.000 ;
    END
  END la_data_in_core[15]
  PIN la_data_in_core[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.130 156.000 609.410 162.000 ;
    END
  END la_data_in_core[16]
  PIN la_data_in_core[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.170 156.000 620.450 162.000 ;
    END
  END la_data_in_core[17]
  PIN la_data_in_core[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 156.000 631.490 162.000 ;
    END
  END la_data_in_core[18]
  PIN la_data_in_core[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.250 156.000 642.530 162.000 ;
    END
  END la_data_in_core[19]
  PIN la_data_in_core[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 156.000 443.810 162.000 ;
    END
  END la_data_in_core[1]
  PIN la_data_in_core[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 156.000 653.570 162.000 ;
    END
  END la_data_in_core[20]
  PIN la_data_in_core[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.330 156.000 664.610 162.000 ;
    END
  END la_data_in_core[21]
  PIN la_data_in_core[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.370 156.000 675.650 162.000 ;
    END
  END la_data_in_core[22]
  PIN la_data_in_core[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.410 156.000 686.690 162.000 ;
    END
  END la_data_in_core[23]
  PIN la_data_in_core[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.450 156.000 697.730 162.000 ;
    END
  END la_data_in_core[24]
  PIN la_data_in_core[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 156.000 708.770 162.000 ;
    END
  END la_data_in_core[25]
  PIN la_data_in_core[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.530 156.000 719.810 162.000 ;
    END
  END la_data_in_core[26]
  PIN la_data_in_core[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.570 156.000 730.850 162.000 ;
    END
  END la_data_in_core[27]
  PIN la_data_in_core[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 156.000 741.890 162.000 ;
    END
  END la_data_in_core[28]
  PIN la_data_in_core[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.650 156.000 752.930 162.000 ;
    END
  END la_data_in_core[29]
  PIN la_data_in_core[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.570 156.000 454.850 162.000 ;
    END
  END la_data_in_core[2]
  PIN la_data_in_core[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.690 156.000 763.970 162.000 ;
    END
  END la_data_in_core[30]
  PIN la_data_in_core[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.730 156.000 775.010 162.000 ;
    END
  END la_data_in_core[31]
  PIN la_data_in_core[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 156.000 786.050 162.000 ;
    END
  END la_data_in_core[32]
  PIN la_data_in_core[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.810 156.000 797.090 162.000 ;
    END
  END la_data_in_core[33]
  PIN la_data_in_core[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.850 156.000 808.130 162.000 ;
    END
  END la_data_in_core[34]
  PIN la_data_in_core[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.890 156.000 819.170 162.000 ;
    END
  END la_data_in_core[35]
  PIN la_data_in_core[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.930 156.000 830.210 162.000 ;
    END
  END la_data_in_core[36]
  PIN la_data_in_core[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.970 156.000 841.250 162.000 ;
    END
  END la_data_in_core[37]
  PIN la_data_in_core[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.010 156.000 852.290 162.000 ;
    END
  END la_data_in_core[38]
  PIN la_data_in_core[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 156.000 863.330 162.000 ;
    END
  END la_data_in_core[39]
  PIN la_data_in_core[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 156.000 465.890 162.000 ;
    END
  END la_data_in_core[3]
  PIN la_data_in_core[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.090 156.000 874.370 162.000 ;
    END
  END la_data_in_core[40]
  PIN la_data_in_core[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.130 156.000 885.410 162.000 ;
    END
  END la_data_in_core[41]
  PIN la_data_in_core[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.170 156.000 896.450 162.000 ;
    END
  END la_data_in_core[42]
  PIN la_data_in_core[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.210 156.000 907.490 162.000 ;
    END
  END la_data_in_core[43]
  PIN la_data_in_core[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.250 156.000 918.530 162.000 ;
    END
  END la_data_in_core[44]
  PIN la_data_in_core[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.290 156.000 929.570 162.000 ;
    END
  END la_data_in_core[45]
  PIN la_data_in_core[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.330 156.000 940.610 162.000 ;
    END
  END la_data_in_core[46]
  PIN la_data_in_core[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.370 156.000 951.650 162.000 ;
    END
  END la_data_in_core[47]
  PIN la_data_in_core[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.410 156.000 962.690 162.000 ;
    END
  END la_data_in_core[48]
  PIN la_data_in_core[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 973.450 156.000 973.730 162.000 ;
    END
  END la_data_in_core[49]
  PIN la_data_in_core[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 156.000 476.930 162.000 ;
    END
  END la_data_in_core[4]
  PIN la_data_in_core[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.490 156.000 984.770 162.000 ;
    END
  END la_data_in_core[50]
  PIN la_data_in_core[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.530 156.000 995.810 162.000 ;
    END
  END la_data_in_core[51]
  PIN la_data_in_core[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1006.570 156.000 1006.850 162.000 ;
    END
  END la_data_in_core[52]
  PIN la_data_in_core[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.610 156.000 1017.890 162.000 ;
    END
  END la_data_in_core[53]
  PIN la_data_in_core[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1028.650 156.000 1028.930 162.000 ;
    END
  END la_data_in_core[54]
  PIN la_data_in_core[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1039.690 156.000 1039.970 162.000 ;
    END
  END la_data_in_core[55]
  PIN la_data_in_core[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.730 156.000 1051.010 162.000 ;
    END
  END la_data_in_core[56]
  PIN la_data_in_core[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.770 156.000 1062.050 162.000 ;
    END
  END la_data_in_core[57]
  PIN la_data_in_core[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.810 156.000 1073.090 162.000 ;
    END
  END la_data_in_core[58]
  PIN la_data_in_core[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1083.850 156.000 1084.130 162.000 ;
    END
  END la_data_in_core[59]
  PIN la_data_in_core[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 156.000 487.970 162.000 ;
    END
  END la_data_in_core[5]
  PIN la_data_in_core[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.890 156.000 1095.170 162.000 ;
    END
  END la_data_in_core[60]
  PIN la_data_in_core[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1105.930 156.000 1106.210 162.000 ;
    END
  END la_data_in_core[61]
  PIN la_data_in_core[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.970 156.000 1117.250 162.000 ;
    END
  END la_data_in_core[62]
  PIN la_data_in_core[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.010 156.000 1128.290 162.000 ;
    END
  END la_data_in_core[63]
  PIN la_data_in_core[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.050 156.000 1139.330 162.000 ;
    END
  END la_data_in_core[64]
  PIN la_data_in_core[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.090 156.000 1150.370 162.000 ;
    END
  END la_data_in_core[65]
  PIN la_data_in_core[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1161.130 156.000 1161.410 162.000 ;
    END
  END la_data_in_core[66]
  PIN la_data_in_core[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.170 156.000 1172.450 162.000 ;
    END
  END la_data_in_core[67]
  PIN la_data_in_core[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1183.210 156.000 1183.490 162.000 ;
    END
  END la_data_in_core[68]
  PIN la_data_in_core[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.250 156.000 1194.530 162.000 ;
    END
  END la_data_in_core[69]
  PIN la_data_in_core[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 156.000 499.010 162.000 ;
    END
  END la_data_in_core[6]
  PIN la_data_in_core[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1205.290 156.000 1205.570 162.000 ;
    END
  END la_data_in_core[70]
  PIN la_data_in_core[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1216.330 156.000 1216.610 162.000 ;
    END
  END la_data_in_core[71]
  PIN la_data_in_core[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.370 156.000 1227.650 162.000 ;
    END
  END la_data_in_core[72]
  PIN la_data_in_core[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1238.410 156.000 1238.690 162.000 ;
    END
  END la_data_in_core[73]
  PIN la_data_in_core[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.450 156.000 1249.730 162.000 ;
    END
  END la_data_in_core[74]
  PIN la_data_in_core[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1260.490 156.000 1260.770 162.000 ;
    END
  END la_data_in_core[75]
  PIN la_data_in_core[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.530 156.000 1271.810 162.000 ;
    END
  END la_data_in_core[76]
  PIN la_data_in_core[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1282.570 156.000 1282.850 162.000 ;
    END
  END la_data_in_core[77]
  PIN la_data_in_core[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1293.610 156.000 1293.890 162.000 ;
    END
  END la_data_in_core[78]
  PIN la_data_in_core[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.650 156.000 1304.930 162.000 ;
    END
  END la_data_in_core[79]
  PIN la_data_in_core[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 156.000 510.050 162.000 ;
    END
  END la_data_in_core[7]
  PIN la_data_in_core[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1315.690 156.000 1315.970 162.000 ;
    END
  END la_data_in_core[80]
  PIN la_data_in_core[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.730 156.000 1327.010 162.000 ;
    END
  END la_data_in_core[81]
  PIN la_data_in_core[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1337.770 156.000 1338.050 162.000 ;
    END
  END la_data_in_core[82]
  PIN la_data_in_core[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1348.810 156.000 1349.090 162.000 ;
    END
  END la_data_in_core[83]
  PIN la_data_in_core[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1359.850 156.000 1360.130 162.000 ;
    END
  END la_data_in_core[84]
  PIN la_data_in_core[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1370.890 156.000 1371.170 162.000 ;
    END
  END la_data_in_core[85]
  PIN la_data_in_core[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.930 156.000 1382.210 162.000 ;
    END
  END la_data_in_core[86]
  PIN la_data_in_core[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1392.970 156.000 1393.250 162.000 ;
    END
  END la_data_in_core[87]
  PIN la_data_in_core[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.010 156.000 1404.290 162.000 ;
    END
  END la_data_in_core[88]
  PIN la_data_in_core[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.050 156.000 1415.330 162.000 ;
    END
  END la_data_in_core[89]
  PIN la_data_in_core[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 156.000 521.090 162.000 ;
    END
  END la_data_in_core[8]
  PIN la_data_in_core[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.090 156.000 1426.370 162.000 ;
    END
  END la_data_in_core[90]
  PIN la_data_in_core[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1437.130 156.000 1437.410 162.000 ;
    END
  END la_data_in_core[91]
  PIN la_data_in_core[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1448.170 156.000 1448.450 162.000 ;
    END
  END la_data_in_core[92]
  PIN la_data_in_core[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1459.210 156.000 1459.490 162.000 ;
    END
  END la_data_in_core[93]
  PIN la_data_in_core[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1470.250 156.000 1470.530 162.000 ;
    END
  END la_data_in_core[94]
  PIN la_data_in_core[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.290 156.000 1481.570 162.000 ;
    END
  END la_data_in_core[95]
  PIN la_data_in_core[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.330 156.000 1492.610 162.000 ;
    END
  END la_data_in_core[96]
  PIN la_data_in_core[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.370 156.000 1503.650 162.000 ;
    END
  END la_data_in_core[97]
  PIN la_data_in_core[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1514.410 156.000 1514.690 162.000 ;
    END
  END la_data_in_core[98]
  PIN la_data_in_core[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1525.450 156.000 1525.730 162.000 ;
    END
  END la_data_in_core[99]
  PIN la_data_in_core[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 156.000 532.130 162.000 ;
    END
  END la_data_in_core[9]
  PIN la_data_in_mprj[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 -2.000 99.730 4.000 ;
    END
  END la_data_in_mprj[0]
  PIN la_data_in_mprj[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1203.450 -2.000 1203.730 4.000 ;
    END
  END la_data_in_mprj[100]
  PIN la_data_in_mprj[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.490 -2.000 1214.770 4.000 ;
    END
  END la_data_in_mprj[101]
  PIN la_data_in_mprj[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.530 -2.000 1225.810 4.000 ;
    END
  END la_data_in_mprj[102]
  PIN la_data_in_mprj[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1236.570 -2.000 1236.850 4.000 ;
    END
  END la_data_in_mprj[103]
  PIN la_data_in_mprj[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.610 -2.000 1247.890 4.000 ;
    END
  END la_data_in_mprj[104]
  PIN la_data_in_mprj[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1258.650 -2.000 1258.930 4.000 ;
    END
  END la_data_in_mprj[105]
  PIN la_data_in_mprj[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.690 -2.000 1269.970 4.000 ;
    END
  END la_data_in_mprj[106]
  PIN la_data_in_mprj[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.730 -2.000 1281.010 4.000 ;
    END
  END la_data_in_mprj[107]
  PIN la_data_in_mprj[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.770 -2.000 1292.050 4.000 ;
    END
  END la_data_in_mprj[108]
  PIN la_data_in_mprj[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1302.810 -2.000 1303.090 4.000 ;
    END
  END la_data_in_mprj[109]
  PIN la_data_in_mprj[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 -2.000 210.130 4.000 ;
    END
  END la_data_in_mprj[10]
  PIN la_data_in_mprj[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.850 -2.000 1314.130 4.000 ;
    END
  END la_data_in_mprj[110]
  PIN la_data_in_mprj[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1324.890 -2.000 1325.170 4.000 ;
    END
  END la_data_in_mprj[111]
  PIN la_data_in_mprj[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.930 -2.000 1336.210 4.000 ;
    END
  END la_data_in_mprj[112]
  PIN la_data_in_mprj[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.970 -2.000 1347.250 4.000 ;
    END
  END la_data_in_mprj[113]
  PIN la_data_in_mprj[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.010 -2.000 1358.290 4.000 ;
    END
  END la_data_in_mprj[114]
  PIN la_data_in_mprj[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1369.050 -2.000 1369.330 4.000 ;
    END
  END la_data_in_mprj[115]
  PIN la_data_in_mprj[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1380.090 -2.000 1380.370 4.000 ;
    END
  END la_data_in_mprj[116]
  PIN la_data_in_mprj[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.130 -2.000 1391.410 4.000 ;
    END
  END la_data_in_mprj[117]
  PIN la_data_in_mprj[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1402.170 -2.000 1402.450 4.000 ;
    END
  END la_data_in_mprj[118]
  PIN la_data_in_mprj[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.210 -2.000 1413.490 4.000 ;
    END
  END la_data_in_mprj[119]
  PIN la_data_in_mprj[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 -2.000 221.170 4.000 ;
    END
  END la_data_in_mprj[11]
  PIN la_data_in_mprj[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1424.250 -2.000 1424.530 4.000 ;
    END
  END la_data_in_mprj[120]
  PIN la_data_in_mprj[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.290 -2.000 1435.570 4.000 ;
    END
  END la_data_in_mprj[121]
  PIN la_data_in_mprj[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1446.330 -2.000 1446.610 4.000 ;
    END
  END la_data_in_mprj[122]
  PIN la_data_in_mprj[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1457.370 -2.000 1457.650 4.000 ;
    END
  END la_data_in_mprj[123]
  PIN la_data_in_mprj[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.410 -2.000 1468.690 4.000 ;
    END
  END la_data_in_mprj[124]
  PIN la_data_in_mprj[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1479.450 -2.000 1479.730 4.000 ;
    END
  END la_data_in_mprj[125]
  PIN la_data_in_mprj[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.490 -2.000 1490.770 4.000 ;
    END
  END la_data_in_mprj[126]
  PIN la_data_in_mprj[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1501.530 -2.000 1501.810 4.000 ;
    END
  END la_data_in_mprj[127]
  PIN la_data_in_mprj[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 -2.000 232.210 4.000 ;
    END
  END la_data_in_mprj[12]
  PIN la_data_in_mprj[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 -2.000 243.250 4.000 ;
    END
  END la_data_in_mprj[13]
  PIN la_data_in_mprj[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 -2.000 254.290 4.000 ;
    END
  END la_data_in_mprj[14]
  PIN la_data_in_mprj[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 -2.000 265.330 4.000 ;
    END
  END la_data_in_mprj[15]
  PIN la_data_in_mprj[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 -2.000 276.370 4.000 ;
    END
  END la_data_in_mprj[16]
  PIN la_data_in_mprj[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 -2.000 287.410 4.000 ;
    END
  END la_data_in_mprj[17]
  PIN la_data_in_mprj[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 -2.000 298.450 4.000 ;
    END
  END la_data_in_mprj[18]
  PIN la_data_in_mprj[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 -2.000 309.490 4.000 ;
    END
  END la_data_in_mprj[19]
  PIN la_data_in_mprj[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 -2.000 110.770 4.000 ;
    END
  END la_data_in_mprj[1]
  PIN la_data_in_mprj[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 -2.000 320.530 4.000 ;
    END
  END la_data_in_mprj[20]
  PIN la_data_in_mprj[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 -2.000 331.570 4.000 ;
    END
  END la_data_in_mprj[21]
  PIN la_data_in_mprj[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 -2.000 342.610 4.000 ;
    END
  END la_data_in_mprj[22]
  PIN la_data_in_mprj[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.370 -2.000 353.650 4.000 ;
    END
  END la_data_in_mprj[23]
  PIN la_data_in_mprj[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 -2.000 364.690 4.000 ;
    END
  END la_data_in_mprj[24]
  PIN la_data_in_mprj[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 -2.000 375.730 4.000 ;
    END
  END la_data_in_mprj[25]
  PIN la_data_in_mprj[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 -2.000 386.770 4.000 ;
    END
  END la_data_in_mprj[26]
  PIN la_data_in_mprj[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 -2.000 397.810 4.000 ;
    END
  END la_data_in_mprj[27]
  PIN la_data_in_mprj[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 -2.000 408.850 4.000 ;
    END
  END la_data_in_mprj[28]
  PIN la_data_in_mprj[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.610 -2.000 419.890 4.000 ;
    END
  END la_data_in_mprj[29]
  PIN la_data_in_mprj[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 -2.000 121.810 4.000 ;
    END
  END la_data_in_mprj[2]
  PIN la_data_in_mprj[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 -2.000 430.930 4.000 ;
    END
  END la_data_in_mprj[30]
  PIN la_data_in_mprj[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 -2.000 441.970 4.000 ;
    END
  END la_data_in_mprj[31]
  PIN la_data_in_mprj[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.730 -2.000 453.010 4.000 ;
    END
  END la_data_in_mprj[32]
  PIN la_data_in_mprj[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 -2.000 464.050 4.000 ;
    END
  END la_data_in_mprj[33]
  PIN la_data_in_mprj[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.810 -2.000 475.090 4.000 ;
    END
  END la_data_in_mprj[34]
  PIN la_data_in_mprj[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 -2.000 486.130 4.000 ;
    END
  END la_data_in_mprj[35]
  PIN la_data_in_mprj[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 -2.000 497.170 4.000 ;
    END
  END la_data_in_mprj[36]
  PIN la_data_in_mprj[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.930 -2.000 508.210 4.000 ;
    END
  END la_data_in_mprj[37]
  PIN la_data_in_mprj[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.970 -2.000 519.250 4.000 ;
    END
  END la_data_in_mprj[38]
  PIN la_data_in_mprj[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 -2.000 530.290 4.000 ;
    END
  END la_data_in_mprj[39]
  PIN la_data_in_mprj[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 -2.000 132.850 4.000 ;
    END
  END la_data_in_mprj[3]
  PIN la_data_in_mprj[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 -2.000 541.330 4.000 ;
    END
  END la_data_in_mprj[40]
  PIN la_data_in_mprj[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 -2.000 552.370 4.000 ;
    END
  END la_data_in_mprj[41]
  PIN la_data_in_mprj[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.130 -2.000 563.410 4.000 ;
    END
  END la_data_in_mprj[42]
  PIN la_data_in_mprj[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.170 -2.000 574.450 4.000 ;
    END
  END la_data_in_mprj[43]
  PIN la_data_in_mprj[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 -2.000 585.490 4.000 ;
    END
  END la_data_in_mprj[44]
  PIN la_data_in_mprj[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 -2.000 596.530 4.000 ;
    END
  END la_data_in_mprj[45]
  PIN la_data_in_mprj[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.290 -2.000 607.570 4.000 ;
    END
  END la_data_in_mprj[46]
  PIN la_data_in_mprj[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 -2.000 618.610 4.000 ;
    END
  END la_data_in_mprj[47]
  PIN la_data_in_mprj[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.370 -2.000 629.650 4.000 ;
    END
  END la_data_in_mprj[48]
  PIN la_data_in_mprj[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.410 -2.000 640.690 4.000 ;
    END
  END la_data_in_mprj[49]
  PIN la_data_in_mprj[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 -2.000 143.890 4.000 ;
    END
  END la_data_in_mprj[4]
  PIN la_data_in_mprj[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.450 -2.000 651.730 4.000 ;
    END
  END la_data_in_mprj[50]
  PIN la_data_in_mprj[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.490 -2.000 662.770 4.000 ;
    END
  END la_data_in_mprj[51]
  PIN la_data_in_mprj[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 -2.000 673.810 4.000 ;
    END
  END la_data_in_mprj[52]
  PIN la_data_in_mprj[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.570 -2.000 684.850 4.000 ;
    END
  END la_data_in_mprj[53]
  PIN la_data_in_mprj[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 -2.000 695.890 4.000 ;
    END
  END la_data_in_mprj[54]
  PIN la_data_in_mprj[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.650 -2.000 706.930 4.000 ;
    END
  END la_data_in_mprj[55]
  PIN la_data_in_mprj[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.690 -2.000 717.970 4.000 ;
    END
  END la_data_in_mprj[56]
  PIN la_data_in_mprj[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.730 -2.000 729.010 4.000 ;
    END
  END la_data_in_mprj[57]
  PIN la_data_in_mprj[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.770 -2.000 740.050 4.000 ;
    END
  END la_data_in_mprj[58]
  PIN la_data_in_mprj[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.810 -2.000 751.090 4.000 ;
    END
  END la_data_in_mprj[59]
  PIN la_data_in_mprj[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 -2.000 154.930 4.000 ;
    END
  END la_data_in_mprj[5]
  PIN la_data_in_mprj[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.850 -2.000 762.130 4.000 ;
    END
  END la_data_in_mprj[60]
  PIN la_data_in_mprj[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 -2.000 773.170 4.000 ;
    END
  END la_data_in_mprj[61]
  PIN la_data_in_mprj[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.930 -2.000 784.210 4.000 ;
    END
  END la_data_in_mprj[62]
  PIN la_data_in_mprj[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.970 -2.000 795.250 4.000 ;
    END
  END la_data_in_mprj[63]
  PIN la_data_in_mprj[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.010 -2.000 806.290 4.000 ;
    END
  END la_data_in_mprj[64]
  PIN la_data_in_mprj[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.050 -2.000 817.330 4.000 ;
    END
  END la_data_in_mprj[65]
  PIN la_data_in_mprj[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.090 -2.000 828.370 4.000 ;
    END
  END la_data_in_mprj[66]
  PIN la_data_in_mprj[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.130 -2.000 839.410 4.000 ;
    END
  END la_data_in_mprj[67]
  PIN la_data_in_mprj[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.170 -2.000 850.450 4.000 ;
    END
  END la_data_in_mprj[68]
  PIN la_data_in_mprj[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.210 -2.000 861.490 4.000 ;
    END
  END la_data_in_mprj[69]
  PIN la_data_in_mprj[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 -2.000 165.970 4.000 ;
    END
  END la_data_in_mprj[6]
  PIN la_data_in_mprj[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.250 -2.000 872.530 4.000 ;
    END
  END la_data_in_mprj[70]
  PIN la_data_in_mprj[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.290 -2.000 883.570 4.000 ;
    END
  END la_data_in_mprj[71]
  PIN la_data_in_mprj[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.330 -2.000 894.610 4.000 ;
    END
  END la_data_in_mprj[72]
  PIN la_data_in_mprj[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.370 -2.000 905.650 4.000 ;
    END
  END la_data_in_mprj[73]
  PIN la_data_in_mprj[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.410 -2.000 916.690 4.000 ;
    END
  END la_data_in_mprj[74]
  PIN la_data_in_mprj[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 -2.000 927.730 4.000 ;
    END
  END la_data_in_mprj[75]
  PIN la_data_in_mprj[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.490 -2.000 938.770 4.000 ;
    END
  END la_data_in_mprj[76]
  PIN la_data_in_mprj[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.530 -2.000 949.810 4.000 ;
    END
  END la_data_in_mprj[77]
  PIN la_data_in_mprj[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.570 -2.000 960.850 4.000 ;
    END
  END la_data_in_mprj[78]
  PIN la_data_in_mprj[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.610 -2.000 971.890 4.000 ;
    END
  END la_data_in_mprj[79]
  PIN la_data_in_mprj[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 -2.000 177.010 4.000 ;
    END
  END la_data_in_mprj[7]
  PIN la_data_in_mprj[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.650 -2.000 982.930 4.000 ;
    END
  END la_data_in_mprj[80]
  PIN la_data_in_mprj[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.690 -2.000 993.970 4.000 ;
    END
  END la_data_in_mprj[81]
  PIN la_data_in_mprj[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.730 -2.000 1005.010 4.000 ;
    END
  END la_data_in_mprj[82]
  PIN la_data_in_mprj[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.770 -2.000 1016.050 4.000 ;
    END
  END la_data_in_mprj[83]
  PIN la_data_in_mprj[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.810 -2.000 1027.090 4.000 ;
    END
  END la_data_in_mprj[84]
  PIN la_data_in_mprj[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.850 -2.000 1038.130 4.000 ;
    END
  END la_data_in_mprj[85]
  PIN la_data_in_mprj[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.890 -2.000 1049.170 4.000 ;
    END
  END la_data_in_mprj[86]
  PIN la_data_in_mprj[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.930 -2.000 1060.210 4.000 ;
    END
  END la_data_in_mprj[87]
  PIN la_data_in_mprj[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.970 -2.000 1071.250 4.000 ;
    END
  END la_data_in_mprj[88]
  PIN la_data_in_mprj[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.010 -2.000 1082.290 4.000 ;
    END
  END la_data_in_mprj[89]
  PIN la_data_in_mprj[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 -2.000 188.050 4.000 ;
    END
  END la_data_in_mprj[8]
  PIN la_data_in_mprj[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.050 -2.000 1093.330 4.000 ;
    END
  END la_data_in_mprj[90]
  PIN la_data_in_mprj[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.090 -2.000 1104.370 4.000 ;
    END
  END la_data_in_mprj[91]
  PIN la_data_in_mprj[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1115.130 -2.000 1115.410 4.000 ;
    END
  END la_data_in_mprj[92]
  PIN la_data_in_mprj[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1126.170 -2.000 1126.450 4.000 ;
    END
  END la_data_in_mprj[93]
  PIN la_data_in_mprj[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.210 -2.000 1137.490 4.000 ;
    END
  END la_data_in_mprj[94]
  PIN la_data_in_mprj[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1148.250 -2.000 1148.530 4.000 ;
    END
  END la_data_in_mprj[95]
  PIN la_data_in_mprj[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.290 -2.000 1159.570 4.000 ;
    END
  END la_data_in_mprj[96]
  PIN la_data_in_mprj[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1170.330 -2.000 1170.610 4.000 ;
    END
  END la_data_in_mprj[97]
  PIN la_data_in_mprj[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.370 -2.000 1181.650 4.000 ;
    END
  END la_data_in_mprj[98]
  PIN la_data_in_mprj[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1192.410 -2.000 1192.690 4.000 ;
    END
  END la_data_in_mprj[99]
  PIN la_data_in_mprj[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 -2.000 199.090 4.000 ;
    END
  END la_data_in_mprj[9]
  PIN la_data_out_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 156.000 436.450 162.000 ;
    END
  END la_data_out_core[0]
  PIN la_data_out_core[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1540.170 156.000 1540.450 162.000 ;
    END
  END la_data_out_core[100]
  PIN la_data_out_core[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.210 156.000 1551.490 162.000 ;
    END
  END la_data_out_core[101]
  PIN la_data_out_core[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1562.250 156.000 1562.530 162.000 ;
    END
  END la_data_out_core[102]
  PIN la_data_out_core[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1573.290 156.000 1573.570 162.000 ;
    END
  END la_data_out_core[103]
  PIN la_data_out_core[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.330 156.000 1584.610 162.000 ;
    END
  END la_data_out_core[104]
  PIN la_data_out_core[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1595.370 156.000 1595.650 162.000 ;
    END
  END la_data_out_core[105]
  PIN la_data_out_core[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1606.410 156.000 1606.690 162.000 ;
    END
  END la_data_out_core[106]
  PIN la_data_out_core[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1617.450 156.000 1617.730 162.000 ;
    END
  END la_data_out_core[107]
  PIN la_data_out_core[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1628.490 156.000 1628.770 162.000 ;
    END
  END la_data_out_core[108]
  PIN la_data_out_core[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.530 156.000 1639.810 162.000 ;
    END
  END la_data_out_core[109]
  PIN la_data_out_core[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.570 156.000 546.850 162.000 ;
    END
  END la_data_out_core[10]
  PIN la_data_out_core[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1650.570 156.000 1650.850 162.000 ;
    END
  END la_data_out_core[110]
  PIN la_data_out_core[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.610 156.000 1661.890 162.000 ;
    END
  END la_data_out_core[111]
  PIN la_data_out_core[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1672.650 156.000 1672.930 162.000 ;
    END
  END la_data_out_core[112]
  PIN la_data_out_core[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1683.690 156.000 1683.970 162.000 ;
    END
  END la_data_out_core[113]
  PIN la_data_out_core[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1694.730 156.000 1695.010 162.000 ;
    END
  END la_data_out_core[114]
  PIN la_data_out_core[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1705.770 156.000 1706.050 162.000 ;
    END
  END la_data_out_core[115]
  PIN la_data_out_core[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.810 156.000 1717.090 162.000 ;
    END
  END la_data_out_core[116]
  PIN la_data_out_core[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1727.850 156.000 1728.130 162.000 ;
    END
  END la_data_out_core[117]
  PIN la_data_out_core[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1738.890 156.000 1739.170 162.000 ;
    END
  END la_data_out_core[118]
  PIN la_data_out_core[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1749.930 156.000 1750.210 162.000 ;
    END
  END la_data_out_core[119]
  PIN la_data_out_core[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.610 156.000 557.890 162.000 ;
    END
  END la_data_out_core[11]
  PIN la_data_out_core[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.970 156.000 1761.250 162.000 ;
    END
  END la_data_out_core[120]
  PIN la_data_out_core[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1772.010 156.000 1772.290 162.000 ;
    END
  END la_data_out_core[121]
  PIN la_data_out_core[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.050 156.000 1783.330 162.000 ;
    END
  END la_data_out_core[122]
  PIN la_data_out_core[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1794.090 156.000 1794.370 162.000 ;
    END
  END la_data_out_core[123]
  PIN la_data_out_core[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.130 156.000 1805.410 162.000 ;
    END
  END la_data_out_core[124]
  PIN la_data_out_core[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.170 156.000 1816.450 162.000 ;
    END
  END la_data_out_core[125]
  PIN la_data_out_core[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1827.210 156.000 1827.490 162.000 ;
    END
  END la_data_out_core[126]
  PIN la_data_out_core[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1838.250 156.000 1838.530 162.000 ;
    END
  END la_data_out_core[127]
  PIN la_data_out_core[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.650 156.000 568.930 162.000 ;
    END
  END la_data_out_core[12]
  PIN la_data_out_core[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 156.000 579.970 162.000 ;
    END
  END la_data_out_core[13]
  PIN la_data_out_core[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 156.000 591.010 162.000 ;
    END
  END la_data_out_core[14]
  PIN la_data_out_core[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.770 156.000 602.050 162.000 ;
    END
  END la_data_out_core[15]
  PIN la_data_out_core[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 156.000 613.090 162.000 ;
    END
  END la_data_out_core[16]
  PIN la_data_out_core[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 156.000 624.130 162.000 ;
    END
  END la_data_out_core[17]
  PIN la_data_out_core[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 156.000 635.170 162.000 ;
    END
  END la_data_out_core[18]
  PIN la_data_out_core[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.930 156.000 646.210 162.000 ;
    END
  END la_data_out_core[19]
  PIN la_data_out_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 156.000 447.490 162.000 ;
    END
  END la_data_out_core[1]
  PIN la_data_out_core[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 156.000 657.250 162.000 ;
    END
  END la_data_out_core[20]
  PIN la_data_out_core[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.010 156.000 668.290 162.000 ;
    END
  END la_data_out_core[21]
  PIN la_data_out_core[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.050 156.000 679.330 162.000 ;
    END
  END la_data_out_core[22]
  PIN la_data_out_core[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 156.000 690.370 162.000 ;
    END
  END la_data_out_core[23]
  PIN la_data_out_core[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.130 156.000 701.410 162.000 ;
    END
  END la_data_out_core[24]
  PIN la_data_out_core[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 156.000 712.450 162.000 ;
    END
  END la_data_out_core[25]
  PIN la_data_out_core[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.210 156.000 723.490 162.000 ;
    END
  END la_data_out_core[26]
  PIN la_data_out_core[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 156.000 734.530 162.000 ;
    END
  END la_data_out_core[27]
  PIN la_data_out_core[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 156.000 745.570 162.000 ;
    END
  END la_data_out_core[28]
  PIN la_data_out_core[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.330 156.000 756.610 162.000 ;
    END
  END la_data_out_core[29]
  PIN la_data_out_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 156.000 458.530 162.000 ;
    END
  END la_data_out_core[2]
  PIN la_data_out_core[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 156.000 767.650 162.000 ;
    END
  END la_data_out_core[30]
  PIN la_data_out_core[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.410 156.000 778.690 162.000 ;
    END
  END la_data_out_core[31]
  PIN la_data_out_core[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 156.000 789.730 162.000 ;
    END
  END la_data_out_core[32]
  PIN la_data_out_core[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.490 156.000 800.770 162.000 ;
    END
  END la_data_out_core[33]
  PIN la_data_out_core[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 156.000 811.810 162.000 ;
    END
  END la_data_out_core[34]
  PIN la_data_out_core[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.570 156.000 822.850 162.000 ;
    END
  END la_data_out_core[35]
  PIN la_data_out_core[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.610 156.000 833.890 162.000 ;
    END
  END la_data_out_core[36]
  PIN la_data_out_core[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.650 156.000 844.930 162.000 ;
    END
  END la_data_out_core[37]
  PIN la_data_out_core[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 156.000 855.970 162.000 ;
    END
  END la_data_out_core[38]
  PIN la_data_out_core[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.730 156.000 867.010 162.000 ;
    END
  END la_data_out_core[39]
  PIN la_data_out_core[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 156.000 469.570 162.000 ;
    END
  END la_data_out_core[3]
  PIN la_data_out_core[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.770 156.000 878.050 162.000 ;
    END
  END la_data_out_core[40]
  PIN la_data_out_core[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 156.000 889.090 162.000 ;
    END
  END la_data_out_core[41]
  PIN la_data_out_core[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.850 156.000 900.130 162.000 ;
    END
  END la_data_out_core[42]
  PIN la_data_out_core[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.890 156.000 911.170 162.000 ;
    END
  END la_data_out_core[43]
  PIN la_data_out_core[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.930 156.000 922.210 162.000 ;
    END
  END la_data_out_core[44]
  PIN la_data_out_core[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.970 156.000 933.250 162.000 ;
    END
  END la_data_out_core[45]
  PIN la_data_out_core[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.010 156.000 944.290 162.000 ;
    END
  END la_data_out_core[46]
  PIN la_data_out_core[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.050 156.000 955.330 162.000 ;
    END
  END la_data_out_core[47]
  PIN la_data_out_core[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 156.000 966.370 162.000 ;
    END
  END la_data_out_core[48]
  PIN la_data_out_core[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.130 156.000 977.410 162.000 ;
    END
  END la_data_out_core[49]
  PIN la_data_out_core[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 156.000 480.610 162.000 ;
    END
  END la_data_out_core[4]
  PIN la_data_out_core[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.170 156.000 988.450 162.000 ;
    END
  END la_data_out_core[50]
  PIN la_data_out_core[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.210 156.000 999.490 162.000 ;
    END
  END la_data_out_core[51]
  PIN la_data_out_core[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1010.250 156.000 1010.530 162.000 ;
    END
  END la_data_out_core[52]
  PIN la_data_out_core[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1021.290 156.000 1021.570 162.000 ;
    END
  END la_data_out_core[53]
  PIN la_data_out_core[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1032.330 156.000 1032.610 162.000 ;
    END
  END la_data_out_core[54]
  PIN la_data_out_core[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.370 156.000 1043.650 162.000 ;
    END
  END la_data_out_core[55]
  PIN la_data_out_core[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.410 156.000 1054.690 162.000 ;
    END
  END la_data_out_core[56]
  PIN la_data_out_core[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.450 156.000 1065.730 162.000 ;
    END
  END la_data_out_core[57]
  PIN la_data_out_core[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.490 156.000 1076.770 162.000 ;
    END
  END la_data_out_core[58]
  PIN la_data_out_core[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.530 156.000 1087.810 162.000 ;
    END
  END la_data_out_core[59]
  PIN la_data_out_core[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 156.000 491.650 162.000 ;
    END
  END la_data_out_core[5]
  PIN la_data_out_core[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.570 156.000 1098.850 162.000 ;
    END
  END la_data_out_core[60]
  PIN la_data_out_core[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.610 156.000 1109.890 162.000 ;
    END
  END la_data_out_core[61]
  PIN la_data_out_core[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.650 156.000 1120.930 162.000 ;
    END
  END la_data_out_core[62]
  PIN la_data_out_core[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.690 156.000 1131.970 162.000 ;
    END
  END la_data_out_core[63]
  PIN la_data_out_core[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1142.730 156.000 1143.010 162.000 ;
    END
  END la_data_out_core[64]
  PIN la_data_out_core[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1153.770 156.000 1154.050 162.000 ;
    END
  END la_data_out_core[65]
  PIN la_data_out_core[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.810 156.000 1165.090 162.000 ;
    END
  END la_data_out_core[66]
  PIN la_data_out_core[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.850 156.000 1176.130 162.000 ;
    END
  END la_data_out_core[67]
  PIN la_data_out_core[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1186.890 156.000 1187.170 162.000 ;
    END
  END la_data_out_core[68]
  PIN la_data_out_core[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.930 156.000 1198.210 162.000 ;
    END
  END la_data_out_core[69]
  PIN la_data_out_core[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 156.000 502.690 162.000 ;
    END
  END la_data_out_core[6]
  PIN la_data_out_core[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.970 156.000 1209.250 162.000 ;
    END
  END la_data_out_core[70]
  PIN la_data_out_core[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.010 156.000 1220.290 162.000 ;
    END
  END la_data_out_core[71]
  PIN la_data_out_core[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.050 156.000 1231.330 162.000 ;
    END
  END la_data_out_core[72]
  PIN la_data_out_core[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.090 156.000 1242.370 162.000 ;
    END
  END la_data_out_core[73]
  PIN la_data_out_core[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1253.130 156.000 1253.410 162.000 ;
    END
  END la_data_out_core[74]
  PIN la_data_out_core[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1264.170 156.000 1264.450 162.000 ;
    END
  END la_data_out_core[75]
  PIN la_data_out_core[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.210 156.000 1275.490 162.000 ;
    END
  END la_data_out_core[76]
  PIN la_data_out_core[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1286.250 156.000 1286.530 162.000 ;
    END
  END la_data_out_core[77]
  PIN la_data_out_core[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.290 156.000 1297.570 162.000 ;
    END
  END la_data_out_core[78]
  PIN la_data_out_core[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.330 156.000 1308.610 162.000 ;
    END
  END la_data_out_core[79]
  PIN la_data_out_core[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.450 156.000 513.730 162.000 ;
    END
  END la_data_out_core[7]
  PIN la_data_out_core[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1319.370 156.000 1319.650 162.000 ;
    END
  END la_data_out_core[80]
  PIN la_data_out_core[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1330.410 156.000 1330.690 162.000 ;
    END
  END la_data_out_core[81]
  PIN la_data_out_core[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1341.450 156.000 1341.730 162.000 ;
    END
  END la_data_out_core[82]
  PIN la_data_out_core[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.490 156.000 1352.770 162.000 ;
    END
  END la_data_out_core[83]
  PIN la_data_out_core[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1363.530 156.000 1363.810 162.000 ;
    END
  END la_data_out_core[84]
  PIN la_data_out_core[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1374.570 156.000 1374.850 162.000 ;
    END
  END la_data_out_core[85]
  PIN la_data_out_core[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.610 156.000 1385.890 162.000 ;
    END
  END la_data_out_core[86]
  PIN la_data_out_core[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1396.650 156.000 1396.930 162.000 ;
    END
  END la_data_out_core[87]
  PIN la_data_out_core[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.690 156.000 1407.970 162.000 ;
    END
  END la_data_out_core[88]
  PIN la_data_out_core[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.730 156.000 1419.010 162.000 ;
    END
  END la_data_out_core[89]
  PIN la_data_out_core[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 156.000 524.770 162.000 ;
    END
  END la_data_out_core[8]
  PIN la_data_out_core[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.770 156.000 1430.050 162.000 ;
    END
  END la_data_out_core[90]
  PIN la_data_out_core[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1440.810 156.000 1441.090 162.000 ;
    END
  END la_data_out_core[91]
  PIN la_data_out_core[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1451.850 156.000 1452.130 162.000 ;
    END
  END la_data_out_core[92]
  PIN la_data_out_core[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.890 156.000 1463.170 162.000 ;
    END
  END la_data_out_core[93]
  PIN la_data_out_core[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.930 156.000 1474.210 162.000 ;
    END
  END la_data_out_core[94]
  PIN la_data_out_core[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.970 156.000 1485.250 162.000 ;
    END
  END la_data_out_core[95]
  PIN la_data_out_core[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1496.010 156.000 1496.290 162.000 ;
    END
  END la_data_out_core[96]
  PIN la_data_out_core[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.050 156.000 1507.330 162.000 ;
    END
  END la_data_out_core[97]
  PIN la_data_out_core[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1518.090 156.000 1518.370 162.000 ;
    END
  END la_data_out_core[98]
  PIN la_data_out_core[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1529.130 156.000 1529.410 162.000 ;
    END
  END la_data_out_core[99]
  PIN la_data_out_core[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 156.000 535.810 162.000 ;
    END
  END la_data_out_core[9]
  PIN la_data_out_mprj[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 -2.000 102.490 4.000 ;
    END
  END la_data_out_mprj[0]
  PIN la_data_out_mprj[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1206.210 -2.000 1206.490 4.000 ;
    END
  END la_data_out_mprj[100]
  PIN la_data_out_mprj[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.250 -2.000 1217.530 4.000 ;
    END
  END la_data_out_mprj[101]
  PIN la_data_out_mprj[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1228.290 -2.000 1228.570 4.000 ;
    END
  END la_data_out_mprj[102]
  PIN la_data_out_mprj[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.330 -2.000 1239.610 4.000 ;
    END
  END la_data_out_mprj[103]
  PIN la_data_out_mprj[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1250.370 -2.000 1250.650 4.000 ;
    END
  END la_data_out_mprj[104]
  PIN la_data_out_mprj[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.410 -2.000 1261.690 4.000 ;
    END
  END la_data_out_mprj[105]
  PIN la_data_out_mprj[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1272.450 -2.000 1272.730 4.000 ;
    END
  END la_data_out_mprj[106]
  PIN la_data_out_mprj[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.490 -2.000 1283.770 4.000 ;
    END
  END la_data_out_mprj[107]
  PIN la_data_out_mprj[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.530 -2.000 1294.810 4.000 ;
    END
  END la_data_out_mprj[108]
  PIN la_data_out_mprj[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1305.570 -2.000 1305.850 4.000 ;
    END
  END la_data_out_mprj[109]
  PIN la_data_out_mprj[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 -2.000 212.890 4.000 ;
    END
  END la_data_out_mprj[10]
  PIN la_data_out_mprj[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1316.610 -2.000 1316.890 4.000 ;
    END
  END la_data_out_mprj[110]
  PIN la_data_out_mprj[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1327.650 -2.000 1327.930 4.000 ;
    END
  END la_data_out_mprj[111]
  PIN la_data_out_mprj[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.690 -2.000 1338.970 4.000 ;
    END
  END la_data_out_mprj[112]
  PIN la_data_out_mprj[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.730 -2.000 1350.010 4.000 ;
    END
  END la_data_out_mprj[113]
  PIN la_data_out_mprj[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1360.770 -2.000 1361.050 4.000 ;
    END
  END la_data_out_mprj[114]
  PIN la_data_out_mprj[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.810 -2.000 1372.090 4.000 ;
    END
  END la_data_out_mprj[115]
  PIN la_data_out_mprj[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1382.850 -2.000 1383.130 4.000 ;
    END
  END la_data_out_mprj[116]
  PIN la_data_out_mprj[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1393.890 -2.000 1394.170 4.000 ;
    END
  END la_data_out_mprj[117]
  PIN la_data_out_mprj[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.930 -2.000 1405.210 4.000 ;
    END
  END la_data_out_mprj[118]
  PIN la_data_out_mprj[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.970 -2.000 1416.250 4.000 ;
    END
  END la_data_out_mprj[119]
  PIN la_data_out_mprj[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 -2.000 223.930 4.000 ;
    END
  END la_data_out_mprj[11]
  PIN la_data_out_mprj[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1427.010 -2.000 1427.290 4.000 ;
    END
  END la_data_out_mprj[120]
  PIN la_data_out_mprj[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.050 -2.000 1438.330 4.000 ;
    END
  END la_data_out_mprj[121]
  PIN la_data_out_mprj[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.090 -2.000 1449.370 4.000 ;
    END
  END la_data_out_mprj[122]
  PIN la_data_out_mprj[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1460.130 -2.000 1460.410 4.000 ;
    END
  END la_data_out_mprj[123]
  PIN la_data_out_mprj[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.170 -2.000 1471.450 4.000 ;
    END
  END la_data_out_mprj[124]
  PIN la_data_out_mprj[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1482.210 -2.000 1482.490 4.000 ;
    END
  END la_data_out_mprj[125]
  PIN la_data_out_mprj[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1493.250 -2.000 1493.530 4.000 ;
    END
  END la_data_out_mprj[126]
  PIN la_data_out_mprj[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1504.290 -2.000 1504.570 4.000 ;
    END
  END la_data_out_mprj[127]
  PIN la_data_out_mprj[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 -2.000 234.970 4.000 ;
    END
  END la_data_out_mprj[12]
  PIN la_data_out_mprj[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 -2.000 246.010 4.000 ;
    END
  END la_data_out_mprj[13]
  PIN la_data_out_mprj[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 -2.000 257.050 4.000 ;
    END
  END la_data_out_mprj[14]
  PIN la_data_out_mprj[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 -2.000 268.090 4.000 ;
    END
  END la_data_out_mprj[15]
  PIN la_data_out_mprj[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 -2.000 279.130 4.000 ;
    END
  END la_data_out_mprj[16]
  PIN la_data_out_mprj[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 -2.000 290.170 4.000 ;
    END
  END la_data_out_mprj[17]
  PIN la_data_out_mprj[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 -2.000 301.210 4.000 ;
    END
  END la_data_out_mprj[18]
  PIN la_data_out_mprj[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 -2.000 312.250 4.000 ;
    END
  END la_data_out_mprj[19]
  PIN la_data_out_mprj[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 -2.000 113.530 4.000 ;
    END
  END la_data_out_mprj[1]
  PIN la_data_out_mprj[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 -2.000 323.290 4.000 ;
    END
  END la_data_out_mprj[20]
  PIN la_data_out_mprj[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 -2.000 334.330 4.000 ;
    END
  END la_data_out_mprj[21]
  PIN la_data_out_mprj[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 -2.000 345.370 4.000 ;
    END
  END la_data_out_mprj[22]
  PIN la_data_out_mprj[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 -2.000 356.410 4.000 ;
    END
  END la_data_out_mprj[23]
  PIN la_data_out_mprj[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 -2.000 367.450 4.000 ;
    END
  END la_data_out_mprj[24]
  PIN la_data_out_mprj[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 -2.000 378.490 4.000 ;
    END
  END la_data_out_mprj[25]
  PIN la_data_out_mprj[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 -2.000 389.530 4.000 ;
    END
  END la_data_out_mprj[26]
  PIN la_data_out_mprj[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 -2.000 400.570 4.000 ;
    END
  END la_data_out_mprj[27]
  PIN la_data_out_mprj[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 -2.000 411.610 4.000 ;
    END
  END la_data_out_mprj[28]
  PIN la_data_out_mprj[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.370 -2.000 422.650 4.000 ;
    END
  END la_data_out_mprj[29]
  PIN la_data_out_mprj[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 -2.000 124.570 4.000 ;
    END
  END la_data_out_mprj[2]
  PIN la_data_out_mprj[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 -2.000 433.690 4.000 ;
    END
  END la_data_out_mprj[30]
  PIN la_data_out_mprj[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 -2.000 444.730 4.000 ;
    END
  END la_data_out_mprj[31]
  PIN la_data_out_mprj[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 -2.000 455.770 4.000 ;
    END
  END la_data_out_mprj[32]
  PIN la_data_out_mprj[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.530 -2.000 466.810 4.000 ;
    END
  END la_data_out_mprj[33]
  PIN la_data_out_mprj[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.570 -2.000 477.850 4.000 ;
    END
  END la_data_out_mprj[34]
  PIN la_data_out_mprj[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 -2.000 488.890 4.000 ;
    END
  END la_data_out_mprj[35]
  PIN la_data_out_mprj[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 -2.000 499.930 4.000 ;
    END
  END la_data_out_mprj[36]
  PIN la_data_out_mprj[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 -2.000 510.970 4.000 ;
    END
  END la_data_out_mprj[37]
  PIN la_data_out_mprj[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 -2.000 522.010 4.000 ;
    END
  END la_data_out_mprj[38]
  PIN la_data_out_mprj[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.770 -2.000 533.050 4.000 ;
    END
  END la_data_out_mprj[39]
  PIN la_data_out_mprj[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 -2.000 135.610 4.000 ;
    END
  END la_data_out_mprj[3]
  PIN la_data_out_mprj[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 -2.000 544.090 4.000 ;
    END
  END la_data_out_mprj[40]
  PIN la_data_out_mprj[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.850 -2.000 555.130 4.000 ;
    END
  END la_data_out_mprj[41]
  PIN la_data_out_mprj[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.890 -2.000 566.170 4.000 ;
    END
  END la_data_out_mprj[42]
  PIN la_data_out_mprj[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.930 -2.000 577.210 4.000 ;
    END
  END la_data_out_mprj[43]
  PIN la_data_out_mprj[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.970 -2.000 588.250 4.000 ;
    END
  END la_data_out_mprj[44]
  PIN la_data_out_mprj[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 -2.000 599.290 4.000 ;
    END
  END la_data_out_mprj[45]
  PIN la_data_out_mprj[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.050 -2.000 610.330 4.000 ;
    END
  END la_data_out_mprj[46]
  PIN la_data_out_mprj[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.090 -2.000 621.370 4.000 ;
    END
  END la_data_out_mprj[47]
  PIN la_data_out_mprj[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 -2.000 632.410 4.000 ;
    END
  END la_data_out_mprj[48]
  PIN la_data_out_mprj[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.170 -2.000 643.450 4.000 ;
    END
  END la_data_out_mprj[49]
  PIN la_data_out_mprj[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 -2.000 146.650 4.000 ;
    END
  END la_data_out_mprj[4]
  PIN la_data_out_mprj[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.210 -2.000 654.490 4.000 ;
    END
  END la_data_out_mprj[50]
  PIN la_data_out_mprj[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.250 -2.000 665.530 4.000 ;
    END
  END la_data_out_mprj[51]
  PIN la_data_out_mprj[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 -2.000 676.570 4.000 ;
    END
  END la_data_out_mprj[52]
  PIN la_data_out_mprj[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.330 -2.000 687.610 4.000 ;
    END
  END la_data_out_mprj[53]
  PIN la_data_out_mprj[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.370 -2.000 698.650 4.000 ;
    END
  END la_data_out_mprj[54]
  PIN la_data_out_mprj[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.410 -2.000 709.690 4.000 ;
    END
  END la_data_out_mprj[55]
  PIN la_data_out_mprj[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.450 -2.000 720.730 4.000 ;
    END
  END la_data_out_mprj[56]
  PIN la_data_out_mprj[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.490 -2.000 731.770 4.000 ;
    END
  END la_data_out_mprj[57]
  PIN la_data_out_mprj[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.530 -2.000 742.810 4.000 ;
    END
  END la_data_out_mprj[58]
  PIN la_data_out_mprj[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 -2.000 753.850 4.000 ;
    END
  END la_data_out_mprj[59]
  PIN la_data_out_mprj[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 -2.000 157.690 4.000 ;
    END
  END la_data_out_mprj[5]
  PIN la_data_out_mprj[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.610 -2.000 764.890 4.000 ;
    END
  END la_data_out_mprj[60]
  PIN la_data_out_mprj[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 -2.000 775.930 4.000 ;
    END
  END la_data_out_mprj[61]
  PIN la_data_out_mprj[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 -2.000 786.970 4.000 ;
    END
  END la_data_out_mprj[62]
  PIN la_data_out_mprj[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 -2.000 798.010 4.000 ;
    END
  END la_data_out_mprj[63]
  PIN la_data_out_mprj[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.770 -2.000 809.050 4.000 ;
    END
  END la_data_out_mprj[64]
  PIN la_data_out_mprj[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.810 -2.000 820.090 4.000 ;
    END
  END la_data_out_mprj[65]
  PIN la_data_out_mprj[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 -2.000 831.130 4.000 ;
    END
  END la_data_out_mprj[66]
  PIN la_data_out_mprj[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.890 -2.000 842.170 4.000 ;
    END
  END la_data_out_mprj[67]
  PIN la_data_out_mprj[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.930 -2.000 853.210 4.000 ;
    END
  END la_data_out_mprj[68]
  PIN la_data_out_mprj[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.970 -2.000 864.250 4.000 ;
    END
  END la_data_out_mprj[69]
  PIN la_data_out_mprj[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 -2.000 168.730 4.000 ;
    END
  END la_data_out_mprj[6]
  PIN la_data_out_mprj[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.010 -2.000 875.290 4.000 ;
    END
  END la_data_out_mprj[70]
  PIN la_data_out_mprj[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.050 -2.000 886.330 4.000 ;
    END
  END la_data_out_mprj[71]
  PIN la_data_out_mprj[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.090 -2.000 897.370 4.000 ;
    END
  END la_data_out_mprj[72]
  PIN la_data_out_mprj[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.130 -2.000 908.410 4.000 ;
    END
  END la_data_out_mprj[73]
  PIN la_data_out_mprj[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.170 -2.000 919.450 4.000 ;
    END
  END la_data_out_mprj[74]
  PIN la_data_out_mprj[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.210 -2.000 930.490 4.000 ;
    END
  END la_data_out_mprj[75]
  PIN la_data_out_mprj[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.250 -2.000 941.530 4.000 ;
    END
  END la_data_out_mprj[76]
  PIN la_data_out_mprj[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.290 -2.000 952.570 4.000 ;
    END
  END la_data_out_mprj[77]
  PIN la_data_out_mprj[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.330 -2.000 963.610 4.000 ;
    END
  END la_data_out_mprj[78]
  PIN la_data_out_mprj[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.370 -2.000 974.650 4.000 ;
    END
  END la_data_out_mprj[79]
  PIN la_data_out_mprj[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 -2.000 179.770 4.000 ;
    END
  END la_data_out_mprj[7]
  PIN la_data_out_mprj[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 -2.000 985.690 4.000 ;
    END
  END la_data_out_mprj[80]
  PIN la_data_out_mprj[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.450 -2.000 996.730 4.000 ;
    END
  END la_data_out_mprj[81]
  PIN la_data_out_mprj[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.490 -2.000 1007.770 4.000 ;
    END
  END la_data_out_mprj[82]
  PIN la_data_out_mprj[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.530 -2.000 1018.810 4.000 ;
    END
  END la_data_out_mprj[83]
  PIN la_data_out_mprj[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.570 -2.000 1029.850 4.000 ;
    END
  END la_data_out_mprj[84]
  PIN la_data_out_mprj[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.610 -2.000 1040.890 4.000 ;
    END
  END la_data_out_mprj[85]
  PIN la_data_out_mprj[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.650 -2.000 1051.930 4.000 ;
    END
  END la_data_out_mprj[86]
  PIN la_data_out_mprj[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 -2.000 1062.970 4.000 ;
    END
  END la_data_out_mprj[87]
  PIN la_data_out_mprj[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.730 -2.000 1074.010 4.000 ;
    END
  END la_data_out_mprj[88]
  PIN la_data_out_mprj[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.770 -2.000 1085.050 4.000 ;
    END
  END la_data_out_mprj[89]
  PIN la_data_out_mprj[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 -2.000 190.810 4.000 ;
    END
  END la_data_out_mprj[8]
  PIN la_data_out_mprj[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.810 -2.000 1096.090 4.000 ;
    END
  END la_data_out_mprj[90]
  PIN la_data_out_mprj[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1106.850 -2.000 1107.130 4.000 ;
    END
  END la_data_out_mprj[91]
  PIN la_data_out_mprj[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.890 -2.000 1118.170 4.000 ;
    END
  END la_data_out_mprj[92]
  PIN la_data_out_mprj[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.930 -2.000 1129.210 4.000 ;
    END
  END la_data_out_mprj[93]
  PIN la_data_out_mprj[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.970 -2.000 1140.250 4.000 ;
    END
  END la_data_out_mprj[94]
  PIN la_data_out_mprj[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1151.010 -2.000 1151.290 4.000 ;
    END
  END la_data_out_mprj[95]
  PIN la_data_out_mprj[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.050 -2.000 1162.330 4.000 ;
    END
  END la_data_out_mprj[96]
  PIN la_data_out_mprj[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.090 -2.000 1173.370 4.000 ;
    END
  END la_data_out_mprj[97]
  PIN la_data_out_mprj[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.130 -2.000 1184.410 4.000 ;
    END
  END la_data_out_mprj[98]
  PIN la_data_out_mprj[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1195.170 -2.000 1195.450 4.000 ;
    END
  END la_data_out_mprj[99]
  PIN la_data_out_mprj[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 -2.000 201.850 4.000 ;
    END
  END la_data_out_mprj[9]
  PIN la_iena_mprj[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 -2.000 105.250 4.000 ;
    END
  END la_iena_mprj[0]
  PIN la_iena_mprj[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.970 -2.000 1209.250 4.000 ;
    END
  END la_iena_mprj[100]
  PIN la_iena_mprj[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.010 -2.000 1220.290 4.000 ;
    END
  END la_iena_mprj[101]
  PIN la_iena_mprj[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.050 -2.000 1231.330 4.000 ;
    END
  END la_iena_mprj[102]
  PIN la_iena_mprj[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.090 -2.000 1242.370 4.000 ;
    END
  END la_iena_mprj[103]
  PIN la_iena_mprj[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1253.130 -2.000 1253.410 4.000 ;
    END
  END la_iena_mprj[104]
  PIN la_iena_mprj[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1264.170 -2.000 1264.450 4.000 ;
    END
  END la_iena_mprj[105]
  PIN la_iena_mprj[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.210 -2.000 1275.490 4.000 ;
    END
  END la_iena_mprj[106]
  PIN la_iena_mprj[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1286.250 -2.000 1286.530 4.000 ;
    END
  END la_iena_mprj[107]
  PIN la_iena_mprj[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.290 -2.000 1297.570 4.000 ;
    END
  END la_iena_mprj[108]
  PIN la_iena_mprj[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.330 -2.000 1308.610 4.000 ;
    END
  END la_iena_mprj[109]
  PIN la_iena_mprj[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 -2.000 215.650 4.000 ;
    END
  END la_iena_mprj[10]
  PIN la_iena_mprj[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1319.370 -2.000 1319.650 4.000 ;
    END
  END la_iena_mprj[110]
  PIN la_iena_mprj[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1330.410 -2.000 1330.690 4.000 ;
    END
  END la_iena_mprj[111]
  PIN la_iena_mprj[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1341.450 -2.000 1341.730 4.000 ;
    END
  END la_iena_mprj[112]
  PIN la_iena_mprj[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.490 -2.000 1352.770 4.000 ;
    END
  END la_iena_mprj[113]
  PIN la_iena_mprj[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1363.530 -2.000 1363.810 4.000 ;
    END
  END la_iena_mprj[114]
  PIN la_iena_mprj[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1374.570 -2.000 1374.850 4.000 ;
    END
  END la_iena_mprj[115]
  PIN la_iena_mprj[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.610 -2.000 1385.890 4.000 ;
    END
  END la_iena_mprj[116]
  PIN la_iena_mprj[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1396.650 -2.000 1396.930 4.000 ;
    END
  END la_iena_mprj[117]
  PIN la_iena_mprj[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.690 -2.000 1407.970 4.000 ;
    END
  END la_iena_mprj[118]
  PIN la_iena_mprj[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.730 -2.000 1419.010 4.000 ;
    END
  END la_iena_mprj[119]
  PIN la_iena_mprj[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 -2.000 226.690 4.000 ;
    END
  END la_iena_mprj[11]
  PIN la_iena_mprj[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.770 -2.000 1430.050 4.000 ;
    END
  END la_iena_mprj[120]
  PIN la_iena_mprj[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1440.810 -2.000 1441.090 4.000 ;
    END
  END la_iena_mprj[121]
  PIN la_iena_mprj[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1451.850 -2.000 1452.130 4.000 ;
    END
  END la_iena_mprj[122]
  PIN la_iena_mprj[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.890 -2.000 1463.170 4.000 ;
    END
  END la_iena_mprj[123]
  PIN la_iena_mprj[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.930 -2.000 1474.210 4.000 ;
    END
  END la_iena_mprj[124]
  PIN la_iena_mprj[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.970 -2.000 1485.250 4.000 ;
    END
  END la_iena_mprj[125]
  PIN la_iena_mprj[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1496.010 -2.000 1496.290 4.000 ;
    END
  END la_iena_mprj[126]
  PIN la_iena_mprj[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.050 -2.000 1507.330 4.000 ;
    END
  END la_iena_mprj[127]
  PIN la_iena_mprj[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 -2.000 237.730 4.000 ;
    END
  END la_iena_mprj[12]
  PIN la_iena_mprj[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 -2.000 248.770 4.000 ;
    END
  END la_iena_mprj[13]
  PIN la_iena_mprj[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 -2.000 259.810 4.000 ;
    END
  END la_iena_mprj[14]
  PIN la_iena_mprj[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 -2.000 270.850 4.000 ;
    END
  END la_iena_mprj[15]
  PIN la_iena_mprj[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 -2.000 281.890 4.000 ;
    END
  END la_iena_mprj[16]
  PIN la_iena_mprj[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 -2.000 292.930 4.000 ;
    END
  END la_iena_mprj[17]
  PIN la_iena_mprj[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 -2.000 303.970 4.000 ;
    END
  END la_iena_mprj[18]
  PIN la_iena_mprj[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 -2.000 315.010 4.000 ;
    END
  END la_iena_mprj[19]
  PIN la_iena_mprj[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 -2.000 116.290 4.000 ;
    END
  END la_iena_mprj[1]
  PIN la_iena_mprj[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 -2.000 326.050 4.000 ;
    END
  END la_iena_mprj[20]
  PIN la_iena_mprj[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 -2.000 337.090 4.000 ;
    END
  END la_iena_mprj[21]
  PIN la_iena_mprj[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 -2.000 348.130 4.000 ;
    END
  END la_iena_mprj[22]
  PIN la_iena_mprj[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 -2.000 359.170 4.000 ;
    END
  END la_iena_mprj[23]
  PIN la_iena_mprj[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 -2.000 370.210 4.000 ;
    END
  END la_iena_mprj[24]
  PIN la_iena_mprj[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 -2.000 381.250 4.000 ;
    END
  END la_iena_mprj[25]
  PIN la_iena_mprj[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 -2.000 392.290 4.000 ;
    END
  END la_iena_mprj[26]
  PIN la_iena_mprj[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 -2.000 403.330 4.000 ;
    END
  END la_iena_mprj[27]
  PIN la_iena_mprj[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 -2.000 414.370 4.000 ;
    END
  END la_iena_mprj[28]
  PIN la_iena_mprj[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 -2.000 425.410 4.000 ;
    END
  END la_iena_mprj[29]
  PIN la_iena_mprj[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 -2.000 127.330 4.000 ;
    END
  END la_iena_mprj[2]
  PIN la_iena_mprj[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 -2.000 436.450 4.000 ;
    END
  END la_iena_mprj[30]
  PIN la_iena_mprj[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 -2.000 447.490 4.000 ;
    END
  END la_iena_mprj[31]
  PIN la_iena_mprj[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 -2.000 458.530 4.000 ;
    END
  END la_iena_mprj[32]
  PIN la_iena_mprj[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 -2.000 469.570 4.000 ;
    END
  END la_iena_mprj[33]
  PIN la_iena_mprj[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 -2.000 480.610 4.000 ;
    END
  END la_iena_mprj[34]
  PIN la_iena_mprj[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 -2.000 491.650 4.000 ;
    END
  END la_iena_mprj[35]
  PIN la_iena_mprj[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 -2.000 502.690 4.000 ;
    END
  END la_iena_mprj[36]
  PIN la_iena_mprj[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.450 -2.000 513.730 4.000 ;
    END
  END la_iena_mprj[37]
  PIN la_iena_mprj[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 -2.000 524.770 4.000 ;
    END
  END la_iena_mprj[38]
  PIN la_iena_mprj[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 -2.000 535.810 4.000 ;
    END
  END la_iena_mprj[39]
  PIN la_iena_mprj[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 -2.000 138.370 4.000 ;
    END
  END la_iena_mprj[3]
  PIN la_iena_mprj[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.570 -2.000 546.850 4.000 ;
    END
  END la_iena_mprj[40]
  PIN la_iena_mprj[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.610 -2.000 557.890 4.000 ;
    END
  END la_iena_mprj[41]
  PIN la_iena_mprj[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.650 -2.000 568.930 4.000 ;
    END
  END la_iena_mprj[42]
  PIN la_iena_mprj[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 -2.000 579.970 4.000 ;
    END
  END la_iena_mprj[43]
  PIN la_iena_mprj[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 -2.000 591.010 4.000 ;
    END
  END la_iena_mprj[44]
  PIN la_iena_mprj[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.770 -2.000 602.050 4.000 ;
    END
  END la_iena_mprj[45]
  PIN la_iena_mprj[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 -2.000 613.090 4.000 ;
    END
  END la_iena_mprj[46]
  PIN la_iena_mprj[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 -2.000 624.130 4.000 ;
    END
  END la_iena_mprj[47]
  PIN la_iena_mprj[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 -2.000 635.170 4.000 ;
    END
  END la_iena_mprj[48]
  PIN la_iena_mprj[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.930 -2.000 646.210 4.000 ;
    END
  END la_iena_mprj[49]
  PIN la_iena_mprj[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 -2.000 149.410 4.000 ;
    END
  END la_iena_mprj[4]
  PIN la_iena_mprj[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 -2.000 657.250 4.000 ;
    END
  END la_iena_mprj[50]
  PIN la_iena_mprj[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.010 -2.000 668.290 4.000 ;
    END
  END la_iena_mprj[51]
  PIN la_iena_mprj[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.050 -2.000 679.330 4.000 ;
    END
  END la_iena_mprj[52]
  PIN la_iena_mprj[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 -2.000 690.370 4.000 ;
    END
  END la_iena_mprj[53]
  PIN la_iena_mprj[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.130 -2.000 701.410 4.000 ;
    END
  END la_iena_mprj[54]
  PIN la_iena_mprj[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 -2.000 712.450 4.000 ;
    END
  END la_iena_mprj[55]
  PIN la_iena_mprj[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.210 -2.000 723.490 4.000 ;
    END
  END la_iena_mprj[56]
  PIN la_iena_mprj[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 -2.000 734.530 4.000 ;
    END
  END la_iena_mprj[57]
  PIN la_iena_mprj[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 -2.000 745.570 4.000 ;
    END
  END la_iena_mprj[58]
  PIN la_iena_mprj[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.330 -2.000 756.610 4.000 ;
    END
  END la_iena_mprj[59]
  PIN la_iena_mprj[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 -2.000 160.450 4.000 ;
    END
  END la_iena_mprj[5]
  PIN la_iena_mprj[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 -2.000 767.650 4.000 ;
    END
  END la_iena_mprj[60]
  PIN la_iena_mprj[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.410 -2.000 778.690 4.000 ;
    END
  END la_iena_mprj[61]
  PIN la_iena_mprj[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 -2.000 789.730 4.000 ;
    END
  END la_iena_mprj[62]
  PIN la_iena_mprj[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.490 -2.000 800.770 4.000 ;
    END
  END la_iena_mprj[63]
  PIN la_iena_mprj[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 -2.000 811.810 4.000 ;
    END
  END la_iena_mprj[64]
  PIN la_iena_mprj[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.570 -2.000 822.850 4.000 ;
    END
  END la_iena_mprj[65]
  PIN la_iena_mprj[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.610 -2.000 833.890 4.000 ;
    END
  END la_iena_mprj[66]
  PIN la_iena_mprj[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.650 -2.000 844.930 4.000 ;
    END
  END la_iena_mprj[67]
  PIN la_iena_mprj[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 -2.000 855.970 4.000 ;
    END
  END la_iena_mprj[68]
  PIN la_iena_mprj[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.730 -2.000 867.010 4.000 ;
    END
  END la_iena_mprj[69]
  PIN la_iena_mprj[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 -2.000 171.490 4.000 ;
    END
  END la_iena_mprj[6]
  PIN la_iena_mprj[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.770 -2.000 878.050 4.000 ;
    END
  END la_iena_mprj[70]
  PIN la_iena_mprj[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 -2.000 889.090 4.000 ;
    END
  END la_iena_mprj[71]
  PIN la_iena_mprj[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.850 -2.000 900.130 4.000 ;
    END
  END la_iena_mprj[72]
  PIN la_iena_mprj[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.890 -2.000 911.170 4.000 ;
    END
  END la_iena_mprj[73]
  PIN la_iena_mprj[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.930 -2.000 922.210 4.000 ;
    END
  END la_iena_mprj[74]
  PIN la_iena_mprj[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.970 -2.000 933.250 4.000 ;
    END
  END la_iena_mprj[75]
  PIN la_iena_mprj[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.010 -2.000 944.290 4.000 ;
    END
  END la_iena_mprj[76]
  PIN la_iena_mprj[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.050 -2.000 955.330 4.000 ;
    END
  END la_iena_mprj[77]
  PIN la_iena_mprj[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 -2.000 966.370 4.000 ;
    END
  END la_iena_mprj[78]
  PIN la_iena_mprj[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.130 -2.000 977.410 4.000 ;
    END
  END la_iena_mprj[79]
  PIN la_iena_mprj[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 -2.000 182.530 4.000 ;
    END
  END la_iena_mprj[7]
  PIN la_iena_mprj[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.170 -2.000 988.450 4.000 ;
    END
  END la_iena_mprj[80]
  PIN la_iena_mprj[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.210 -2.000 999.490 4.000 ;
    END
  END la_iena_mprj[81]
  PIN la_iena_mprj[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1010.250 -2.000 1010.530 4.000 ;
    END
  END la_iena_mprj[82]
  PIN la_iena_mprj[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1021.290 -2.000 1021.570 4.000 ;
    END
  END la_iena_mprj[83]
  PIN la_iena_mprj[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1032.330 -2.000 1032.610 4.000 ;
    END
  END la_iena_mprj[84]
  PIN la_iena_mprj[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.370 -2.000 1043.650 4.000 ;
    END
  END la_iena_mprj[85]
  PIN la_iena_mprj[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.410 -2.000 1054.690 4.000 ;
    END
  END la_iena_mprj[86]
  PIN la_iena_mprj[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.450 -2.000 1065.730 4.000 ;
    END
  END la_iena_mprj[87]
  PIN la_iena_mprj[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.490 -2.000 1076.770 4.000 ;
    END
  END la_iena_mprj[88]
  PIN la_iena_mprj[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.530 -2.000 1087.810 4.000 ;
    END
  END la_iena_mprj[89]
  PIN la_iena_mprj[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 -2.000 193.570 4.000 ;
    END
  END la_iena_mprj[8]
  PIN la_iena_mprj[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.570 -2.000 1098.850 4.000 ;
    END
  END la_iena_mprj[90]
  PIN la_iena_mprj[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.610 -2.000 1109.890 4.000 ;
    END
  END la_iena_mprj[91]
  PIN la_iena_mprj[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.650 -2.000 1120.930 4.000 ;
    END
  END la_iena_mprj[92]
  PIN la_iena_mprj[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.690 -2.000 1131.970 4.000 ;
    END
  END la_iena_mprj[93]
  PIN la_iena_mprj[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1142.730 -2.000 1143.010 4.000 ;
    END
  END la_iena_mprj[94]
  PIN la_iena_mprj[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1153.770 -2.000 1154.050 4.000 ;
    END
  END la_iena_mprj[95]
  PIN la_iena_mprj[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.810 -2.000 1165.090 4.000 ;
    END
  END la_iena_mprj[96]
  PIN la_iena_mprj[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.850 -2.000 1176.130 4.000 ;
    END
  END la_iena_mprj[97]
  PIN la_iena_mprj[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1186.890 -2.000 1187.170 4.000 ;
    END
  END la_iena_mprj[98]
  PIN la_iena_mprj[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.930 -2.000 1198.210 4.000 ;
    END
  END la_iena_mprj[99]
  PIN la_iena_mprj[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 -2.000 204.610 4.000 ;
    END
  END la_iena_mprj[9]
  PIN la_oenb_core[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 156.000 440.130 162.000 ;
    END
  END la_oenb_core[0]
  PIN la_oenb_core[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1543.850 156.000 1544.130 162.000 ;
    END
  END la_oenb_core[100]
  PIN la_oenb_core[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1554.890 156.000 1555.170 162.000 ;
    END
  END la_oenb_core[101]
  PIN la_oenb_core[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.930 156.000 1566.210 162.000 ;
    END
  END la_oenb_core[102]
  PIN la_oenb_core[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1576.970 156.000 1577.250 162.000 ;
    END
  END la_oenb_core[103]
  PIN la_oenb_core[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.010 156.000 1588.290 162.000 ;
    END
  END la_oenb_core[104]
  PIN la_oenb_core[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1599.050 156.000 1599.330 162.000 ;
    END
  END la_oenb_core[105]
  PIN la_oenb_core[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.090 156.000 1610.370 162.000 ;
    END
  END la_oenb_core[106]
  PIN la_oenb_core[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.130 156.000 1621.410 162.000 ;
    END
  END la_oenb_core[107]
  PIN la_oenb_core[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1632.170 156.000 1632.450 162.000 ;
    END
  END la_oenb_core[108]
  PIN la_oenb_core[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1643.210 156.000 1643.490 162.000 ;
    END
  END la_oenb_core[109]
  PIN la_oenb_core[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.250 156.000 550.530 162.000 ;
    END
  END la_oenb_core[10]
  PIN la_oenb_core[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1654.250 156.000 1654.530 162.000 ;
    END
  END la_oenb_core[110]
  PIN la_oenb_core[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1665.290 156.000 1665.570 162.000 ;
    END
  END la_oenb_core[111]
  PIN la_oenb_core[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1676.330 156.000 1676.610 162.000 ;
    END
  END la_oenb_core[112]
  PIN la_oenb_core[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.370 156.000 1687.650 162.000 ;
    END
  END la_oenb_core[113]
  PIN la_oenb_core[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1698.410 156.000 1698.690 162.000 ;
    END
  END la_oenb_core[114]
  PIN la_oenb_core[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.450 156.000 1709.730 162.000 ;
    END
  END la_oenb_core[115]
  PIN la_oenb_core[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1720.490 156.000 1720.770 162.000 ;
    END
  END la_oenb_core[116]
  PIN la_oenb_core[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1731.530 156.000 1731.810 162.000 ;
    END
  END la_oenb_core[117]
  PIN la_oenb_core[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1742.570 156.000 1742.850 162.000 ;
    END
  END la_oenb_core[118]
  PIN la_oenb_core[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1753.610 156.000 1753.890 162.000 ;
    END
  END la_oenb_core[119]
  PIN la_oenb_core[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.290 156.000 561.570 162.000 ;
    END
  END la_oenb_core[11]
  PIN la_oenb_core[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.650 156.000 1764.930 162.000 ;
    END
  END la_oenb_core[120]
  PIN la_oenb_core[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1775.690 156.000 1775.970 162.000 ;
    END
  END la_oenb_core[121]
  PIN la_oenb_core[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1786.730 156.000 1787.010 162.000 ;
    END
  END la_oenb_core[122]
  PIN la_oenb_core[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1797.770 156.000 1798.050 162.000 ;
    END
  END la_oenb_core[123]
  PIN la_oenb_core[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1808.810 156.000 1809.090 162.000 ;
    END
  END la_oenb_core[124]
  PIN la_oenb_core[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1819.850 156.000 1820.130 162.000 ;
    END
  END la_oenb_core[125]
  PIN la_oenb_core[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1830.890 156.000 1831.170 162.000 ;
    END
  END la_oenb_core[126]
  PIN la_oenb_core[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1841.930 156.000 1842.210 162.000 ;
    END
  END la_oenb_core[127]
  PIN la_oenb_core[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.330 156.000 572.610 162.000 ;
    END
  END la_oenb_core[12]
  PIN la_oenb_core[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.370 156.000 583.650 162.000 ;
    END
  END la_oenb_core[13]
  PIN la_oenb_core[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 156.000 594.690 162.000 ;
    END
  END la_oenb_core[14]
  PIN la_oenb_core[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 156.000 605.730 162.000 ;
    END
  END la_oenb_core[15]
  PIN la_oenb_core[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.490 156.000 616.770 162.000 ;
    END
  END la_oenb_core[16]
  PIN la_oenb_core[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 156.000 627.810 162.000 ;
    END
  END la_oenb_core[17]
  PIN la_oenb_core[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 156.000 638.850 162.000 ;
    END
  END la_oenb_core[18]
  PIN la_oenb_core[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 156.000 649.890 162.000 ;
    END
  END la_oenb_core[19]
  PIN la_oenb_core[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 156.000 451.170 162.000 ;
    END
  END la_oenb_core[1]
  PIN la_oenb_core[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 156.000 660.930 162.000 ;
    END
  END la_oenb_core[20]
  PIN la_oenb_core[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.690 156.000 671.970 162.000 ;
    END
  END la_oenb_core[21]
  PIN la_oenb_core[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 156.000 683.010 162.000 ;
    END
  END la_oenb_core[22]
  PIN la_oenb_core[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.770 156.000 694.050 162.000 ;
    END
  END la_oenb_core[23]
  PIN la_oenb_core[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.810 156.000 705.090 162.000 ;
    END
  END la_oenb_core[24]
  PIN la_oenb_core[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 156.000 716.130 162.000 ;
    END
  END la_oenb_core[25]
  PIN la_oenb_core[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.890 156.000 727.170 162.000 ;
    END
  END la_oenb_core[26]
  PIN la_oenb_core[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.930 156.000 738.210 162.000 ;
    END
  END la_oenb_core[27]
  PIN la_oenb_core[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.970 156.000 749.250 162.000 ;
    END
  END la_oenb_core[28]
  PIN la_oenb_core[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 156.000 760.290 162.000 ;
    END
  END la_oenb_core[29]
  PIN la_oenb_core[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.930 156.000 462.210 162.000 ;
    END
  END la_oenb_core[2]
  PIN la_oenb_core[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.050 156.000 771.330 162.000 ;
    END
  END la_oenb_core[30]
  PIN la_oenb_core[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.090 156.000 782.370 162.000 ;
    END
  END la_oenb_core[31]
  PIN la_oenb_core[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.130 156.000 793.410 162.000 ;
    END
  END la_oenb_core[32]
  PIN la_oenb_core[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.170 156.000 804.450 162.000 ;
    END
  END la_oenb_core[33]
  PIN la_oenb_core[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.210 156.000 815.490 162.000 ;
    END
  END la_oenb_core[34]
  PIN la_oenb_core[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.250 156.000 826.530 162.000 ;
    END
  END la_oenb_core[35]
  PIN la_oenb_core[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 156.000 837.570 162.000 ;
    END
  END la_oenb_core[36]
  PIN la_oenb_core[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.330 156.000 848.610 162.000 ;
    END
  END la_oenb_core[37]
  PIN la_oenb_core[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.370 156.000 859.650 162.000 ;
    END
  END la_oenb_core[38]
  PIN la_oenb_core[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.410 156.000 870.690 162.000 ;
    END
  END la_oenb_core[39]
  PIN la_oenb_core[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.970 156.000 473.250 162.000 ;
    END
  END la_oenb_core[3]
  PIN la_oenb_core[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.450 156.000 881.730 162.000 ;
    END
  END la_oenb_core[40]
  PIN la_oenb_core[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.490 156.000 892.770 162.000 ;
    END
  END la_oenb_core[41]
  PIN la_oenb_core[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.530 156.000 903.810 162.000 ;
    END
  END la_oenb_core[42]
  PIN la_oenb_core[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 156.000 914.850 162.000 ;
    END
  END la_oenb_core[43]
  PIN la_oenb_core[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 925.610 156.000 925.890 162.000 ;
    END
  END la_oenb_core[44]
  PIN la_oenb_core[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.650 156.000 936.930 162.000 ;
    END
  END la_oenb_core[45]
  PIN la_oenb_core[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.690 156.000 947.970 162.000 ;
    END
  END la_oenb_core[46]
  PIN la_oenb_core[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.730 156.000 959.010 162.000 ;
    END
  END la_oenb_core[47]
  PIN la_oenb_core[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.770 156.000 970.050 162.000 ;
    END
  END la_oenb_core[48]
  PIN la_oenb_core[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.810 156.000 981.090 162.000 ;
    END
  END la_oenb_core[49]
  PIN la_oenb_core[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.010 156.000 484.290 162.000 ;
    END
  END la_oenb_core[4]
  PIN la_oenb_core[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.850 156.000 992.130 162.000 ;
    END
  END la_oenb_core[50]
  PIN la_oenb_core[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.890 156.000 1003.170 162.000 ;
    END
  END la_oenb_core[51]
  PIN la_oenb_core[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.930 156.000 1014.210 162.000 ;
    END
  END la_oenb_core[52]
  PIN la_oenb_core[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.970 156.000 1025.250 162.000 ;
    END
  END la_oenb_core[53]
  PIN la_oenb_core[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.010 156.000 1036.290 162.000 ;
    END
  END la_oenb_core[54]
  PIN la_oenb_core[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.050 156.000 1047.330 162.000 ;
    END
  END la_oenb_core[55]
  PIN la_oenb_core[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.090 156.000 1058.370 162.000 ;
    END
  END la_oenb_core[56]
  PIN la_oenb_core[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.130 156.000 1069.410 162.000 ;
    END
  END la_oenb_core[57]
  PIN la_oenb_core[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.170 156.000 1080.450 162.000 ;
    END
  END la_oenb_core[58]
  PIN la_oenb_core[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.210 156.000 1091.490 162.000 ;
    END
  END la_oenb_core[59]
  PIN la_oenb_core[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.050 156.000 495.330 162.000 ;
    END
  END la_oenb_core[5]
  PIN la_oenb_core[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.250 156.000 1102.530 162.000 ;
    END
  END la_oenb_core[60]
  PIN la_oenb_core[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.290 156.000 1113.570 162.000 ;
    END
  END la_oenb_core[61]
  PIN la_oenb_core[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.330 156.000 1124.610 162.000 ;
    END
  END la_oenb_core[62]
  PIN la_oenb_core[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1135.370 156.000 1135.650 162.000 ;
    END
  END la_oenb_core[63]
  PIN la_oenb_core[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.410 156.000 1146.690 162.000 ;
    END
  END la_oenb_core[64]
  PIN la_oenb_core[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1157.450 156.000 1157.730 162.000 ;
    END
  END la_oenb_core[65]
  PIN la_oenb_core[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.490 156.000 1168.770 162.000 ;
    END
  END la_oenb_core[66]
  PIN la_oenb_core[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.530 156.000 1179.810 162.000 ;
    END
  END la_oenb_core[67]
  PIN la_oenb_core[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.570 156.000 1190.850 162.000 ;
    END
  END la_oenb_core[68]
  PIN la_oenb_core[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.610 156.000 1201.890 162.000 ;
    END
  END la_oenb_core[69]
  PIN la_oenb_core[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 156.000 506.370 162.000 ;
    END
  END la_oenb_core[6]
  PIN la_oenb_core[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1212.650 156.000 1212.930 162.000 ;
    END
  END la_oenb_core[70]
  PIN la_oenb_core[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.690 156.000 1223.970 162.000 ;
    END
  END la_oenb_core[71]
  PIN la_oenb_core[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1234.730 156.000 1235.010 162.000 ;
    END
  END la_oenb_core[72]
  PIN la_oenb_core[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1245.770 156.000 1246.050 162.000 ;
    END
  END la_oenb_core[73]
  PIN la_oenb_core[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1256.810 156.000 1257.090 162.000 ;
    END
  END la_oenb_core[74]
  PIN la_oenb_core[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.850 156.000 1268.130 162.000 ;
    END
  END la_oenb_core[75]
  PIN la_oenb_core[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.890 156.000 1279.170 162.000 ;
    END
  END la_oenb_core[76]
  PIN la_oenb_core[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1289.930 156.000 1290.210 162.000 ;
    END
  END la_oenb_core[77]
  PIN la_oenb_core[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1300.970 156.000 1301.250 162.000 ;
    END
  END la_oenb_core[78]
  PIN la_oenb_core[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1312.010 156.000 1312.290 162.000 ;
    END
  END la_oenb_core[79]
  PIN la_oenb_core[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.130 156.000 517.410 162.000 ;
    END
  END la_oenb_core[7]
  PIN la_oenb_core[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.050 156.000 1323.330 162.000 ;
    END
  END la_oenb_core[80]
  PIN la_oenb_core[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1334.090 156.000 1334.370 162.000 ;
    END
  END la_oenb_core[81]
  PIN la_oenb_core[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1345.130 156.000 1345.410 162.000 ;
    END
  END la_oenb_core[82]
  PIN la_oenb_core[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.170 156.000 1356.450 162.000 ;
    END
  END la_oenb_core[83]
  PIN la_oenb_core[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.210 156.000 1367.490 162.000 ;
    END
  END la_oenb_core[84]
  PIN la_oenb_core[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.250 156.000 1378.530 162.000 ;
    END
  END la_oenb_core[85]
  PIN la_oenb_core[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1389.290 156.000 1389.570 162.000 ;
    END
  END la_oenb_core[86]
  PIN la_oenb_core[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.330 156.000 1400.610 162.000 ;
    END
  END la_oenb_core[87]
  PIN la_oenb_core[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1411.370 156.000 1411.650 162.000 ;
    END
  END la_oenb_core[88]
  PIN la_oenb_core[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1422.410 156.000 1422.690 162.000 ;
    END
  END la_oenb_core[89]
  PIN la_oenb_core[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 156.000 528.450 162.000 ;
    END
  END la_oenb_core[8]
  PIN la_oenb_core[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1433.450 156.000 1433.730 162.000 ;
    END
  END la_oenb_core[90]
  PIN la_oenb_core[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.490 156.000 1444.770 162.000 ;
    END
  END la_oenb_core[91]
  PIN la_oenb_core[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.530 156.000 1455.810 162.000 ;
    END
  END la_oenb_core[92]
  PIN la_oenb_core[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1466.570 156.000 1466.850 162.000 ;
    END
  END la_oenb_core[93]
  PIN la_oenb_core[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1477.610 156.000 1477.890 162.000 ;
    END
  END la_oenb_core[94]
  PIN la_oenb_core[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1488.650 156.000 1488.930 162.000 ;
    END
  END la_oenb_core[95]
  PIN la_oenb_core[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1499.690 156.000 1499.970 162.000 ;
    END
  END la_oenb_core[96]
  PIN la_oenb_core[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1510.730 156.000 1511.010 162.000 ;
    END
  END la_oenb_core[97]
  PIN la_oenb_core[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.770 156.000 1522.050 162.000 ;
    END
  END la_oenb_core[98]
  PIN la_oenb_core[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1532.810 156.000 1533.090 162.000 ;
    END
  END la_oenb_core[99]
  PIN la_oenb_core[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 156.000 539.490 162.000 ;
    END
  END la_oenb_core[9]
  PIN la_oenb_mprj[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 -2.000 108.010 4.000 ;
    END
  END la_oenb_mprj[0]
  PIN la_oenb_mprj[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1211.730 -2.000 1212.010 4.000 ;
    END
  END la_oenb_mprj[100]
  PIN la_oenb_mprj[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1222.770 -2.000 1223.050 4.000 ;
    END
  END la_oenb_mprj[101]
  PIN la_oenb_mprj[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.810 -2.000 1234.090 4.000 ;
    END
  END la_oenb_mprj[102]
  PIN la_oenb_mprj[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1244.850 -2.000 1245.130 4.000 ;
    END
  END la_oenb_mprj[103]
  PIN la_oenb_mprj[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.890 -2.000 1256.170 4.000 ;
    END
  END la_oenb_mprj[104]
  PIN la_oenb_mprj[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.930 -2.000 1267.210 4.000 ;
    END
  END la_oenb_mprj[105]
  PIN la_oenb_mprj[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1277.970 -2.000 1278.250 4.000 ;
    END
  END la_oenb_mprj[106]
  PIN la_oenb_mprj[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1289.010 -2.000 1289.290 4.000 ;
    END
  END la_oenb_mprj[107]
  PIN la_oenb_mprj[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1300.050 -2.000 1300.330 4.000 ;
    END
  END la_oenb_mprj[108]
  PIN la_oenb_mprj[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1311.090 -2.000 1311.370 4.000 ;
    END
  END la_oenb_mprj[109]
  PIN la_oenb_mprj[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 -2.000 218.410 4.000 ;
    END
  END la_oenb_mprj[10]
  PIN la_oenb_mprj[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1322.130 -2.000 1322.410 4.000 ;
    END
  END la_oenb_mprj[110]
  PIN la_oenb_mprj[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.170 -2.000 1333.450 4.000 ;
    END
  END la_oenb_mprj[111]
  PIN la_oenb_mprj[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.210 -2.000 1344.490 4.000 ;
    END
  END la_oenb_mprj[112]
  PIN la_oenb_mprj[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.250 -2.000 1355.530 4.000 ;
    END
  END la_oenb_mprj[113]
  PIN la_oenb_mprj[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1366.290 -2.000 1366.570 4.000 ;
    END
  END la_oenb_mprj[114]
  PIN la_oenb_mprj[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1377.330 -2.000 1377.610 4.000 ;
    END
  END la_oenb_mprj[115]
  PIN la_oenb_mprj[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1388.370 -2.000 1388.650 4.000 ;
    END
  END la_oenb_mprj[116]
  PIN la_oenb_mprj[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1399.410 -2.000 1399.690 4.000 ;
    END
  END la_oenb_mprj[117]
  PIN la_oenb_mprj[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.450 -2.000 1410.730 4.000 ;
    END
  END la_oenb_mprj[118]
  PIN la_oenb_mprj[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.490 -2.000 1421.770 4.000 ;
    END
  END la_oenb_mprj[119]
  PIN la_oenb_mprj[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 -2.000 229.450 4.000 ;
    END
  END la_oenb_mprj[11]
  PIN la_oenb_mprj[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.530 -2.000 1432.810 4.000 ;
    END
  END la_oenb_mprj[120]
  PIN la_oenb_mprj[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1443.570 -2.000 1443.850 4.000 ;
    END
  END la_oenb_mprj[121]
  PIN la_oenb_mprj[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1454.610 -2.000 1454.890 4.000 ;
    END
  END la_oenb_mprj[122]
  PIN la_oenb_mprj[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.650 -2.000 1465.930 4.000 ;
    END
  END la_oenb_mprj[123]
  PIN la_oenb_mprj[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1476.690 -2.000 1476.970 4.000 ;
    END
  END la_oenb_mprj[124]
  PIN la_oenb_mprj[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1487.730 -2.000 1488.010 4.000 ;
    END
  END la_oenb_mprj[125]
  PIN la_oenb_mprj[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1498.770 -2.000 1499.050 4.000 ;
    END
  END la_oenb_mprj[126]
  PIN la_oenb_mprj[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1509.810 -2.000 1510.090 4.000 ;
    END
  END la_oenb_mprj[127]
  PIN la_oenb_mprj[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 -2.000 240.490 4.000 ;
    END
  END la_oenb_mprj[12]
  PIN la_oenb_mprj[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 -2.000 251.530 4.000 ;
    END
  END la_oenb_mprj[13]
  PIN la_oenb_mprj[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 -2.000 262.570 4.000 ;
    END
  END la_oenb_mprj[14]
  PIN la_oenb_mprj[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 -2.000 273.610 4.000 ;
    END
  END la_oenb_mprj[15]
  PIN la_oenb_mprj[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 -2.000 284.650 4.000 ;
    END
  END la_oenb_mprj[16]
  PIN la_oenb_mprj[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 -2.000 295.690 4.000 ;
    END
  END la_oenb_mprj[17]
  PIN la_oenb_mprj[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 -2.000 306.730 4.000 ;
    END
  END la_oenb_mprj[18]
  PIN la_oenb_mprj[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 -2.000 317.770 4.000 ;
    END
  END la_oenb_mprj[19]
  PIN la_oenb_mprj[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 -2.000 119.050 4.000 ;
    END
  END la_oenb_mprj[1]
  PIN la_oenb_mprj[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 -2.000 328.810 4.000 ;
    END
  END la_oenb_mprj[20]
  PIN la_oenb_mprj[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 -2.000 339.850 4.000 ;
    END
  END la_oenb_mprj[21]
  PIN la_oenb_mprj[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 -2.000 350.890 4.000 ;
    END
  END la_oenb_mprj[22]
  PIN la_oenb_mprj[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 -2.000 361.930 4.000 ;
    END
  END la_oenb_mprj[23]
  PIN la_oenb_mprj[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 -2.000 372.970 4.000 ;
    END
  END la_oenb_mprj[24]
  PIN la_oenb_mprj[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.730 -2.000 384.010 4.000 ;
    END
  END la_oenb_mprj[25]
  PIN la_oenb_mprj[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 -2.000 395.050 4.000 ;
    END
  END la_oenb_mprj[26]
  PIN la_oenb_mprj[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 -2.000 406.090 4.000 ;
    END
  END la_oenb_mprj[27]
  PIN la_oenb_mprj[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 -2.000 417.130 4.000 ;
    END
  END la_oenb_mprj[28]
  PIN la_oenb_mprj[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 -2.000 428.170 4.000 ;
    END
  END la_oenb_mprj[29]
  PIN la_oenb_mprj[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 -2.000 130.090 4.000 ;
    END
  END la_oenb_mprj[2]
  PIN la_oenb_mprj[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 -2.000 439.210 4.000 ;
    END
  END la_oenb_mprj[30]
  PIN la_oenb_mprj[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 -2.000 450.250 4.000 ;
    END
  END la_oenb_mprj[31]
  PIN la_oenb_mprj[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 -2.000 461.290 4.000 ;
    END
  END la_oenb_mprj[32]
  PIN la_oenb_mprj[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.050 -2.000 472.330 4.000 ;
    END
  END la_oenb_mprj[33]
  PIN la_oenb_mprj[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 -2.000 483.370 4.000 ;
    END
  END la_oenb_mprj[34]
  PIN la_oenb_mprj[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.130 -2.000 494.410 4.000 ;
    END
  END la_oenb_mprj[35]
  PIN la_oenb_mprj[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 -2.000 505.450 4.000 ;
    END
  END la_oenb_mprj[36]
  PIN la_oenb_mprj[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 -2.000 516.490 4.000 ;
    END
  END la_oenb_mprj[37]
  PIN la_oenb_mprj[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.250 -2.000 527.530 4.000 ;
    END
  END la_oenb_mprj[38]
  PIN la_oenb_mprj[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 -2.000 538.570 4.000 ;
    END
  END la_oenb_mprj[39]
  PIN la_oenb_mprj[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 -2.000 141.130 4.000 ;
    END
  END la_oenb_mprj[3]
  PIN la_oenb_mprj[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.330 -2.000 549.610 4.000 ;
    END
  END la_oenb_mprj[40]
  PIN la_oenb_mprj[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 -2.000 560.650 4.000 ;
    END
  END la_oenb_mprj[41]
  PIN la_oenb_mprj[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 -2.000 571.690 4.000 ;
    END
  END la_oenb_mprj[42]
  PIN la_oenb_mprj[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.450 -2.000 582.730 4.000 ;
    END
  END la_oenb_mprj[43]
  PIN la_oenb_mprj[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.490 -2.000 593.770 4.000 ;
    END
  END la_oenb_mprj[44]
  PIN la_oenb_mprj[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 -2.000 604.810 4.000 ;
    END
  END la_oenb_mprj[45]
  PIN la_oenb_mprj[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.570 -2.000 615.850 4.000 ;
    END
  END la_oenb_mprj[46]
  PIN la_oenb_mprj[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.610 -2.000 626.890 4.000 ;
    END
  END la_oenb_mprj[47]
  PIN la_oenb_mprj[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 -2.000 637.930 4.000 ;
    END
  END la_oenb_mprj[48]
  PIN la_oenb_mprj[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.690 -2.000 648.970 4.000 ;
    END
  END la_oenb_mprj[49]
  PIN la_oenb_mprj[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 -2.000 152.170 4.000 ;
    END
  END la_oenb_mprj[4]
  PIN la_oenb_mprj[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.730 -2.000 660.010 4.000 ;
    END
  END la_oenb_mprj[50]
  PIN la_oenb_mprj[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.770 -2.000 671.050 4.000 ;
    END
  END la_oenb_mprj[51]
  PIN la_oenb_mprj[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 -2.000 682.090 4.000 ;
    END
  END la_oenb_mprj[52]
  PIN la_oenb_mprj[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.850 -2.000 693.130 4.000 ;
    END
  END la_oenb_mprj[53]
  PIN la_oenb_mprj[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 -2.000 704.170 4.000 ;
    END
  END la_oenb_mprj[54]
  PIN la_oenb_mprj[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 -2.000 715.210 4.000 ;
    END
  END la_oenb_mprj[55]
  PIN la_oenb_mprj[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.970 -2.000 726.250 4.000 ;
    END
  END la_oenb_mprj[56]
  PIN la_oenb_mprj[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 -2.000 737.290 4.000 ;
    END
  END la_oenb_mprj[57]
  PIN la_oenb_mprj[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.050 -2.000 748.330 4.000 ;
    END
  END la_oenb_mprj[58]
  PIN la_oenb_mprj[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 -2.000 759.370 4.000 ;
    END
  END la_oenb_mprj[59]
  PIN la_oenb_mprj[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 -2.000 163.210 4.000 ;
    END
  END la_oenb_mprj[5]
  PIN la_oenb_mprj[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.130 -2.000 770.410 4.000 ;
    END
  END la_oenb_mprj[60]
  PIN la_oenb_mprj[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.170 -2.000 781.450 4.000 ;
    END
  END la_oenb_mprj[61]
  PIN la_oenb_mprj[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 -2.000 792.490 4.000 ;
    END
  END la_oenb_mprj[62]
  PIN la_oenb_mprj[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.250 -2.000 803.530 4.000 ;
    END
  END la_oenb_mprj[63]
  PIN la_oenb_mprj[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 -2.000 814.570 4.000 ;
    END
  END la_oenb_mprj[64]
  PIN la_oenb_mprj[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.330 -2.000 825.610 4.000 ;
    END
  END la_oenb_mprj[65]
  PIN la_oenb_mprj[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.370 -2.000 836.650 4.000 ;
    END
  END la_oenb_mprj[66]
  PIN la_oenb_mprj[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.410 -2.000 847.690 4.000 ;
    END
  END la_oenb_mprj[67]
  PIN la_oenb_mprj[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.450 -2.000 858.730 4.000 ;
    END
  END la_oenb_mprj[68]
  PIN la_oenb_mprj[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 -2.000 869.770 4.000 ;
    END
  END la_oenb_mprj[69]
  PIN la_oenb_mprj[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 -2.000 174.250 4.000 ;
    END
  END la_oenb_mprj[6]
  PIN la_oenb_mprj[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.530 -2.000 880.810 4.000 ;
    END
  END la_oenb_mprj[70]
  PIN la_oenb_mprj[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.570 -2.000 891.850 4.000 ;
    END
  END la_oenb_mprj[71]
  PIN la_oenb_mprj[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.610 -2.000 902.890 4.000 ;
    END
  END la_oenb_mprj[72]
  PIN la_oenb_mprj[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.650 -2.000 913.930 4.000 ;
    END
  END la_oenb_mprj[73]
  PIN la_oenb_mprj[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.690 -2.000 924.970 4.000 ;
    END
  END la_oenb_mprj[74]
  PIN la_oenb_mprj[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.730 -2.000 936.010 4.000 ;
    END
  END la_oenb_mprj[75]
  PIN la_oenb_mprj[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.770 -2.000 947.050 4.000 ;
    END
  END la_oenb_mprj[76]
  PIN la_oenb_mprj[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.810 -2.000 958.090 4.000 ;
    END
  END la_oenb_mprj[77]
  PIN la_oenb_mprj[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.850 -2.000 969.130 4.000 ;
    END
  END la_oenb_mprj[78]
  PIN la_oenb_mprj[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.890 -2.000 980.170 4.000 ;
    END
  END la_oenb_mprj[79]
  PIN la_oenb_mprj[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 -2.000 185.290 4.000 ;
    END
  END la_oenb_mprj[7]
  PIN la_oenb_mprj[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.930 -2.000 991.210 4.000 ;
    END
  END la_oenb_mprj[80]
  PIN la_oenb_mprj[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.970 -2.000 1002.250 4.000 ;
    END
  END la_oenb_mprj[81]
  PIN la_oenb_mprj[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.010 -2.000 1013.290 4.000 ;
    END
  END la_oenb_mprj[82]
  PIN la_oenb_mprj[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.050 -2.000 1024.330 4.000 ;
    END
  END la_oenb_mprj[83]
  PIN la_oenb_mprj[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1035.090 -2.000 1035.370 4.000 ;
    END
  END la_oenb_mprj[84]
  PIN la_oenb_mprj[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.130 -2.000 1046.410 4.000 ;
    END
  END la_oenb_mprj[85]
  PIN la_oenb_mprj[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1057.170 -2.000 1057.450 4.000 ;
    END
  END la_oenb_mprj[86]
  PIN la_oenb_mprj[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1068.210 -2.000 1068.490 4.000 ;
    END
  END la_oenb_mprj[87]
  PIN la_oenb_mprj[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.250 -2.000 1079.530 4.000 ;
    END
  END la_oenb_mprj[88]
  PIN la_oenb_mprj[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.290 -2.000 1090.570 4.000 ;
    END
  END la_oenb_mprj[89]
  PIN la_oenb_mprj[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 -2.000 196.330 4.000 ;
    END
  END la_oenb_mprj[8]
  PIN la_oenb_mprj[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.330 -2.000 1101.610 4.000 ;
    END
  END la_oenb_mprj[90]
  PIN la_oenb_mprj[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1112.370 -2.000 1112.650 4.000 ;
    END
  END la_oenb_mprj[91]
  PIN la_oenb_mprj[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.410 -2.000 1123.690 4.000 ;
    END
  END la_oenb_mprj[92]
  PIN la_oenb_mprj[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.450 -2.000 1134.730 4.000 ;
    END
  END la_oenb_mprj[93]
  PIN la_oenb_mprj[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.490 -2.000 1145.770 4.000 ;
    END
  END la_oenb_mprj[94]
  PIN la_oenb_mprj[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.530 -2.000 1156.810 4.000 ;
    END
  END la_oenb_mprj[95]
  PIN la_oenb_mprj[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1167.570 -2.000 1167.850 4.000 ;
    END
  END la_oenb_mprj[96]
  PIN la_oenb_mprj[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.610 -2.000 1178.890 4.000 ;
    END
  END la_oenb_mprj[97]
  PIN la_oenb_mprj[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1189.650 -2.000 1189.930 4.000 ;
    END
  END la_oenb_mprj[98]
  PIN la_oenb_mprj[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1200.690 -2.000 1200.970 4.000 ;
    END
  END la_oenb_mprj[99]
  PIN la_oenb_mprj[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 -2.000 207.370 4.000 ;
    END
  END la_oenb_mprj[9]
  PIN mprj_ack_i_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1512.570 -2.000 1512.850 4.000 ;
    END
  END mprj_ack_i_core
  PIN mprj_ack_i_user
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 156.000 50.050 162.000 ;
    END
  END mprj_ack_i_user
  PIN mprj_adr_o_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.610 -2.000 1523.890 4.000 ;
    END
  END mprj_adr_o_core[0]
  PIN mprj_adr_o_core[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1617.450 -2.000 1617.730 4.000 ;
    END
  END mprj_adr_o_core[10]
  PIN mprj_adr_o_core[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1625.730 -2.000 1626.010 4.000 ;
    END
  END mprj_adr_o_core[11]
  PIN mprj_adr_o_core[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1634.010 -2.000 1634.290 4.000 ;
    END
  END mprj_adr_o_core[12]
  PIN mprj_adr_o_core[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1642.290 -2.000 1642.570 4.000 ;
    END
  END mprj_adr_o_core[13]
  PIN mprj_adr_o_core[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1650.570 -2.000 1650.850 4.000 ;
    END
  END mprj_adr_o_core[14]
  PIN mprj_adr_o_core[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.850 -2.000 1659.130 4.000 ;
    END
  END mprj_adr_o_core[15]
  PIN mprj_adr_o_core[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1667.130 -2.000 1667.410 4.000 ;
    END
  END mprj_adr_o_core[16]
  PIN mprj_adr_o_core[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.410 -2.000 1675.690 4.000 ;
    END
  END mprj_adr_o_core[17]
  PIN mprj_adr_o_core[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1683.690 -2.000 1683.970 4.000 ;
    END
  END mprj_adr_o_core[18]
  PIN mprj_adr_o_core[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.970 -2.000 1692.250 4.000 ;
    END
  END mprj_adr_o_core[19]
  PIN mprj_adr_o_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1534.650 -2.000 1534.930 4.000 ;
    END
  END mprj_adr_o_core[1]
  PIN mprj_adr_o_core[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1700.250 -2.000 1700.530 4.000 ;
    END
  END mprj_adr_o_core[20]
  PIN mprj_adr_o_core[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1708.530 -2.000 1708.810 4.000 ;
    END
  END mprj_adr_o_core[21]
  PIN mprj_adr_o_core[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.810 -2.000 1717.090 4.000 ;
    END
  END mprj_adr_o_core[22]
  PIN mprj_adr_o_core[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1725.090 -2.000 1725.370 4.000 ;
    END
  END mprj_adr_o_core[23]
  PIN mprj_adr_o_core[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1733.370 -2.000 1733.650 4.000 ;
    END
  END mprj_adr_o_core[24]
  PIN mprj_adr_o_core[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1741.650 -2.000 1741.930 4.000 ;
    END
  END mprj_adr_o_core[25]
  PIN mprj_adr_o_core[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1749.930 -2.000 1750.210 4.000 ;
    END
  END mprj_adr_o_core[26]
  PIN mprj_adr_o_core[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.210 -2.000 1758.490 4.000 ;
    END
  END mprj_adr_o_core[27]
  PIN mprj_adr_o_core[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1766.490 -2.000 1766.770 4.000 ;
    END
  END mprj_adr_o_core[28]
  PIN mprj_adr_o_core[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1774.770 -2.000 1775.050 4.000 ;
    END
  END mprj_adr_o_core[29]
  PIN mprj_adr_o_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.690 -2.000 1545.970 4.000 ;
    END
  END mprj_adr_o_core[2]
  PIN mprj_adr_o_core[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.050 -2.000 1783.330 4.000 ;
    END
  END mprj_adr_o_core[30]
  PIN mprj_adr_o_core[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1791.330 -2.000 1791.610 4.000 ;
    END
  END mprj_adr_o_core[31]
  PIN mprj_adr_o_core[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1556.730 -2.000 1557.010 4.000 ;
    END
  END mprj_adr_o_core[3]
  PIN mprj_adr_o_core[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1567.770 -2.000 1568.050 4.000 ;
    END
  END mprj_adr_o_core[4]
  PIN mprj_adr_o_core[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1576.050 -2.000 1576.330 4.000 ;
    END
  END mprj_adr_o_core[5]
  PIN mprj_adr_o_core[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.330 -2.000 1584.610 4.000 ;
    END
  END mprj_adr_o_core[6]
  PIN mprj_adr_o_core[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.610 -2.000 1592.890 4.000 ;
    END
  END mprj_adr_o_core[7]
  PIN mprj_adr_o_core[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1600.890 -2.000 1601.170 4.000 ;
    END
  END mprj_adr_o_core[8]
  PIN mprj_adr_o_core[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1609.170 -2.000 1609.450 4.000 ;
    END
  END mprj_adr_o_core[9]
  PIN mprj_adr_o_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 156.000 64.770 162.000 ;
    END
  END mprj_adr_o_user[0]
  PIN mprj_adr_o_user[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 156.000 189.890 162.000 ;
    END
  END mprj_adr_o_user[10]
  PIN mprj_adr_o_user[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 156.000 200.930 162.000 ;
    END
  END mprj_adr_o_user[11]
  PIN mprj_adr_o_user[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 156.000 211.970 162.000 ;
    END
  END mprj_adr_o_user[12]
  PIN mprj_adr_o_user[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 156.000 223.010 162.000 ;
    END
  END mprj_adr_o_user[13]
  PIN mprj_adr_o_user[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 156.000 234.050 162.000 ;
    END
  END mprj_adr_o_user[14]
  PIN mprj_adr_o_user[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 156.000 245.090 162.000 ;
    END
  END mprj_adr_o_user[15]
  PIN mprj_adr_o_user[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 156.000 256.130 162.000 ;
    END
  END mprj_adr_o_user[16]
  PIN mprj_adr_o_user[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 156.000 267.170 162.000 ;
    END
  END mprj_adr_o_user[17]
  PIN mprj_adr_o_user[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 156.000 278.210 162.000 ;
    END
  END mprj_adr_o_user[18]
  PIN mprj_adr_o_user[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 156.000 289.250 162.000 ;
    END
  END mprj_adr_o_user[19]
  PIN mprj_adr_o_user[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 156.000 79.490 162.000 ;
    END
  END mprj_adr_o_user[1]
  PIN mprj_adr_o_user[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 156.000 300.290 162.000 ;
    END
  END mprj_adr_o_user[20]
  PIN mprj_adr_o_user[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 156.000 311.330 162.000 ;
    END
  END mprj_adr_o_user[21]
  PIN mprj_adr_o_user[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 156.000 322.370 162.000 ;
    END
  END mprj_adr_o_user[22]
  PIN mprj_adr_o_user[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 156.000 333.410 162.000 ;
    END
  END mprj_adr_o_user[23]
  PIN mprj_adr_o_user[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 156.000 344.450 162.000 ;
    END
  END mprj_adr_o_user[24]
  PIN mprj_adr_o_user[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 156.000 355.490 162.000 ;
    END
  END mprj_adr_o_user[25]
  PIN mprj_adr_o_user[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 156.000 366.530 162.000 ;
    END
  END mprj_adr_o_user[26]
  PIN mprj_adr_o_user[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 156.000 377.570 162.000 ;
    END
  END mprj_adr_o_user[27]
  PIN mprj_adr_o_user[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 156.000 388.610 162.000 ;
    END
  END mprj_adr_o_user[28]
  PIN mprj_adr_o_user[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 156.000 399.650 162.000 ;
    END
  END mprj_adr_o_user[29]
  PIN mprj_adr_o_user[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 156.000 94.210 162.000 ;
    END
  END mprj_adr_o_user[2]
  PIN mprj_adr_o_user[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 156.000 410.690 162.000 ;
    END
  END mprj_adr_o_user[30]
  PIN mprj_adr_o_user[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 156.000 421.730 162.000 ;
    END
  END mprj_adr_o_user[31]
  PIN mprj_adr_o_user[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 156.000 108.930 162.000 ;
    END
  END mprj_adr_o_user[3]
  PIN mprj_adr_o_user[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 156.000 123.650 162.000 ;
    END
  END mprj_adr_o_user[4]
  PIN mprj_adr_o_user[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 156.000 134.690 162.000 ;
    END
  END mprj_adr_o_user[5]
  PIN mprj_adr_o_user[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 156.000 145.730 162.000 ;
    END
  END mprj_adr_o_user[6]
  PIN mprj_adr_o_user[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 156.000 156.770 162.000 ;
    END
  END mprj_adr_o_user[7]
  PIN mprj_adr_o_user[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 156.000 167.810 162.000 ;
    END
  END mprj_adr_o_user[8]
  PIN mprj_adr_o_user[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 156.000 178.850 162.000 ;
    END
  END mprj_adr_o_user[9]
  PIN mprj_cyc_o_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.330 -2.000 1515.610 4.000 ;
    END
  END mprj_cyc_o_core
  PIN mprj_cyc_o_user
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 156.000 53.730 162.000 ;
    END
  END mprj_cyc_o_user
  PIN mprj_dat_i_core[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.370 -2.000 1526.650 4.000 ;
    END
  END mprj_dat_i_core[0]
  PIN mprj_dat_i_core[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1620.210 -2.000 1620.490 4.000 ;
    END
  END mprj_dat_i_core[10]
  PIN mprj_dat_i_core[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1628.490 -2.000 1628.770 4.000 ;
    END
  END mprj_dat_i_core[11]
  PIN mprj_dat_i_core[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1636.770 -2.000 1637.050 4.000 ;
    END
  END mprj_dat_i_core[12]
  PIN mprj_dat_i_core[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.050 -2.000 1645.330 4.000 ;
    END
  END mprj_dat_i_core[13]
  PIN mprj_dat_i_core[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1653.330 -2.000 1653.610 4.000 ;
    END
  END mprj_dat_i_core[14]
  PIN mprj_dat_i_core[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.610 -2.000 1661.890 4.000 ;
    END
  END mprj_dat_i_core[15]
  PIN mprj_dat_i_core[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1669.890 -2.000 1670.170 4.000 ;
    END
  END mprj_dat_i_core[16]
  PIN mprj_dat_i_core[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1678.170 -2.000 1678.450 4.000 ;
    END
  END mprj_dat_i_core[17]
  PIN mprj_dat_i_core[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1686.450 -2.000 1686.730 4.000 ;
    END
  END mprj_dat_i_core[18]
  PIN mprj_dat_i_core[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1694.730 -2.000 1695.010 4.000 ;
    END
  END mprj_dat_i_core[19]
  PIN mprj_dat_i_core[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1537.410 -2.000 1537.690 4.000 ;
    END
  END mprj_dat_i_core[1]
  PIN mprj_dat_i_core[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.010 -2.000 1703.290 4.000 ;
    END
  END mprj_dat_i_core[20]
  PIN mprj_dat_i_core[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1711.290 -2.000 1711.570 4.000 ;
    END
  END mprj_dat_i_core[21]
  PIN mprj_dat_i_core[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1719.570 -2.000 1719.850 4.000 ;
    END
  END mprj_dat_i_core[22]
  PIN mprj_dat_i_core[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1727.850 -2.000 1728.130 4.000 ;
    END
  END mprj_dat_i_core[23]
  PIN mprj_dat_i_core[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1736.130 -2.000 1736.410 4.000 ;
    END
  END mprj_dat_i_core[24]
  PIN mprj_dat_i_core[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1744.410 -2.000 1744.690 4.000 ;
    END
  END mprj_dat_i_core[25]
  PIN mprj_dat_i_core[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.690 -2.000 1752.970 4.000 ;
    END
  END mprj_dat_i_core[26]
  PIN mprj_dat_i_core[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.970 -2.000 1761.250 4.000 ;
    END
  END mprj_dat_i_core[27]
  PIN mprj_dat_i_core[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1769.250 -2.000 1769.530 4.000 ;
    END
  END mprj_dat_i_core[28]
  PIN mprj_dat_i_core[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1777.530 -2.000 1777.810 4.000 ;
    END
  END mprj_dat_i_core[29]
  PIN mprj_dat_i_core[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.450 -2.000 1548.730 4.000 ;
    END
  END mprj_dat_i_core[2]
  PIN mprj_dat_i_core[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1785.810 -2.000 1786.090 4.000 ;
    END
  END mprj_dat_i_core[30]
  PIN mprj_dat_i_core[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1794.090 -2.000 1794.370 4.000 ;
    END
  END mprj_dat_i_core[31]
  PIN mprj_dat_i_core[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1559.490 -2.000 1559.770 4.000 ;
    END
  END mprj_dat_i_core[3]
  PIN mprj_dat_i_core[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1570.530 -2.000 1570.810 4.000 ;
    END
  END mprj_dat_i_core[4]
  PIN mprj_dat_i_core[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1578.810 -2.000 1579.090 4.000 ;
    END
  END mprj_dat_i_core[5]
  PIN mprj_dat_i_core[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1587.090 -2.000 1587.370 4.000 ;
    END
  END mprj_dat_i_core[6]
  PIN mprj_dat_i_core[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1595.370 -2.000 1595.650 4.000 ;
    END
  END mprj_dat_i_core[7]
  PIN mprj_dat_i_core[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.650 -2.000 1603.930 4.000 ;
    END
  END mprj_dat_i_core[8]
  PIN mprj_dat_i_core[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1611.930 -2.000 1612.210 4.000 ;
    END
  END mprj_dat_i_core[9]
  PIN mprj_dat_i_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 156.000 68.450 162.000 ;
    END
  END mprj_dat_i_user[0]
  PIN mprj_dat_i_user[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 156.000 193.570 162.000 ;
    END
  END mprj_dat_i_user[10]
  PIN mprj_dat_i_user[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 156.000 204.610 162.000 ;
    END
  END mprj_dat_i_user[11]
  PIN mprj_dat_i_user[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 156.000 215.650 162.000 ;
    END
  END mprj_dat_i_user[12]
  PIN mprj_dat_i_user[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 156.000 226.690 162.000 ;
    END
  END mprj_dat_i_user[13]
  PIN mprj_dat_i_user[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 156.000 237.730 162.000 ;
    END
  END mprj_dat_i_user[14]
  PIN mprj_dat_i_user[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 156.000 248.770 162.000 ;
    END
  END mprj_dat_i_user[15]
  PIN mprj_dat_i_user[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 156.000 259.810 162.000 ;
    END
  END mprj_dat_i_user[16]
  PIN mprj_dat_i_user[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 156.000 270.850 162.000 ;
    END
  END mprj_dat_i_user[17]
  PIN mprj_dat_i_user[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 156.000 281.890 162.000 ;
    END
  END mprj_dat_i_user[18]
  PIN mprj_dat_i_user[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 156.000 292.930 162.000 ;
    END
  END mprj_dat_i_user[19]
  PIN mprj_dat_i_user[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 156.000 83.170 162.000 ;
    END
  END mprj_dat_i_user[1]
  PIN mprj_dat_i_user[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 156.000 303.970 162.000 ;
    END
  END mprj_dat_i_user[20]
  PIN mprj_dat_i_user[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 156.000 315.010 162.000 ;
    END
  END mprj_dat_i_user[21]
  PIN mprj_dat_i_user[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 156.000 326.050 162.000 ;
    END
  END mprj_dat_i_user[22]
  PIN mprj_dat_i_user[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 156.000 337.090 162.000 ;
    END
  END mprj_dat_i_user[23]
  PIN mprj_dat_i_user[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 156.000 348.130 162.000 ;
    END
  END mprj_dat_i_user[24]
  PIN mprj_dat_i_user[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 156.000 359.170 162.000 ;
    END
  END mprj_dat_i_user[25]
  PIN mprj_dat_i_user[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 156.000 370.210 162.000 ;
    END
  END mprj_dat_i_user[26]
  PIN mprj_dat_i_user[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 156.000 381.250 162.000 ;
    END
  END mprj_dat_i_user[27]
  PIN mprj_dat_i_user[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 156.000 392.290 162.000 ;
    END
  END mprj_dat_i_user[28]
  PIN mprj_dat_i_user[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 156.000 403.330 162.000 ;
    END
  END mprj_dat_i_user[29]
  PIN mprj_dat_i_user[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 156.000 97.890 162.000 ;
    END
  END mprj_dat_i_user[2]
  PIN mprj_dat_i_user[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 156.000 414.370 162.000 ;
    END
  END mprj_dat_i_user[30]
  PIN mprj_dat_i_user[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 156.000 425.410 162.000 ;
    END
  END mprj_dat_i_user[31]
  PIN mprj_dat_i_user[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 156.000 112.610 162.000 ;
    END
  END mprj_dat_i_user[3]
  PIN mprj_dat_i_user[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 156.000 127.330 162.000 ;
    END
  END mprj_dat_i_user[4]
  PIN mprj_dat_i_user[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 156.000 138.370 162.000 ;
    END
  END mprj_dat_i_user[5]
  PIN mprj_dat_i_user[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 156.000 149.410 162.000 ;
    END
  END mprj_dat_i_user[6]
  PIN mprj_dat_i_user[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 156.000 160.450 162.000 ;
    END
  END mprj_dat_i_user[7]
  PIN mprj_dat_i_user[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 156.000 171.490 162.000 ;
    END
  END mprj_dat_i_user[8]
  PIN mprj_dat_i_user[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 156.000 182.530 162.000 ;
    END
  END mprj_dat_i_user[9]
  PIN mprj_dat_o_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1529.130 -2.000 1529.410 4.000 ;
    END
  END mprj_dat_o_core[0]
  PIN mprj_dat_o_core[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.970 -2.000 1623.250 4.000 ;
    END
  END mprj_dat_o_core[10]
  PIN mprj_dat_o_core[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1631.250 -2.000 1631.530 4.000 ;
    END
  END mprj_dat_o_core[11]
  PIN mprj_dat_o_core[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.530 -2.000 1639.810 4.000 ;
    END
  END mprj_dat_o_core[12]
  PIN mprj_dat_o_core[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1647.810 -2.000 1648.090 4.000 ;
    END
  END mprj_dat_o_core[13]
  PIN mprj_dat_o_core[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1656.090 -2.000 1656.370 4.000 ;
    END
  END mprj_dat_o_core[14]
  PIN mprj_dat_o_core[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1664.370 -2.000 1664.650 4.000 ;
    END
  END mprj_dat_o_core[15]
  PIN mprj_dat_o_core[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1672.650 -2.000 1672.930 4.000 ;
    END
  END mprj_dat_o_core[16]
  PIN mprj_dat_o_core[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1680.930 -2.000 1681.210 4.000 ;
    END
  END mprj_dat_o_core[17]
  PIN mprj_dat_o_core[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1689.210 -2.000 1689.490 4.000 ;
    END
  END mprj_dat_o_core[18]
  PIN mprj_dat_o_core[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.490 -2.000 1697.770 4.000 ;
    END
  END mprj_dat_o_core[19]
  PIN mprj_dat_o_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1540.170 -2.000 1540.450 4.000 ;
    END
  END mprj_dat_o_core[1]
  PIN mprj_dat_o_core[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1705.770 -2.000 1706.050 4.000 ;
    END
  END mprj_dat_o_core[20]
  PIN mprj_dat_o_core[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1714.050 -2.000 1714.330 4.000 ;
    END
  END mprj_dat_o_core[21]
  PIN mprj_dat_o_core[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.330 -2.000 1722.610 4.000 ;
    END
  END mprj_dat_o_core[22]
  PIN mprj_dat_o_core[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1730.610 -2.000 1730.890 4.000 ;
    END
  END mprj_dat_o_core[23]
  PIN mprj_dat_o_core[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1738.890 -2.000 1739.170 4.000 ;
    END
  END mprj_dat_o_core[24]
  PIN mprj_dat_o_core[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1747.170 -2.000 1747.450 4.000 ;
    END
  END mprj_dat_o_core[25]
  PIN mprj_dat_o_core[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1755.450 -2.000 1755.730 4.000 ;
    END
  END mprj_dat_o_core[26]
  PIN mprj_dat_o_core[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1763.730 -2.000 1764.010 4.000 ;
    END
  END mprj_dat_o_core[27]
  PIN mprj_dat_o_core[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1772.010 -2.000 1772.290 4.000 ;
    END
  END mprj_dat_o_core[28]
  PIN mprj_dat_o_core[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1780.290 -2.000 1780.570 4.000 ;
    END
  END mprj_dat_o_core[29]
  PIN mprj_dat_o_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.210 -2.000 1551.490 4.000 ;
    END
  END mprj_dat_o_core[2]
  PIN mprj_dat_o_core[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1788.570 -2.000 1788.850 4.000 ;
    END
  END mprj_dat_o_core[30]
  PIN mprj_dat_o_core[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1796.850 -2.000 1797.130 4.000 ;
    END
  END mprj_dat_o_core[31]
  PIN mprj_dat_o_core[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1562.250 -2.000 1562.530 4.000 ;
    END
  END mprj_dat_o_core[3]
  PIN mprj_dat_o_core[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1573.290 -2.000 1573.570 4.000 ;
    END
  END mprj_dat_o_core[4]
  PIN mprj_dat_o_core[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.570 -2.000 1581.850 4.000 ;
    END
  END mprj_dat_o_core[5]
  PIN mprj_dat_o_core[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1589.850 -2.000 1590.130 4.000 ;
    END
  END mprj_dat_o_core[6]
  PIN mprj_dat_o_core[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.130 -2.000 1598.410 4.000 ;
    END
  END mprj_dat_o_core[7]
  PIN mprj_dat_o_core[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1606.410 -2.000 1606.690 4.000 ;
    END
  END mprj_dat_o_core[8]
  PIN mprj_dat_o_core[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1614.690 -2.000 1614.970 4.000 ;
    END
  END mprj_dat_o_core[9]
  PIN mprj_dat_o_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 156.000 72.130 162.000 ;
    END
  END mprj_dat_o_user[0]
  PIN mprj_dat_o_user[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 156.000 197.250 162.000 ;
    END
  END mprj_dat_o_user[10]
  PIN mprj_dat_o_user[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 156.000 208.290 162.000 ;
    END
  END mprj_dat_o_user[11]
  PIN mprj_dat_o_user[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 156.000 219.330 162.000 ;
    END
  END mprj_dat_o_user[12]
  PIN mprj_dat_o_user[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 156.000 230.370 162.000 ;
    END
  END mprj_dat_o_user[13]
  PIN mprj_dat_o_user[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 156.000 241.410 162.000 ;
    END
  END mprj_dat_o_user[14]
  PIN mprj_dat_o_user[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 156.000 252.450 162.000 ;
    END
  END mprj_dat_o_user[15]
  PIN mprj_dat_o_user[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 156.000 263.490 162.000 ;
    END
  END mprj_dat_o_user[16]
  PIN mprj_dat_o_user[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 156.000 274.530 162.000 ;
    END
  END mprj_dat_o_user[17]
  PIN mprj_dat_o_user[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 156.000 285.570 162.000 ;
    END
  END mprj_dat_o_user[18]
  PIN mprj_dat_o_user[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 156.000 296.610 162.000 ;
    END
  END mprj_dat_o_user[19]
  PIN mprj_dat_o_user[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 156.000 86.850 162.000 ;
    END
  END mprj_dat_o_user[1]
  PIN mprj_dat_o_user[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 156.000 307.650 162.000 ;
    END
  END mprj_dat_o_user[20]
  PIN mprj_dat_o_user[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 156.000 318.690 162.000 ;
    END
  END mprj_dat_o_user[21]
  PIN mprj_dat_o_user[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 156.000 329.730 162.000 ;
    END
  END mprj_dat_o_user[22]
  PIN mprj_dat_o_user[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 156.000 340.770 162.000 ;
    END
  END mprj_dat_o_user[23]
  PIN mprj_dat_o_user[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 156.000 351.810 162.000 ;
    END
  END mprj_dat_o_user[24]
  PIN mprj_dat_o_user[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 156.000 362.850 162.000 ;
    END
  END mprj_dat_o_user[25]
  PIN mprj_dat_o_user[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 156.000 373.890 162.000 ;
    END
  END mprj_dat_o_user[26]
  PIN mprj_dat_o_user[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 156.000 384.930 162.000 ;
    END
  END mprj_dat_o_user[27]
  PIN mprj_dat_o_user[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 156.000 395.970 162.000 ;
    END
  END mprj_dat_o_user[28]
  PIN mprj_dat_o_user[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.730 156.000 407.010 162.000 ;
    END
  END mprj_dat_o_user[29]
  PIN mprj_dat_o_user[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 156.000 101.570 162.000 ;
    END
  END mprj_dat_o_user[2]
  PIN mprj_dat_o_user[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 156.000 418.050 162.000 ;
    END
  END mprj_dat_o_user[30]
  PIN mprj_dat_o_user[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 156.000 429.090 162.000 ;
    END
  END mprj_dat_o_user[31]
  PIN mprj_dat_o_user[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 156.000 116.290 162.000 ;
    END
  END mprj_dat_o_user[3]
  PIN mprj_dat_o_user[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 156.000 131.010 162.000 ;
    END
  END mprj_dat_o_user[4]
  PIN mprj_dat_o_user[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 156.000 142.050 162.000 ;
    END
  END mprj_dat_o_user[5]
  PIN mprj_dat_o_user[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 156.000 153.090 162.000 ;
    END
  END mprj_dat_o_user[6]
  PIN mprj_dat_o_user[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 156.000 164.130 162.000 ;
    END
  END mprj_dat_o_user[7]
  PIN mprj_dat_o_user[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 156.000 175.170 162.000 ;
    END
  END mprj_dat_o_user[8]
  PIN mprj_dat_o_user[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 156.000 186.210 162.000 ;
    END
  END mprj_dat_o_user[9]
  PIN mprj_iena_wb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.610 -2.000 1799.890 4.000 ;
    END
  END mprj_iena_wb
  PIN mprj_sel_o_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1531.890 -2.000 1532.170 4.000 ;
    END
  END mprj_sel_o_core[0]
  PIN mprj_sel_o_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.930 -2.000 1543.210 4.000 ;
    END
  END mprj_sel_o_core[1]
  PIN mprj_sel_o_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1553.970 -2.000 1554.250 4.000 ;
    END
  END mprj_sel_o_core[2]
  PIN mprj_sel_o_core[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.010 -2.000 1565.290 4.000 ;
    END
  END mprj_sel_o_core[3]
  PIN mprj_sel_o_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 156.000 75.810 162.000 ;
    END
  END mprj_sel_o_user[0]
  PIN mprj_sel_o_user[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 156.000 90.530 162.000 ;
    END
  END mprj_sel_o_user[1]
  PIN mprj_sel_o_user[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 156.000 105.250 162.000 ;
    END
  END mprj_sel_o_user[2]
  PIN mprj_sel_o_user[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 156.000 119.970 162.000 ;
    END
  END mprj_sel_o_user[3]
  PIN mprj_stb_o_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1518.090 -2.000 1518.370 4.000 ;
    END
  END mprj_stb_o_core
  PIN mprj_stb_o_user
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 156.000 57.410 162.000 ;
    END
  END mprj_stb_o_user
  PIN mprj_we_o_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1520.850 -2.000 1521.130 4.000 ;
    END
  END mprj_we_o_core
  PIN mprj_we_o_user
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 156.000 61.090 162.000 ;
    END
  END mprj_we_o_user
  PIN user1_vcc_powergood
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 42.880 1902.000 43.480 ;
    END
  END user1_vcc_powergood
  PIN user1_vdd_powergood
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 55.120 1902.000 55.720 ;
    END
  END user1_vdd_powergood
  PIN user2_vcc_powergood
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 67.360 1902.000 67.960 ;
    END
  END user2_vcc_powergood
  PIN user2_vdd_powergood
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 79.600 1902.000 80.200 ;
    END
  END user2_vdd_powergood
  PIN user_clock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 156.000 42.690 162.000 ;
    END
  END user_clock
  PIN user_clock2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.610 156.000 1845.890 162.000 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 91.840 1902.000 92.440 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 104.080 1902.000 104.680 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 116.320 1902.000 116.920 ;
    END
  END user_irq[2]
  PIN user_irq_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1849.290 156.000 1849.570 162.000 ;
    END
  END user_irq_core[0]
  PIN user_irq_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1852.970 156.000 1853.250 162.000 ;
    END
  END user_irq_core[1]
  PIN user_irq_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1856.650 156.000 1856.930 162.000 ;
    END
  END user_irq_core[2]
  PIN user_irq_ena[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 128.560 1902.000 129.160 ;
    END
  END user_irq_ena[0]
  PIN user_irq_ena[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 140.800 1902.000 141.400 ;
    END
  END user_irq_ena[1]
  PIN user_irq_ena[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 153.040 1902.000 153.640 ;
    END
  END user_irq_ena[2]
  PIN user_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 156.000 46.370 162.000 ;
    END
  END user_reset
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 25.070 5.200 25.970 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 100.320 5.200 101.220 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 175.570 5.200 176.470 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 250.820 5.200 251.720 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 326.070 5.200 326.970 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 401.320 5.200 402.220 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 476.570 5.200 477.470 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 551.820 5.200 552.720 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 627.070 5.200 627.970 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 702.320 5.200 703.220 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 777.570 5.200 778.470 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 852.820 5.200 853.720 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 928.070 5.200 928.970 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1003.320 5.200 1004.220 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1078.570 5.200 1079.470 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1153.820 5.200 1154.720 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1229.070 5.200 1229.970 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1304.320 5.200 1305.220 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1379.570 5.200 1380.470 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1454.820 5.200 1455.720 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1530.070 5.200 1530.970 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1605.320 5.200 1606.220 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1680.570 5.200 1681.470 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1755.820 5.200 1756.720 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1831.070 5.200 1831.970 152.560 ;
    END
  END vccd
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 706.420 5.200 707.320 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 781.670 5.200 782.570 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 856.920 5.200 857.820 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 932.170 5.200 933.070 152.560 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 334.270 5.200 335.170 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 384.270 5.200 385.170 152.560 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1279.070 5.200 1279.970 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1354.320 5.200 1355.220 152.560 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1283.070 5.200 1283.970 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.320 5.200 1359.220 152.560 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1315.970 5.200 1316.870 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1391.220 5.200 1392.120 152.560 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1319.970 5.200 1320.870 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1395.220 5.200 1396.120 152.560 ;
    END
  END vssa2
  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 61.970 5.200 62.870 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 137.220 5.200 138.120 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 212.470 5.200 213.370 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 287.720 5.200 288.620 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 362.970 5.200 363.870 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 438.220 5.200 439.120 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 513.470 5.200 514.370 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 588.720 5.200 589.620 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 663.970 5.200 664.870 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 739.220 5.200 740.120 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 814.470 5.200 815.370 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 889.720 5.200 890.620 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 964.970 5.200 965.870 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1040.220 5.200 1041.120 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1115.470 5.200 1116.370 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1190.720 5.200 1191.620 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1265.970 5.200 1266.870 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1341.220 5.200 1342.120 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1416.470 5.200 1417.370 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.720 5.200 1492.620 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1566.970 5.200 1567.870 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1642.220 5.200 1643.120 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1717.470 5.200 1718.370 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1792.720 5.200 1793.620 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1867.970 5.200 1868.870 152.560 ;
    END
  END vssd
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 743.320 5.200 744.220 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.570 5.200 819.470 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 893.820 5.200 894.720 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 969.070 5.200 969.970 152.560 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 355.170 5.200 356.070 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.170 5.200 406.070 152.560 ;
    END
  END vssd2
  OBS
      LAYER nwell ;
        RECT 5.330 148.185 1894.470 151.015 ;
        RECT 5.330 142.745 1894.470 145.575 ;
        RECT 5.330 137.305 1894.470 140.135 ;
        RECT 5.330 131.865 1894.470 134.695 ;
        RECT 5.330 126.425 1894.470 129.255 ;
        RECT 5.330 120.985 1894.470 123.815 ;
        RECT 5.330 115.545 1894.470 118.375 ;
        RECT 5.330 110.105 1894.470 112.935 ;
        RECT 5.330 104.665 1894.470 107.495 ;
        RECT 5.330 99.225 1894.470 102.055 ;
        RECT 5.330 93.785 1894.470 96.615 ;
        RECT 5.330 88.345 1894.470 91.175 ;
        RECT 5.330 82.905 1894.470 85.735 ;
        RECT 5.330 77.465 668.570 80.295 ;
        RECT 5.330 72.025 668.570 74.855 ;
        RECT 5.330 66.585 668.570 69.415 ;
        RECT 5.330 61.145 668.570 63.975 ;
        RECT 5.330 56.930 668.570 58.535 ;
        RECT 5.330 55.705 320.350 56.930 ;
        RECT 5.330 50.265 320.350 53.095 ;
        RECT 5.330 44.825 320.350 47.655 ;
        RECT 5.330 39.385 320.350 42.215 ;
        RECT 5.330 33.945 320.350 36.775 ;
        RECT 5.330 28.505 320.350 31.335 ;
        RECT 5.330 23.065 1894.470 25.895 ;
        RECT 5.330 17.625 1894.470 20.455 ;
        RECT 5.330 12.185 1894.470 15.015 ;
        RECT 5.330 6.745 1894.470 9.575 ;
      LAYER li1 ;
        RECT 5.520 5.355 1894.280 152.405 ;
      LAYER met1 ;
        RECT 131.030 160.000 711.920 160.040 ;
        RECT 724.430 160.000 738.370 160.040 ;
        RECT 5.520 0.040 1894.280 160.000 ;
      LAYER met2 ;
        RECT 25.180 155.720 42.130 159.790 ;
        RECT 42.970 155.720 45.810 159.790 ;
        RECT 46.650 155.720 49.490 159.790 ;
        RECT 50.330 155.720 53.170 159.790 ;
        RECT 54.010 155.720 56.850 159.790 ;
        RECT 57.690 155.720 60.530 159.790 ;
        RECT 61.370 155.720 64.210 159.790 ;
        RECT 65.050 155.720 67.890 159.790 ;
        RECT 68.730 155.720 71.570 159.790 ;
        RECT 72.410 155.720 75.250 159.790 ;
        RECT 76.090 155.720 78.930 159.790 ;
        RECT 79.770 155.720 82.610 159.790 ;
        RECT 83.450 155.720 86.290 159.790 ;
        RECT 87.130 155.720 89.970 159.790 ;
        RECT 90.810 155.720 93.650 159.790 ;
        RECT 94.490 155.720 97.330 159.790 ;
        RECT 98.170 155.720 101.010 159.790 ;
        RECT 101.850 155.720 104.690 159.790 ;
        RECT 105.530 155.720 108.370 159.790 ;
        RECT 109.210 155.720 112.050 159.790 ;
        RECT 112.890 155.720 115.730 159.790 ;
        RECT 116.570 155.720 119.410 159.790 ;
        RECT 120.250 155.720 123.090 159.790 ;
        RECT 123.930 155.720 126.770 159.790 ;
        RECT 127.610 155.720 130.450 159.790 ;
        RECT 131.290 155.720 134.130 159.790 ;
        RECT 134.970 155.720 137.810 159.790 ;
        RECT 138.650 155.720 141.490 159.790 ;
        RECT 142.330 155.720 145.170 159.790 ;
        RECT 146.010 155.720 148.850 159.790 ;
        RECT 149.690 155.720 152.530 159.790 ;
        RECT 153.370 155.720 156.210 159.790 ;
        RECT 157.050 155.720 159.890 159.790 ;
        RECT 160.730 155.720 163.570 159.790 ;
        RECT 164.410 155.720 167.250 159.790 ;
        RECT 168.090 155.720 170.930 159.790 ;
        RECT 171.770 155.720 174.610 159.790 ;
        RECT 175.450 155.720 178.290 159.790 ;
        RECT 179.130 155.720 181.970 159.790 ;
        RECT 182.810 155.720 185.650 159.790 ;
        RECT 186.490 155.720 189.330 159.790 ;
        RECT 190.170 155.720 193.010 159.790 ;
        RECT 193.850 155.720 196.690 159.790 ;
        RECT 197.530 155.720 200.370 159.790 ;
        RECT 201.210 155.720 204.050 159.790 ;
        RECT 204.890 155.720 207.730 159.790 ;
        RECT 208.570 155.720 211.410 159.790 ;
        RECT 212.250 155.720 215.090 159.790 ;
        RECT 215.930 155.720 218.770 159.790 ;
        RECT 219.610 155.720 222.450 159.790 ;
        RECT 223.290 155.720 226.130 159.790 ;
        RECT 226.970 155.720 229.810 159.790 ;
        RECT 230.650 155.720 233.490 159.790 ;
        RECT 234.330 155.720 237.170 159.790 ;
        RECT 238.010 155.720 240.850 159.790 ;
        RECT 241.690 155.720 244.530 159.790 ;
        RECT 245.370 155.720 248.210 159.790 ;
        RECT 249.050 155.720 251.890 159.790 ;
        RECT 252.730 155.720 255.570 159.790 ;
        RECT 256.410 155.720 259.250 159.790 ;
        RECT 260.090 155.720 262.930 159.790 ;
        RECT 263.770 155.720 266.610 159.790 ;
        RECT 267.450 155.720 270.290 159.790 ;
        RECT 271.130 155.720 273.970 159.790 ;
        RECT 274.810 155.720 277.650 159.790 ;
        RECT 278.490 155.720 281.330 159.790 ;
        RECT 282.170 155.720 285.010 159.790 ;
        RECT 285.850 155.720 288.690 159.790 ;
        RECT 289.530 155.720 292.370 159.790 ;
        RECT 293.210 155.720 296.050 159.790 ;
        RECT 296.890 155.720 299.730 159.790 ;
        RECT 300.570 155.720 303.410 159.790 ;
        RECT 304.250 155.720 307.090 159.790 ;
        RECT 307.930 155.720 310.770 159.790 ;
        RECT 311.610 155.720 314.450 159.790 ;
        RECT 315.290 155.720 318.130 159.790 ;
        RECT 318.970 155.720 321.810 159.790 ;
        RECT 322.650 155.720 325.490 159.790 ;
        RECT 326.330 155.720 329.170 159.790 ;
        RECT 330.010 155.720 332.850 159.790 ;
        RECT 333.690 155.720 336.530 159.790 ;
        RECT 337.370 155.720 340.210 159.790 ;
        RECT 341.050 155.720 343.890 159.790 ;
        RECT 344.730 155.720 347.570 159.790 ;
        RECT 348.410 155.720 351.250 159.790 ;
        RECT 352.090 155.720 354.930 159.790 ;
        RECT 355.770 155.720 358.610 159.790 ;
        RECT 359.450 155.720 362.290 159.790 ;
        RECT 363.130 155.720 365.970 159.790 ;
        RECT 366.810 155.720 369.650 159.790 ;
        RECT 370.490 155.720 373.330 159.790 ;
        RECT 374.170 155.720 377.010 159.790 ;
        RECT 377.850 155.720 380.690 159.790 ;
        RECT 381.530 155.720 384.370 159.790 ;
        RECT 385.210 155.720 388.050 159.790 ;
        RECT 388.890 155.720 391.730 159.790 ;
        RECT 392.570 155.720 395.410 159.790 ;
        RECT 396.250 155.720 399.090 159.790 ;
        RECT 399.930 155.720 402.770 159.790 ;
        RECT 403.610 155.720 406.450 159.790 ;
        RECT 407.290 155.720 410.130 159.790 ;
        RECT 410.970 155.720 413.810 159.790 ;
        RECT 414.650 155.720 417.490 159.790 ;
        RECT 418.330 155.720 421.170 159.790 ;
        RECT 422.010 155.720 424.850 159.790 ;
        RECT 425.690 155.720 428.530 159.790 ;
        RECT 429.370 155.720 432.210 159.790 ;
        RECT 433.050 155.720 435.890 159.790 ;
        RECT 436.730 155.720 439.570 159.790 ;
        RECT 440.410 155.720 443.250 159.790 ;
        RECT 444.090 155.720 446.930 159.790 ;
        RECT 447.770 155.720 450.610 159.790 ;
        RECT 451.450 155.720 454.290 159.790 ;
        RECT 455.130 155.720 457.970 159.790 ;
        RECT 458.810 155.720 461.650 159.790 ;
        RECT 462.490 155.720 465.330 159.790 ;
        RECT 466.170 155.720 469.010 159.790 ;
        RECT 469.850 155.720 472.690 159.790 ;
        RECT 473.530 155.720 476.370 159.790 ;
        RECT 477.210 155.720 480.050 159.790 ;
        RECT 480.890 155.720 483.730 159.790 ;
        RECT 484.570 155.720 487.410 159.790 ;
        RECT 488.250 155.720 491.090 159.790 ;
        RECT 491.930 155.720 494.770 159.790 ;
        RECT 495.610 155.720 498.450 159.790 ;
        RECT 499.290 155.720 502.130 159.790 ;
        RECT 502.970 155.720 505.810 159.790 ;
        RECT 506.650 155.720 509.490 159.790 ;
        RECT 510.330 155.720 513.170 159.790 ;
        RECT 514.010 155.720 516.850 159.790 ;
        RECT 517.690 155.720 520.530 159.790 ;
        RECT 521.370 155.720 524.210 159.790 ;
        RECT 525.050 155.720 527.890 159.790 ;
        RECT 528.730 155.720 531.570 159.790 ;
        RECT 532.410 155.720 535.250 159.790 ;
        RECT 536.090 155.720 538.930 159.790 ;
        RECT 539.770 155.720 542.610 159.790 ;
        RECT 543.450 155.720 546.290 159.790 ;
        RECT 547.130 155.720 549.970 159.790 ;
        RECT 550.810 155.720 553.650 159.790 ;
        RECT 554.490 155.720 557.330 159.790 ;
        RECT 558.170 155.720 561.010 159.790 ;
        RECT 561.850 155.720 564.690 159.790 ;
        RECT 565.530 155.720 568.370 159.790 ;
        RECT 569.210 155.720 572.050 159.790 ;
        RECT 572.890 155.720 575.730 159.790 ;
        RECT 576.570 155.720 579.410 159.790 ;
        RECT 580.250 155.720 583.090 159.790 ;
        RECT 583.930 155.720 586.770 159.790 ;
        RECT 587.610 155.720 590.450 159.790 ;
        RECT 591.290 155.720 594.130 159.790 ;
        RECT 594.970 155.720 597.810 159.790 ;
        RECT 598.650 155.720 601.490 159.790 ;
        RECT 602.330 155.720 605.170 159.790 ;
        RECT 606.010 155.720 608.850 159.790 ;
        RECT 609.690 155.720 612.530 159.790 ;
        RECT 613.370 155.720 616.210 159.790 ;
        RECT 617.050 155.720 619.890 159.790 ;
        RECT 620.730 155.720 623.570 159.790 ;
        RECT 624.410 155.720 627.250 159.790 ;
        RECT 628.090 155.720 630.930 159.790 ;
        RECT 631.770 155.720 634.610 159.790 ;
        RECT 635.450 155.720 638.290 159.790 ;
        RECT 639.130 155.720 641.970 159.790 ;
        RECT 642.810 155.720 645.650 159.790 ;
        RECT 646.490 155.720 649.330 159.790 ;
        RECT 650.170 155.720 653.010 159.790 ;
        RECT 653.850 155.720 656.690 159.790 ;
        RECT 657.530 155.720 660.370 159.790 ;
        RECT 661.210 155.720 664.050 159.790 ;
        RECT 664.890 155.720 667.730 159.790 ;
        RECT 668.570 155.720 671.410 159.790 ;
        RECT 672.250 155.720 675.090 159.790 ;
        RECT 675.930 155.720 678.770 159.790 ;
        RECT 679.610 155.720 682.450 159.790 ;
        RECT 683.290 155.720 686.130 159.790 ;
        RECT 686.970 155.720 689.810 159.790 ;
        RECT 690.650 155.720 693.490 159.790 ;
        RECT 694.330 155.720 697.170 159.790 ;
        RECT 698.010 155.720 700.850 159.790 ;
        RECT 701.690 155.720 704.530 159.790 ;
        RECT 705.370 155.720 708.210 159.790 ;
        RECT 709.050 155.720 711.890 159.790 ;
        RECT 712.730 155.720 715.570 159.790 ;
        RECT 716.410 155.720 719.250 159.790 ;
        RECT 720.090 155.720 722.930 159.790 ;
        RECT 723.770 155.720 726.610 159.790 ;
        RECT 727.450 155.720 730.290 159.790 ;
        RECT 731.130 155.720 733.970 159.790 ;
        RECT 734.810 155.720 737.650 159.790 ;
        RECT 738.490 155.720 741.330 159.790 ;
        RECT 742.170 155.720 745.010 159.790 ;
        RECT 745.850 155.720 748.690 159.790 ;
        RECT 749.530 155.720 752.370 159.790 ;
        RECT 753.210 155.720 756.050 159.790 ;
        RECT 756.890 155.720 759.730 159.790 ;
        RECT 760.570 155.720 763.410 159.790 ;
        RECT 764.250 155.720 767.090 159.790 ;
        RECT 767.930 155.720 770.770 159.790 ;
        RECT 771.610 155.720 774.450 159.790 ;
        RECT 775.290 155.720 778.130 159.790 ;
        RECT 778.970 155.720 781.810 159.790 ;
        RECT 782.650 155.720 785.490 159.790 ;
        RECT 786.330 155.720 789.170 159.790 ;
        RECT 790.010 155.720 792.850 159.790 ;
        RECT 793.690 155.720 796.530 159.790 ;
        RECT 797.370 155.720 800.210 159.790 ;
        RECT 801.050 155.720 803.890 159.790 ;
        RECT 804.730 155.720 807.570 159.790 ;
        RECT 808.410 155.720 811.250 159.790 ;
        RECT 812.090 155.720 814.930 159.790 ;
        RECT 815.770 155.720 818.610 159.790 ;
        RECT 819.450 155.720 822.290 159.790 ;
        RECT 823.130 155.720 825.970 159.790 ;
        RECT 826.810 155.720 829.650 159.790 ;
        RECT 830.490 155.720 833.330 159.790 ;
        RECT 834.170 155.720 837.010 159.790 ;
        RECT 837.850 155.720 840.690 159.790 ;
        RECT 841.530 155.720 844.370 159.790 ;
        RECT 845.210 155.720 848.050 159.790 ;
        RECT 848.890 155.720 851.730 159.790 ;
        RECT 852.570 155.720 855.410 159.790 ;
        RECT 856.250 155.720 859.090 159.790 ;
        RECT 859.930 155.720 862.770 159.790 ;
        RECT 863.610 155.720 866.450 159.790 ;
        RECT 867.290 155.720 870.130 159.790 ;
        RECT 870.970 155.720 873.810 159.790 ;
        RECT 874.650 155.720 877.490 159.790 ;
        RECT 878.330 155.720 881.170 159.790 ;
        RECT 882.010 155.720 884.850 159.790 ;
        RECT 885.690 155.720 888.530 159.790 ;
        RECT 889.370 155.720 892.210 159.790 ;
        RECT 893.050 155.720 895.890 159.790 ;
        RECT 896.730 155.720 899.570 159.790 ;
        RECT 900.410 155.720 903.250 159.790 ;
        RECT 904.090 155.720 906.930 159.790 ;
        RECT 907.770 155.720 910.610 159.790 ;
        RECT 911.450 155.720 914.290 159.790 ;
        RECT 915.130 155.720 917.970 159.790 ;
        RECT 918.810 155.720 921.650 159.790 ;
        RECT 922.490 155.720 925.330 159.790 ;
        RECT 926.170 155.720 929.010 159.790 ;
        RECT 929.850 155.720 932.690 159.790 ;
        RECT 933.530 155.720 936.370 159.790 ;
        RECT 937.210 155.720 940.050 159.790 ;
        RECT 940.890 155.720 943.730 159.790 ;
        RECT 944.570 155.720 947.410 159.790 ;
        RECT 948.250 155.720 951.090 159.790 ;
        RECT 951.930 155.720 954.770 159.790 ;
        RECT 955.610 155.720 958.450 159.790 ;
        RECT 959.290 155.720 962.130 159.790 ;
        RECT 962.970 155.720 965.810 159.790 ;
        RECT 966.650 155.720 969.490 159.790 ;
        RECT 970.330 155.720 973.170 159.790 ;
        RECT 974.010 155.720 976.850 159.790 ;
        RECT 977.690 155.720 980.530 159.790 ;
        RECT 981.370 155.720 984.210 159.790 ;
        RECT 985.050 155.720 987.890 159.790 ;
        RECT 988.730 155.720 991.570 159.790 ;
        RECT 992.410 155.720 995.250 159.790 ;
        RECT 996.090 155.720 998.930 159.790 ;
        RECT 999.770 155.720 1002.610 159.790 ;
        RECT 1003.450 155.720 1006.290 159.790 ;
        RECT 1007.130 155.720 1009.970 159.790 ;
        RECT 1010.810 155.720 1013.650 159.790 ;
        RECT 1014.490 155.720 1017.330 159.790 ;
        RECT 1018.170 155.720 1021.010 159.790 ;
        RECT 1021.850 155.720 1024.690 159.790 ;
        RECT 1025.530 155.720 1028.370 159.790 ;
        RECT 1029.210 155.720 1032.050 159.790 ;
        RECT 1032.890 155.720 1035.730 159.790 ;
        RECT 1036.570 155.720 1039.410 159.790 ;
        RECT 1040.250 155.720 1043.090 159.790 ;
        RECT 1043.930 155.720 1046.770 159.790 ;
        RECT 1047.610 155.720 1050.450 159.790 ;
        RECT 1051.290 155.720 1054.130 159.790 ;
        RECT 1054.970 155.720 1057.810 159.790 ;
        RECT 1058.650 155.720 1061.490 159.790 ;
        RECT 1062.330 155.720 1065.170 159.790 ;
        RECT 1066.010 155.720 1068.850 159.790 ;
        RECT 1069.690 155.720 1072.530 159.790 ;
        RECT 1073.370 155.720 1076.210 159.790 ;
        RECT 1077.050 155.720 1079.890 159.790 ;
        RECT 1080.730 155.720 1083.570 159.790 ;
        RECT 1084.410 155.720 1087.250 159.790 ;
        RECT 1088.090 155.720 1090.930 159.790 ;
        RECT 1091.770 155.720 1094.610 159.790 ;
        RECT 1095.450 155.720 1098.290 159.790 ;
        RECT 1099.130 155.720 1101.970 159.790 ;
        RECT 1102.810 155.720 1105.650 159.790 ;
        RECT 1106.490 155.720 1109.330 159.790 ;
        RECT 1110.170 155.720 1113.010 159.790 ;
        RECT 1113.850 155.720 1116.690 159.790 ;
        RECT 1117.530 155.720 1120.370 159.790 ;
        RECT 1121.210 155.720 1124.050 159.790 ;
        RECT 1124.890 155.720 1127.730 159.790 ;
        RECT 1128.570 155.720 1131.410 159.790 ;
        RECT 1132.250 155.720 1135.090 159.790 ;
        RECT 1135.930 155.720 1138.770 159.790 ;
        RECT 1139.610 155.720 1142.450 159.790 ;
        RECT 1143.290 155.720 1146.130 159.790 ;
        RECT 1146.970 155.720 1149.810 159.790 ;
        RECT 1150.650 155.720 1153.490 159.790 ;
        RECT 1154.330 155.720 1157.170 159.790 ;
        RECT 1158.010 155.720 1160.850 159.790 ;
        RECT 1161.690 155.720 1164.530 159.790 ;
        RECT 1165.370 155.720 1168.210 159.790 ;
        RECT 1169.050 155.720 1171.890 159.790 ;
        RECT 1172.730 155.720 1175.570 159.790 ;
        RECT 1176.410 155.720 1179.250 159.790 ;
        RECT 1180.090 155.720 1182.930 159.790 ;
        RECT 1183.770 155.720 1186.610 159.790 ;
        RECT 1187.450 155.720 1190.290 159.790 ;
        RECT 1191.130 155.720 1193.970 159.790 ;
        RECT 1194.810 155.720 1197.650 159.790 ;
        RECT 1198.490 155.720 1201.330 159.790 ;
        RECT 1202.170 155.720 1205.010 159.790 ;
        RECT 1205.850 155.720 1208.690 159.790 ;
        RECT 1209.530 155.720 1212.370 159.790 ;
        RECT 1213.210 155.720 1216.050 159.790 ;
        RECT 1216.890 155.720 1219.730 159.790 ;
        RECT 1220.570 155.720 1223.410 159.790 ;
        RECT 1224.250 155.720 1227.090 159.790 ;
        RECT 1227.930 155.720 1230.770 159.790 ;
        RECT 1231.610 155.720 1234.450 159.790 ;
        RECT 1235.290 155.720 1238.130 159.790 ;
        RECT 1238.970 155.720 1241.810 159.790 ;
        RECT 1242.650 155.720 1245.490 159.790 ;
        RECT 1246.330 155.720 1249.170 159.790 ;
        RECT 1250.010 155.720 1252.850 159.790 ;
        RECT 1253.690 155.720 1256.530 159.790 ;
        RECT 1257.370 155.720 1260.210 159.790 ;
        RECT 1261.050 155.720 1263.890 159.790 ;
        RECT 1264.730 155.720 1267.570 159.790 ;
        RECT 1268.410 155.720 1271.250 159.790 ;
        RECT 1272.090 155.720 1274.930 159.790 ;
        RECT 1275.770 155.720 1278.610 159.790 ;
        RECT 1279.450 155.720 1282.290 159.790 ;
        RECT 1283.130 155.720 1285.970 159.790 ;
        RECT 1286.810 155.720 1289.650 159.790 ;
        RECT 1290.490 155.720 1293.330 159.790 ;
        RECT 1294.170 155.720 1297.010 159.790 ;
        RECT 1297.850 155.720 1300.690 159.790 ;
        RECT 1301.530 155.720 1304.370 159.790 ;
        RECT 1305.210 155.720 1308.050 159.790 ;
        RECT 1308.890 155.720 1311.730 159.790 ;
        RECT 1312.570 155.720 1315.410 159.790 ;
        RECT 1316.250 155.720 1319.090 159.790 ;
        RECT 1319.930 155.720 1322.770 159.790 ;
        RECT 1323.610 155.720 1326.450 159.790 ;
        RECT 1327.290 155.720 1330.130 159.790 ;
        RECT 1330.970 155.720 1333.810 159.790 ;
        RECT 1334.650 155.720 1337.490 159.790 ;
        RECT 1338.330 155.720 1341.170 159.790 ;
        RECT 1342.010 155.720 1344.850 159.790 ;
        RECT 1345.690 155.720 1348.530 159.790 ;
        RECT 1349.370 155.720 1352.210 159.790 ;
        RECT 1353.050 155.720 1355.890 159.790 ;
        RECT 1356.730 155.720 1359.570 159.790 ;
        RECT 1360.410 155.720 1363.250 159.790 ;
        RECT 1364.090 155.720 1366.930 159.790 ;
        RECT 1367.770 155.720 1370.610 159.790 ;
        RECT 1371.450 155.720 1374.290 159.790 ;
        RECT 1375.130 155.720 1377.970 159.790 ;
        RECT 1378.810 155.720 1381.650 159.790 ;
        RECT 1382.490 155.720 1385.330 159.790 ;
        RECT 1386.170 155.720 1389.010 159.790 ;
        RECT 1389.850 155.720 1392.690 159.790 ;
        RECT 1393.530 155.720 1396.370 159.790 ;
        RECT 1397.210 155.720 1400.050 159.790 ;
        RECT 1400.890 155.720 1403.730 159.790 ;
        RECT 1404.570 155.720 1407.410 159.790 ;
        RECT 1408.250 155.720 1411.090 159.790 ;
        RECT 1411.930 155.720 1414.770 159.790 ;
        RECT 1415.610 155.720 1418.450 159.790 ;
        RECT 1419.290 155.720 1422.130 159.790 ;
        RECT 1422.970 155.720 1425.810 159.790 ;
        RECT 1426.650 155.720 1429.490 159.790 ;
        RECT 1430.330 155.720 1433.170 159.790 ;
        RECT 1434.010 155.720 1436.850 159.790 ;
        RECT 1437.690 155.720 1440.530 159.790 ;
        RECT 1441.370 155.720 1444.210 159.790 ;
        RECT 1445.050 155.720 1447.890 159.790 ;
        RECT 1448.730 155.720 1451.570 159.790 ;
        RECT 1452.410 155.720 1455.250 159.790 ;
        RECT 1456.090 155.720 1458.930 159.790 ;
        RECT 1459.770 155.720 1462.610 159.790 ;
        RECT 1463.450 155.720 1466.290 159.790 ;
        RECT 1467.130 155.720 1469.970 159.790 ;
        RECT 1470.810 155.720 1473.650 159.790 ;
        RECT 1474.490 155.720 1477.330 159.790 ;
        RECT 1478.170 155.720 1481.010 159.790 ;
        RECT 1481.850 155.720 1484.690 159.790 ;
        RECT 1485.530 155.720 1488.370 159.790 ;
        RECT 1489.210 155.720 1492.050 159.790 ;
        RECT 1492.890 155.720 1495.730 159.790 ;
        RECT 1496.570 155.720 1499.410 159.790 ;
        RECT 1500.250 155.720 1503.090 159.790 ;
        RECT 1503.930 155.720 1506.770 159.790 ;
        RECT 1507.610 155.720 1510.450 159.790 ;
        RECT 1511.290 155.720 1514.130 159.790 ;
        RECT 1514.970 155.720 1517.810 159.790 ;
        RECT 1518.650 155.720 1521.490 159.790 ;
        RECT 1522.330 155.720 1525.170 159.790 ;
        RECT 1526.010 155.720 1528.850 159.790 ;
        RECT 1529.690 155.720 1532.530 159.790 ;
        RECT 1533.370 155.720 1536.210 159.790 ;
        RECT 1537.050 155.720 1539.890 159.790 ;
        RECT 1540.730 155.720 1543.570 159.790 ;
        RECT 1544.410 155.720 1547.250 159.790 ;
        RECT 1548.090 155.720 1550.930 159.790 ;
        RECT 1551.770 155.720 1554.610 159.790 ;
        RECT 1555.450 155.720 1558.290 159.790 ;
        RECT 1559.130 155.720 1561.970 159.790 ;
        RECT 1562.810 155.720 1565.650 159.790 ;
        RECT 1566.490 155.720 1569.330 159.790 ;
        RECT 1570.170 155.720 1573.010 159.790 ;
        RECT 1573.850 155.720 1576.690 159.790 ;
        RECT 1577.530 155.720 1580.370 159.790 ;
        RECT 1581.210 155.720 1584.050 159.790 ;
        RECT 1584.890 155.720 1587.730 159.790 ;
        RECT 1588.570 155.720 1591.410 159.790 ;
        RECT 1592.250 155.720 1595.090 159.790 ;
        RECT 1595.930 155.720 1598.770 159.790 ;
        RECT 1599.610 155.720 1602.450 159.790 ;
        RECT 1603.290 155.720 1606.130 159.790 ;
        RECT 1606.970 155.720 1609.810 159.790 ;
        RECT 1610.650 155.720 1613.490 159.790 ;
        RECT 1614.330 155.720 1617.170 159.790 ;
        RECT 1618.010 155.720 1620.850 159.790 ;
        RECT 1621.690 155.720 1624.530 159.790 ;
        RECT 1625.370 155.720 1628.210 159.790 ;
        RECT 1629.050 155.720 1631.890 159.790 ;
        RECT 1632.730 155.720 1635.570 159.790 ;
        RECT 1636.410 155.720 1639.250 159.790 ;
        RECT 1640.090 155.720 1642.930 159.790 ;
        RECT 1643.770 155.720 1646.610 159.790 ;
        RECT 1647.450 155.720 1650.290 159.790 ;
        RECT 1651.130 155.720 1653.970 159.790 ;
        RECT 1654.810 155.720 1657.650 159.790 ;
        RECT 1658.490 155.720 1661.330 159.790 ;
        RECT 1662.170 155.720 1665.010 159.790 ;
        RECT 1665.850 155.720 1668.690 159.790 ;
        RECT 1669.530 155.720 1672.370 159.790 ;
        RECT 1673.210 155.720 1676.050 159.790 ;
        RECT 1676.890 155.720 1679.730 159.790 ;
        RECT 1680.570 155.720 1683.410 159.790 ;
        RECT 1684.250 155.720 1687.090 159.790 ;
        RECT 1687.930 155.720 1690.770 159.790 ;
        RECT 1691.610 155.720 1694.450 159.790 ;
        RECT 1695.290 155.720 1698.130 159.790 ;
        RECT 1698.970 155.720 1701.810 159.790 ;
        RECT 1702.650 155.720 1705.490 159.790 ;
        RECT 1706.330 155.720 1709.170 159.790 ;
        RECT 1710.010 155.720 1712.850 159.790 ;
        RECT 1713.690 155.720 1716.530 159.790 ;
        RECT 1717.370 155.720 1720.210 159.790 ;
        RECT 1721.050 155.720 1723.890 159.790 ;
        RECT 1724.730 155.720 1727.570 159.790 ;
        RECT 1728.410 155.720 1731.250 159.790 ;
        RECT 1732.090 155.720 1734.930 159.790 ;
        RECT 1735.770 155.720 1738.610 159.790 ;
        RECT 1739.450 155.720 1742.290 159.790 ;
        RECT 1743.130 155.720 1745.970 159.790 ;
        RECT 1746.810 155.720 1749.650 159.790 ;
        RECT 1750.490 155.720 1753.330 159.790 ;
        RECT 1754.170 155.720 1757.010 159.790 ;
        RECT 1757.850 155.720 1760.690 159.790 ;
        RECT 1761.530 155.720 1764.370 159.790 ;
        RECT 1765.210 155.720 1768.050 159.790 ;
        RECT 1768.890 155.720 1771.730 159.790 ;
        RECT 1772.570 155.720 1775.410 159.790 ;
        RECT 1776.250 155.720 1779.090 159.790 ;
        RECT 1779.930 155.720 1782.770 159.790 ;
        RECT 1783.610 155.720 1786.450 159.790 ;
        RECT 1787.290 155.720 1790.130 159.790 ;
        RECT 1790.970 155.720 1793.810 159.790 ;
        RECT 1794.650 155.720 1797.490 159.790 ;
        RECT 1798.330 155.720 1801.170 159.790 ;
        RECT 1802.010 155.720 1804.850 159.790 ;
        RECT 1805.690 155.720 1808.530 159.790 ;
        RECT 1809.370 155.720 1812.210 159.790 ;
        RECT 1813.050 155.720 1815.890 159.790 ;
        RECT 1816.730 155.720 1819.570 159.790 ;
        RECT 1820.410 155.720 1823.250 159.790 ;
        RECT 1824.090 155.720 1826.930 159.790 ;
        RECT 1827.770 155.720 1830.610 159.790 ;
        RECT 1831.450 155.720 1834.290 159.790 ;
        RECT 1835.130 155.720 1837.970 159.790 ;
        RECT 1838.810 155.720 1841.650 159.790 ;
        RECT 1842.490 155.720 1845.330 159.790 ;
        RECT 1846.170 155.720 1849.010 159.790 ;
        RECT 1849.850 155.720 1852.690 159.790 ;
        RECT 1853.530 155.720 1856.370 159.790 ;
        RECT 1857.210 155.720 1891.890 159.790 ;
        RECT 25.180 4.280 1891.890 155.720 ;
        RECT 25.180 0.010 99.170 4.280 ;
        RECT 100.010 0.010 101.930 4.280 ;
        RECT 102.770 0.010 104.690 4.280 ;
        RECT 105.530 0.010 107.450 4.280 ;
        RECT 108.290 0.010 110.210 4.280 ;
        RECT 111.050 0.010 112.970 4.280 ;
        RECT 113.810 0.010 115.730 4.280 ;
        RECT 116.570 0.010 118.490 4.280 ;
        RECT 119.330 0.010 121.250 4.280 ;
        RECT 122.090 0.010 124.010 4.280 ;
        RECT 124.850 0.010 126.770 4.280 ;
        RECT 127.610 0.010 129.530 4.280 ;
        RECT 130.370 0.010 132.290 4.280 ;
        RECT 133.130 0.010 135.050 4.280 ;
        RECT 135.890 0.010 137.810 4.280 ;
        RECT 138.650 0.010 140.570 4.280 ;
        RECT 141.410 0.010 143.330 4.280 ;
        RECT 144.170 0.010 146.090 4.280 ;
        RECT 146.930 0.010 148.850 4.280 ;
        RECT 149.690 0.010 151.610 4.280 ;
        RECT 152.450 0.010 154.370 4.280 ;
        RECT 155.210 0.010 157.130 4.280 ;
        RECT 157.970 0.010 159.890 4.280 ;
        RECT 160.730 0.010 162.650 4.280 ;
        RECT 163.490 0.010 165.410 4.280 ;
        RECT 166.250 0.010 168.170 4.280 ;
        RECT 169.010 0.010 170.930 4.280 ;
        RECT 171.770 0.010 173.690 4.280 ;
        RECT 174.530 0.010 176.450 4.280 ;
        RECT 177.290 0.010 179.210 4.280 ;
        RECT 180.050 0.010 181.970 4.280 ;
        RECT 182.810 0.010 184.730 4.280 ;
        RECT 185.570 0.010 187.490 4.280 ;
        RECT 188.330 0.010 190.250 4.280 ;
        RECT 191.090 0.010 193.010 4.280 ;
        RECT 193.850 0.010 195.770 4.280 ;
        RECT 196.610 0.010 198.530 4.280 ;
        RECT 199.370 0.010 201.290 4.280 ;
        RECT 202.130 0.010 204.050 4.280 ;
        RECT 204.890 0.010 206.810 4.280 ;
        RECT 207.650 0.010 209.570 4.280 ;
        RECT 210.410 0.010 212.330 4.280 ;
        RECT 213.170 0.010 215.090 4.280 ;
        RECT 215.930 0.010 217.850 4.280 ;
        RECT 218.690 0.010 220.610 4.280 ;
        RECT 221.450 0.010 223.370 4.280 ;
        RECT 224.210 0.010 226.130 4.280 ;
        RECT 226.970 0.010 228.890 4.280 ;
        RECT 229.730 0.010 231.650 4.280 ;
        RECT 232.490 0.010 234.410 4.280 ;
        RECT 235.250 0.010 237.170 4.280 ;
        RECT 238.010 0.010 239.930 4.280 ;
        RECT 240.770 0.010 242.690 4.280 ;
        RECT 243.530 0.010 245.450 4.280 ;
        RECT 246.290 0.010 248.210 4.280 ;
        RECT 249.050 0.010 250.970 4.280 ;
        RECT 251.810 0.010 253.730 4.280 ;
        RECT 254.570 0.010 256.490 4.280 ;
        RECT 257.330 0.010 259.250 4.280 ;
        RECT 260.090 0.010 262.010 4.280 ;
        RECT 262.850 0.010 264.770 4.280 ;
        RECT 265.610 0.010 267.530 4.280 ;
        RECT 268.370 0.010 270.290 4.280 ;
        RECT 271.130 0.010 273.050 4.280 ;
        RECT 273.890 0.010 275.810 4.280 ;
        RECT 276.650 0.010 278.570 4.280 ;
        RECT 279.410 0.010 281.330 4.280 ;
        RECT 282.170 0.010 284.090 4.280 ;
        RECT 284.930 0.010 286.850 4.280 ;
        RECT 287.690 0.010 289.610 4.280 ;
        RECT 290.450 0.010 292.370 4.280 ;
        RECT 293.210 0.010 295.130 4.280 ;
        RECT 295.970 0.010 297.890 4.280 ;
        RECT 298.730 0.010 300.650 4.280 ;
        RECT 301.490 0.010 303.410 4.280 ;
        RECT 304.250 0.010 306.170 4.280 ;
        RECT 307.010 0.010 308.930 4.280 ;
        RECT 309.770 0.010 311.690 4.280 ;
        RECT 312.530 0.010 314.450 4.280 ;
        RECT 315.290 0.010 317.210 4.280 ;
        RECT 318.050 0.010 319.970 4.280 ;
        RECT 320.810 0.010 322.730 4.280 ;
        RECT 323.570 0.010 325.490 4.280 ;
        RECT 326.330 0.010 328.250 4.280 ;
        RECT 329.090 0.010 331.010 4.280 ;
        RECT 331.850 0.010 333.770 4.280 ;
        RECT 334.610 0.010 336.530 4.280 ;
        RECT 337.370 0.010 339.290 4.280 ;
        RECT 340.130 0.010 342.050 4.280 ;
        RECT 342.890 0.010 344.810 4.280 ;
        RECT 345.650 0.010 347.570 4.280 ;
        RECT 348.410 0.010 350.330 4.280 ;
        RECT 351.170 0.010 353.090 4.280 ;
        RECT 353.930 0.010 355.850 4.280 ;
        RECT 356.690 0.010 358.610 4.280 ;
        RECT 359.450 0.010 361.370 4.280 ;
        RECT 362.210 0.010 364.130 4.280 ;
        RECT 364.970 0.010 366.890 4.280 ;
        RECT 367.730 0.010 369.650 4.280 ;
        RECT 370.490 0.010 372.410 4.280 ;
        RECT 373.250 0.010 375.170 4.280 ;
        RECT 376.010 0.010 377.930 4.280 ;
        RECT 378.770 0.010 380.690 4.280 ;
        RECT 381.530 0.010 383.450 4.280 ;
        RECT 384.290 0.010 386.210 4.280 ;
        RECT 387.050 0.010 388.970 4.280 ;
        RECT 389.810 0.010 391.730 4.280 ;
        RECT 392.570 0.010 394.490 4.280 ;
        RECT 395.330 0.010 397.250 4.280 ;
        RECT 398.090 0.010 400.010 4.280 ;
        RECT 400.850 0.010 402.770 4.280 ;
        RECT 403.610 0.010 405.530 4.280 ;
        RECT 406.370 0.010 408.290 4.280 ;
        RECT 409.130 0.010 411.050 4.280 ;
        RECT 411.890 0.010 413.810 4.280 ;
        RECT 414.650 0.010 416.570 4.280 ;
        RECT 417.410 0.010 419.330 4.280 ;
        RECT 420.170 0.010 422.090 4.280 ;
        RECT 422.930 0.010 424.850 4.280 ;
        RECT 425.690 0.010 427.610 4.280 ;
        RECT 428.450 0.010 430.370 4.280 ;
        RECT 431.210 0.010 433.130 4.280 ;
        RECT 433.970 0.010 435.890 4.280 ;
        RECT 436.730 0.010 438.650 4.280 ;
        RECT 439.490 0.010 441.410 4.280 ;
        RECT 442.250 0.010 444.170 4.280 ;
        RECT 445.010 0.010 446.930 4.280 ;
        RECT 447.770 0.010 449.690 4.280 ;
        RECT 450.530 0.010 452.450 4.280 ;
        RECT 453.290 0.010 455.210 4.280 ;
        RECT 456.050 0.010 457.970 4.280 ;
        RECT 458.810 0.010 460.730 4.280 ;
        RECT 461.570 0.010 463.490 4.280 ;
        RECT 464.330 0.010 466.250 4.280 ;
        RECT 467.090 0.010 469.010 4.280 ;
        RECT 469.850 0.010 471.770 4.280 ;
        RECT 472.610 0.010 474.530 4.280 ;
        RECT 475.370 0.010 477.290 4.280 ;
        RECT 478.130 0.010 480.050 4.280 ;
        RECT 480.890 0.010 482.810 4.280 ;
        RECT 483.650 0.010 485.570 4.280 ;
        RECT 486.410 0.010 488.330 4.280 ;
        RECT 489.170 0.010 491.090 4.280 ;
        RECT 491.930 0.010 493.850 4.280 ;
        RECT 494.690 0.010 496.610 4.280 ;
        RECT 497.450 0.010 499.370 4.280 ;
        RECT 500.210 0.010 502.130 4.280 ;
        RECT 502.970 0.010 504.890 4.280 ;
        RECT 505.730 0.010 507.650 4.280 ;
        RECT 508.490 0.010 510.410 4.280 ;
        RECT 511.250 0.010 513.170 4.280 ;
        RECT 514.010 0.010 515.930 4.280 ;
        RECT 516.770 0.010 518.690 4.280 ;
        RECT 519.530 0.010 521.450 4.280 ;
        RECT 522.290 0.010 524.210 4.280 ;
        RECT 525.050 0.010 526.970 4.280 ;
        RECT 527.810 0.010 529.730 4.280 ;
        RECT 530.570 0.010 532.490 4.280 ;
        RECT 533.330 0.010 535.250 4.280 ;
        RECT 536.090 0.010 538.010 4.280 ;
        RECT 538.850 0.010 540.770 4.280 ;
        RECT 541.610 0.010 543.530 4.280 ;
        RECT 544.370 0.010 546.290 4.280 ;
        RECT 547.130 0.010 549.050 4.280 ;
        RECT 549.890 0.010 551.810 4.280 ;
        RECT 552.650 0.010 554.570 4.280 ;
        RECT 555.410 0.010 557.330 4.280 ;
        RECT 558.170 0.010 560.090 4.280 ;
        RECT 560.930 0.010 562.850 4.280 ;
        RECT 563.690 0.010 565.610 4.280 ;
        RECT 566.450 0.010 568.370 4.280 ;
        RECT 569.210 0.010 571.130 4.280 ;
        RECT 571.970 0.010 573.890 4.280 ;
        RECT 574.730 0.010 576.650 4.280 ;
        RECT 577.490 0.010 579.410 4.280 ;
        RECT 580.250 0.010 582.170 4.280 ;
        RECT 583.010 0.010 584.930 4.280 ;
        RECT 585.770 0.010 587.690 4.280 ;
        RECT 588.530 0.010 590.450 4.280 ;
        RECT 591.290 0.010 593.210 4.280 ;
        RECT 594.050 0.010 595.970 4.280 ;
        RECT 596.810 0.010 598.730 4.280 ;
        RECT 599.570 0.010 601.490 4.280 ;
        RECT 602.330 0.010 604.250 4.280 ;
        RECT 605.090 0.010 607.010 4.280 ;
        RECT 607.850 0.010 609.770 4.280 ;
        RECT 610.610 0.010 612.530 4.280 ;
        RECT 613.370 0.010 615.290 4.280 ;
        RECT 616.130 0.010 618.050 4.280 ;
        RECT 618.890 0.010 620.810 4.280 ;
        RECT 621.650 0.010 623.570 4.280 ;
        RECT 624.410 0.010 626.330 4.280 ;
        RECT 627.170 0.010 629.090 4.280 ;
        RECT 629.930 0.010 631.850 4.280 ;
        RECT 632.690 0.010 634.610 4.280 ;
        RECT 635.450 0.010 637.370 4.280 ;
        RECT 638.210 0.010 640.130 4.280 ;
        RECT 640.970 0.010 642.890 4.280 ;
        RECT 643.730 0.010 645.650 4.280 ;
        RECT 646.490 0.010 648.410 4.280 ;
        RECT 649.250 0.010 651.170 4.280 ;
        RECT 652.010 0.010 653.930 4.280 ;
        RECT 654.770 0.010 656.690 4.280 ;
        RECT 657.530 0.010 659.450 4.280 ;
        RECT 660.290 0.010 662.210 4.280 ;
        RECT 663.050 0.010 664.970 4.280 ;
        RECT 665.810 0.010 667.730 4.280 ;
        RECT 668.570 0.010 670.490 4.280 ;
        RECT 671.330 0.010 673.250 4.280 ;
        RECT 674.090 0.010 676.010 4.280 ;
        RECT 676.850 0.010 678.770 4.280 ;
        RECT 679.610 0.010 681.530 4.280 ;
        RECT 682.370 0.010 684.290 4.280 ;
        RECT 685.130 0.010 687.050 4.280 ;
        RECT 687.890 0.010 689.810 4.280 ;
        RECT 690.650 0.010 692.570 4.280 ;
        RECT 693.410 0.010 695.330 4.280 ;
        RECT 696.170 0.010 698.090 4.280 ;
        RECT 698.930 0.010 700.850 4.280 ;
        RECT 701.690 0.010 703.610 4.280 ;
        RECT 704.450 0.010 706.370 4.280 ;
        RECT 707.210 0.010 709.130 4.280 ;
        RECT 709.970 0.010 711.890 4.280 ;
        RECT 712.730 0.010 714.650 4.280 ;
        RECT 715.490 0.010 717.410 4.280 ;
        RECT 718.250 0.010 720.170 4.280 ;
        RECT 721.010 0.010 722.930 4.280 ;
        RECT 723.770 0.010 725.690 4.280 ;
        RECT 726.530 0.010 728.450 4.280 ;
        RECT 729.290 0.010 731.210 4.280 ;
        RECT 732.050 0.010 733.970 4.280 ;
        RECT 734.810 0.010 736.730 4.280 ;
        RECT 737.570 0.010 739.490 4.280 ;
        RECT 740.330 0.010 742.250 4.280 ;
        RECT 743.090 0.010 745.010 4.280 ;
        RECT 745.850 0.010 747.770 4.280 ;
        RECT 748.610 0.010 750.530 4.280 ;
        RECT 751.370 0.010 753.290 4.280 ;
        RECT 754.130 0.010 756.050 4.280 ;
        RECT 756.890 0.010 758.810 4.280 ;
        RECT 759.650 0.010 761.570 4.280 ;
        RECT 762.410 0.010 764.330 4.280 ;
        RECT 765.170 0.010 767.090 4.280 ;
        RECT 767.930 0.010 769.850 4.280 ;
        RECT 770.690 0.010 772.610 4.280 ;
        RECT 773.450 0.010 775.370 4.280 ;
        RECT 776.210 0.010 778.130 4.280 ;
        RECT 778.970 0.010 780.890 4.280 ;
        RECT 781.730 0.010 783.650 4.280 ;
        RECT 784.490 0.010 786.410 4.280 ;
        RECT 787.250 0.010 789.170 4.280 ;
        RECT 790.010 0.010 791.930 4.280 ;
        RECT 792.770 0.010 794.690 4.280 ;
        RECT 795.530 0.010 797.450 4.280 ;
        RECT 798.290 0.010 800.210 4.280 ;
        RECT 801.050 0.010 802.970 4.280 ;
        RECT 803.810 0.010 805.730 4.280 ;
        RECT 806.570 0.010 808.490 4.280 ;
        RECT 809.330 0.010 811.250 4.280 ;
        RECT 812.090 0.010 814.010 4.280 ;
        RECT 814.850 0.010 816.770 4.280 ;
        RECT 817.610 0.010 819.530 4.280 ;
        RECT 820.370 0.010 822.290 4.280 ;
        RECT 823.130 0.010 825.050 4.280 ;
        RECT 825.890 0.010 827.810 4.280 ;
        RECT 828.650 0.010 830.570 4.280 ;
        RECT 831.410 0.010 833.330 4.280 ;
        RECT 834.170 0.010 836.090 4.280 ;
        RECT 836.930 0.010 838.850 4.280 ;
        RECT 839.690 0.010 841.610 4.280 ;
        RECT 842.450 0.010 844.370 4.280 ;
        RECT 845.210 0.010 847.130 4.280 ;
        RECT 847.970 0.010 849.890 4.280 ;
        RECT 850.730 0.010 852.650 4.280 ;
        RECT 853.490 0.010 855.410 4.280 ;
        RECT 856.250 0.010 858.170 4.280 ;
        RECT 859.010 0.010 860.930 4.280 ;
        RECT 861.770 0.010 863.690 4.280 ;
        RECT 864.530 0.010 866.450 4.280 ;
        RECT 867.290 0.010 869.210 4.280 ;
        RECT 870.050 0.010 871.970 4.280 ;
        RECT 872.810 0.010 874.730 4.280 ;
        RECT 875.570 0.010 877.490 4.280 ;
        RECT 878.330 0.010 880.250 4.280 ;
        RECT 881.090 0.010 883.010 4.280 ;
        RECT 883.850 0.010 885.770 4.280 ;
        RECT 886.610 0.010 888.530 4.280 ;
        RECT 889.370 0.010 891.290 4.280 ;
        RECT 892.130 0.010 894.050 4.280 ;
        RECT 894.890 0.010 896.810 4.280 ;
        RECT 897.650 0.010 899.570 4.280 ;
        RECT 900.410 0.010 902.330 4.280 ;
        RECT 903.170 0.010 905.090 4.280 ;
        RECT 905.930 0.010 907.850 4.280 ;
        RECT 908.690 0.010 910.610 4.280 ;
        RECT 911.450 0.010 913.370 4.280 ;
        RECT 914.210 0.010 916.130 4.280 ;
        RECT 916.970 0.010 918.890 4.280 ;
        RECT 919.730 0.010 921.650 4.280 ;
        RECT 922.490 0.010 924.410 4.280 ;
        RECT 925.250 0.010 927.170 4.280 ;
        RECT 928.010 0.010 929.930 4.280 ;
        RECT 930.770 0.010 932.690 4.280 ;
        RECT 933.530 0.010 935.450 4.280 ;
        RECT 936.290 0.010 938.210 4.280 ;
        RECT 939.050 0.010 940.970 4.280 ;
        RECT 941.810 0.010 943.730 4.280 ;
        RECT 944.570 0.010 946.490 4.280 ;
        RECT 947.330 0.010 949.250 4.280 ;
        RECT 950.090 0.010 952.010 4.280 ;
        RECT 952.850 0.010 954.770 4.280 ;
        RECT 955.610 0.010 957.530 4.280 ;
        RECT 958.370 0.010 960.290 4.280 ;
        RECT 961.130 0.010 963.050 4.280 ;
        RECT 963.890 0.010 965.810 4.280 ;
        RECT 966.650 0.010 968.570 4.280 ;
        RECT 969.410 0.010 971.330 4.280 ;
        RECT 972.170 0.010 974.090 4.280 ;
        RECT 974.930 0.010 976.850 4.280 ;
        RECT 977.690 0.010 979.610 4.280 ;
        RECT 980.450 0.010 982.370 4.280 ;
        RECT 983.210 0.010 985.130 4.280 ;
        RECT 985.970 0.010 987.890 4.280 ;
        RECT 988.730 0.010 990.650 4.280 ;
        RECT 991.490 0.010 993.410 4.280 ;
        RECT 994.250 0.010 996.170 4.280 ;
        RECT 997.010 0.010 998.930 4.280 ;
        RECT 999.770 0.010 1001.690 4.280 ;
        RECT 1002.530 0.010 1004.450 4.280 ;
        RECT 1005.290 0.010 1007.210 4.280 ;
        RECT 1008.050 0.010 1009.970 4.280 ;
        RECT 1010.810 0.010 1012.730 4.280 ;
        RECT 1013.570 0.010 1015.490 4.280 ;
        RECT 1016.330 0.010 1018.250 4.280 ;
        RECT 1019.090 0.010 1021.010 4.280 ;
        RECT 1021.850 0.010 1023.770 4.280 ;
        RECT 1024.610 0.010 1026.530 4.280 ;
        RECT 1027.370 0.010 1029.290 4.280 ;
        RECT 1030.130 0.010 1032.050 4.280 ;
        RECT 1032.890 0.010 1034.810 4.280 ;
        RECT 1035.650 0.010 1037.570 4.280 ;
        RECT 1038.410 0.010 1040.330 4.280 ;
        RECT 1041.170 0.010 1043.090 4.280 ;
        RECT 1043.930 0.010 1045.850 4.280 ;
        RECT 1046.690 0.010 1048.610 4.280 ;
        RECT 1049.450 0.010 1051.370 4.280 ;
        RECT 1052.210 0.010 1054.130 4.280 ;
        RECT 1054.970 0.010 1056.890 4.280 ;
        RECT 1057.730 0.010 1059.650 4.280 ;
        RECT 1060.490 0.010 1062.410 4.280 ;
        RECT 1063.250 0.010 1065.170 4.280 ;
        RECT 1066.010 0.010 1067.930 4.280 ;
        RECT 1068.770 0.010 1070.690 4.280 ;
        RECT 1071.530 0.010 1073.450 4.280 ;
        RECT 1074.290 0.010 1076.210 4.280 ;
        RECT 1077.050 0.010 1078.970 4.280 ;
        RECT 1079.810 0.010 1081.730 4.280 ;
        RECT 1082.570 0.010 1084.490 4.280 ;
        RECT 1085.330 0.010 1087.250 4.280 ;
        RECT 1088.090 0.010 1090.010 4.280 ;
        RECT 1090.850 0.010 1092.770 4.280 ;
        RECT 1093.610 0.010 1095.530 4.280 ;
        RECT 1096.370 0.010 1098.290 4.280 ;
        RECT 1099.130 0.010 1101.050 4.280 ;
        RECT 1101.890 0.010 1103.810 4.280 ;
        RECT 1104.650 0.010 1106.570 4.280 ;
        RECT 1107.410 0.010 1109.330 4.280 ;
        RECT 1110.170 0.010 1112.090 4.280 ;
        RECT 1112.930 0.010 1114.850 4.280 ;
        RECT 1115.690 0.010 1117.610 4.280 ;
        RECT 1118.450 0.010 1120.370 4.280 ;
        RECT 1121.210 0.010 1123.130 4.280 ;
        RECT 1123.970 0.010 1125.890 4.280 ;
        RECT 1126.730 0.010 1128.650 4.280 ;
        RECT 1129.490 0.010 1131.410 4.280 ;
        RECT 1132.250 0.010 1134.170 4.280 ;
        RECT 1135.010 0.010 1136.930 4.280 ;
        RECT 1137.770 0.010 1139.690 4.280 ;
        RECT 1140.530 0.010 1142.450 4.280 ;
        RECT 1143.290 0.010 1145.210 4.280 ;
        RECT 1146.050 0.010 1147.970 4.280 ;
        RECT 1148.810 0.010 1150.730 4.280 ;
        RECT 1151.570 0.010 1153.490 4.280 ;
        RECT 1154.330 0.010 1156.250 4.280 ;
        RECT 1157.090 0.010 1159.010 4.280 ;
        RECT 1159.850 0.010 1161.770 4.280 ;
        RECT 1162.610 0.010 1164.530 4.280 ;
        RECT 1165.370 0.010 1167.290 4.280 ;
        RECT 1168.130 0.010 1170.050 4.280 ;
        RECT 1170.890 0.010 1172.810 4.280 ;
        RECT 1173.650 0.010 1175.570 4.280 ;
        RECT 1176.410 0.010 1178.330 4.280 ;
        RECT 1179.170 0.010 1181.090 4.280 ;
        RECT 1181.930 0.010 1183.850 4.280 ;
        RECT 1184.690 0.010 1186.610 4.280 ;
        RECT 1187.450 0.010 1189.370 4.280 ;
        RECT 1190.210 0.010 1192.130 4.280 ;
        RECT 1192.970 0.010 1194.890 4.280 ;
        RECT 1195.730 0.010 1197.650 4.280 ;
        RECT 1198.490 0.010 1200.410 4.280 ;
        RECT 1201.250 0.010 1203.170 4.280 ;
        RECT 1204.010 0.010 1205.930 4.280 ;
        RECT 1206.770 0.010 1208.690 4.280 ;
        RECT 1209.530 0.010 1211.450 4.280 ;
        RECT 1212.290 0.010 1214.210 4.280 ;
        RECT 1215.050 0.010 1216.970 4.280 ;
        RECT 1217.810 0.010 1219.730 4.280 ;
        RECT 1220.570 0.010 1222.490 4.280 ;
        RECT 1223.330 0.010 1225.250 4.280 ;
        RECT 1226.090 0.010 1228.010 4.280 ;
        RECT 1228.850 0.010 1230.770 4.280 ;
        RECT 1231.610 0.010 1233.530 4.280 ;
        RECT 1234.370 0.010 1236.290 4.280 ;
        RECT 1237.130 0.010 1239.050 4.280 ;
        RECT 1239.890 0.010 1241.810 4.280 ;
        RECT 1242.650 0.010 1244.570 4.280 ;
        RECT 1245.410 0.010 1247.330 4.280 ;
        RECT 1248.170 0.010 1250.090 4.280 ;
        RECT 1250.930 0.010 1252.850 4.280 ;
        RECT 1253.690 0.010 1255.610 4.280 ;
        RECT 1256.450 0.010 1258.370 4.280 ;
        RECT 1259.210 0.010 1261.130 4.280 ;
        RECT 1261.970 0.010 1263.890 4.280 ;
        RECT 1264.730 0.010 1266.650 4.280 ;
        RECT 1267.490 0.010 1269.410 4.280 ;
        RECT 1270.250 0.010 1272.170 4.280 ;
        RECT 1273.010 0.010 1274.930 4.280 ;
        RECT 1275.770 0.010 1277.690 4.280 ;
        RECT 1278.530 0.010 1280.450 4.280 ;
        RECT 1281.290 0.010 1283.210 4.280 ;
        RECT 1284.050 0.010 1285.970 4.280 ;
        RECT 1286.810 0.010 1288.730 4.280 ;
        RECT 1289.570 0.010 1291.490 4.280 ;
        RECT 1292.330 0.010 1294.250 4.280 ;
        RECT 1295.090 0.010 1297.010 4.280 ;
        RECT 1297.850 0.010 1299.770 4.280 ;
        RECT 1300.610 0.010 1302.530 4.280 ;
        RECT 1303.370 0.010 1305.290 4.280 ;
        RECT 1306.130 0.010 1308.050 4.280 ;
        RECT 1308.890 0.010 1310.810 4.280 ;
        RECT 1311.650 0.010 1313.570 4.280 ;
        RECT 1314.410 0.010 1316.330 4.280 ;
        RECT 1317.170 0.010 1319.090 4.280 ;
        RECT 1319.930 0.010 1321.850 4.280 ;
        RECT 1322.690 0.010 1324.610 4.280 ;
        RECT 1325.450 0.010 1327.370 4.280 ;
        RECT 1328.210 0.010 1330.130 4.280 ;
        RECT 1330.970 0.010 1332.890 4.280 ;
        RECT 1333.730 0.010 1335.650 4.280 ;
        RECT 1336.490 0.010 1338.410 4.280 ;
        RECT 1339.250 0.010 1341.170 4.280 ;
        RECT 1342.010 0.010 1343.930 4.280 ;
        RECT 1344.770 0.010 1346.690 4.280 ;
        RECT 1347.530 0.010 1349.450 4.280 ;
        RECT 1350.290 0.010 1352.210 4.280 ;
        RECT 1353.050 0.010 1354.970 4.280 ;
        RECT 1355.810 0.010 1357.730 4.280 ;
        RECT 1358.570 0.010 1360.490 4.280 ;
        RECT 1361.330 0.010 1363.250 4.280 ;
        RECT 1364.090 0.010 1366.010 4.280 ;
        RECT 1366.850 0.010 1368.770 4.280 ;
        RECT 1369.610 0.010 1371.530 4.280 ;
        RECT 1372.370 0.010 1374.290 4.280 ;
        RECT 1375.130 0.010 1377.050 4.280 ;
        RECT 1377.890 0.010 1379.810 4.280 ;
        RECT 1380.650 0.010 1382.570 4.280 ;
        RECT 1383.410 0.010 1385.330 4.280 ;
        RECT 1386.170 0.010 1388.090 4.280 ;
        RECT 1388.930 0.010 1390.850 4.280 ;
        RECT 1391.690 0.010 1393.610 4.280 ;
        RECT 1394.450 0.010 1396.370 4.280 ;
        RECT 1397.210 0.010 1399.130 4.280 ;
        RECT 1399.970 0.010 1401.890 4.280 ;
        RECT 1402.730 0.010 1404.650 4.280 ;
        RECT 1405.490 0.010 1407.410 4.280 ;
        RECT 1408.250 0.010 1410.170 4.280 ;
        RECT 1411.010 0.010 1412.930 4.280 ;
        RECT 1413.770 0.010 1415.690 4.280 ;
        RECT 1416.530 0.010 1418.450 4.280 ;
        RECT 1419.290 0.010 1421.210 4.280 ;
        RECT 1422.050 0.010 1423.970 4.280 ;
        RECT 1424.810 0.010 1426.730 4.280 ;
        RECT 1427.570 0.010 1429.490 4.280 ;
        RECT 1430.330 0.010 1432.250 4.280 ;
        RECT 1433.090 0.010 1435.010 4.280 ;
        RECT 1435.850 0.010 1437.770 4.280 ;
        RECT 1438.610 0.010 1440.530 4.280 ;
        RECT 1441.370 0.010 1443.290 4.280 ;
        RECT 1444.130 0.010 1446.050 4.280 ;
        RECT 1446.890 0.010 1448.810 4.280 ;
        RECT 1449.650 0.010 1451.570 4.280 ;
        RECT 1452.410 0.010 1454.330 4.280 ;
        RECT 1455.170 0.010 1457.090 4.280 ;
        RECT 1457.930 0.010 1459.850 4.280 ;
        RECT 1460.690 0.010 1462.610 4.280 ;
        RECT 1463.450 0.010 1465.370 4.280 ;
        RECT 1466.210 0.010 1468.130 4.280 ;
        RECT 1468.970 0.010 1470.890 4.280 ;
        RECT 1471.730 0.010 1473.650 4.280 ;
        RECT 1474.490 0.010 1476.410 4.280 ;
        RECT 1477.250 0.010 1479.170 4.280 ;
        RECT 1480.010 0.010 1481.930 4.280 ;
        RECT 1482.770 0.010 1484.690 4.280 ;
        RECT 1485.530 0.010 1487.450 4.280 ;
        RECT 1488.290 0.010 1490.210 4.280 ;
        RECT 1491.050 0.010 1492.970 4.280 ;
        RECT 1493.810 0.010 1495.730 4.280 ;
        RECT 1496.570 0.010 1498.490 4.280 ;
        RECT 1499.330 0.010 1501.250 4.280 ;
        RECT 1502.090 0.010 1504.010 4.280 ;
        RECT 1504.850 0.010 1506.770 4.280 ;
        RECT 1507.610 0.010 1509.530 4.280 ;
        RECT 1510.370 0.010 1512.290 4.280 ;
        RECT 1513.130 0.010 1515.050 4.280 ;
        RECT 1515.890 0.010 1517.810 4.280 ;
        RECT 1518.650 0.010 1520.570 4.280 ;
        RECT 1521.410 0.010 1523.330 4.280 ;
        RECT 1524.170 0.010 1526.090 4.280 ;
        RECT 1526.930 0.010 1528.850 4.280 ;
        RECT 1529.690 0.010 1531.610 4.280 ;
        RECT 1532.450 0.010 1534.370 4.280 ;
        RECT 1535.210 0.010 1537.130 4.280 ;
        RECT 1537.970 0.010 1539.890 4.280 ;
        RECT 1540.730 0.010 1542.650 4.280 ;
        RECT 1543.490 0.010 1545.410 4.280 ;
        RECT 1546.250 0.010 1548.170 4.280 ;
        RECT 1549.010 0.010 1550.930 4.280 ;
        RECT 1551.770 0.010 1553.690 4.280 ;
        RECT 1554.530 0.010 1556.450 4.280 ;
        RECT 1557.290 0.010 1559.210 4.280 ;
        RECT 1560.050 0.010 1561.970 4.280 ;
        RECT 1562.810 0.010 1564.730 4.280 ;
        RECT 1565.570 0.010 1567.490 4.280 ;
        RECT 1568.330 0.010 1570.250 4.280 ;
        RECT 1571.090 0.010 1573.010 4.280 ;
        RECT 1573.850 0.010 1575.770 4.280 ;
        RECT 1576.610 0.010 1578.530 4.280 ;
        RECT 1579.370 0.010 1581.290 4.280 ;
        RECT 1582.130 0.010 1584.050 4.280 ;
        RECT 1584.890 0.010 1586.810 4.280 ;
        RECT 1587.650 0.010 1589.570 4.280 ;
        RECT 1590.410 0.010 1592.330 4.280 ;
        RECT 1593.170 0.010 1595.090 4.280 ;
        RECT 1595.930 0.010 1597.850 4.280 ;
        RECT 1598.690 0.010 1600.610 4.280 ;
        RECT 1601.450 0.010 1603.370 4.280 ;
        RECT 1604.210 0.010 1606.130 4.280 ;
        RECT 1606.970 0.010 1608.890 4.280 ;
        RECT 1609.730 0.010 1611.650 4.280 ;
        RECT 1612.490 0.010 1614.410 4.280 ;
        RECT 1615.250 0.010 1617.170 4.280 ;
        RECT 1618.010 0.010 1619.930 4.280 ;
        RECT 1620.770 0.010 1622.690 4.280 ;
        RECT 1623.530 0.010 1625.450 4.280 ;
        RECT 1626.290 0.010 1628.210 4.280 ;
        RECT 1629.050 0.010 1630.970 4.280 ;
        RECT 1631.810 0.010 1633.730 4.280 ;
        RECT 1634.570 0.010 1636.490 4.280 ;
        RECT 1637.330 0.010 1639.250 4.280 ;
        RECT 1640.090 0.010 1642.010 4.280 ;
        RECT 1642.850 0.010 1644.770 4.280 ;
        RECT 1645.610 0.010 1647.530 4.280 ;
        RECT 1648.370 0.010 1650.290 4.280 ;
        RECT 1651.130 0.010 1653.050 4.280 ;
        RECT 1653.890 0.010 1655.810 4.280 ;
        RECT 1656.650 0.010 1658.570 4.280 ;
        RECT 1659.410 0.010 1661.330 4.280 ;
        RECT 1662.170 0.010 1664.090 4.280 ;
        RECT 1664.930 0.010 1666.850 4.280 ;
        RECT 1667.690 0.010 1669.610 4.280 ;
        RECT 1670.450 0.010 1672.370 4.280 ;
        RECT 1673.210 0.010 1675.130 4.280 ;
        RECT 1675.970 0.010 1677.890 4.280 ;
        RECT 1678.730 0.010 1680.650 4.280 ;
        RECT 1681.490 0.010 1683.410 4.280 ;
        RECT 1684.250 0.010 1686.170 4.280 ;
        RECT 1687.010 0.010 1688.930 4.280 ;
        RECT 1689.770 0.010 1691.690 4.280 ;
        RECT 1692.530 0.010 1694.450 4.280 ;
        RECT 1695.290 0.010 1697.210 4.280 ;
        RECT 1698.050 0.010 1699.970 4.280 ;
        RECT 1700.810 0.010 1702.730 4.280 ;
        RECT 1703.570 0.010 1705.490 4.280 ;
        RECT 1706.330 0.010 1708.250 4.280 ;
        RECT 1709.090 0.010 1711.010 4.280 ;
        RECT 1711.850 0.010 1713.770 4.280 ;
        RECT 1714.610 0.010 1716.530 4.280 ;
        RECT 1717.370 0.010 1719.290 4.280 ;
        RECT 1720.130 0.010 1722.050 4.280 ;
        RECT 1722.890 0.010 1724.810 4.280 ;
        RECT 1725.650 0.010 1727.570 4.280 ;
        RECT 1728.410 0.010 1730.330 4.280 ;
        RECT 1731.170 0.010 1733.090 4.280 ;
        RECT 1733.930 0.010 1735.850 4.280 ;
        RECT 1736.690 0.010 1738.610 4.280 ;
        RECT 1739.450 0.010 1741.370 4.280 ;
        RECT 1742.210 0.010 1744.130 4.280 ;
        RECT 1744.970 0.010 1746.890 4.280 ;
        RECT 1747.730 0.010 1749.650 4.280 ;
        RECT 1750.490 0.010 1752.410 4.280 ;
        RECT 1753.250 0.010 1755.170 4.280 ;
        RECT 1756.010 0.010 1757.930 4.280 ;
        RECT 1758.770 0.010 1760.690 4.280 ;
        RECT 1761.530 0.010 1763.450 4.280 ;
        RECT 1764.290 0.010 1766.210 4.280 ;
        RECT 1767.050 0.010 1768.970 4.280 ;
        RECT 1769.810 0.010 1771.730 4.280 ;
        RECT 1772.570 0.010 1774.490 4.280 ;
        RECT 1775.330 0.010 1777.250 4.280 ;
        RECT 1778.090 0.010 1780.010 4.280 ;
        RECT 1780.850 0.010 1782.770 4.280 ;
        RECT 1783.610 0.010 1785.530 4.280 ;
        RECT 1786.370 0.010 1788.290 4.280 ;
        RECT 1789.130 0.010 1791.050 4.280 ;
        RECT 1791.890 0.010 1793.810 4.280 ;
        RECT 1794.650 0.010 1796.570 4.280 ;
        RECT 1797.410 0.010 1799.330 4.280 ;
        RECT 1800.170 0.010 1891.890 4.280 ;
      LAYER met3 ;
        RECT 25.130 154.040 1896.000 159.625 ;
        RECT 25.130 152.640 1895.600 154.040 ;
        RECT 25.130 141.800 1896.000 152.640 ;
        RECT 25.130 140.400 1895.600 141.800 ;
        RECT 25.130 129.560 1896.000 140.400 ;
        RECT 25.130 128.160 1895.600 129.560 ;
        RECT 25.130 117.320 1896.000 128.160 ;
        RECT 25.130 115.920 1895.600 117.320 ;
        RECT 25.130 105.080 1896.000 115.920 ;
        RECT 25.130 103.680 1895.600 105.080 ;
        RECT 25.130 92.840 1896.000 103.680 ;
        RECT 25.130 91.440 1895.600 92.840 ;
        RECT 25.130 80.600 1896.000 91.440 ;
        RECT 25.130 79.200 1895.600 80.600 ;
        RECT 25.130 68.360 1896.000 79.200 ;
        RECT 25.130 66.960 1895.600 68.360 ;
        RECT 25.130 56.120 1896.000 66.960 ;
        RECT 25.130 54.720 1895.600 56.120 ;
        RECT 25.130 43.880 1896.000 54.720 ;
        RECT 25.130 42.480 1895.600 43.880 ;
        RECT 25.130 31.640 1896.000 42.480 ;
        RECT 25.130 30.240 1895.600 31.640 ;
        RECT 25.130 19.400 1896.000 30.240 ;
        RECT 25.130 18.000 1895.600 19.400 ;
        RECT 25.130 7.160 1896.000 18.000 ;
        RECT 25.130 5.760 1895.600 7.160 ;
        RECT 25.130 0.175 1896.000 5.760 ;
      LAYER met4 ;
        RECT 289.175 4.800 325.670 146.025 ;
        RECT 327.370 4.800 333.870 146.025 ;
        RECT 335.570 4.800 354.770 146.025 ;
        RECT 356.470 4.800 362.570 146.025 ;
        RECT 364.270 4.800 383.870 146.025 ;
        RECT 385.570 4.800 400.920 146.025 ;
        RECT 402.620 4.800 404.770 146.025 ;
        RECT 406.470 4.800 437.820 146.025 ;
        RECT 439.520 4.800 476.170 146.025 ;
        RECT 477.870 4.800 513.070 146.025 ;
        RECT 514.770 4.800 551.420 146.025 ;
        RECT 553.120 4.800 588.320 146.025 ;
        RECT 590.020 4.800 626.670 146.025 ;
        RECT 628.370 4.800 663.570 146.025 ;
        RECT 665.270 4.800 701.920 146.025 ;
        RECT 703.620 4.800 706.020 146.025 ;
        RECT 707.720 4.800 738.820 146.025 ;
        RECT 740.520 4.800 742.920 146.025 ;
        RECT 744.620 4.800 777.170 146.025 ;
        RECT 778.870 4.800 781.270 146.025 ;
        RECT 782.970 4.800 814.070 146.025 ;
        RECT 815.770 4.800 818.170 146.025 ;
        RECT 819.870 4.800 852.420 146.025 ;
        RECT 854.120 4.800 856.520 146.025 ;
        RECT 858.220 4.800 889.320 146.025 ;
        RECT 891.020 4.800 893.420 146.025 ;
        RECT 895.120 4.800 927.670 146.025 ;
        RECT 929.370 4.800 931.770 146.025 ;
        RECT 933.470 4.800 964.570 146.025 ;
        RECT 966.270 4.800 968.670 146.025 ;
        RECT 970.370 4.800 1002.920 146.025 ;
        RECT 1004.620 4.800 1039.820 146.025 ;
        RECT 1041.520 4.800 1078.170 146.025 ;
        RECT 1079.870 4.800 1115.070 146.025 ;
        RECT 1116.770 4.800 1153.420 146.025 ;
        RECT 1155.120 4.800 1190.320 146.025 ;
        RECT 1192.020 4.800 1228.670 146.025 ;
        RECT 1230.370 4.800 1265.570 146.025 ;
        RECT 1267.270 4.800 1278.670 146.025 ;
        RECT 1280.370 4.800 1282.670 146.025 ;
        RECT 1284.370 4.800 1303.920 146.025 ;
        RECT 1305.620 4.800 1315.570 146.025 ;
        RECT 1317.270 4.800 1319.570 146.025 ;
        RECT 1321.270 4.800 1340.820 146.025 ;
        RECT 1342.520 4.800 1353.920 146.025 ;
        RECT 1355.620 4.800 1357.920 146.025 ;
        RECT 1359.620 4.800 1379.170 146.025 ;
        RECT 1380.870 4.800 1390.820 146.025 ;
        RECT 1392.520 4.800 1394.820 146.025 ;
        RECT 1396.520 4.800 1416.070 146.025 ;
        RECT 1417.770 4.800 1454.420 146.025 ;
        RECT 1456.120 4.800 1491.320 146.025 ;
        RECT 1493.020 4.800 1529.670 146.025 ;
        RECT 1531.370 4.800 1566.570 146.025 ;
        RECT 1568.270 4.800 1604.920 146.025 ;
        RECT 1606.620 4.800 1641.820 146.025 ;
        RECT 1643.520 4.800 1680.170 146.025 ;
        RECT 1681.870 4.800 1691.585 146.025 ;
        RECT 289.175 0.175 1691.585 4.800 ;
  END
END mgmt_protect
END LIBRARY

