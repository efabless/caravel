VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gpio_logic_high
  CLASS BLOCK ;
  FOREIGN gpio_logic_high ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.000 BY 16.000 ;
  PIN gpio_logic1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3.000 8.200 7.000 8.800 ;
    END
  END gpio_logic1
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.300 -0.240 1.700 13.840 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 -0.240 5.400 13.840 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT -0.190 12.185 7.090 13.790 ;
        RECT -0.190 6.745 7.090 9.575 ;
        RECT -0.190 1.305 7.090 4.135 ;
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 3.360 -0.055 3.480 0.055 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
      LAYER li1 ;
        RECT 0.000 0.085 6.900 13.685 ;
      LAYER li1 ;
        RECT 0.000 -0.085 6.900 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.240 6.900 13.840 ;
      LAYER met2 ;
        RECT 0.390 0.000 5.310 13.840 ;
        RECT 4.090 -0.240 5.310 0.000 ;
      LAYER met3 ;
        RECT 0.300 9.200 5.400 13.765 ;
        RECT 0.300 7.800 2.600 9.200 ;
        RECT 0.300 0.000 5.400 7.800 ;
        RECT 4.000 -0.165 5.400 0.000 ;
  END
END gpio_logic_high
END LIBRARY

