magic
tech sky130A
magscale 1 2
timestamp 1623523101
<< viali >>
rect 18797 221 18831 255
<< metal1 >>
rect 0 1114 19964 1136
rect 0 1062 174 1114
rect 226 1062 8174 1114
rect 8226 1062 16174 1114
rect 16226 1062 19964 1114
rect 0 1040 19964 1062
rect 0 570 19964 592
rect 0 518 4174 570
rect 4226 518 12174 570
rect 12226 518 19964 570
rect 0 496 19964 518
rect 18782 252 18788 264
rect 18743 224 18788 252
rect 18782 212 18788 224
rect 18840 212 18846 264
rect 0 26 19964 48
rect 0 -26 174 26
rect 226 -26 8174 26
rect 8226 -26 16174 26
rect 16226 -26 19964 26
rect 0 -48 19964 -26
<< via1 >>
rect 174 1062 226 1114
rect 8174 1062 8226 1114
rect 16174 1062 16226 1114
rect 4174 518 4226 570
rect 12174 518 12226 570
rect 18788 255 18840 264
rect 18788 221 18797 255
rect 18797 221 18831 255
rect 18831 221 18840 255
rect 18788 212 18840 221
rect 174 -26 226 26
rect 8174 -26 8226 26
rect 16174 -26 16226 26
<< metal2 >>
rect 170 1114 230 1136
rect 170 1062 174 1114
rect 226 1062 230 1114
rect 170 380 230 1062
rect 4170 960 4230 1136
rect 4170 904 4172 960
rect 4228 904 4230 960
rect 4066 776 4122 785
rect 4066 711 4122 720
rect 170 324 172 380
rect 228 324 230 380
rect 170 26 230 324
rect 4080 241 4108 711
rect 4170 570 4230 904
rect 4170 518 4174 570
rect 4226 518 4230 570
rect 4066 232 4122 241
rect 4066 167 4122 176
rect 170 -26 174 26
rect 226 -26 230 26
rect 170 -48 230 -26
rect 4170 -48 4230 518
rect 8170 1114 8230 1136
rect 8170 1062 8174 1114
rect 8226 1062 8230 1114
rect 8170 380 8230 1062
rect 8170 324 8172 380
rect 8228 324 8230 380
rect 8170 26 8230 324
rect 8170 -26 8174 26
rect 8226 -26 8230 26
rect 8170 -48 8230 -26
rect 12170 960 12230 1136
rect 12170 904 12172 960
rect 12228 904 12230 960
rect 12170 570 12230 904
rect 12170 518 12174 570
rect 12226 518 12230 570
rect 12170 -48 12230 518
rect 16170 1114 16230 1136
rect 16170 1062 16174 1114
rect 16226 1062 16230 1114
rect 16170 380 16230 1062
rect 16170 324 16172 380
rect 16228 324 16230 380
rect 16170 26 16230 324
rect 18788 264 18840 270
rect 18786 232 18788 241
rect 18840 232 18842 241
rect 18786 167 18842 176
rect 16170 -26 16174 26
rect 16226 -26 16230 26
rect 16170 -48 16230 -26
<< via2 >>
rect 4172 904 4228 960
rect 4066 720 4122 776
rect 172 324 228 380
rect 4066 176 4122 232
rect 8172 324 8228 380
rect 12172 904 12228 960
rect 16172 324 16228 380
rect 18786 212 18788 232
rect 18788 212 18840 232
rect 18840 212 18842 232
rect 18786 176 18842 212
<< metal3 >>
rect 0 960 19964 977
rect 0 904 4172 960
rect 4228 904 12172 960
rect 12228 904 19964 960
rect 0 887 19964 904
rect 0 778 800 808
rect 4061 778 4127 781
rect 0 776 4127 778
rect 0 720 4066 776
rect 4122 720 4127 776
rect 0 718 4127 720
rect 0 688 800 718
rect 4061 715 4127 718
rect 0 380 19964 397
rect 0 324 172 380
rect 228 324 8172 380
rect 8228 324 16172 380
rect 16228 324 19964 380
rect 0 307 19964 324
rect 4061 234 4127 237
rect 18781 234 18847 237
rect 4061 232 18847 234
rect 4061 176 4066 232
rect 4122 176 18786 232
rect 18842 176 18847 232
rect 4061 174 18847 176
rect 4061 171 4127 174
rect 18781 171 18847 174
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623438133
transform 1 0 0 0 -1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1623438133
transform 1 0 0 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623438133
transform 1 0 276 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1623438133
transform 1 0 276 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1623438133
transform 1 0 1380 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1623438133
transform 1 0 1380 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623438133
transform 1 0 2668 0 -1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_11
timestamp 1623438133
transform 1 0 2668 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623438133
transform 1 0 2484 0 -1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_30
timestamp 1623438133
transform 1 0 2760 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_27
timestamp 1623438133
transform 1 0 2484 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_30
timestamp 1623438133
transform 1 0 2760 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_42
timestamp 1623438133
transform 1 0 3864 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_42
timestamp 1623438133
transform 1 0 3864 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_5
timestamp 1623438133
transform 1 0 5336 0 -1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_12
timestamp 1623438133
transform 1 0 5336 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623438133
transform 1 0 4968 0 -1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_59
timestamp 1623438133
transform 1 0 5428 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_54
timestamp 1623438133
transform 1 0 4968 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_59
timestamp 1623438133
transform 1 0 5428 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_71
timestamp 1623438133
transform 1 0 6532 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_71
timestamp 1623438133
transform 1 0 6532 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_6
timestamp 1623438133
transform 1 0 8004 0 -1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_13
timestamp 1623438133
transform 1 0 8004 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83
timestamp 1623438133
transform 1 0 7636 0 -1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_88
timestamp 1623438133
transform 1 0 8096 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_83
timestamp 1623438133
transform 1 0 7636 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_88
timestamp 1623438133
transform 1 0 8096 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_100
timestamp 1623438133
transform 1 0 9200 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_100
timestamp 1623438133
transform 1 0 9200 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112
timestamp 1623438133
transform 1 0 10304 0 -1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_112
timestamp 1623438133
transform 1 0 10304 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_7
timestamp 1623438133
transform 1 0 10672 0 -1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_14
timestamp 1623438133
transform 1 0 10672 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_117
timestamp 1623438133
transform 1 0 10764 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_117
timestamp 1623438133
transform 1 0 10764 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_129
timestamp 1623438133
transform 1 0 11868 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1623438133
transform 1 0 12972 0 -1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_129
timestamp 1623438133
transform 1 0 11868 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_141
timestamp 1623438133
transform 1 0 12972 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_8
timestamp 1623438133
transform 1 0 13340 0 -1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_15
timestamp 1623438133
transform 1 0 13340 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_146
timestamp 1623438133
transform 1 0 13432 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_146
timestamp 1623438133
transform 1 0 13432 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_158
timestamp 1623438133
transform 1 0 14536 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_158
timestamp 1623438133
transform 1 0 14536 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_9
timestamp 1623438133
transform 1 0 16008 0 -1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_16
timestamp 1623438133
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_170
timestamp 1623438133
transform 1 0 15640 0 -1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_175
timestamp 1623438133
transform 1 0 16100 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_170
timestamp 1623438133
transform 1 0 15640 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_175
timestamp 1623438133
transform 1 0 16100 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1623438133
transform 1 0 17204 0 -1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_187
timestamp 1623438133
transform 1 0 17204 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  inst $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623438133
transform 1 0 18768 0 -1 544
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_10
timestamp 1623438133
transform 1 0 18676 0 -1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_17
timestamp 1623438133
transform 1 0 18676 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_199
timestamp 1623438133
transform 1 0 18308 0 -1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_199
timestamp 1623438133
transform 1 0 18308 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_204 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623438133
transform 1 0 18768 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1623438133
transform -1 0 19964 0 -1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1623438133
transform -1 0 19964 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_207 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623438133
transform 1 0 19044 0 -1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_213 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623438133
transform 1 0 19596 0 -1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_212
timestamp 1623438133
transform 1 0 19504 0 1 544
box -38 -48 222 592
<< labels >>
rlabel metal3 s 0 688 800 808 6 HI
port 0 nsew signal tristate
rlabel metal2 s 16170 -48 16230 1136 6 vccd2
port 1 nsew power bidirectional
rlabel metal2 s 8170 -48 8230 1136 6 vccd2
port 2 nsew power bidirectional
rlabel metal2 s 170 -48 230 1136 6 vccd2
port 3 nsew power bidirectional
rlabel metal3 s 0 307 19964 397 6 vccd2
port 4 nsew power bidirectional
rlabel metal2 s 12170 -48 12230 1136 6 vssd2
port 5 nsew ground bidirectional
rlabel metal2 s 4170 -48 4230 1136 6 vssd2
port 6 nsew ground bidirectional
rlabel metal3 s 0 887 19964 977 6 vssd2
port 7 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 1400
<< end >>
