VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gpio_signal_buffering_alt
  CLASS BLOCK ;
  FOREIGN gpio_signal_buffering_alt ;
  ORIGIN 0.000 0.000 ;
  SIZE 3588.000 BY 5188.000 ;
  PIN mgmt_io_in_unbuf[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3381.660 3606.800 3381.860 3608.390 ;
      LAYER mcon ;
        RECT 3381.690 3607.300 3381.860 3608.390 ;
      LAYER met1 ;
        RECT 3370.780 3608.085 3370.920 3641.605 ;
        RECT 3370.780 3607.765 3371.040 3608.085 ;
        RECT 3381.640 3607.240 3381.900 3608.450 ;
      LAYER via ;
        RECT 3370.780 3607.795 3371.040 3608.055 ;
        RECT 3381.640 3607.300 3381.900 3608.390 ;
      LAYER met2 ;
        RECT 3370.750 3607.935 3371.070 3608.055 ;
        RECT 3381.610 3607.935 3381.930 3608.390 ;
        RECT 3370.330 3607.795 3381.930 3607.935 ;
        RECT 3381.610 3607.300 3381.930 3607.795 ;
    END
  END mgmt_io_in_unbuf[6]
  PIN mgmt_io_out_buf[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.560 3606.895 3385.770 3607.065 ;
        RECT 3384.410 3606.810 3385.290 3606.895 ;
        RECT 3384.410 3606.225 3384.580 3606.810 ;
        RECT 3383.560 3606.055 3384.580 3606.225 ;
        RECT 3384.410 3605.385 3384.580 3606.055 ;
        RECT 3383.560 3605.215 3384.580 3605.385 ;
        RECT 3384.410 3604.545 3384.580 3605.215 ;
        RECT 3383.560 3604.375 3384.580 3604.545 ;
        RECT 3385.120 3606.225 3385.290 3606.810 ;
        RECT 3385.120 3606.055 3385.770 3606.225 ;
        RECT 3385.120 3605.385 3385.290 3606.055 ;
        RECT 3385.120 3605.215 3385.770 3605.385 ;
        RECT 3385.120 3604.545 3385.290 3605.215 ;
        RECT 3385.120 3604.375 3385.770 3604.545 ;
      LAYER met1 ;
        RECT 3370.220 3638.535 3370.360 3640.605 ;
        RECT 3370.220 3638.395 3370.640 3638.535 ;
        RECT 3370.500 3607.115 3370.640 3638.395 ;
        RECT 3370.500 3606.795 3370.760 3607.115 ;
        RECT 3384.350 3606.760 3385.320 3607.020 ;
      LAYER via ;
        RECT 3370.500 3606.825 3370.760 3607.085 ;
        RECT 3384.410 3606.760 3385.260 3607.020 ;
      LAYER met2 ;
        RECT 3370.470 3606.965 3370.790 3607.085 ;
        RECT 3384.410 3606.965 3385.260 3607.050 ;
        RECT 3370.330 3606.825 3385.260 3606.965 ;
        RECT 3384.410 3606.730 3385.260 3606.825 ;
    END
  END mgmt_io_out_buf[6]
  PIN mgmt_io_in_unbuf[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3381.660 2230.700 3381.860 2232.290 ;
      LAYER mcon ;
        RECT 3381.690 2231.200 3381.860 2232.290 ;
      LAYER met1 ;
        RECT 3369.800 2231.985 3369.940 2281.275 ;
        RECT 3369.800 2231.665 3370.060 2231.985 ;
        RECT 3381.640 2231.140 3381.900 2232.350 ;
      LAYER via ;
        RECT 3369.800 2231.695 3370.060 2231.955 ;
        RECT 3381.640 2231.200 3381.900 2232.290 ;
      LAYER met2 ;
        RECT 3369.770 2231.835 3370.090 2231.955 ;
        RECT 3381.610 2231.835 3381.930 2232.290 ;
        RECT 3365.990 2231.695 3381.930 2231.835 ;
        RECT 3381.610 2231.200 3381.930 2231.695 ;
    END
  END mgmt_io_in_unbuf[5]
  PIN mgmt_io_in_unbuf[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3381.660 2224.720 3381.860 2226.310 ;
      LAYER mcon ;
        RECT 3381.690 2225.220 3381.860 2226.310 ;
      LAYER met1 ;
        RECT 3368.680 2226.005 3368.820 2279.275 ;
        RECT 3368.680 2225.685 3368.940 2226.005 ;
        RECT 3381.640 2225.160 3381.900 2226.370 ;
      LAYER via ;
        RECT 3368.680 2225.715 3368.940 2225.975 ;
        RECT 3381.640 2225.220 3381.900 2226.310 ;
      LAYER met2 ;
        RECT 3368.650 2225.855 3368.970 2225.975 ;
        RECT 3381.610 2225.855 3381.930 2226.310 ;
        RECT 3365.990 2225.715 3381.930 2225.855 ;
        RECT 3381.610 2225.220 3381.930 2225.715 ;
    END
  END mgmt_io_in_unbuf[4]
  PIN mgmt_io_in_unbuf[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3381.660 2218.740 3381.860 2220.330 ;
      LAYER mcon ;
        RECT 3381.690 2219.240 3381.860 2220.330 ;
      LAYER met1 ;
        RECT 3367.560 2220.025 3367.700 2277.275 ;
        RECT 3367.560 2219.705 3367.820 2220.025 ;
        RECT 3381.640 2219.180 3381.900 2220.390 ;
      LAYER via ;
        RECT 3367.560 2219.735 3367.820 2219.995 ;
        RECT 3381.640 2219.240 3381.900 2220.330 ;
      LAYER met2 ;
        RECT 3367.530 2219.875 3367.850 2219.995 ;
        RECT 3381.610 2219.875 3381.930 2220.330 ;
        RECT 3365.990 2219.735 3381.930 2219.875 ;
        RECT 3381.610 2219.240 3381.930 2219.735 ;
    END
  END mgmt_io_in_unbuf[3]
  PIN mgmt_io_in_unbuf[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3381.660 2212.760 3381.860 2214.350 ;
      LAYER mcon ;
        RECT 3381.690 2213.260 3381.860 2214.350 ;
      LAYER met1 ;
        RECT 3366.440 2214.045 3366.580 2275.275 ;
        RECT 3366.440 2213.725 3366.700 2214.045 ;
        RECT 3381.640 2213.200 3381.900 2214.410 ;
      LAYER via ;
        RECT 3366.440 2213.755 3366.700 2214.015 ;
        RECT 3381.640 2213.260 3381.900 2214.350 ;
      LAYER met2 ;
        RECT 3366.410 2213.895 3366.730 2214.015 ;
        RECT 3381.610 2213.895 3381.930 2214.350 ;
        RECT 3365.990 2213.755 3381.930 2213.895 ;
        RECT 3381.610 2213.260 3381.930 2213.755 ;
    END
  END mgmt_io_in_unbuf[2]
  PIN mgmt_io_in_unbuf[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3381.660 2206.780 3381.860 2208.370 ;
      LAYER mcon ;
        RECT 3381.690 2207.280 3381.860 2208.370 ;
      LAYER met1 ;
        RECT 3365.320 2208.065 3365.460 2273.275 ;
        RECT 3365.320 2207.745 3365.580 2208.065 ;
        RECT 3381.640 2207.220 3381.900 2208.430 ;
      LAYER via ;
        RECT 3365.320 2207.775 3365.580 2208.035 ;
        RECT 3381.640 2207.280 3381.900 2208.370 ;
      LAYER met2 ;
        RECT 3365.290 2207.915 3365.610 2208.035 ;
        RECT 3381.610 2207.915 3381.930 2208.370 ;
        RECT 3364.865 2207.775 3381.930 2207.915 ;
        RECT 3381.610 2207.280 3381.930 2207.775 ;
    END
  END mgmt_io_in_unbuf[1]
  PIN mgmt_io_in_unbuf[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3381.660 2200.800 3381.860 2202.390 ;
      LAYER mcon ;
        RECT 3381.690 2201.300 3381.860 2202.390 ;
      LAYER met1 ;
        RECT 3364.200 2202.085 3364.340 2271.275 ;
        RECT 3364.200 2201.765 3364.460 2202.085 ;
        RECT 3381.640 2201.240 3381.900 2202.450 ;
      LAYER via ;
        RECT 3364.200 2201.795 3364.460 2202.055 ;
        RECT 3381.640 2201.300 3381.900 2202.390 ;
      LAYER met2 ;
        RECT 3364.170 2201.935 3364.490 2202.055 ;
        RECT 3381.610 2201.935 3381.930 2202.390 ;
        RECT 3363.750 2201.795 3381.930 2201.935 ;
        RECT 3381.610 2201.300 3381.930 2201.795 ;
    END
  END mgmt_io_in_unbuf[0]
  PIN mgmt_io_out_buf[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.560 2200.895 3385.770 2201.065 ;
        RECT 3384.410 2200.810 3385.290 2200.895 ;
        RECT 3384.410 2200.225 3384.580 2200.810 ;
        RECT 3383.560 2200.055 3384.580 2200.225 ;
        RECT 3384.410 2199.385 3384.580 2200.055 ;
        RECT 3383.560 2199.215 3384.580 2199.385 ;
        RECT 3384.410 2198.545 3384.580 2199.215 ;
        RECT 3383.560 2198.375 3384.580 2198.545 ;
        RECT 3385.120 2200.225 3385.290 2200.810 ;
        RECT 3385.120 2200.055 3385.770 2200.225 ;
        RECT 3385.120 2199.385 3385.290 2200.055 ;
        RECT 3385.120 2199.215 3385.770 2199.385 ;
        RECT 3385.120 2198.545 3385.290 2199.215 ;
        RECT 3385.120 2198.375 3385.770 2198.545 ;
      LAYER met1 ;
        RECT 3363.640 2267.635 3363.780 2270.275 ;
        RECT 3363.640 2267.495 3364.060 2267.635 ;
        RECT 3363.920 2201.115 3364.060 2267.495 ;
        RECT 3363.920 2200.795 3364.180 2201.115 ;
        RECT 3384.350 2200.760 3385.320 2201.020 ;
      LAYER via ;
        RECT 3363.920 2200.825 3364.180 2201.085 ;
        RECT 3384.410 2200.760 3385.260 2201.020 ;
      LAYER met2 ;
        RECT 3363.890 2200.965 3364.210 2201.085 ;
        RECT 3384.410 2200.965 3385.260 2201.050 ;
        RECT 3363.750 2200.825 3385.260 2200.965 ;
        RECT 3384.410 2200.730 3385.260 2200.825 ;
    END
  END mgmt_io_out_buf[0]
  PIN mgmt_io_out_buf[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.560 2206.875 3385.770 2207.045 ;
        RECT 3384.410 2206.790 3385.290 2206.875 ;
        RECT 3384.410 2206.205 3384.580 2206.790 ;
        RECT 3383.560 2206.035 3384.580 2206.205 ;
        RECT 3384.410 2205.365 3384.580 2206.035 ;
        RECT 3383.560 2205.195 3384.580 2205.365 ;
        RECT 3384.410 2204.525 3384.580 2205.195 ;
        RECT 3383.560 2204.355 3384.580 2204.525 ;
        RECT 3385.120 2206.205 3385.290 2206.790 ;
        RECT 3385.120 2206.035 3385.770 2206.205 ;
        RECT 3385.120 2205.365 3385.290 2206.035 ;
        RECT 3385.120 2205.195 3385.770 2205.365 ;
        RECT 3385.120 2204.525 3385.290 2205.195 ;
        RECT 3385.120 2204.355 3385.770 2204.525 ;
      LAYER met1 ;
        RECT 3364.760 2269.660 3364.900 2272.275 ;
        RECT 3364.760 2269.520 3365.180 2269.660 ;
        RECT 3365.040 2207.095 3365.180 2269.520 ;
        RECT 3365.040 2206.775 3365.300 2207.095 ;
        RECT 3384.350 2206.740 3385.320 2207.000 ;
      LAYER via ;
        RECT 3365.040 2206.805 3365.300 2207.065 ;
        RECT 3384.410 2206.740 3385.260 2207.000 ;
      LAYER met2 ;
        RECT 3365.010 2206.945 3365.330 2207.065 ;
        RECT 3384.410 2206.945 3385.260 2207.030 ;
        RECT 3364.865 2206.805 3385.260 2206.945 ;
        RECT 3384.410 2206.710 3385.260 2206.805 ;
    END
  END mgmt_io_out_buf[1]
  PIN mgmt_io_out_buf[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.560 2212.855 3385.770 2213.025 ;
        RECT 3384.410 2212.770 3385.290 2212.855 ;
        RECT 3384.410 2212.185 3384.580 2212.770 ;
        RECT 3383.560 2212.015 3384.580 2212.185 ;
        RECT 3384.410 2211.345 3384.580 2212.015 ;
        RECT 3383.560 2211.175 3384.580 2211.345 ;
        RECT 3384.410 2210.505 3384.580 2211.175 ;
        RECT 3383.560 2210.335 3384.580 2210.505 ;
        RECT 3385.120 2212.185 3385.290 2212.770 ;
        RECT 3385.120 2212.015 3385.770 2212.185 ;
        RECT 3385.120 2211.345 3385.290 2212.015 ;
        RECT 3385.120 2211.175 3385.770 2211.345 ;
        RECT 3385.120 2210.505 3385.290 2211.175 ;
        RECT 3385.120 2210.335 3385.770 2210.505 ;
      LAYER met1 ;
        RECT 3365.880 2271.665 3366.020 2274.275 ;
        RECT 3365.880 2271.525 3366.300 2271.665 ;
        RECT 3366.160 2213.075 3366.300 2271.525 ;
        RECT 3366.160 2212.755 3366.420 2213.075 ;
        RECT 3384.350 2212.720 3385.320 2212.980 ;
      LAYER via ;
        RECT 3366.160 2212.785 3366.420 2213.045 ;
        RECT 3384.410 2212.720 3385.260 2212.980 ;
      LAYER met2 ;
        RECT 3366.130 2212.925 3366.450 2213.045 ;
        RECT 3384.410 2212.925 3385.260 2213.010 ;
        RECT 3365.990 2212.785 3385.260 2212.925 ;
        RECT 3384.410 2212.690 3385.260 2212.785 ;
    END
  END mgmt_io_out_buf[2]
  PIN mgmt_io_out_buf[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.560 2218.835 3385.770 2219.005 ;
        RECT 3384.410 2218.750 3385.290 2218.835 ;
        RECT 3384.410 2218.165 3384.580 2218.750 ;
        RECT 3383.560 2217.995 3384.580 2218.165 ;
        RECT 3384.410 2217.325 3384.580 2217.995 ;
        RECT 3383.560 2217.155 3384.580 2217.325 ;
        RECT 3384.410 2216.485 3384.580 2217.155 ;
        RECT 3383.560 2216.315 3384.580 2216.485 ;
        RECT 3385.120 2218.165 3385.290 2218.750 ;
        RECT 3385.120 2217.995 3385.770 2218.165 ;
        RECT 3385.120 2217.325 3385.290 2217.995 ;
        RECT 3385.120 2217.155 3385.770 2217.325 ;
        RECT 3385.120 2216.485 3385.290 2217.155 ;
        RECT 3385.120 2216.315 3385.770 2216.485 ;
      LAYER met1 ;
        RECT 3367.000 2273.895 3367.140 2276.275 ;
        RECT 3367.000 2273.755 3367.420 2273.895 ;
        RECT 3367.280 2219.055 3367.420 2273.755 ;
        RECT 3367.280 2218.735 3367.540 2219.055 ;
        RECT 3384.350 2218.700 3385.320 2218.960 ;
      LAYER via ;
        RECT 3367.280 2218.765 3367.540 2219.025 ;
        RECT 3384.410 2218.700 3385.260 2218.960 ;
      LAYER met2 ;
        RECT 3367.250 2218.905 3367.570 2219.025 ;
        RECT 3384.410 2218.905 3385.260 2218.990 ;
        RECT 3365.990 2218.765 3385.260 2218.905 ;
        RECT 3384.410 2218.670 3385.260 2218.765 ;
    END
  END mgmt_io_out_buf[3]
  PIN mgmt_io_out_buf[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.560 2224.815 3385.770 2224.985 ;
        RECT 3384.410 2224.730 3385.290 2224.815 ;
        RECT 3384.410 2224.145 3384.580 2224.730 ;
        RECT 3383.560 2223.975 3384.580 2224.145 ;
        RECT 3384.410 2223.305 3384.580 2223.975 ;
        RECT 3383.560 2223.135 3384.580 2223.305 ;
        RECT 3384.410 2222.465 3384.580 2223.135 ;
        RECT 3383.560 2222.295 3384.580 2222.465 ;
        RECT 3385.120 2224.145 3385.290 2224.730 ;
        RECT 3385.120 2223.975 3385.770 2224.145 ;
        RECT 3385.120 2223.305 3385.290 2223.975 ;
        RECT 3385.120 2223.135 3385.770 2223.305 ;
        RECT 3385.120 2222.465 3385.290 2223.135 ;
        RECT 3385.120 2222.295 3385.770 2222.465 ;
      LAYER met1 ;
        RECT 3368.120 2275.655 3368.260 2278.275 ;
        RECT 3368.120 2275.515 3368.540 2275.655 ;
        RECT 3368.400 2225.035 3368.540 2275.515 ;
        RECT 3368.400 2224.715 3368.660 2225.035 ;
        RECT 3384.350 2224.680 3385.320 2224.940 ;
      LAYER via ;
        RECT 3368.400 2224.745 3368.660 2225.005 ;
        RECT 3384.410 2224.680 3385.260 2224.940 ;
      LAYER met2 ;
        RECT 3368.370 2224.885 3368.690 2225.005 ;
        RECT 3384.410 2224.885 3385.260 2224.970 ;
        RECT 3365.990 2224.745 3385.260 2224.885 ;
        RECT 3384.410 2224.650 3385.260 2224.745 ;
    END
  END mgmt_io_out_buf[4]
  PIN mgmt_io_out_buf[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.560 2230.795 3385.770 2230.965 ;
        RECT 3384.410 2230.710 3385.290 2230.795 ;
        RECT 3384.410 2230.125 3384.580 2230.710 ;
        RECT 3383.560 2229.955 3384.580 2230.125 ;
        RECT 3384.410 2229.285 3384.580 2229.955 ;
        RECT 3383.560 2229.115 3384.580 2229.285 ;
        RECT 3384.410 2228.445 3384.580 2229.115 ;
        RECT 3383.560 2228.275 3384.580 2228.445 ;
        RECT 3385.120 2230.125 3385.290 2230.710 ;
        RECT 3385.120 2229.955 3385.770 2230.125 ;
        RECT 3385.120 2229.285 3385.290 2229.955 ;
        RECT 3385.120 2229.115 3385.770 2229.285 ;
        RECT 3385.120 2228.445 3385.290 2229.115 ;
        RECT 3385.120 2228.275 3385.770 2228.445 ;
      LAYER met1 ;
        RECT 3369.240 2277.665 3369.380 2280.275 ;
        RECT 3369.240 2277.525 3369.660 2277.665 ;
        RECT 3369.520 2231.015 3369.660 2277.525 ;
        RECT 3369.520 2230.695 3369.780 2231.015 ;
        RECT 3384.350 2230.660 3385.320 2230.920 ;
      LAYER via ;
        RECT 3369.520 2230.725 3369.780 2230.985 ;
        RECT 3384.410 2230.660 3385.260 2230.920 ;
      LAYER met2 ;
        RECT 3369.490 2230.865 3369.810 2230.985 ;
        RECT 3384.410 2230.865 3385.260 2230.950 ;
        RECT 3365.990 2230.725 3385.260 2230.865 ;
        RECT 3384.410 2230.630 3385.260 2230.725 ;
    END
  END mgmt_io_out_buf[5]
  PIN mgmt_io_out_unbuf[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.750 2196.660 3384.950 2197.760 ;
      LAYER mcon ;
        RECT 3384.750 2196.670 3384.920 2197.760 ;
      LAYER met1 ;
        RECT 3363.940 2196.930 3364.200 2197.250 ;
        RECT 3364.060 1188.225 3364.200 2196.930 ;
        RECT 3384.700 2196.610 3384.960 2197.820 ;
        RECT 3363.780 1188.085 3364.200 1188.225 ;
        RECT 3363.780 1185.250 3363.920 1188.085 ;
      LAYER via ;
        RECT 3363.940 2196.960 3364.200 2197.220 ;
        RECT 3384.700 2196.670 3384.960 2197.760 ;
      LAYER met2 ;
        RECT 3363.910 2197.100 3364.230 2197.220 ;
        RECT 3384.670 2197.100 3384.990 2197.760 ;
        RECT 3363.750 2196.960 3384.990 2197.100 ;
        RECT 3384.670 2196.670 3384.990 2196.960 ;
    END
  END mgmt_io_out_unbuf[0]
  PIN mgmt_io_out_unbuf[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.750 2202.640 3384.950 2203.740 ;
      LAYER mcon ;
        RECT 3384.750 2202.650 3384.920 2203.740 ;
      LAYER met1 ;
        RECT 3365.060 2202.910 3365.320 2203.230 ;
        RECT 3365.180 1186.500 3365.320 2202.910 ;
        RECT 3384.700 2202.590 3384.960 2203.800 ;
        RECT 3364.900 1186.360 3365.320 1186.500 ;
        RECT 3364.900 1183.250 3365.040 1186.360 ;
      LAYER via ;
        RECT 3365.060 2202.940 3365.320 2203.200 ;
        RECT 3384.700 2202.650 3384.960 2203.740 ;
      LAYER met2 ;
        RECT 3365.030 2203.080 3365.350 2203.200 ;
        RECT 3384.670 2203.080 3384.990 2203.740 ;
        RECT 3364.900 2202.940 3384.990 2203.080 ;
        RECT 3384.670 2202.650 3384.990 2202.940 ;
    END
  END mgmt_io_out_unbuf[1]
  PIN mgmt_io_out_unbuf[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.750 2208.620 3384.950 2209.720 ;
      LAYER mcon ;
        RECT 3384.750 2208.630 3384.920 2209.720 ;
      LAYER met1 ;
        RECT 3366.180 2208.890 3366.440 2209.210 ;
        RECT 3366.300 1184.485 3366.440 2208.890 ;
        RECT 3384.700 2208.570 3384.960 2209.780 ;
        RECT 3366.020 1184.345 3366.440 1184.485 ;
        RECT 3366.020 1181.250 3366.160 1184.345 ;
      LAYER via ;
        RECT 3366.180 2208.920 3366.440 2209.180 ;
        RECT 3384.700 2208.630 3384.960 2209.720 ;
      LAYER met2 ;
        RECT 3366.150 2209.060 3366.470 2209.180 ;
        RECT 3384.670 2209.060 3384.990 2209.720 ;
        RECT 3365.990 2208.920 3384.990 2209.060 ;
        RECT 3384.670 2208.630 3384.990 2208.920 ;
    END
  END mgmt_io_out_unbuf[2]
  PIN mgmt_io_out_unbuf[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.750 2214.600 3384.950 2215.700 ;
      LAYER mcon ;
        RECT 3384.750 2214.610 3384.920 2215.700 ;
      LAYER met1 ;
        RECT 3367.300 2214.870 3367.560 2215.190 ;
        RECT 3367.420 1182.440 3367.560 2214.870 ;
        RECT 3384.700 2214.550 3384.960 2215.760 ;
        RECT 3367.140 1182.300 3367.560 1182.440 ;
        RECT 3367.140 1179.250 3367.280 1182.300 ;
      LAYER via ;
        RECT 3367.300 2214.900 3367.560 2215.160 ;
        RECT 3384.700 2214.610 3384.960 2215.700 ;
      LAYER met2 ;
        RECT 3367.270 2215.040 3367.590 2215.160 ;
        RECT 3384.670 2215.040 3384.990 2215.700 ;
        RECT 3365.990 2214.900 3384.990 2215.040 ;
        RECT 3384.670 2214.610 3384.990 2214.900 ;
    END
  END mgmt_io_out_unbuf[3]
  PIN mgmt_io_out_unbuf[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.750 2220.580 3384.950 2221.680 ;
      LAYER mcon ;
        RECT 3384.750 2220.590 3384.920 2221.680 ;
      LAYER met1 ;
        RECT 3368.420 2220.850 3368.680 2221.170 ;
        RECT 3368.540 1180.470 3368.680 2220.850 ;
        RECT 3384.700 2220.530 3384.960 2221.740 ;
        RECT 3368.260 1180.330 3368.680 1180.470 ;
        RECT 3368.260 1177.250 3368.400 1180.330 ;
      LAYER via ;
        RECT 3368.420 2220.880 3368.680 2221.140 ;
        RECT 3384.700 2220.590 3384.960 2221.680 ;
      LAYER met2 ;
        RECT 3368.390 2221.020 3368.710 2221.140 ;
        RECT 3384.670 2221.020 3384.990 2221.680 ;
        RECT 3365.990 2220.880 3384.990 2221.020 ;
        RECT 3384.670 2220.590 3384.990 2220.880 ;
    END
  END mgmt_io_out_unbuf[4]
  PIN mgmt_io_out_unbuf[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.750 2226.560 3384.950 2227.660 ;
      LAYER mcon ;
        RECT 3384.750 2226.570 3384.920 2227.660 ;
      LAYER met1 ;
        RECT 3369.540 2226.830 3369.800 2227.150 ;
        RECT 3369.660 1178.500 3369.800 2226.830 ;
        RECT 3384.700 2226.510 3384.960 2227.720 ;
        RECT 3369.380 1178.360 3369.800 1178.500 ;
        RECT 3369.380 1175.250 3369.520 1178.360 ;
      LAYER via ;
        RECT 3369.540 2226.860 3369.800 2227.120 ;
        RECT 3384.700 2226.570 3384.960 2227.660 ;
      LAYER met2 ;
        RECT 3369.510 2227.000 3369.830 2227.120 ;
        RECT 3384.670 2227.000 3384.990 2227.660 ;
        RECT 3365.990 2226.860 3384.990 2227.000 ;
        RECT 3384.670 2226.570 3384.990 2226.860 ;
    END
  END mgmt_io_out_unbuf[5]
  PIN mgmt_io_out_unbuf[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.750 2232.540 3384.950 2233.640 ;
      LAYER mcon ;
        RECT 3384.750 2232.550 3384.920 2233.640 ;
      LAYER met1 ;
        RECT 3370.660 2232.810 3370.920 2233.130 ;
        RECT 3370.780 1176.490 3370.920 2232.810 ;
        RECT 3384.700 2232.490 3384.960 2233.700 ;
        RECT 3370.500 1176.350 3370.920 1176.490 ;
        RECT 3370.500 1173.250 3370.640 1176.350 ;
      LAYER via ;
        RECT 3370.660 2232.840 3370.920 2233.100 ;
        RECT 3384.700 2232.550 3384.960 2233.640 ;
      LAYER met2 ;
        RECT 3370.630 2232.980 3370.950 2233.100 ;
        RECT 3384.670 2232.980 3384.990 2233.640 ;
        RECT 3365.990 2232.840 3384.990 2232.980 ;
        RECT 3384.670 2232.550 3384.990 2232.840 ;
    END
  END mgmt_io_out_unbuf[6]
  PIN mgmt_io_in_buf[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3380.840 2235.895 3381.490 2236.065 ;
        RECT 3381.320 2235.225 3381.490 2235.895 ;
        RECT 3380.840 2235.055 3381.490 2235.225 ;
        RECT 3381.320 2234.385 3381.490 2235.055 ;
        RECT 3380.840 2234.215 3381.490 2234.385 ;
        RECT 3381.320 2233.630 3381.490 2234.215 ;
        RECT 3382.030 2235.895 3383.050 2236.065 ;
        RECT 3382.030 2235.225 3382.200 2235.895 ;
        RECT 3382.030 2235.055 3383.050 2235.225 ;
        RECT 3382.030 2234.385 3382.200 2235.055 ;
        RECT 3382.030 2234.215 3383.050 2234.385 ;
        RECT 3382.030 2233.630 3382.200 2234.215 ;
        RECT 3381.320 2233.545 3382.200 2233.630 ;
        RECT 3380.840 2233.375 3383.050 2233.545 ;
      LAYER mcon ;
        RECT 3381.350 2233.460 3382.200 2233.630 ;
      LAYER met1 ;
        RECT 3370.940 2233.430 3371.200 2233.750 ;
        RECT 3371.060 1172.250 3371.200 2233.430 ;
        RECT 3381.290 2233.410 3382.260 2233.670 ;
      LAYER via ;
        RECT 3370.940 2233.460 3371.200 2233.720 ;
        RECT 3381.350 2233.410 3382.200 2233.670 ;
      LAYER met2 ;
        RECT 3370.910 2233.600 3371.230 2233.720 ;
        RECT 3381.350 2233.600 3382.200 2233.700 ;
        RECT 3365.990 2233.460 3382.200 2233.600 ;
        RECT 3381.350 2233.380 3382.200 2233.460 ;
    END
  END mgmt_io_in_buf[6]
  PIN mgmt_io_in_buf[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3380.840 2229.915 3381.490 2230.085 ;
        RECT 3381.320 2229.245 3381.490 2229.915 ;
        RECT 3380.840 2229.075 3381.490 2229.245 ;
        RECT 3381.320 2228.405 3381.490 2229.075 ;
        RECT 3380.840 2228.235 3381.490 2228.405 ;
        RECT 3381.320 2227.650 3381.490 2228.235 ;
        RECT 3382.030 2229.915 3383.050 2230.085 ;
        RECT 3382.030 2229.245 3382.200 2229.915 ;
        RECT 3382.030 2229.075 3383.050 2229.245 ;
        RECT 3382.030 2228.405 3382.200 2229.075 ;
        RECT 3382.030 2228.235 3383.050 2228.405 ;
        RECT 3382.030 2227.650 3382.200 2228.235 ;
        RECT 3381.320 2227.565 3382.200 2227.650 ;
        RECT 3380.840 2227.395 3383.050 2227.565 ;
      LAYER mcon ;
        RECT 3381.350 2227.480 3382.200 2227.650 ;
      LAYER met1 ;
        RECT 3369.820 2227.450 3370.080 2227.770 ;
        RECT 3369.940 1174.250 3370.080 2227.450 ;
        RECT 3381.290 2227.430 3382.260 2227.690 ;
      LAYER via ;
        RECT 3369.820 2227.480 3370.080 2227.740 ;
        RECT 3381.350 2227.430 3382.200 2227.690 ;
      LAYER met2 ;
        RECT 3369.790 2227.620 3370.110 2227.740 ;
        RECT 3381.350 2227.620 3382.200 2227.720 ;
        RECT 3365.990 2227.480 3382.200 2227.620 ;
        RECT 3381.350 2227.400 3382.200 2227.480 ;
    END
  END mgmt_io_in_buf[5]
  PIN mgmt_io_in_buf[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3380.840 2223.935 3381.490 2224.105 ;
        RECT 3381.320 2223.265 3381.490 2223.935 ;
        RECT 3380.840 2223.095 3381.490 2223.265 ;
        RECT 3381.320 2222.425 3381.490 2223.095 ;
        RECT 3380.840 2222.255 3381.490 2222.425 ;
        RECT 3381.320 2221.670 3381.490 2222.255 ;
        RECT 3382.030 2223.935 3383.050 2224.105 ;
        RECT 3382.030 2223.265 3382.200 2223.935 ;
        RECT 3382.030 2223.095 3383.050 2223.265 ;
        RECT 3382.030 2222.425 3382.200 2223.095 ;
        RECT 3382.030 2222.255 3383.050 2222.425 ;
        RECT 3382.030 2221.670 3382.200 2222.255 ;
        RECT 3381.320 2221.585 3382.200 2221.670 ;
        RECT 3380.840 2221.415 3383.050 2221.585 ;
      LAYER mcon ;
        RECT 3381.350 2221.500 3382.200 2221.670 ;
      LAYER met1 ;
        RECT 3368.700 2221.470 3368.960 2221.790 ;
        RECT 3368.820 1176.250 3368.960 2221.470 ;
        RECT 3381.290 2221.450 3382.260 2221.710 ;
      LAYER via ;
        RECT 3368.700 2221.500 3368.960 2221.760 ;
        RECT 3381.350 2221.450 3382.200 2221.710 ;
      LAYER met2 ;
        RECT 3368.670 2221.640 3368.990 2221.760 ;
        RECT 3381.350 2221.640 3382.200 2221.740 ;
        RECT 3365.990 2221.500 3382.200 2221.640 ;
        RECT 3381.350 2221.420 3382.200 2221.500 ;
    END
  END mgmt_io_in_buf[4]
  PIN mgmt_io_in_buf[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3380.840 2217.955 3381.490 2218.125 ;
        RECT 3381.320 2217.285 3381.490 2217.955 ;
        RECT 3380.840 2217.115 3381.490 2217.285 ;
        RECT 3381.320 2216.445 3381.490 2217.115 ;
        RECT 3380.840 2216.275 3381.490 2216.445 ;
        RECT 3381.320 2215.690 3381.490 2216.275 ;
        RECT 3382.030 2217.955 3383.050 2218.125 ;
        RECT 3382.030 2217.285 3382.200 2217.955 ;
        RECT 3382.030 2217.115 3383.050 2217.285 ;
        RECT 3382.030 2216.445 3382.200 2217.115 ;
        RECT 3382.030 2216.275 3383.050 2216.445 ;
        RECT 3382.030 2215.690 3382.200 2216.275 ;
        RECT 3381.320 2215.605 3382.200 2215.690 ;
        RECT 3380.840 2215.435 3383.050 2215.605 ;
      LAYER mcon ;
        RECT 3381.350 2215.520 3382.200 2215.690 ;
      LAYER met1 ;
        RECT 3367.580 2215.490 3367.840 2215.810 ;
        RECT 3367.700 1178.250 3367.840 2215.490 ;
        RECT 3381.290 2215.470 3382.260 2215.730 ;
      LAYER via ;
        RECT 3367.580 2215.520 3367.840 2215.780 ;
        RECT 3381.350 2215.470 3382.200 2215.730 ;
      LAYER met2 ;
        RECT 3367.550 2215.660 3367.870 2215.780 ;
        RECT 3381.350 2215.660 3382.200 2215.760 ;
        RECT 3365.990 2215.520 3382.200 2215.660 ;
        RECT 3381.350 2215.440 3382.200 2215.520 ;
    END
  END mgmt_io_in_buf[3]
  PIN mgmt_io_in_buf[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3380.840 2211.975 3381.490 2212.145 ;
        RECT 3381.320 2211.305 3381.490 2211.975 ;
        RECT 3380.840 2211.135 3381.490 2211.305 ;
        RECT 3381.320 2210.465 3381.490 2211.135 ;
        RECT 3380.840 2210.295 3381.490 2210.465 ;
        RECT 3381.320 2209.710 3381.490 2210.295 ;
        RECT 3382.030 2211.975 3383.050 2212.145 ;
        RECT 3382.030 2211.305 3382.200 2211.975 ;
        RECT 3382.030 2211.135 3383.050 2211.305 ;
        RECT 3382.030 2210.465 3382.200 2211.135 ;
        RECT 3382.030 2210.295 3383.050 2210.465 ;
        RECT 3382.030 2209.710 3382.200 2210.295 ;
        RECT 3381.320 2209.625 3382.200 2209.710 ;
        RECT 3380.840 2209.455 3383.050 2209.625 ;
      LAYER mcon ;
        RECT 3381.350 2209.540 3382.200 2209.710 ;
      LAYER met1 ;
        RECT 3366.460 2209.510 3366.720 2209.830 ;
        RECT 3366.580 1180.250 3366.720 2209.510 ;
        RECT 3381.290 2209.490 3382.260 2209.750 ;
      LAYER via ;
        RECT 3366.460 2209.540 3366.720 2209.800 ;
        RECT 3381.350 2209.490 3382.200 2209.750 ;
      LAYER met2 ;
        RECT 3366.430 2209.680 3366.750 2209.800 ;
        RECT 3381.350 2209.680 3382.200 2209.780 ;
        RECT 3365.990 2209.540 3382.200 2209.680 ;
        RECT 3381.350 2209.460 3382.200 2209.540 ;
    END
  END mgmt_io_in_buf[2]
  PIN mgmt_io_in_buf[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3380.840 2205.995 3381.490 2206.165 ;
        RECT 3381.320 2205.325 3381.490 2205.995 ;
        RECT 3380.840 2205.155 3381.490 2205.325 ;
        RECT 3381.320 2204.485 3381.490 2205.155 ;
        RECT 3380.840 2204.315 3381.490 2204.485 ;
        RECT 3381.320 2203.730 3381.490 2204.315 ;
        RECT 3382.030 2205.995 3383.050 2206.165 ;
        RECT 3382.030 2205.325 3382.200 2205.995 ;
        RECT 3382.030 2205.155 3383.050 2205.325 ;
        RECT 3382.030 2204.485 3382.200 2205.155 ;
        RECT 3382.030 2204.315 3383.050 2204.485 ;
        RECT 3382.030 2203.730 3382.200 2204.315 ;
        RECT 3381.320 2203.645 3382.200 2203.730 ;
        RECT 3380.840 2203.475 3383.050 2203.645 ;
      LAYER mcon ;
        RECT 3381.350 2203.560 3382.200 2203.730 ;
      LAYER met1 ;
        RECT 3365.340 2203.530 3365.600 2203.850 ;
        RECT 3365.460 1182.250 3365.600 2203.530 ;
        RECT 3381.290 2203.510 3382.260 2203.770 ;
      LAYER via ;
        RECT 3365.340 2203.560 3365.600 2203.820 ;
        RECT 3381.350 2203.510 3382.200 2203.770 ;
      LAYER met2 ;
        RECT 3365.310 2203.700 3365.630 2203.820 ;
        RECT 3381.350 2203.700 3382.200 2203.800 ;
        RECT 3364.900 2203.560 3382.200 2203.700 ;
        RECT 3381.350 2203.480 3382.200 2203.560 ;
    END
  END mgmt_io_in_buf[1]
  PIN mgmt_io_in_buf[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3380.840 2200.015 3381.490 2200.185 ;
        RECT 3381.320 2199.345 3381.490 2200.015 ;
        RECT 3380.840 2199.175 3381.490 2199.345 ;
        RECT 3381.320 2198.505 3381.490 2199.175 ;
        RECT 3380.840 2198.335 3381.490 2198.505 ;
        RECT 3381.320 2197.750 3381.490 2198.335 ;
        RECT 3382.030 2200.015 3383.050 2200.185 ;
        RECT 3382.030 2199.345 3382.200 2200.015 ;
        RECT 3382.030 2199.175 3383.050 2199.345 ;
        RECT 3382.030 2198.505 3382.200 2199.175 ;
        RECT 3382.030 2198.335 3383.050 2198.505 ;
        RECT 3382.030 2197.750 3382.200 2198.335 ;
        RECT 3381.320 2197.665 3382.200 2197.750 ;
        RECT 3380.840 2197.495 3383.050 2197.665 ;
      LAYER mcon ;
        RECT 3381.350 2197.580 3382.200 2197.750 ;
      LAYER met1 ;
        RECT 3364.220 2197.550 3364.480 2197.870 ;
        RECT 3364.340 1184.250 3364.480 2197.550 ;
        RECT 3381.290 2197.530 3382.260 2197.790 ;
      LAYER via ;
        RECT 3364.220 2197.580 3364.480 2197.840 ;
        RECT 3381.350 2197.530 3382.200 2197.790 ;
      LAYER met2 ;
        RECT 3364.190 2197.720 3364.510 2197.840 ;
        RECT 3381.350 2197.720 3382.200 2197.820 ;
        RECT 3363.750 2197.580 3382.200 2197.720 ;
        RECT 3381.350 2197.500 3382.200 2197.580 ;
    END
  END mgmt_io_in_buf[0]
  PIN mgmt_io_out_buf[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.225 3013.485 204.435 3013.655 ;
        RECT 202.705 3013.400 203.585 3013.485 ;
        RECT 202.705 3012.815 202.875 3013.400 ;
        RECT 202.225 3012.645 202.875 3012.815 ;
        RECT 202.705 3011.975 202.875 3012.645 ;
        RECT 202.225 3011.805 202.875 3011.975 ;
        RECT 202.705 3011.135 202.875 3011.805 ;
        RECT 202.225 3010.965 202.875 3011.135 ;
        RECT 203.415 3012.815 203.585 3013.400 ;
        RECT 203.415 3012.645 204.435 3012.815 ;
        RECT 203.415 3011.975 203.585 3012.645 ;
        RECT 203.415 3011.805 204.435 3011.975 ;
        RECT 203.415 3011.135 203.585 3011.805 ;
        RECT 203.415 3010.965 204.435 3011.135 ;
      LAYER mcon ;
        RECT 202.735 3013.400 203.585 3013.570 ;
      LAYER met1 ;
        RECT 218.315 3059.235 218.455 3061.780 ;
        RECT 218.035 3059.095 218.455 3059.235 ;
        RECT 218.035 3013.705 218.175 3059.095 ;
        RECT 202.675 3013.350 203.645 3013.610 ;
        RECT 217.915 3013.385 218.175 3013.705 ;
      LAYER via ;
        RECT 202.735 3013.350 203.585 3013.610 ;
        RECT 217.915 3013.415 218.175 3013.675 ;
      LAYER met2 ;
        RECT 202.735 3013.555 203.585 3013.640 ;
        RECT 217.885 3013.555 218.205 3013.675 ;
        RECT 202.735 3013.415 221.600 3013.555 ;
        RECT 202.735 3013.320 203.585 3013.415 ;
    END
  END mgmt_io_out_buf[7]
  PIN mgmt_io_out_buf[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.225 3007.505 204.435 3007.675 ;
        RECT 202.705 3007.420 203.585 3007.505 ;
        RECT 202.705 3006.835 202.875 3007.420 ;
        RECT 202.225 3006.665 202.875 3006.835 ;
        RECT 202.705 3005.995 202.875 3006.665 ;
        RECT 202.225 3005.825 202.875 3005.995 ;
        RECT 202.705 3005.155 202.875 3005.825 ;
        RECT 202.225 3004.985 202.875 3005.155 ;
        RECT 203.415 3006.835 203.585 3007.420 ;
        RECT 203.415 3006.665 204.435 3006.835 ;
        RECT 203.415 3005.995 203.585 3006.665 ;
        RECT 203.415 3005.825 204.435 3005.995 ;
        RECT 203.415 3005.155 203.585 3005.825 ;
        RECT 203.415 3004.985 204.435 3005.155 ;
      LAYER mcon ;
        RECT 202.735 3007.420 203.585 3007.590 ;
      LAYER met1 ;
        RECT 219.435 3057.210 219.575 3059.780 ;
        RECT 219.155 3057.070 219.575 3057.210 ;
        RECT 219.155 3007.725 219.295 3057.070 ;
        RECT 202.675 3007.370 203.645 3007.630 ;
        RECT 219.035 3007.405 219.295 3007.725 ;
      LAYER via ;
        RECT 202.735 3007.370 203.585 3007.630 ;
        RECT 219.035 3007.435 219.295 3007.695 ;
      LAYER met2 ;
        RECT 202.735 3007.575 203.585 3007.660 ;
        RECT 219.005 3007.575 219.325 3007.695 ;
        RECT 202.735 3007.435 221.600 3007.575 ;
        RECT 202.735 3007.340 203.585 3007.435 ;
    END
  END mgmt_io_out_buf[8]
  PIN mgmt_io_out_buf[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.225 3001.525 204.435 3001.695 ;
        RECT 202.705 3001.440 203.585 3001.525 ;
        RECT 202.705 3000.855 202.875 3001.440 ;
        RECT 202.225 3000.685 202.875 3000.855 ;
        RECT 202.705 3000.015 202.875 3000.685 ;
        RECT 202.225 2999.845 202.875 3000.015 ;
        RECT 202.705 2999.175 202.875 2999.845 ;
        RECT 202.225 2999.005 202.875 2999.175 ;
        RECT 203.415 3000.855 203.585 3001.440 ;
        RECT 203.415 3000.685 204.435 3000.855 ;
        RECT 203.415 3000.015 203.585 3000.685 ;
        RECT 203.415 2999.845 204.435 3000.015 ;
        RECT 203.415 2999.175 203.585 2999.845 ;
        RECT 203.415 2999.005 204.435 2999.175 ;
      LAYER mcon ;
        RECT 202.735 3001.440 203.585 3001.610 ;
      LAYER met1 ;
        RECT 220.555 3055.155 220.695 3057.780 ;
        RECT 220.275 3055.015 220.695 3055.155 ;
        RECT 220.275 3001.745 220.415 3055.015 ;
        RECT 202.675 3001.390 203.645 3001.650 ;
        RECT 220.155 3001.425 220.415 3001.745 ;
      LAYER via ;
        RECT 202.735 3001.390 203.585 3001.650 ;
        RECT 220.155 3001.455 220.415 3001.715 ;
      LAYER met2 ;
        RECT 202.735 3001.595 203.585 3001.680 ;
        RECT 220.125 3001.595 220.445 3001.715 ;
        RECT 202.735 3001.455 221.600 3001.595 ;
        RECT 202.735 3001.360 203.585 3001.455 ;
    END
  END mgmt_io_out_buf[9]
  PIN mgmt_io_out_buf[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.225 2995.545 204.435 2995.715 ;
        RECT 202.705 2995.460 203.585 2995.545 ;
        RECT 202.705 2994.875 202.875 2995.460 ;
        RECT 202.225 2994.705 202.875 2994.875 ;
        RECT 202.705 2994.035 202.875 2994.705 ;
        RECT 202.225 2993.865 202.875 2994.035 ;
        RECT 202.705 2993.195 202.875 2993.865 ;
        RECT 202.225 2993.025 202.875 2993.195 ;
        RECT 203.415 2994.875 203.585 2995.460 ;
        RECT 203.415 2994.705 204.435 2994.875 ;
        RECT 203.415 2994.035 203.585 2994.705 ;
        RECT 203.415 2993.865 204.435 2994.035 ;
        RECT 203.415 2993.195 203.585 2993.865 ;
        RECT 203.415 2993.025 204.435 2993.195 ;
      LAYER mcon ;
        RECT 202.735 2995.460 203.585 2995.630 ;
      LAYER met1 ;
        RECT 221.675 3053.175 221.815 3055.780 ;
        RECT 221.395 3053.035 221.815 3053.175 ;
        RECT 221.395 2995.765 221.535 3053.035 ;
        RECT 202.675 2995.410 203.645 2995.670 ;
        RECT 221.275 2995.445 221.535 2995.765 ;
      LAYER via ;
        RECT 202.735 2995.410 203.585 2995.670 ;
        RECT 221.275 2995.475 221.535 2995.735 ;
      LAYER met2 ;
        RECT 202.735 2995.615 203.585 2995.700 ;
        RECT 221.245 2995.615 221.565 2995.735 ;
        RECT 202.735 2995.475 221.605 2995.615 ;
        RECT 202.735 2995.380 203.585 2995.475 ;
    END
  END mgmt_io_out_buf[10]
  PIN mgmt_io_out_buf[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.225 2989.565 204.435 2989.735 ;
        RECT 202.705 2989.480 203.585 2989.565 ;
        RECT 202.705 2988.895 202.875 2989.480 ;
        RECT 202.225 2988.725 202.875 2988.895 ;
        RECT 202.705 2988.055 202.875 2988.725 ;
        RECT 202.225 2987.885 202.875 2988.055 ;
        RECT 202.705 2987.215 202.875 2987.885 ;
        RECT 202.225 2987.045 202.875 2987.215 ;
        RECT 203.415 2988.895 203.585 2989.480 ;
        RECT 203.415 2988.725 204.435 2988.895 ;
        RECT 203.415 2988.055 203.585 2988.725 ;
        RECT 203.415 2987.885 204.435 2988.055 ;
        RECT 203.415 2987.215 203.585 2987.885 ;
        RECT 203.415 2987.045 204.435 2987.215 ;
      LAYER mcon ;
        RECT 202.735 2989.480 203.585 2989.650 ;
      LAYER met1 ;
        RECT 222.795 3051.110 222.935 3053.780 ;
        RECT 222.515 3050.970 222.935 3051.110 ;
        RECT 222.515 2989.785 222.655 3050.970 ;
        RECT 202.675 2989.430 203.645 2989.690 ;
        RECT 222.395 2989.465 222.655 2989.785 ;
      LAYER via ;
        RECT 202.735 2989.430 203.585 2989.690 ;
        RECT 222.395 2989.495 222.655 2989.755 ;
      LAYER met2 ;
        RECT 202.735 2989.635 203.585 2989.720 ;
        RECT 222.365 2989.635 222.685 2989.755 ;
        RECT 202.735 2989.495 222.720 2989.635 ;
        RECT 202.735 2989.400 203.585 2989.495 ;
    END
  END mgmt_io_out_buf[11]
  PIN mgmt_io_in_unbuf[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 206.135 2989.470 206.335 2991.060 ;
      LAYER mcon ;
        RECT 206.135 2989.970 206.305 2991.060 ;
      LAYER met1 ;
        RECT 206.095 2989.910 206.355 2991.120 ;
        RECT 222.235 2990.755 222.375 3054.780 ;
        RECT 222.115 2990.435 222.375 2990.755 ;
      LAYER via ;
        RECT 206.095 2989.970 206.355 2991.060 ;
        RECT 222.115 2990.465 222.375 2990.725 ;
      LAYER met2 ;
        RECT 206.065 2990.605 206.385 2991.060 ;
        RECT 222.085 2990.605 222.405 2990.725 ;
        RECT 206.065 2990.465 222.720 2990.605 ;
        RECT 206.065 2989.970 206.385 2990.465 ;
    END
  END mgmt_io_in_unbuf[11]
  PIN mgmt_io_in_unbuf[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 206.135 2995.450 206.335 2997.040 ;
      LAYER mcon ;
        RECT 206.135 2995.950 206.305 2997.040 ;
      LAYER met1 ;
        RECT 206.095 2995.890 206.355 2997.100 ;
        RECT 221.115 2996.735 221.255 3056.780 ;
        RECT 220.995 2996.415 221.255 2996.735 ;
      LAYER via ;
        RECT 206.095 2995.950 206.355 2997.040 ;
        RECT 220.995 2996.445 221.255 2996.705 ;
      LAYER met2 ;
        RECT 206.065 2996.585 206.385 2997.040 ;
        RECT 220.965 2996.585 221.285 2996.705 ;
        RECT 206.065 2996.445 221.605 2996.585 ;
        RECT 206.065 2995.950 206.385 2996.445 ;
    END
  END mgmt_io_in_unbuf[10]
  PIN mgmt_io_in_unbuf[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 206.135 3001.430 206.335 3003.020 ;
      LAYER mcon ;
        RECT 206.135 3001.930 206.305 3003.020 ;
      LAYER met1 ;
        RECT 206.095 3001.870 206.355 3003.080 ;
        RECT 219.995 3002.715 220.135 3058.780 ;
        RECT 219.875 3002.395 220.135 3002.715 ;
      LAYER via ;
        RECT 206.095 3001.930 206.355 3003.020 ;
        RECT 219.875 3002.425 220.135 3002.685 ;
      LAYER met2 ;
        RECT 206.065 3002.565 206.385 3003.020 ;
        RECT 219.845 3002.565 220.165 3002.685 ;
        RECT 206.065 3002.425 221.600 3002.565 ;
        RECT 206.065 3001.930 206.385 3002.425 ;
    END
  END mgmt_io_in_unbuf[9]
  PIN mgmt_io_in_unbuf[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 206.135 3007.410 206.335 3009.000 ;
      LAYER mcon ;
        RECT 206.135 3007.910 206.305 3009.000 ;
      LAYER met1 ;
        RECT 206.095 3007.850 206.355 3009.060 ;
        RECT 218.875 3008.695 219.015 3060.780 ;
        RECT 218.755 3008.375 219.015 3008.695 ;
      LAYER via ;
        RECT 206.095 3007.910 206.355 3009.000 ;
        RECT 218.755 3008.405 219.015 3008.665 ;
      LAYER met2 ;
        RECT 206.065 3008.545 206.385 3009.000 ;
        RECT 218.725 3008.545 219.045 3008.665 ;
        RECT 206.065 3008.405 221.600 3008.545 ;
        RECT 206.065 3007.910 206.385 3008.405 ;
    END
  END mgmt_io_in_unbuf[8]
  PIN mgmt_io_in_unbuf[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 206.135 3013.390 206.335 3014.980 ;
      LAYER mcon ;
        RECT 206.135 3013.890 206.305 3014.980 ;
      LAYER met1 ;
        RECT 206.095 3013.830 206.355 3015.040 ;
        RECT 217.755 3014.675 217.895 3062.780 ;
        RECT 217.635 3014.355 217.895 3014.675 ;
      LAYER via ;
        RECT 206.095 3013.890 206.355 3014.980 ;
        RECT 217.635 3014.385 217.895 3014.645 ;
      LAYER met2 ;
        RECT 206.065 3014.525 206.385 3014.980 ;
        RECT 217.605 3014.525 217.925 3014.645 ;
        RECT 206.065 3014.385 221.600 3014.525 ;
        RECT 206.065 3013.890 206.385 3014.385 ;
    END
  END mgmt_io_in_unbuf[7]
  PIN mgmt_io_out_buf[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.335 1695.680 204.545 1695.850 ;
        RECT 202.815 1695.595 203.695 1695.680 ;
        RECT 202.815 1695.010 202.985 1695.595 ;
        RECT 202.335 1694.840 202.985 1695.010 ;
        RECT 202.815 1694.170 202.985 1694.840 ;
        RECT 202.335 1694.000 202.985 1694.170 ;
        RECT 202.815 1693.330 202.985 1694.000 ;
        RECT 202.335 1693.160 202.985 1693.330 ;
        RECT 203.525 1695.010 203.695 1695.595 ;
        RECT 203.525 1694.840 204.545 1695.010 ;
        RECT 203.525 1694.170 203.695 1694.840 ;
        RECT 203.525 1694.000 204.545 1694.170 ;
        RECT 203.525 1693.330 203.695 1694.000 ;
        RECT 203.525 1693.160 204.545 1693.330 ;
      LAYER mcon ;
        RECT 202.845 1695.595 203.695 1695.765 ;
      LAYER met1 ;
        RECT 223.775 1769.515 223.915 1772.650 ;
        RECT 223.495 1769.375 223.915 1769.515 ;
        RECT 223.495 1695.900 223.635 1769.375 ;
        RECT 202.785 1695.545 203.755 1695.805 ;
        RECT 223.375 1695.580 223.635 1695.900 ;
      LAYER via ;
        RECT 202.845 1695.545 203.695 1695.805 ;
        RECT 223.375 1695.610 223.635 1695.870 ;
      LAYER met2 ;
        RECT 202.845 1695.750 203.695 1695.835 ;
        RECT 223.345 1695.750 223.665 1695.870 ;
        RECT 202.845 1695.610 223.840 1695.750 ;
        RECT 202.845 1695.515 203.695 1695.610 ;
    END
  END mgmt_io_out_buf[12]
  PIN mgmt_io_out_buf[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.335 1689.700 204.545 1689.870 ;
        RECT 202.815 1689.615 203.695 1689.700 ;
        RECT 202.815 1689.030 202.985 1689.615 ;
        RECT 202.335 1688.860 202.985 1689.030 ;
        RECT 202.815 1688.190 202.985 1688.860 ;
        RECT 202.335 1688.020 202.985 1688.190 ;
        RECT 202.815 1687.350 202.985 1688.020 ;
        RECT 202.335 1687.180 202.985 1687.350 ;
        RECT 203.525 1689.030 203.695 1689.615 ;
        RECT 203.525 1688.860 204.545 1689.030 ;
        RECT 203.525 1688.190 203.695 1688.860 ;
        RECT 203.525 1688.020 204.545 1688.190 ;
        RECT 203.525 1687.350 203.695 1688.020 ;
        RECT 203.525 1687.180 204.545 1687.350 ;
      LAYER mcon ;
        RECT 202.845 1689.615 203.695 1689.785 ;
      LAYER met1 ;
        RECT 224.895 1767.530 225.035 1770.650 ;
        RECT 224.615 1767.390 225.035 1767.530 ;
        RECT 224.615 1689.920 224.755 1767.390 ;
        RECT 202.785 1689.565 203.755 1689.825 ;
        RECT 224.495 1689.600 224.755 1689.920 ;
      LAYER via ;
        RECT 202.845 1689.565 203.695 1689.825 ;
        RECT 224.495 1689.630 224.755 1689.890 ;
      LAYER met2 ;
        RECT 202.845 1689.770 203.695 1689.855 ;
        RECT 224.465 1689.770 224.785 1689.890 ;
        RECT 202.845 1689.630 224.910 1689.770 ;
        RECT 202.845 1689.535 203.695 1689.630 ;
    END
  END mgmt_io_out_buf[13]
  PIN mgmt_io_out_buf[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.335 1683.720 204.545 1683.890 ;
        RECT 202.815 1683.635 203.695 1683.720 ;
        RECT 202.815 1683.050 202.985 1683.635 ;
        RECT 202.335 1682.880 202.985 1683.050 ;
        RECT 202.815 1682.210 202.985 1682.880 ;
        RECT 202.335 1682.040 202.985 1682.210 ;
        RECT 202.815 1681.370 202.985 1682.040 ;
        RECT 202.335 1681.200 202.985 1681.370 ;
        RECT 203.525 1683.050 203.695 1683.635 ;
        RECT 203.525 1682.880 204.545 1683.050 ;
        RECT 203.525 1682.210 203.695 1682.880 ;
        RECT 203.525 1682.040 204.545 1682.210 ;
        RECT 203.525 1681.370 203.695 1682.040 ;
        RECT 203.525 1681.200 204.545 1681.370 ;
      LAYER mcon ;
        RECT 202.845 1683.635 203.695 1683.805 ;
      LAYER met1 ;
        RECT 226.015 1765.600 226.155 1768.650 ;
        RECT 225.735 1765.460 226.155 1765.600 ;
        RECT 225.735 1683.940 225.875 1765.460 ;
        RECT 202.785 1683.585 203.755 1683.845 ;
        RECT 225.615 1683.620 225.875 1683.940 ;
      LAYER via ;
        RECT 202.845 1683.585 203.695 1683.845 ;
        RECT 225.615 1683.650 225.875 1683.910 ;
      LAYER met2 ;
        RECT 202.845 1683.790 203.695 1683.875 ;
        RECT 225.585 1683.790 225.905 1683.910 ;
        RECT 202.845 1683.650 225.975 1683.790 ;
        RECT 202.845 1683.555 203.695 1683.650 ;
    END
  END mgmt_io_out_buf[14]
  PIN mgmt_io_out_buf[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.335 1677.740 204.545 1677.910 ;
        RECT 202.815 1677.655 203.695 1677.740 ;
        RECT 202.815 1677.070 202.985 1677.655 ;
        RECT 202.335 1676.900 202.985 1677.070 ;
        RECT 202.815 1676.230 202.985 1676.900 ;
        RECT 202.335 1676.060 202.985 1676.230 ;
        RECT 202.815 1675.390 202.985 1676.060 ;
        RECT 202.335 1675.220 202.985 1675.390 ;
        RECT 203.525 1677.070 203.695 1677.655 ;
        RECT 203.525 1676.900 204.545 1677.070 ;
        RECT 203.525 1676.230 203.695 1676.900 ;
        RECT 203.525 1676.060 204.545 1676.230 ;
        RECT 203.525 1675.390 203.695 1676.060 ;
        RECT 203.525 1675.220 204.545 1675.390 ;
      LAYER mcon ;
        RECT 202.845 1677.655 203.695 1677.825 ;
      LAYER met1 ;
        RECT 227.135 1763.525 227.275 1766.650 ;
        RECT 226.855 1763.385 227.275 1763.525 ;
        RECT 226.855 1677.960 226.995 1763.385 ;
        RECT 202.785 1677.605 203.755 1677.865 ;
        RECT 226.735 1677.640 226.995 1677.960 ;
      LAYER via ;
        RECT 202.845 1677.605 203.695 1677.865 ;
        RECT 226.735 1677.670 226.995 1677.930 ;
      LAYER met2 ;
        RECT 202.845 1677.810 203.695 1677.895 ;
        RECT 226.705 1677.810 227.025 1677.930 ;
        RECT 202.845 1677.670 227.100 1677.810 ;
        RECT 202.845 1677.575 203.695 1677.670 ;
    END
  END mgmt_io_out_buf[15]
  PIN mgmt_io_in_unbuf[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 206.245 1677.645 206.445 1679.235 ;
      LAYER mcon ;
        RECT 206.245 1678.145 206.415 1679.235 ;
      LAYER met1 ;
        RECT 206.205 1678.085 206.465 1679.295 ;
        RECT 226.575 1678.930 226.715 1767.650 ;
        RECT 226.455 1678.610 226.715 1678.930 ;
      LAYER via ;
        RECT 206.205 1678.145 206.465 1679.235 ;
        RECT 226.455 1678.640 226.715 1678.900 ;
      LAYER met2 ;
        RECT 206.175 1678.780 206.495 1679.235 ;
        RECT 226.425 1678.780 226.745 1678.900 ;
        RECT 206.175 1678.640 227.100 1678.780 ;
        RECT 206.175 1678.145 206.495 1678.640 ;
    END
  END mgmt_io_in_unbuf[15]
  PIN mgmt_io_in_unbuf[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 206.245 1683.625 206.445 1685.215 ;
      LAYER mcon ;
        RECT 206.245 1684.125 206.415 1685.215 ;
      LAYER met1 ;
        RECT 206.205 1684.065 206.465 1685.275 ;
        RECT 225.455 1684.790 225.595 1769.650 ;
        RECT 225.335 1684.470 225.595 1684.790 ;
      LAYER via ;
        RECT 206.205 1684.125 206.465 1685.215 ;
        RECT 225.335 1684.500 225.595 1684.760 ;
      LAYER met2 ;
        RECT 206.175 1684.760 206.495 1685.215 ;
        RECT 206.175 1684.620 225.975 1684.760 ;
        RECT 206.175 1684.125 206.495 1684.620 ;
        RECT 225.305 1684.500 225.625 1684.620 ;
    END
  END mgmt_io_in_unbuf[14]
  PIN mgmt_io_in_unbuf[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 206.245 1689.605 206.445 1691.195 ;
      LAYER mcon ;
        RECT 206.245 1690.105 206.415 1691.195 ;
      LAYER met1 ;
        RECT 206.205 1690.045 206.465 1691.255 ;
        RECT 224.335 1690.890 224.475 1771.650 ;
        RECT 224.215 1690.570 224.475 1690.890 ;
      LAYER via ;
        RECT 206.205 1690.105 206.465 1691.195 ;
        RECT 224.215 1690.600 224.475 1690.860 ;
      LAYER met2 ;
        RECT 206.175 1690.740 206.495 1691.195 ;
        RECT 224.185 1690.740 224.505 1690.860 ;
        RECT 206.175 1690.600 224.910 1690.740 ;
        RECT 206.175 1690.105 206.495 1690.600 ;
    END
  END mgmt_io_in_unbuf[13]
  PIN mgmt_io_in_unbuf[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 206.245 1695.585 206.445 1697.175 ;
      LAYER mcon ;
        RECT 206.245 1696.085 206.415 1697.175 ;
      LAYER met1 ;
        RECT 206.205 1696.025 206.465 1697.235 ;
        RECT 223.215 1696.870 223.355 1773.650 ;
        RECT 223.095 1696.550 223.355 1696.870 ;
      LAYER via ;
        RECT 206.205 1696.085 206.465 1697.175 ;
        RECT 223.095 1696.580 223.355 1696.840 ;
      LAYER met2 ;
        RECT 206.175 1696.720 206.495 1697.175 ;
        RECT 223.065 1696.720 223.385 1696.840 ;
        RECT 206.175 1696.580 223.840 1696.720 ;
        RECT 206.175 1696.085 206.495 1696.580 ;
    END
  END mgmt_io_in_unbuf[12]
  PIN mgmt_io_out_buf[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 760.135 216.390 760.305 216.870 ;
        RECT 760.975 216.390 761.145 216.870 ;
        RECT 761.815 216.390 761.985 216.870 ;
        RECT 762.655 216.390 762.825 216.870 ;
        RECT 760.135 216.220 762.825 216.390 ;
        RECT 760.135 215.680 760.390 216.220 ;
        RECT 760.135 215.510 762.825 215.680 ;
        RECT 760.135 214.660 760.305 215.510 ;
        RECT 760.975 214.660 761.145 215.510 ;
        RECT 761.815 214.660 761.985 215.510 ;
        RECT 762.655 214.660 762.825 215.510 ;
      LAYER mcon ;
        RECT 760.220 215.510 760.390 216.360 ;
      LAYER met1 ;
        RECT 655.755 225.380 659.600 225.520 ;
        RECT 760.190 225.380 760.510 225.500 ;
        RECT 659.460 225.240 760.510 225.380 ;
        RECT 760.170 215.450 760.430 216.420 ;
      LAYER via ;
        RECT 760.220 225.240 760.480 225.500 ;
        RECT 760.170 215.510 760.430 216.360 ;
      LAYER met2 ;
        RECT 760.220 225.530 760.360 232.345 ;
        RECT 760.220 225.210 760.480 225.530 ;
        RECT 760.220 216.360 760.360 225.210 ;
        RECT 760.140 215.510 760.460 216.360 ;
    END
  END mgmt_io_out_buf[16]
  PIN mgmt_io_out_buf[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 766.115 216.390 766.285 216.870 ;
        RECT 766.955 216.390 767.125 216.870 ;
        RECT 767.795 216.390 767.965 216.870 ;
        RECT 768.635 216.390 768.805 216.870 ;
        RECT 766.115 216.220 768.805 216.390 ;
        RECT 766.115 215.680 766.370 216.220 ;
        RECT 766.115 215.510 768.805 215.680 ;
        RECT 766.115 214.660 766.285 215.510 ;
        RECT 766.955 214.660 767.125 215.510 ;
        RECT 767.795 214.660 767.965 215.510 ;
        RECT 768.635 214.660 768.805 215.510 ;
      LAYER mcon ;
        RECT 766.200 215.510 766.370 216.360 ;
      LAYER met1 ;
        RECT 657.755 224.540 661.640 224.680 ;
        RECT 766.170 224.540 766.490 224.660 ;
        RECT 661.500 224.400 766.490 224.540 ;
        RECT 766.150 215.450 766.410 216.420 ;
      LAYER via ;
        RECT 766.200 224.400 766.460 224.660 ;
        RECT 766.150 215.510 766.410 216.360 ;
      LAYER met2 ;
        RECT 766.200 224.690 766.340 232.345 ;
        RECT 766.200 224.370 766.460 224.690 ;
        RECT 766.200 216.360 766.340 224.370 ;
        RECT 766.120 215.510 766.440 216.360 ;
    END
  END mgmt_io_out_buf[17]
  PIN mgmt_io_out_buf[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 772.095 216.390 772.265 216.870 ;
        RECT 772.935 216.390 773.105 216.870 ;
        RECT 773.775 216.390 773.945 216.870 ;
        RECT 774.615 216.390 774.785 216.870 ;
        RECT 772.095 216.220 774.785 216.390 ;
        RECT 772.095 215.680 772.350 216.220 ;
        RECT 772.095 215.510 774.785 215.680 ;
        RECT 772.095 214.660 772.265 215.510 ;
        RECT 772.935 214.660 773.105 215.510 ;
        RECT 773.775 214.660 773.945 215.510 ;
        RECT 774.615 214.660 774.785 215.510 ;
      LAYER mcon ;
        RECT 772.180 215.510 772.350 216.360 ;
      LAYER met1 ;
        RECT 659.755 223.700 663.635 223.840 ;
        RECT 772.150 223.700 772.470 223.820 ;
        RECT 663.495 223.560 772.470 223.700 ;
        RECT 772.130 215.450 772.390 216.420 ;
      LAYER via ;
        RECT 772.180 223.560 772.440 223.820 ;
        RECT 772.130 215.510 772.390 216.360 ;
      LAYER met2 ;
        RECT 772.180 223.850 772.320 232.345 ;
        RECT 772.180 223.530 772.440 223.850 ;
        RECT 772.180 216.360 772.320 223.530 ;
        RECT 772.100 215.510 772.420 216.360 ;
    END
  END mgmt_io_out_buf[18]
  PIN mgmt_io_out_buf[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 778.075 216.390 778.245 216.870 ;
        RECT 778.915 216.390 779.085 216.870 ;
        RECT 779.755 216.390 779.925 216.870 ;
        RECT 780.595 216.390 780.765 216.870 ;
        RECT 778.075 216.220 780.765 216.390 ;
        RECT 778.075 215.680 778.330 216.220 ;
        RECT 778.075 215.510 780.765 215.680 ;
        RECT 778.075 214.660 778.245 215.510 ;
        RECT 778.915 214.660 779.085 215.510 ;
        RECT 779.755 214.660 779.925 215.510 ;
        RECT 780.595 214.660 780.765 215.510 ;
      LAYER mcon ;
        RECT 778.160 215.510 778.330 216.360 ;
      LAYER met1 ;
        RECT 661.755 222.860 665.585 223.000 ;
        RECT 778.130 222.860 778.450 222.980 ;
        RECT 665.445 222.720 778.450 222.860 ;
        RECT 778.110 215.450 778.370 216.420 ;
      LAYER via ;
        RECT 778.160 222.720 778.420 222.980 ;
        RECT 778.110 215.510 778.370 216.360 ;
      LAYER met2 ;
        RECT 778.160 223.010 778.300 232.345 ;
        RECT 778.160 222.690 778.420 223.010 ;
        RECT 778.160 216.360 778.300 222.690 ;
        RECT 778.080 215.510 778.400 216.360 ;
    END
  END mgmt_io_out_buf[19]
  PIN mgmt_io_in_unbuf[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 783.220 212.760 784.320 212.960 ;
      LAYER mcon ;
        RECT 783.230 212.790 784.320 212.960 ;
      LAYER met1 ;
        RECT 783.490 222.580 783.810 222.700 ;
        RECT 662.615 222.440 783.810 222.580 ;
        RECT 783.170 212.750 784.380 213.010 ;
      LAYER via ;
        RECT 783.520 222.440 783.780 222.700 ;
        RECT 783.230 212.750 784.320 213.010 ;
      LAYER met2 ;
        RECT 783.520 222.730 783.660 232.345 ;
        RECT 783.520 222.410 783.780 222.730 ;
        RECT 783.520 213.040 783.660 222.410 ;
        RECT 783.230 212.720 784.320 213.040 ;
    END
  END mgmt_io_in_unbuf[19]
  PIN mgmt_io_in_unbuf[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 777.240 212.760 778.340 212.960 ;
      LAYER mcon ;
        RECT 777.250 212.790 778.340 212.960 ;
      LAYER met1 ;
        RECT 777.510 223.420 777.830 223.540 ;
        RECT 660.615 223.280 777.830 223.420 ;
        RECT 777.190 212.750 778.400 213.010 ;
      LAYER via ;
        RECT 777.540 223.280 777.800 223.540 ;
        RECT 777.250 212.750 778.340 213.010 ;
      LAYER met2 ;
        RECT 777.540 223.570 777.680 232.345 ;
        RECT 777.540 223.250 777.800 223.570 ;
        RECT 777.540 213.040 777.680 223.250 ;
        RECT 777.250 212.720 778.340 213.040 ;
    END
  END mgmt_io_in_unbuf[18]
  PIN mgmt_io_in_unbuf[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 771.260 212.760 772.360 212.960 ;
      LAYER mcon ;
        RECT 771.270 212.790 772.360 212.960 ;
      LAYER met1 ;
        RECT 771.530 224.260 771.850 224.380 ;
        RECT 658.615 224.120 771.850 224.260 ;
        RECT 771.210 212.750 772.420 213.010 ;
      LAYER via ;
        RECT 771.560 224.120 771.820 224.380 ;
        RECT 771.270 212.750 772.360 213.010 ;
      LAYER met2 ;
        RECT 771.560 224.410 771.700 232.345 ;
        RECT 771.560 224.090 771.820 224.410 ;
        RECT 771.560 213.040 771.700 224.090 ;
        RECT 771.270 212.720 772.360 213.040 ;
    END
  END mgmt_io_in_unbuf[17]
  PIN mgmt_io_in_unbuf[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 765.280 212.760 766.380 212.960 ;
      LAYER mcon ;
        RECT 765.290 212.790 766.380 212.960 ;
      LAYER met1 ;
        RECT 765.550 225.100 765.870 225.220 ;
        RECT 656.615 224.960 765.870 225.100 ;
        RECT 765.230 212.750 766.440 213.010 ;
      LAYER via ;
        RECT 765.580 224.960 765.840 225.220 ;
        RECT 765.290 212.750 766.380 213.010 ;
      LAYER met2 ;
        RECT 765.580 225.250 765.720 232.345 ;
        RECT 765.580 224.930 765.840 225.250 ;
        RECT 765.580 213.040 765.720 224.930 ;
        RECT 765.290 212.720 766.380 213.040 ;
    END
  END mgmt_io_in_unbuf[16]
  PIN mgmt_io_oeb_buf[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 784.055 216.390 784.225 216.870 ;
        RECT 784.895 216.390 785.065 216.870 ;
        RECT 785.735 216.390 785.905 216.870 ;
        RECT 786.575 216.390 786.745 216.870 ;
        RECT 784.055 216.220 786.745 216.390 ;
        RECT 784.055 215.680 784.310 216.220 ;
        RECT 784.055 215.510 786.745 215.680 ;
        RECT 784.055 214.660 784.225 215.510 ;
        RECT 784.895 214.660 785.065 215.510 ;
        RECT 785.735 214.660 785.905 215.510 ;
        RECT 786.575 214.660 786.745 215.510 ;
      LAYER mcon ;
        RECT 784.140 215.510 784.310 216.360 ;
      LAYER met1 ;
        RECT 784.110 222.020 784.430 222.140 ;
        RECT 663.615 221.880 784.430 222.020 ;
        RECT 784.090 215.450 784.350 216.420 ;
      LAYER via ;
        RECT 784.140 221.880 784.400 222.140 ;
        RECT 784.090 215.510 784.350 216.360 ;
      LAYER met2 ;
        RECT 784.140 222.170 784.280 232.345 ;
        RECT 784.140 221.850 784.400 222.170 ;
        RECT 784.140 216.360 784.280 221.850 ;
        RECT 784.060 215.510 784.380 216.360 ;
    END
  END mgmt_io_oeb_buf[0]
  PIN mgmt_io_oeb_buf[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 790.035 213.300 790.205 214.150 ;
        RECT 790.875 213.300 791.045 214.150 ;
        RECT 791.715 213.300 791.885 214.150 ;
        RECT 792.555 213.300 792.725 214.150 ;
        RECT 790.035 213.130 792.725 213.300 ;
        RECT 790.035 212.590 790.290 213.130 ;
        RECT 790.035 212.420 792.725 212.590 ;
        RECT 790.035 211.940 790.205 212.420 ;
        RECT 790.875 211.940 791.045 212.420 ;
        RECT 791.715 211.940 791.885 212.420 ;
        RECT 792.555 211.940 792.725 212.420 ;
      LAYER mcon ;
        RECT 790.120 212.450 790.290 213.300 ;
      LAYER met1 ;
        RECT 789.470 221.460 789.790 221.580 ;
        RECT 664.615 221.320 789.790 221.460 ;
        RECT 790.080 212.390 790.340 213.360 ;
      LAYER via ;
        RECT 789.500 221.320 789.760 221.580 ;
        RECT 790.080 212.450 790.340 213.300 ;
      LAYER met2 ;
        RECT 789.500 221.610 789.640 232.345 ;
        RECT 789.500 221.290 789.760 221.610 ;
        RECT 789.500 214.240 789.640 221.290 ;
        RECT 789.500 214.100 790.275 214.240 ;
        RECT 790.135 213.300 790.275 214.100 ;
        RECT 790.050 212.450 790.370 213.300 ;
    END
  END mgmt_io_oeb_buf[1]
  PIN mgmt_io_oeb_buf[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 790.035 216.390 790.205 216.870 ;
        RECT 790.875 216.390 791.045 216.870 ;
        RECT 791.715 216.390 791.885 216.870 ;
        RECT 792.555 216.390 792.725 216.870 ;
        RECT 790.035 216.220 792.725 216.390 ;
        RECT 790.035 215.680 790.290 216.220 ;
        RECT 790.035 215.510 792.725 215.680 ;
        RECT 790.035 214.660 790.205 215.510 ;
        RECT 790.875 214.660 791.045 215.510 ;
        RECT 791.715 214.660 791.885 215.510 ;
        RECT 792.555 214.660 792.725 215.510 ;
      LAYER mcon ;
        RECT 790.120 215.510 790.290 216.360 ;
      LAYER met1 ;
        RECT 790.090 220.900 790.410 221.020 ;
        RECT 665.615 220.760 790.410 220.900 ;
        RECT 790.070 215.450 790.330 216.420 ;
      LAYER via ;
        RECT 790.120 220.760 790.380 221.020 ;
        RECT 790.070 215.510 790.330 216.360 ;
      LAYER met2 ;
        RECT 790.120 221.050 790.260 232.345 ;
        RECT 790.120 220.730 790.380 221.050 ;
        RECT 790.120 216.360 790.260 220.730 ;
        RECT 790.040 215.510 790.360 216.360 ;
    END
  END mgmt_io_oeb_buf[2]
  PIN mgmt_io_oeb_unbuf[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2270.340 215.850 2271.930 216.050 ;
      LAYER mcon ;
        RECT 2270.840 215.850 2271.930 216.020 ;
      LAYER met1 ;
        RECT 2271.305 221.040 2416.200 221.180 ;
        RECT 2271.305 220.920 2271.625 221.040 ;
        RECT 2270.780 215.810 2271.990 216.070 ;
        RECT 2416.060 211.780 2416.200 221.040 ;
        RECT 3377.640 212.245 3377.780 1156.450 ;
        RECT 2537.220 212.105 3377.780 212.245 ;
        RECT 2537.220 211.780 2537.360 212.105 ;
        RECT 2416.060 211.640 2537.360 211.780 ;
      LAYER via ;
        RECT 2271.335 220.920 2271.595 221.180 ;
        RECT 2270.840 215.810 2271.930 216.070 ;
      LAYER met2 ;
        RECT 2271.335 221.210 2271.475 232.485 ;
        RECT 2271.335 220.890 2271.595 221.210 ;
        RECT 2271.335 216.100 2271.475 220.890 ;
        RECT 2270.840 215.780 2271.930 216.100 ;
    END
  END mgmt_io_oeb_unbuf[2]
  PIN mgmt_io_oeb_unbuf[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2270.340 212.760 2271.440 212.960 ;
      LAYER mcon ;
        RECT 2270.340 212.790 2271.430 212.960 ;
      LAYER met1 ;
        RECT 2270.335 221.600 2417.040 221.740 ;
        RECT 2270.335 221.480 2270.655 221.600 ;
        RECT 2270.280 212.750 2271.490 213.010 ;
        RECT 2416.900 212.060 2417.040 221.600 ;
        RECT 3376.800 212.740 3376.940 1155.450 ;
        RECT 2536.380 212.600 3376.940 212.740 ;
        RECT 2536.380 212.060 2536.520 212.600 ;
        RECT 2416.900 211.920 2536.520 212.060 ;
      LAYER via ;
        RECT 2270.365 221.480 2270.625 221.740 ;
        RECT 2270.340 212.750 2271.430 213.010 ;
      LAYER met2 ;
        RECT 2270.365 221.770 2270.505 232.485 ;
        RECT 2270.365 221.450 2270.625 221.770 ;
        RECT 2270.365 214.170 2270.505 221.450 ;
        RECT 2270.365 214.030 2271.140 214.170 ;
        RECT 2271.000 213.040 2271.140 214.030 ;
        RECT 2270.340 212.720 2271.430 213.040 ;
    END
  END mgmt_io_oeb_unbuf[1]
  PIN mgmt_io_oeb_unbuf[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2264.360 215.850 2265.950 216.050 ;
      LAYER mcon ;
        RECT 2264.860 215.850 2265.950 216.020 ;
      LAYER met1 ;
        RECT 2265.205 222.160 2417.880 222.300 ;
        RECT 2265.205 222.040 2265.525 222.160 ;
        RECT 2264.800 215.810 2266.010 216.070 ;
        RECT 2417.740 212.340 2417.880 222.160 ;
        RECT 3375.960 213.300 3376.100 1154.440 ;
        RECT 2535.540 213.160 3376.100 213.300 ;
        RECT 2535.540 212.340 2535.680 213.160 ;
        RECT 2417.740 212.200 2535.680 212.340 ;
      LAYER via ;
        RECT 2265.235 222.040 2265.495 222.300 ;
        RECT 2264.860 215.810 2265.950 216.070 ;
      LAYER met2 ;
        RECT 2265.355 222.330 2265.495 232.485 ;
        RECT 2265.235 222.010 2265.495 222.330 ;
        RECT 2265.355 216.100 2265.495 222.010 ;
        RECT 2264.860 215.780 2265.950 216.100 ;
    END
  END mgmt_io_oeb_unbuf[0]
  PIN mgmt_io_in_buf[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2261.935 213.300 2262.105 214.150 ;
        RECT 2262.775 213.300 2262.945 214.150 ;
        RECT 2263.615 213.300 2263.785 214.150 ;
        RECT 2264.455 213.300 2264.625 214.150 ;
        RECT 2261.935 213.130 2264.625 213.300 ;
        RECT 2264.370 212.590 2264.625 213.130 ;
        RECT 2261.935 212.420 2264.625 212.590 ;
        RECT 2261.935 211.940 2262.105 212.420 ;
        RECT 2262.775 211.940 2262.945 212.420 ;
        RECT 2263.615 211.940 2263.785 212.420 ;
        RECT 2264.455 211.940 2264.625 212.420 ;
      LAYER mcon ;
        RECT 2264.370 212.450 2264.540 213.300 ;
      LAYER met1 ;
        RECT 2264.355 222.720 2418.720 222.860 ;
        RECT 2264.355 222.600 2264.675 222.720 ;
        RECT 2264.320 212.390 2264.580 213.360 ;
        RECT 2418.580 212.620 2418.720 222.720 ;
        RECT 3375.120 213.860 3375.260 1153.450 ;
        RECT 2534.700 213.720 3375.260 213.860 ;
        RECT 2534.700 212.620 2534.840 213.720 ;
        RECT 2418.580 212.480 2534.840 212.620 ;
      LAYER via ;
        RECT 2264.385 222.600 2264.645 222.860 ;
        RECT 2264.320 212.450 2264.580 213.300 ;
      LAYER met2 ;
        RECT 2264.385 222.890 2264.525 232.485 ;
        RECT 2264.385 222.570 2264.645 222.890 ;
        RECT 2264.385 213.300 2264.525 222.570 ;
        RECT 2264.290 212.450 2264.610 213.300 ;
    END
  END mgmt_io_in_buf[19]
  PIN mgmt_io_in_buf[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2255.955 213.300 2256.125 214.150 ;
        RECT 2256.795 213.300 2256.965 214.150 ;
        RECT 2257.635 213.300 2257.805 214.150 ;
        RECT 2258.475 213.300 2258.645 214.150 ;
        RECT 2255.955 213.130 2258.645 213.300 ;
        RECT 2258.390 212.590 2258.645 213.130 ;
        RECT 2255.955 212.420 2258.645 212.590 ;
        RECT 2255.955 211.940 2256.125 212.420 ;
        RECT 2256.795 211.940 2256.965 212.420 ;
        RECT 2257.635 211.940 2257.805 212.420 ;
        RECT 2258.475 211.940 2258.645 212.420 ;
      LAYER mcon ;
        RECT 2258.390 212.450 2258.560 213.300 ;
      LAYER met1 ;
        RECT 2258.375 223.560 2419.840 223.700 ;
        RECT 2258.375 223.440 2258.695 223.560 ;
        RECT 2258.340 212.390 2258.600 213.360 ;
        RECT 2419.695 213.180 2419.835 223.560 ;
        RECT 3374.000 214.700 3374.140 1151.450 ;
        RECT 2533.580 214.560 3374.140 214.700 ;
        RECT 2533.580 213.180 2533.720 214.560 ;
        RECT 2419.695 213.040 2533.720 213.180 ;
      LAYER via ;
        RECT 2258.405 223.440 2258.665 223.700 ;
        RECT 2258.340 212.450 2258.600 213.300 ;
      LAYER met2 ;
        RECT 2258.405 223.730 2258.545 232.485 ;
        RECT 2258.405 223.410 2258.665 223.730 ;
        RECT 2258.405 213.300 2258.545 223.410 ;
        RECT 2258.310 212.450 2258.630 213.300 ;
    END
  END mgmt_io_in_buf[18]
  PIN mgmt_io_in_buf[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2249.975 213.300 2250.145 214.150 ;
        RECT 2250.815 213.300 2250.985 214.150 ;
        RECT 2251.655 213.300 2251.825 214.150 ;
        RECT 2252.495 213.300 2252.665 214.150 ;
        RECT 2249.975 213.130 2252.665 213.300 ;
        RECT 2252.410 212.590 2252.665 213.130 ;
        RECT 2249.975 212.420 2252.665 212.590 ;
        RECT 2249.975 211.940 2250.145 212.420 ;
        RECT 2250.815 211.940 2250.985 212.420 ;
        RECT 2251.655 211.940 2251.825 212.420 ;
        RECT 2252.495 211.940 2252.665 212.420 ;
      LAYER mcon ;
        RECT 2252.410 212.450 2252.580 213.300 ;
      LAYER met1 ;
        RECT 2252.395 224.400 2420.960 224.540 ;
        RECT 2252.395 224.280 2252.715 224.400 ;
        RECT 2420.820 213.740 2420.960 224.400 ;
        RECT 3372.880 215.540 3373.020 1149.440 ;
        RECT 2532.460 215.400 3373.020 215.540 ;
        RECT 2532.460 213.740 2532.600 215.400 ;
        RECT 2420.820 213.600 2532.600 213.740 ;
        RECT 2252.360 212.390 2252.620 213.360 ;
      LAYER via ;
        RECT 2252.425 224.280 2252.685 224.540 ;
        RECT 2252.360 212.450 2252.620 213.300 ;
      LAYER met2 ;
        RECT 2252.425 224.570 2252.565 232.485 ;
        RECT 2252.425 224.250 2252.685 224.570 ;
        RECT 2252.425 213.300 2252.565 224.250 ;
        RECT 2252.330 212.450 2252.650 213.300 ;
    END
  END mgmt_io_in_buf[17]
  PIN mgmt_io_in_buf[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2243.995 213.300 2244.165 214.150 ;
        RECT 2244.835 213.300 2245.005 214.150 ;
        RECT 2245.675 213.300 2245.845 214.150 ;
        RECT 2246.515 213.300 2246.685 214.150 ;
        RECT 2243.995 213.130 2246.685 213.300 ;
        RECT 2246.430 212.590 2246.685 213.130 ;
        RECT 2243.995 212.420 2246.685 212.590 ;
        RECT 2243.995 211.940 2244.165 212.420 ;
        RECT 2244.835 211.940 2245.005 212.420 ;
        RECT 2245.675 211.940 2245.845 212.420 ;
        RECT 2246.515 211.940 2246.685 212.420 ;
      LAYER mcon ;
        RECT 2246.430 212.450 2246.600 213.300 ;
      LAYER met1 ;
        RECT 2246.415 225.240 2422.080 225.380 ;
        RECT 2246.415 225.120 2246.735 225.240 ;
        RECT 2421.940 214.300 2422.080 225.240 ;
        RECT 3371.760 216.380 3371.900 1147.440 ;
        RECT 2531.340 216.240 3371.900 216.380 ;
        RECT 2531.340 214.300 2531.480 216.240 ;
        RECT 2421.940 214.160 2531.480 214.300 ;
        RECT 2246.380 212.390 2246.640 213.360 ;
      LAYER via ;
        RECT 2246.445 225.120 2246.705 225.380 ;
        RECT 2246.380 212.450 2246.640 213.300 ;
      LAYER met2 ;
        RECT 2246.445 225.410 2246.585 232.485 ;
        RECT 2246.445 225.090 2246.705 225.410 ;
        RECT 2246.445 213.300 2246.585 225.090 ;
        RECT 2246.350 212.450 2246.670 213.300 ;
    END
  END mgmt_io_in_buf[16]
  PIN mgmt_io_out_unbuf[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2240.440 215.850 2242.030 216.050 ;
      LAYER mcon ;
        RECT 2240.940 215.850 2242.030 216.020 ;
      LAYER met1 ;
        RECT 3371.200 1143.040 3371.340 1146.440 ;
        RECT 3371.200 1142.900 3371.620 1143.040 ;
        RECT 2241.405 225.520 2422.360 225.660 ;
        RECT 2241.405 225.400 2241.725 225.520 ;
        RECT 2240.880 215.810 2242.090 216.070 ;
        RECT 2422.220 214.580 2422.360 225.520 ;
        RECT 3371.480 216.660 3371.620 1142.900 ;
        RECT 2531.060 216.520 3371.620 216.660 ;
        RECT 2531.060 214.580 2531.200 216.520 ;
        RECT 2422.220 214.440 2531.200 214.580 ;
      LAYER via ;
        RECT 2241.435 225.400 2241.695 225.660 ;
        RECT 2240.940 215.810 2242.030 216.070 ;
      LAYER met2 ;
        RECT 2241.435 225.690 2241.575 232.485 ;
        RECT 2241.435 225.370 2241.695 225.690 ;
        RECT 2241.435 216.100 2241.575 225.370 ;
        RECT 2240.940 215.780 2242.030 216.100 ;
    END
  END mgmt_io_out_unbuf[16]
  PIN mgmt_io_out_unbuf[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2246.420 215.850 2248.010 216.050 ;
      LAYER mcon ;
        RECT 2246.920 215.850 2248.010 216.020 ;
      LAYER met1 ;
        RECT 3372.320 1145.005 3372.460 1148.450 ;
        RECT 3372.320 1144.865 3372.740 1145.005 ;
        RECT 2247.385 224.680 2421.240 224.820 ;
        RECT 2247.385 224.560 2247.705 224.680 ;
        RECT 2246.860 215.810 2248.070 216.070 ;
        RECT 2421.100 214.020 2421.240 224.680 ;
        RECT 3372.600 215.820 3372.740 1144.865 ;
        RECT 2532.180 215.680 3372.740 215.820 ;
        RECT 2532.180 214.020 2532.320 215.680 ;
        RECT 2421.100 213.880 2532.320 214.020 ;
      LAYER via ;
        RECT 2247.415 224.560 2247.675 224.820 ;
        RECT 2246.920 215.810 2248.010 216.070 ;
      LAYER met2 ;
        RECT 2247.415 224.850 2247.555 232.485 ;
        RECT 2247.415 224.530 2247.675 224.850 ;
        RECT 2247.415 216.100 2247.555 224.530 ;
        RECT 2246.920 215.780 2248.010 216.100 ;
    END
  END mgmt_io_out_unbuf[17]
  PIN mgmt_io_out_unbuf[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2252.400 215.850 2253.990 216.050 ;
      LAYER mcon ;
        RECT 2252.900 215.850 2253.990 216.020 ;
      LAYER met1 ;
        RECT 3373.440 1146.985 3373.580 1150.440 ;
        RECT 3373.440 1146.845 3373.860 1146.985 ;
        RECT 2253.245 223.840 2420.120 223.980 ;
        RECT 2253.245 223.720 2253.565 223.840 ;
        RECT 2252.840 215.810 2254.050 216.070 ;
        RECT 2419.980 213.460 2420.120 223.840 ;
        RECT 3373.720 214.980 3373.860 1146.845 ;
        RECT 2533.300 214.840 3373.860 214.980 ;
        RECT 2533.300 213.460 2533.440 214.840 ;
        RECT 2419.980 213.320 2533.440 213.460 ;
      LAYER via ;
        RECT 2253.275 223.720 2253.535 223.980 ;
        RECT 2252.900 215.810 2253.990 216.070 ;
      LAYER met2 ;
        RECT 2253.395 224.010 2253.535 232.485 ;
        RECT 2253.275 223.690 2253.535 224.010 ;
        RECT 2253.395 216.100 2253.535 223.690 ;
        RECT 2252.900 215.780 2253.990 216.100 ;
    END
  END mgmt_io_out_unbuf[18]
  PIN mgmt_io_out_unbuf[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2258.380 215.850 2259.970 216.050 ;
      LAYER mcon ;
        RECT 2258.880 215.850 2259.970 216.020 ;
      LAYER met1 ;
        RECT 3374.560 1148.980 3374.700 1152.450 ;
        RECT 3374.560 1148.840 3374.980 1148.980 ;
        RECT 2259.345 223.000 2419.000 223.140 ;
        RECT 2259.345 222.880 2259.665 223.000 ;
        RECT 2258.820 215.810 2260.030 216.070 ;
        RECT 2418.860 212.900 2419.000 223.000 ;
        RECT 3374.840 214.140 3374.980 1148.840 ;
        RECT 2534.420 214.000 3374.980 214.140 ;
        RECT 2534.420 212.900 2534.560 214.000 ;
        RECT 2418.860 212.760 2534.560 212.900 ;
      LAYER via ;
        RECT 2259.375 222.880 2259.635 223.140 ;
        RECT 2258.880 215.810 2259.970 216.070 ;
      LAYER met2 ;
        RECT 2259.375 223.170 2259.515 232.485 ;
        RECT 2259.375 222.850 2259.635 223.170 ;
        RECT 2259.375 216.100 2259.515 222.850 ;
        RECT 2258.880 215.780 2259.970 216.100 ;
    END
  END mgmt_io_out_unbuf[19]
  PIN mgmt_io_out_unbuf[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2150.740 215.850 2152.330 216.050 ;
      LAYER mcon ;
        RECT 2151.240 215.850 2152.330 216.020 ;
      LAYER met1 ;
        RECT 2151.705 238.120 2439.160 238.260 ;
        RECT 2151.705 238.000 2152.025 238.120 ;
        RECT 2439.020 222.980 2439.160 238.120 ;
        RECT 3354.680 229.260 3354.820 1116.750 ;
        RECT 2514.260 229.120 3354.820 229.260 ;
        RECT 2514.260 222.980 2514.400 229.120 ;
        RECT 2439.020 222.840 2514.400 222.980 ;
        RECT 2151.180 215.810 2152.390 216.070 ;
      LAYER via ;
        RECT 2151.735 238.000 2151.995 238.260 ;
        RECT 2151.240 215.810 2152.330 216.070 ;
      LAYER met2 ;
        RECT 2151.735 238.290 2151.875 238.365 ;
        RECT 2151.735 237.970 2151.995 238.290 ;
        RECT 2151.735 216.100 2151.875 237.970 ;
        RECT 2151.240 215.780 2152.330 216.100 ;
    END
  END mgmt_io_out_unbuf[15]
  PIN mgmt_io_out_unbuf[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2156.720 215.850 2158.310 216.050 ;
      LAYER mcon ;
        RECT 2157.220 215.850 2158.310 216.020 ;
      LAYER met1 ;
        RECT 2157.685 237.280 2438.040 237.420 ;
        RECT 2157.685 237.160 2158.005 237.280 ;
        RECT 2437.900 222.420 2438.040 237.280 ;
        RECT 3355.800 228.420 3355.940 1118.700 ;
        RECT 2515.380 228.280 3355.940 228.420 ;
        RECT 2515.380 222.420 2515.520 228.280 ;
        RECT 2437.900 222.280 2515.520 222.420 ;
        RECT 2157.160 215.810 2158.370 216.070 ;
      LAYER via ;
        RECT 2157.715 237.160 2157.975 237.420 ;
        RECT 2157.220 215.810 2158.310 216.070 ;
      LAYER met2 ;
        RECT 2157.715 237.450 2157.855 237.575 ;
        RECT 2157.715 237.130 2157.975 237.450 ;
        RECT 2157.715 216.100 2157.855 237.130 ;
        RECT 2157.220 215.780 2158.310 216.100 ;
    END
  END mgmt_io_out_unbuf[14]
  PIN mgmt_io_out_unbuf[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2162.700 215.850 2164.290 216.050 ;
      LAYER mcon ;
        RECT 2163.200 215.850 2164.290 216.020 ;
      LAYER met1 ;
        RECT 2163.665 236.440 2436.920 236.580 ;
        RECT 2163.665 236.320 2163.985 236.440 ;
        RECT 2436.780 221.860 2436.920 236.440 ;
        RECT 3356.920 227.580 3357.060 1120.690 ;
        RECT 2516.500 227.440 3357.060 227.580 ;
        RECT 2516.500 221.860 2516.640 227.440 ;
        RECT 2436.780 221.720 2516.640 221.860 ;
        RECT 2163.140 215.810 2164.350 216.070 ;
      LAYER via ;
        RECT 2163.695 236.320 2163.955 236.580 ;
        RECT 2163.200 215.810 2164.290 216.070 ;
      LAYER met2 ;
        RECT 2163.695 236.610 2163.835 236.720 ;
        RECT 2163.695 236.290 2163.955 236.610 ;
        RECT 2163.695 216.100 2163.835 236.290 ;
        RECT 2163.200 215.780 2164.290 216.100 ;
    END
  END mgmt_io_out_unbuf[13]
  PIN mgmt_io_out_unbuf[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2168.680 215.850 2170.270 216.050 ;
      LAYER mcon ;
        RECT 2169.180 215.850 2170.270 216.020 ;
      LAYER met1 ;
        RECT 2169.645 235.600 2435.800 235.740 ;
        RECT 2169.645 235.480 2169.965 235.600 ;
        RECT 2435.660 221.300 2435.800 235.600 ;
        RECT 3358.040 226.740 3358.180 1122.710 ;
        RECT 2517.620 226.600 3358.180 226.740 ;
        RECT 2517.620 221.300 2517.760 226.600 ;
        RECT 2435.660 221.160 2517.760 221.300 ;
        RECT 2169.120 215.810 2170.330 216.070 ;
      LAYER via ;
        RECT 2169.675 235.480 2169.935 235.740 ;
        RECT 2169.180 215.810 2170.270 216.070 ;
      LAYER met2 ;
        RECT 2169.675 235.770 2169.815 235.930 ;
        RECT 2169.675 235.450 2169.935 235.770 ;
        RECT 2169.675 216.100 2169.815 235.450 ;
        RECT 2169.180 215.780 2170.270 216.100 ;
    END
  END mgmt_io_out_unbuf[12]
  PIN mgmt_io_out_unbuf[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2174.660 215.850 2176.250 216.050 ;
      LAYER mcon ;
        RECT 2175.160 215.850 2176.250 216.020 ;
      LAYER met1 ;
        RECT 2175.625 234.760 2434.680 234.900 ;
        RECT 2175.625 234.640 2175.945 234.760 ;
        RECT 2434.540 220.740 2434.680 234.760 ;
        RECT 3359.160 225.900 3359.300 1124.680 ;
        RECT 2518.740 225.760 3359.300 225.900 ;
        RECT 2518.740 220.740 2518.880 225.760 ;
        RECT 2434.540 220.600 2518.880 220.740 ;
        RECT 2175.100 215.810 2176.310 216.070 ;
      LAYER via ;
        RECT 2175.655 234.640 2175.915 234.900 ;
        RECT 2175.160 215.810 2176.250 216.070 ;
      LAYER met2 ;
        RECT 2175.655 234.930 2175.795 235.010 ;
        RECT 2175.655 234.610 2175.915 234.930 ;
        RECT 2175.655 216.100 2175.795 234.610 ;
        RECT 2175.160 215.780 2176.250 216.100 ;
    END
  END mgmt_io_out_unbuf[11]
  PIN mgmt_io_out_unbuf[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2180.640 215.850 2182.230 216.050 ;
      LAYER mcon ;
        RECT 2181.140 215.850 2182.230 216.020 ;
      LAYER met1 ;
        RECT 2181.485 233.920 2433.560 234.060 ;
        RECT 2181.485 233.800 2181.805 233.920 ;
        RECT 2433.420 220.180 2433.560 233.920 ;
        RECT 3360.280 225.060 3360.420 1126.700 ;
        RECT 2519.860 224.920 3360.420 225.060 ;
        RECT 2519.860 220.180 2520.000 224.920 ;
        RECT 2433.420 220.040 2520.000 220.180 ;
        RECT 2181.080 215.810 2182.290 216.070 ;
      LAYER via ;
        RECT 2181.515 233.800 2181.775 234.060 ;
        RECT 2181.140 215.810 2182.230 216.070 ;
      LAYER met2 ;
        RECT 2181.635 234.090 2181.775 234.200 ;
        RECT 2181.515 233.770 2181.775 234.090 ;
        RECT 2181.635 216.100 2181.775 233.770 ;
        RECT 2181.140 215.780 2182.230 216.100 ;
    END
  END mgmt_io_out_unbuf[10]
  PIN mgmt_io_out_unbuf[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2186.620 215.850 2188.210 216.050 ;
      LAYER mcon ;
        RECT 2187.120 215.850 2188.210 216.020 ;
      LAYER met1 ;
        RECT 2187.585 233.080 2432.440 233.220 ;
        RECT 2187.585 232.960 2187.905 233.080 ;
        RECT 2432.300 219.620 2432.440 233.080 ;
        RECT 3361.400 224.220 3361.540 1128.690 ;
        RECT 2520.980 224.080 3361.540 224.220 ;
        RECT 2520.980 219.620 2521.120 224.080 ;
        RECT 2432.300 219.480 2521.120 219.620 ;
        RECT 2187.060 215.810 2188.270 216.070 ;
      LAYER via ;
        RECT 2187.615 232.960 2187.875 233.220 ;
        RECT 2187.120 215.810 2188.210 216.070 ;
      LAYER met2 ;
        RECT 2187.615 233.250 2187.755 233.365 ;
        RECT 2187.615 232.930 2187.875 233.250 ;
        RECT 2187.615 216.100 2187.755 232.930 ;
        RECT 2187.120 215.780 2188.210 216.100 ;
    END
  END mgmt_io_out_unbuf[9]
  PIN mgmt_io_out_unbuf[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2192.600 215.850 2194.190 216.050 ;
      LAYER mcon ;
        RECT 2193.100 215.850 2194.190 216.020 ;
      LAYER met1 ;
        RECT 2193.445 232.240 2431.320 232.380 ;
        RECT 2193.445 232.120 2193.765 232.240 ;
        RECT 2431.180 219.060 2431.320 232.240 ;
        RECT 3362.520 223.380 3362.660 1130.690 ;
        RECT 2522.100 223.240 3362.660 223.380 ;
        RECT 2522.100 219.060 2522.240 223.240 ;
        RECT 2431.180 218.920 2522.240 219.060 ;
        RECT 2193.040 215.810 2194.250 216.070 ;
      LAYER via ;
        RECT 2193.475 232.120 2193.735 232.380 ;
        RECT 2193.100 215.810 2194.190 216.070 ;
      LAYER met2 ;
        RECT 2193.595 232.410 2193.735 232.485 ;
        RECT 2193.475 232.090 2193.735 232.410 ;
        RECT 2193.595 216.100 2193.735 232.090 ;
        RECT 2193.100 215.780 2194.190 216.100 ;
    END
  END mgmt_io_out_unbuf[8]
  PIN mgmt_io_out_unbuf[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2198.580 215.850 2200.170 216.050 ;
      LAYER mcon ;
        RECT 2199.080 215.850 2200.170 216.020 ;
      LAYER met1 ;
        RECT 2199.545 231.400 2430.200 231.540 ;
        RECT 2199.545 231.280 2199.865 231.400 ;
        RECT 2430.060 218.500 2430.200 231.400 ;
        RECT 3363.640 222.540 3363.780 1132.690 ;
        RECT 2523.220 222.400 3363.780 222.540 ;
        RECT 2523.220 218.500 2523.360 222.400 ;
        RECT 2430.060 218.360 2523.360 218.500 ;
        RECT 2199.020 215.810 2200.230 216.070 ;
      LAYER via ;
        RECT 2199.575 231.280 2199.835 231.540 ;
        RECT 2199.080 215.810 2200.170 216.070 ;
      LAYER met2 ;
        RECT 2199.575 231.570 2199.715 232.485 ;
        RECT 2199.575 231.250 2199.835 231.570 ;
        RECT 2199.575 216.100 2199.715 231.250 ;
        RECT 2199.080 215.780 2200.170 216.100 ;
    END
  END mgmt_io_out_unbuf[7]
  PIN mgmt_io_in_buf[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2202.135 213.300 2202.305 214.150 ;
        RECT 2202.975 213.300 2203.145 214.150 ;
        RECT 2203.815 213.300 2203.985 214.150 ;
        RECT 2204.655 213.300 2204.825 214.150 ;
        RECT 2202.135 213.130 2204.825 213.300 ;
        RECT 2204.570 212.590 2204.825 213.130 ;
        RECT 2202.135 212.420 2204.825 212.590 ;
        RECT 2202.135 211.940 2202.305 212.420 ;
        RECT 2202.975 211.940 2203.145 212.420 ;
        RECT 2203.815 211.940 2203.985 212.420 ;
        RECT 2204.655 211.940 2204.825 212.420 ;
      LAYER mcon ;
        RECT 2204.570 212.450 2204.740 213.300 ;
      LAYER met1 ;
        RECT 3364.200 1130.145 3364.340 1133.680 ;
        RECT 3363.920 1130.005 3364.340 1130.145 ;
        RECT 2204.555 231.120 2429.920 231.260 ;
        RECT 2204.555 231.000 2204.875 231.120 ;
        RECT 2429.780 218.220 2429.920 231.120 ;
        RECT 3363.920 222.260 3364.060 1130.005 ;
        RECT 2523.500 222.120 3364.060 222.260 ;
        RECT 2523.500 218.220 2523.640 222.120 ;
        RECT 2429.780 218.080 2523.640 218.220 ;
        RECT 2204.520 212.390 2204.780 213.360 ;
      LAYER via ;
        RECT 2204.585 231.000 2204.845 231.260 ;
        RECT 2204.520 212.450 2204.780 213.300 ;
      LAYER met2 ;
        RECT 2204.585 231.290 2204.725 232.485 ;
        RECT 2204.585 230.970 2204.845 231.290 ;
        RECT 2204.585 213.300 2204.725 230.970 ;
        RECT 2204.490 212.450 2204.810 213.300 ;
    END
  END mgmt_io_in_buf[7]
  PIN mgmt_io_in_buf[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2196.155 213.300 2196.325 214.150 ;
        RECT 2196.995 213.300 2197.165 214.150 ;
        RECT 2197.835 213.300 2198.005 214.150 ;
        RECT 2198.675 213.300 2198.845 214.150 ;
        RECT 2196.155 213.130 2198.845 213.300 ;
        RECT 2198.590 212.590 2198.845 213.130 ;
        RECT 2196.155 212.420 2198.845 212.590 ;
        RECT 2196.155 211.940 2196.325 212.420 ;
        RECT 2196.995 211.940 2197.165 212.420 ;
        RECT 2197.835 211.940 2198.005 212.420 ;
        RECT 2198.675 211.940 2198.845 212.420 ;
      LAYER mcon ;
        RECT 2198.590 212.450 2198.760 213.300 ;
      LAYER met1 ;
        RECT 3363.080 1128.270 3363.220 1131.680 ;
        RECT 3362.800 1128.130 3363.220 1128.270 ;
        RECT 2198.575 231.960 2431.040 232.100 ;
        RECT 2198.575 231.840 2198.895 231.960 ;
        RECT 2430.900 218.780 2431.040 231.960 ;
        RECT 3362.800 223.100 3362.940 1128.130 ;
        RECT 2522.380 222.960 3362.940 223.100 ;
        RECT 2522.380 218.780 2522.520 222.960 ;
        RECT 2430.900 218.640 2522.520 218.780 ;
        RECT 2198.540 212.390 2198.800 213.360 ;
      LAYER via ;
        RECT 2198.605 231.840 2198.865 232.100 ;
        RECT 2198.540 212.450 2198.800 213.300 ;
      LAYER met2 ;
        RECT 2198.605 232.130 2198.745 232.485 ;
        RECT 2198.605 231.810 2198.865 232.130 ;
        RECT 2198.605 213.300 2198.745 231.810 ;
        RECT 2198.510 212.450 2198.830 213.300 ;
    END
  END mgmt_io_in_buf[8]
  PIN mgmt_io_in_buf[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2190.175 213.300 2190.345 214.150 ;
        RECT 2191.015 213.300 2191.185 214.150 ;
        RECT 2191.855 213.300 2192.025 214.150 ;
        RECT 2192.695 213.300 2192.865 214.150 ;
        RECT 2190.175 213.130 2192.865 213.300 ;
        RECT 2192.610 212.590 2192.865 213.130 ;
        RECT 2190.175 212.420 2192.865 212.590 ;
        RECT 2190.175 211.940 2190.345 212.420 ;
        RECT 2191.015 211.940 2191.185 212.420 ;
        RECT 2191.855 211.940 2192.025 212.420 ;
        RECT 2192.695 211.940 2192.865 212.420 ;
      LAYER mcon ;
        RECT 2192.610 212.450 2192.780 213.300 ;
      LAYER met1 ;
        RECT 3361.960 1126.275 3362.100 1129.710 ;
        RECT 3361.680 1126.135 3362.100 1126.275 ;
        RECT 2192.595 232.800 2432.160 232.940 ;
        RECT 2192.595 232.680 2192.915 232.800 ;
        RECT 2432.020 219.340 2432.160 232.800 ;
        RECT 3361.680 223.940 3361.820 1126.135 ;
        RECT 2521.260 223.800 3361.820 223.940 ;
        RECT 2521.260 219.340 2521.400 223.800 ;
        RECT 2432.020 219.200 2521.400 219.340 ;
        RECT 2192.560 212.390 2192.820 213.360 ;
      LAYER via ;
        RECT 2192.625 232.680 2192.885 232.940 ;
        RECT 2192.560 212.450 2192.820 213.300 ;
      LAYER met2 ;
        RECT 2192.625 232.970 2192.765 233.010 ;
        RECT 2192.625 232.650 2192.885 232.970 ;
        RECT 2192.625 213.300 2192.765 232.650 ;
        RECT 2192.530 212.450 2192.850 213.300 ;
    END
  END mgmt_io_in_buf[9]
  PIN mgmt_io_in_buf[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2184.195 213.300 2184.365 214.150 ;
        RECT 2185.035 213.300 2185.205 214.150 ;
        RECT 2185.875 213.300 2186.045 214.150 ;
        RECT 2186.715 213.300 2186.885 214.150 ;
        RECT 2184.195 213.130 2186.885 213.300 ;
        RECT 2186.630 212.590 2186.885 213.130 ;
        RECT 2184.195 212.420 2186.885 212.590 ;
        RECT 2184.195 211.940 2184.365 212.420 ;
        RECT 2185.035 211.940 2185.205 212.420 ;
        RECT 2185.875 211.940 2186.045 212.420 ;
        RECT 2186.715 211.940 2186.885 212.420 ;
      LAYER mcon ;
        RECT 2186.630 212.450 2186.800 213.300 ;
      LAYER met1 ;
        RECT 3360.840 1124.165 3360.980 1127.680 ;
        RECT 3360.560 1124.025 3360.980 1124.165 ;
        RECT 2186.615 233.640 2433.280 233.780 ;
        RECT 2186.615 233.520 2186.935 233.640 ;
        RECT 2433.140 219.900 2433.280 233.640 ;
        RECT 3360.560 224.780 3360.700 1124.025 ;
        RECT 2520.140 224.640 3360.700 224.780 ;
        RECT 2520.140 219.900 2520.280 224.640 ;
        RECT 2433.140 219.760 2520.280 219.900 ;
        RECT 2186.580 212.390 2186.840 213.360 ;
      LAYER via ;
        RECT 2186.645 233.520 2186.905 233.780 ;
        RECT 2186.580 212.450 2186.840 213.300 ;
      LAYER met2 ;
        RECT 2186.645 233.810 2186.785 233.870 ;
        RECT 2186.645 233.490 2186.905 233.810 ;
        RECT 2186.645 213.300 2186.785 233.490 ;
        RECT 2186.550 212.450 2186.870 213.300 ;
    END
  END mgmt_io_in_buf[10]
  PIN mgmt_io_in_buf[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2178.215 213.300 2178.385 214.150 ;
        RECT 2179.055 213.300 2179.225 214.150 ;
        RECT 2179.895 213.300 2180.065 214.150 ;
        RECT 2180.735 213.300 2180.905 214.150 ;
        RECT 2178.215 213.130 2180.905 213.300 ;
        RECT 2180.650 212.590 2180.905 213.130 ;
        RECT 2178.215 212.420 2180.905 212.590 ;
        RECT 2178.215 211.940 2178.385 212.420 ;
        RECT 2179.055 211.940 2179.225 212.420 ;
        RECT 2179.895 211.940 2180.065 212.420 ;
        RECT 2180.735 211.940 2180.905 212.420 ;
      LAYER mcon ;
        RECT 2180.650 212.450 2180.820 213.300 ;
      LAYER met1 ;
        RECT 3359.720 1122.215 3359.860 1125.700 ;
        RECT 3359.440 1122.075 3359.860 1122.215 ;
        RECT 2180.635 234.480 2434.400 234.620 ;
        RECT 2180.635 234.360 2180.955 234.480 ;
        RECT 2434.260 220.460 2434.400 234.480 ;
        RECT 3359.440 225.620 3359.580 1122.075 ;
        RECT 2519.020 225.480 3359.580 225.620 ;
        RECT 2519.020 220.460 2519.160 225.480 ;
        RECT 2434.260 220.320 2519.160 220.460 ;
        RECT 2180.600 212.390 2180.860 213.360 ;
      LAYER via ;
        RECT 2180.665 234.360 2180.925 234.620 ;
        RECT 2180.600 212.450 2180.860 213.300 ;
      LAYER met2 ;
        RECT 2180.665 234.650 2180.805 234.705 ;
        RECT 2180.665 234.330 2180.925 234.650 ;
        RECT 2180.665 213.300 2180.805 234.330 ;
        RECT 2180.570 212.450 2180.890 213.300 ;
    END
  END mgmt_io_in_buf[11]
  PIN mgmt_io_in_buf[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2172.235 213.300 2172.405 214.150 ;
        RECT 2173.075 213.300 2173.245 214.150 ;
        RECT 2173.915 213.300 2174.085 214.150 ;
        RECT 2174.755 213.300 2174.925 214.150 ;
        RECT 2172.235 213.130 2174.925 213.300 ;
        RECT 2174.670 212.590 2174.925 213.130 ;
        RECT 2172.235 212.420 2174.925 212.590 ;
        RECT 2172.235 211.940 2172.405 212.420 ;
        RECT 2173.075 211.940 2173.245 212.420 ;
        RECT 2173.915 211.940 2174.085 212.420 ;
        RECT 2174.755 211.940 2174.925 212.420 ;
      LAYER mcon ;
        RECT 2174.670 212.450 2174.840 213.300 ;
      LAYER met1 ;
        RECT 3358.600 1120.330 3358.740 1123.720 ;
        RECT 3358.320 1120.190 3358.740 1120.330 ;
        RECT 2174.655 235.320 2435.520 235.460 ;
        RECT 2174.655 235.200 2174.975 235.320 ;
        RECT 2435.380 221.020 2435.520 235.320 ;
        RECT 3358.320 226.460 3358.460 1120.190 ;
        RECT 2517.900 226.320 3358.460 226.460 ;
        RECT 2517.900 221.020 2518.040 226.320 ;
        RECT 2435.380 220.880 2518.040 221.020 ;
        RECT 2174.620 212.390 2174.880 213.360 ;
      LAYER via ;
        RECT 2174.685 235.200 2174.945 235.460 ;
        RECT 2174.620 212.450 2174.880 213.300 ;
      LAYER met2 ;
        RECT 2174.685 235.490 2174.825 235.530 ;
        RECT 2174.685 235.170 2174.945 235.490 ;
        RECT 2174.685 213.300 2174.825 235.170 ;
        RECT 2174.590 212.450 2174.910 213.300 ;
    END
  END mgmt_io_in_buf[12]
  PIN mgmt_io_in_buf[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2166.255 213.300 2166.425 214.150 ;
        RECT 2167.095 213.300 2167.265 214.150 ;
        RECT 2167.935 213.300 2168.105 214.150 ;
        RECT 2168.775 213.300 2168.945 214.150 ;
        RECT 2166.255 213.130 2168.945 213.300 ;
        RECT 2168.690 212.590 2168.945 213.130 ;
        RECT 2166.255 212.420 2168.945 212.590 ;
        RECT 2166.255 211.940 2166.425 212.420 ;
        RECT 2167.095 211.940 2167.265 212.420 ;
        RECT 2167.935 211.940 2168.105 212.420 ;
        RECT 2168.775 211.940 2168.945 212.420 ;
      LAYER mcon ;
        RECT 2168.690 212.450 2168.860 213.300 ;
      LAYER met1 ;
        RECT 3357.480 1118.210 3357.620 1121.740 ;
        RECT 3357.200 1118.070 3357.620 1118.210 ;
        RECT 2168.675 236.160 2436.640 236.300 ;
        RECT 2168.675 236.040 2168.995 236.160 ;
        RECT 2436.500 221.580 2436.640 236.160 ;
        RECT 3357.200 227.300 3357.340 1118.070 ;
        RECT 2516.780 227.160 3357.340 227.300 ;
        RECT 2516.780 221.580 2516.920 227.160 ;
        RECT 2436.500 221.440 2516.920 221.580 ;
        RECT 2168.640 212.390 2168.900 213.360 ;
      LAYER via ;
        RECT 2168.705 236.040 2168.965 236.300 ;
        RECT 2168.640 212.450 2168.900 213.300 ;
      LAYER met2 ;
        RECT 2168.705 236.330 2168.845 236.400 ;
        RECT 2168.705 236.010 2168.965 236.330 ;
        RECT 2168.705 213.300 2168.845 236.010 ;
        RECT 2168.610 212.450 2168.930 213.300 ;
    END
  END mgmt_io_in_buf[13]
  PIN mgmt_io_in_buf[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2160.275 213.300 2160.445 214.150 ;
        RECT 2161.115 213.300 2161.285 214.150 ;
        RECT 2161.955 213.300 2162.125 214.150 ;
        RECT 2162.795 213.300 2162.965 214.150 ;
        RECT 2160.275 213.130 2162.965 213.300 ;
        RECT 2162.710 212.590 2162.965 213.130 ;
        RECT 2160.275 212.420 2162.965 212.590 ;
        RECT 2160.275 211.940 2160.445 212.420 ;
        RECT 2161.115 211.940 2161.285 212.420 ;
        RECT 2161.955 211.940 2162.125 212.420 ;
        RECT 2162.795 211.940 2162.965 212.420 ;
      LAYER mcon ;
        RECT 2162.710 212.450 2162.880 213.300 ;
      LAYER met1 ;
        RECT 3356.360 1116.205 3356.500 1119.690 ;
        RECT 3356.080 1116.065 3356.500 1116.205 ;
        RECT 2162.695 237.000 2437.760 237.140 ;
        RECT 2162.695 236.880 2163.015 237.000 ;
        RECT 2437.620 222.140 2437.760 237.000 ;
        RECT 3356.080 228.140 3356.220 1116.065 ;
        RECT 2515.660 228.000 3356.220 228.140 ;
        RECT 2515.660 222.140 2515.800 228.000 ;
        RECT 2437.620 222.000 2515.800 222.140 ;
        RECT 2162.660 212.390 2162.920 213.360 ;
      LAYER via ;
        RECT 2162.725 236.880 2162.985 237.140 ;
        RECT 2162.660 212.450 2162.920 213.300 ;
      LAYER met2 ;
        RECT 2162.725 237.170 2162.865 237.225 ;
        RECT 2162.725 236.850 2162.985 237.170 ;
        RECT 2162.725 213.300 2162.865 236.850 ;
        RECT 2162.630 212.450 2162.950 213.300 ;
    END
  END mgmt_io_in_buf[14]
  PIN mgmt_io_in_buf[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2154.295 213.300 2154.465 214.150 ;
        RECT 2155.135 213.300 2155.305 214.150 ;
        RECT 2155.975 213.300 2156.145 214.150 ;
        RECT 2156.815 213.300 2156.985 214.150 ;
        RECT 2154.295 213.130 2156.985 213.300 ;
        RECT 2156.730 212.590 2156.985 213.130 ;
        RECT 2154.295 212.420 2156.985 212.590 ;
        RECT 2154.295 211.940 2154.465 212.420 ;
        RECT 2155.135 211.940 2155.305 212.420 ;
        RECT 2155.975 211.940 2156.145 212.420 ;
        RECT 2156.815 211.940 2156.985 212.420 ;
      LAYER mcon ;
        RECT 2156.730 212.450 2156.900 213.300 ;
      LAYER met1 ;
        RECT 3355.240 1114.280 3355.380 1117.730 ;
        RECT 3354.960 1114.140 3355.380 1114.280 ;
        RECT 2156.715 237.840 2438.880 237.980 ;
        RECT 2156.715 237.720 2157.035 237.840 ;
        RECT 2438.740 222.700 2438.880 237.840 ;
        RECT 3354.960 228.980 3355.100 1114.140 ;
        RECT 2514.540 228.840 3355.100 228.980 ;
        RECT 2514.540 222.700 2514.680 228.840 ;
        RECT 2438.740 222.560 2514.680 222.700 ;
        RECT 2156.680 212.390 2156.940 213.360 ;
      LAYER via ;
        RECT 2156.745 237.720 2157.005 237.980 ;
        RECT 2156.680 212.450 2156.940 213.300 ;
      LAYER met2 ;
        RECT 2156.745 238.010 2156.885 238.085 ;
        RECT 2156.745 237.690 2157.005 238.010 ;
        RECT 2156.745 213.300 2156.885 237.690 ;
        RECT 2156.650 212.450 2156.970 213.300 ;
    END
  END mgmt_io_in_buf[15]
  PIN vssd
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 3380.500 2238.065 3380.670 2238.235 ;
        RECT 3385.940 2238.065 3386.110 2238.235 ;
      LAYER li1 ;
        RECT 3380.500 2237.835 3380.670 2237.920 ;
        RECT 3379.955 2237.775 3380.670 2237.835 ;
        RECT 3379.955 2237.605 3380.500 2237.775 ;
      LAYER li1 ;
        RECT 3385.940 2237.605 3386.110 2237.775 ;
      LAYER li1 ;
        RECT 3379.955 2236.250 3380.670 2237.605 ;
      LAYER li1 ;
        RECT 3385.940 2237.145 3386.110 2237.315 ;
        RECT 3385.940 2236.685 3386.110 2236.855 ;
      LAYER li1 ;
        RECT 3379.125 2235.910 3380.670 2236.250 ;
      LAYER li1 ;
        RECT 3385.940 2236.225 3386.110 2236.395 ;
      LAYER li1 ;
        RECT 3379.955 2232.490 3380.670 2235.910 ;
      LAYER li1 ;
        RECT 3385.940 2235.765 3386.110 2235.935 ;
        RECT 3385.940 2235.305 3386.110 2235.475 ;
        RECT 3385.940 2234.845 3386.110 2235.015 ;
        RECT 3385.940 2234.385 3386.110 2234.555 ;
        RECT 3385.940 2233.925 3386.110 2234.095 ;
        RECT 3385.940 2233.465 3386.110 2233.635 ;
        RECT 3385.940 2233.005 3386.110 2233.175 ;
        RECT 3385.940 2232.545 3386.110 2232.715 ;
      LAYER li1 ;
        RECT 3380.500 2232.400 3380.670 2232.490 ;
      LAYER li1 ;
        RECT 3380.500 2232.085 3380.670 2232.255 ;
        RECT 3385.940 2232.085 3386.110 2232.255 ;
        RECT 3380.500 2231.625 3380.670 2231.795 ;
        RECT 3385.940 2231.625 3386.110 2231.795 ;
        RECT 3380.500 2231.165 3380.670 2231.335 ;
        RECT 3385.940 2231.165 3386.110 2231.335 ;
        RECT 3380.500 2230.705 3380.670 2230.875 ;
        RECT 3385.940 2230.705 3386.110 2230.875 ;
        RECT 3380.500 2230.245 3380.670 2230.415 ;
        RECT 3385.940 2230.245 3386.110 2230.415 ;
        RECT 3380.500 2229.785 3380.670 2229.955 ;
        RECT 3385.940 2229.785 3386.110 2229.955 ;
        RECT 3380.500 2229.325 3380.670 2229.495 ;
        RECT 3385.940 2229.325 3386.110 2229.495 ;
        RECT 3380.500 2228.865 3380.670 2229.035 ;
        RECT 3385.940 2228.865 3386.110 2229.035 ;
        RECT 3380.500 2228.405 3380.670 2228.575 ;
        RECT 3385.940 2228.405 3386.110 2228.575 ;
        RECT 3380.500 2227.945 3380.670 2228.115 ;
        RECT 3385.940 2227.945 3386.110 2228.115 ;
        RECT 3380.500 2227.485 3380.670 2227.655 ;
        RECT 3385.940 2227.485 3386.110 2227.655 ;
        RECT 3380.500 2227.025 3380.670 2227.195 ;
        RECT 3385.940 2227.025 3386.110 2227.195 ;
        RECT 3380.500 2226.565 3380.670 2226.735 ;
        RECT 3385.940 2226.565 3386.110 2226.735 ;
        RECT 3380.500 2226.105 3380.670 2226.275 ;
        RECT 3385.940 2226.105 3386.110 2226.275 ;
        RECT 3380.500 2225.645 3380.670 2225.815 ;
        RECT 3385.940 2225.645 3386.110 2225.815 ;
        RECT 3380.500 2225.185 3380.670 2225.355 ;
        RECT 3385.940 2225.185 3386.110 2225.355 ;
        RECT 3380.500 2224.725 3380.670 2224.895 ;
        RECT 3385.940 2224.725 3386.110 2224.895 ;
        RECT 3380.500 2224.265 3380.670 2224.435 ;
        RECT 3385.940 2224.265 3386.110 2224.435 ;
        RECT 3380.500 2223.805 3380.670 2223.975 ;
        RECT 3385.940 2223.805 3386.110 2223.975 ;
        RECT 3380.500 2223.345 3380.670 2223.515 ;
        RECT 3385.940 2223.345 3386.110 2223.515 ;
        RECT 3380.500 2222.885 3380.670 2223.055 ;
        RECT 3385.940 2222.885 3386.110 2223.055 ;
        RECT 3380.500 2222.425 3380.670 2222.595 ;
        RECT 3385.940 2222.425 3386.110 2222.595 ;
        RECT 3380.500 2221.965 3380.670 2222.135 ;
        RECT 3385.940 2221.965 3386.110 2222.135 ;
        RECT 3380.500 2221.505 3380.670 2221.675 ;
        RECT 3385.940 2221.505 3386.110 2221.675 ;
        RECT 3380.500 2221.045 3380.670 2221.215 ;
        RECT 3385.940 2221.045 3386.110 2221.215 ;
        RECT 3380.500 2220.585 3380.670 2220.755 ;
        RECT 3385.940 2220.585 3386.110 2220.755 ;
        RECT 3380.500 2220.125 3380.670 2220.295 ;
        RECT 3385.940 2220.125 3386.110 2220.295 ;
        RECT 3380.500 2219.665 3380.670 2219.835 ;
        RECT 3385.940 2219.665 3386.110 2219.835 ;
        RECT 3380.500 2219.205 3380.670 2219.375 ;
        RECT 3385.940 2219.205 3386.110 2219.375 ;
        RECT 3380.500 2218.745 3380.670 2218.915 ;
        RECT 3385.940 2218.745 3386.110 2218.915 ;
        RECT 3380.500 2218.285 3380.670 2218.455 ;
        RECT 3385.940 2218.285 3386.110 2218.455 ;
        RECT 3380.500 2217.825 3380.670 2217.995 ;
        RECT 3385.940 2217.825 3386.110 2217.995 ;
        RECT 3380.500 2217.365 3380.670 2217.535 ;
        RECT 3385.940 2217.365 3386.110 2217.535 ;
        RECT 3380.500 2216.905 3380.670 2217.075 ;
        RECT 3385.940 2216.905 3386.110 2217.075 ;
        RECT 3380.500 2216.445 3380.670 2216.615 ;
        RECT 3385.940 2216.445 3386.110 2216.615 ;
        RECT 3380.500 2215.985 3380.670 2216.155 ;
        RECT 3385.940 2215.985 3386.110 2216.155 ;
        RECT 3380.500 2215.525 3380.670 2215.695 ;
        RECT 3385.940 2215.525 3386.110 2215.695 ;
        RECT 3380.500 2215.065 3380.670 2215.235 ;
        RECT 3385.940 2215.065 3386.110 2215.235 ;
        RECT 3380.500 2214.605 3380.670 2214.775 ;
        RECT 3385.940 2214.605 3386.110 2214.775 ;
        RECT 3380.500 2214.145 3380.670 2214.315 ;
        RECT 3385.940 2214.145 3386.110 2214.315 ;
        RECT 3380.500 2213.685 3380.670 2213.855 ;
        RECT 3385.940 2213.685 3386.110 2213.855 ;
        RECT 3380.500 2213.225 3380.670 2213.395 ;
        RECT 3385.940 2213.225 3386.110 2213.395 ;
        RECT 3380.500 2212.765 3380.670 2212.935 ;
        RECT 3385.940 2212.765 3386.110 2212.935 ;
        RECT 3380.500 2212.305 3380.670 2212.475 ;
        RECT 3385.940 2212.305 3386.110 2212.475 ;
        RECT 3380.500 2211.845 3380.670 2212.015 ;
        RECT 3385.940 2211.845 3386.110 2212.015 ;
        RECT 3380.500 2211.385 3380.670 2211.555 ;
        RECT 3385.940 2211.385 3386.110 2211.555 ;
        RECT 3380.500 2210.925 3380.670 2211.095 ;
        RECT 3385.940 2210.925 3386.110 2211.095 ;
        RECT 3380.500 2210.465 3380.670 2210.635 ;
        RECT 3385.940 2210.465 3386.110 2210.635 ;
        RECT 3380.500 2210.005 3380.670 2210.175 ;
        RECT 3385.940 2210.005 3386.110 2210.175 ;
        RECT 3380.500 2209.545 3380.670 2209.715 ;
        RECT 3385.940 2209.545 3386.110 2209.715 ;
        RECT 3380.500 2209.085 3380.670 2209.255 ;
        RECT 3385.940 2209.085 3386.110 2209.255 ;
        RECT 3380.500 2208.625 3380.670 2208.795 ;
        RECT 3385.940 2208.625 3386.110 2208.795 ;
        RECT 3380.500 2208.165 3380.670 2208.335 ;
        RECT 3385.940 2208.165 3386.110 2208.335 ;
        RECT 3380.500 2207.705 3380.670 2207.875 ;
        RECT 3385.940 2207.705 3386.110 2207.875 ;
        RECT 3380.500 2207.245 3380.670 2207.415 ;
        RECT 3385.940 2207.245 3386.110 2207.415 ;
        RECT 3380.500 2206.785 3380.670 2206.955 ;
        RECT 3385.940 2206.785 3386.110 2206.955 ;
        RECT 3380.500 2206.325 3380.670 2206.495 ;
        RECT 3385.940 2206.325 3386.110 2206.495 ;
        RECT 3380.500 2205.865 3380.670 2206.035 ;
        RECT 3385.940 2205.865 3386.110 2206.035 ;
        RECT 3380.500 2205.405 3380.670 2205.575 ;
        RECT 3385.940 2205.405 3386.110 2205.575 ;
        RECT 3380.500 2204.945 3380.670 2205.115 ;
        RECT 3385.940 2204.945 3386.110 2205.115 ;
        RECT 3380.500 2204.485 3380.670 2204.655 ;
        RECT 3385.940 2204.485 3386.110 2204.655 ;
        RECT 3380.500 2204.025 3380.670 2204.195 ;
        RECT 3385.940 2204.025 3386.110 2204.195 ;
        RECT 3380.500 2203.565 3380.670 2203.735 ;
        RECT 3385.940 2203.565 3386.110 2203.735 ;
        RECT 3380.500 2203.105 3380.670 2203.275 ;
        RECT 3385.940 2203.105 3386.110 2203.275 ;
        RECT 3380.500 2202.645 3380.670 2202.815 ;
        RECT 3385.940 2202.645 3386.110 2202.815 ;
        RECT 3380.500 2202.185 3380.670 2202.355 ;
        RECT 3385.940 2202.185 3386.110 2202.355 ;
        RECT 3380.500 2201.725 3380.670 2201.895 ;
        RECT 3385.940 2201.725 3386.110 2201.895 ;
        RECT 3380.500 2201.265 3380.670 2201.435 ;
        RECT 3385.940 2201.265 3386.110 2201.435 ;
        RECT 3380.500 2200.805 3380.670 2200.975 ;
        RECT 3385.940 2200.805 3386.110 2200.975 ;
        RECT 3380.500 2200.345 3380.670 2200.515 ;
        RECT 3385.940 2200.345 3386.110 2200.515 ;
        RECT 3380.500 2199.885 3380.670 2200.055 ;
        RECT 3385.940 2199.885 3386.110 2200.055 ;
        RECT 3380.500 2199.425 3380.670 2199.595 ;
        RECT 3385.940 2199.425 3386.110 2199.595 ;
        RECT 3380.500 2198.965 3380.670 2199.135 ;
        RECT 3385.940 2198.965 3386.110 2199.135 ;
        RECT 3380.500 2198.505 3380.670 2198.675 ;
        RECT 3385.940 2198.505 3386.110 2198.675 ;
        RECT 3380.500 2198.045 3380.670 2198.215 ;
        RECT 3385.940 2198.045 3386.110 2198.215 ;
        RECT 3380.500 2197.585 3380.670 2197.755 ;
        RECT 3385.940 2197.585 3386.110 2197.755 ;
        RECT 3380.500 2197.125 3380.670 2197.295 ;
        RECT 3385.940 2197.125 3386.110 2197.295 ;
        RECT 3380.500 2196.665 3380.670 2196.835 ;
        RECT 3385.940 2196.665 3386.110 2196.835 ;
        RECT 3380.500 2196.205 3380.670 2196.375 ;
        RECT 3385.940 2196.205 3386.110 2196.375 ;
      LAYER mcon ;
        RECT 3380.500 2237.145 3380.670 2237.315 ;
        RECT 3380.500 2236.685 3380.670 2236.855 ;
        RECT 3380.500 2236.225 3380.670 2236.395 ;
        RECT 3380.500 2235.765 3380.670 2235.935 ;
        RECT 3380.500 2235.305 3380.670 2235.475 ;
        RECT 3380.500 2234.845 3380.670 2235.015 ;
        RECT 3380.500 2234.385 3380.670 2234.555 ;
        RECT 3380.500 2233.925 3380.670 2234.095 ;
        RECT 3380.500 2233.465 3380.670 2233.635 ;
        RECT 3380.500 2233.005 3380.670 2233.175 ;
        RECT 3380.500 2232.545 3380.670 2232.715 ;
      LAYER met1 ;
        RECT 3380.345 2196.060 3380.825 2242.390 ;
        RECT 3385.785 2196.060 3386.265 2242.380 ;
      LAYER via ;
        RECT 3380.425 2240.475 3380.725 2242.260 ;
        RECT 3385.835 2240.475 3386.135 2242.260 ;
      LAYER met2 ;
        RECT 3380.365 2240.435 3380.795 2242.300 ;
        RECT 3385.790 2240.435 3386.220 2242.300 ;
      LAYER via2 ;
        RECT 3380.425 2240.475 3380.725 2242.260 ;
        RECT 3385.835 2240.475 3386.135 2242.260 ;
      LAYER met3 ;
        RECT 3380.350 2240.440 3387.875 2242.305 ;
    END
    PORT
      LAYER li1 ;
        RECT 3380.500 3608.185 3380.670 3608.355 ;
        RECT 3385.940 3608.185 3386.110 3608.355 ;
        RECT 3380.500 3607.725 3380.670 3607.895 ;
        RECT 3385.940 3607.725 3386.110 3607.895 ;
        RECT 3380.500 3607.265 3380.670 3607.435 ;
        RECT 3385.940 3607.265 3386.110 3607.435 ;
        RECT 3380.500 3606.805 3380.670 3606.975 ;
        RECT 3385.940 3606.805 3386.110 3606.975 ;
        RECT 3380.500 3606.345 3380.670 3606.515 ;
        RECT 3385.940 3606.345 3386.110 3606.515 ;
        RECT 3380.500 3605.885 3380.670 3606.055 ;
        RECT 3385.940 3605.885 3386.110 3606.055 ;
        RECT 3380.500 3605.425 3380.670 3605.595 ;
        RECT 3385.940 3605.425 3386.110 3605.595 ;
        RECT 3380.500 3604.965 3380.670 3605.135 ;
        RECT 3385.940 3604.965 3386.110 3605.135 ;
        RECT 3380.500 3604.505 3380.670 3604.675 ;
        RECT 3385.940 3604.505 3386.110 3604.675 ;
        RECT 3380.500 3604.045 3380.670 3604.215 ;
        RECT 3385.940 3604.045 3386.110 3604.215 ;
        RECT 3380.500 3603.585 3380.670 3603.755 ;
        RECT 3385.940 3603.585 3386.110 3603.755 ;
        RECT 3380.500 3603.125 3380.670 3603.295 ;
        RECT 3385.940 3603.125 3386.110 3603.295 ;
        RECT 3380.500 3602.665 3380.670 3602.835 ;
        RECT 3385.940 3602.665 3386.110 3602.835 ;
        RECT 3380.500 3602.205 3380.670 3602.375 ;
        RECT 3385.940 3602.205 3386.110 3602.375 ;
      LAYER met1 ;
        RECT 3380.345 3602.060 3380.825 3624.410 ;
        RECT 3385.785 3602.060 3386.265 3624.470 ;
      LAYER via ;
        RECT 3380.465 3622.480 3380.765 3624.265 ;
        RECT 3385.875 3622.480 3386.175 3624.265 ;
      LAYER met2 ;
        RECT 3380.405 3622.440 3380.835 3624.305 ;
        RECT 3385.830 3622.440 3386.260 3624.305 ;
      LAYER via2 ;
        RECT 3380.465 3622.480 3380.765 3624.265 ;
        RECT 3385.875 3622.480 3386.175 3624.265 ;
      LAYER met3 ;
        RECT 3380.390 3622.445 3387.915 3624.310 ;
    END
    PORT
      LAYER li1 ;
        RECT 671.130 217.755 671.470 218.585 ;
        RECT 677.110 217.755 677.450 218.585 ;
        RECT 683.090 217.755 683.430 218.585 ;
        RECT 689.070 217.755 689.410 218.585 ;
        RECT 712.990 217.755 713.330 218.585 ;
        RECT 718.970 217.755 719.310 218.585 ;
        RECT 724.950 217.755 725.290 218.585 ;
        RECT 790.730 217.755 791.070 218.585 ;
        RECT 669.545 217.210 674.890 217.755 ;
        RECT 675.525 217.210 680.870 217.755 ;
        RECT 681.505 217.210 686.850 217.755 ;
        RECT 687.485 217.210 692.830 217.755 ;
        RECT 711.405 217.210 716.750 217.755 ;
        RECT 717.385 217.210 722.730 217.755 ;
        RECT 723.365 217.210 728.710 217.755 ;
        RECT 789.145 217.210 794.490 217.755 ;
      LAYER li1 ;
        RECT 669.145 217.040 669.315 217.210 ;
      LAYER li1 ;
        RECT 669.460 217.040 669.605 217.210 ;
        RECT 669.775 217.040 674.980 217.210 ;
      LAYER li1 ;
        RECT 675.125 217.040 675.295 217.210 ;
      LAYER li1 ;
        RECT 675.440 217.040 675.585 217.210 ;
        RECT 675.755 217.040 680.960 217.210 ;
      LAYER li1 ;
        RECT 681.105 217.040 681.275 217.210 ;
      LAYER li1 ;
        RECT 681.420 217.040 681.565 217.210 ;
        RECT 681.735 217.040 686.940 217.210 ;
      LAYER li1 ;
        RECT 687.085 217.040 687.255 217.210 ;
      LAYER li1 ;
        RECT 687.400 217.040 687.545 217.210 ;
        RECT 687.715 217.040 692.920 217.210 ;
      LAYER li1 ;
        RECT 693.065 217.040 693.235 217.210 ;
        RECT 693.525 217.040 693.695 217.210 ;
        RECT 693.985 217.040 694.155 217.210 ;
        RECT 694.445 217.040 694.615 217.210 ;
        RECT 694.905 217.040 695.075 217.210 ;
        RECT 695.365 217.040 695.535 217.210 ;
        RECT 695.825 217.040 695.995 217.210 ;
        RECT 696.285 217.040 696.455 217.210 ;
        RECT 696.745 217.040 696.915 217.210 ;
        RECT 697.205 217.040 697.375 217.210 ;
        RECT 697.665 217.040 697.835 217.210 ;
        RECT 698.125 217.040 698.295 217.210 ;
        RECT 698.585 217.040 698.755 217.210 ;
        RECT 699.045 217.040 699.215 217.210 ;
        RECT 699.505 217.040 699.675 217.210 ;
        RECT 699.965 217.040 700.135 217.210 ;
        RECT 700.425 217.040 700.595 217.210 ;
        RECT 700.885 217.040 701.055 217.210 ;
        RECT 701.345 217.040 701.515 217.210 ;
        RECT 701.805 217.040 701.975 217.210 ;
        RECT 702.265 217.040 702.435 217.210 ;
        RECT 702.725 217.040 702.895 217.210 ;
        RECT 703.185 217.040 703.355 217.210 ;
        RECT 703.645 217.040 703.815 217.210 ;
        RECT 704.105 217.040 704.275 217.210 ;
        RECT 704.565 217.040 704.735 217.210 ;
        RECT 705.025 217.040 705.195 217.210 ;
        RECT 705.485 217.040 705.655 217.210 ;
        RECT 705.945 217.040 706.115 217.210 ;
        RECT 706.405 217.040 706.575 217.210 ;
        RECT 706.865 217.040 707.035 217.210 ;
        RECT 707.325 217.040 707.495 217.210 ;
        RECT 707.785 217.040 707.955 217.210 ;
        RECT 708.245 217.040 708.415 217.210 ;
        RECT 708.705 217.040 708.875 217.210 ;
        RECT 709.165 217.040 709.335 217.210 ;
        RECT 709.625 217.040 709.795 217.210 ;
        RECT 710.085 217.040 710.255 217.210 ;
        RECT 710.545 217.040 710.715 217.210 ;
        RECT 711.005 217.040 711.175 217.210 ;
      LAYER li1 ;
        RECT 711.320 217.040 711.465 217.210 ;
        RECT 711.635 217.040 716.840 217.210 ;
      LAYER li1 ;
        RECT 716.985 217.040 717.155 217.210 ;
      LAYER li1 ;
        RECT 717.300 217.040 717.445 217.210 ;
        RECT 717.615 217.040 722.820 217.210 ;
      LAYER li1 ;
        RECT 722.965 217.040 723.135 217.210 ;
      LAYER li1 ;
        RECT 723.280 217.040 728.800 217.210 ;
      LAYER li1 ;
        RECT 728.945 217.040 729.115 217.210 ;
        RECT 758.845 217.040 759.015 217.210 ;
        RECT 759.305 217.040 759.475 217.210 ;
        RECT 759.765 217.040 759.935 217.210 ;
        RECT 760.225 217.040 760.395 217.210 ;
        RECT 760.685 217.040 760.855 217.210 ;
        RECT 761.145 217.040 761.315 217.210 ;
        RECT 761.605 217.040 761.775 217.210 ;
        RECT 762.065 217.040 762.235 217.210 ;
        RECT 762.525 217.040 762.695 217.210 ;
        RECT 762.985 217.040 763.155 217.210 ;
        RECT 763.445 217.040 763.615 217.210 ;
        RECT 763.905 217.040 764.075 217.210 ;
        RECT 764.365 217.040 764.535 217.210 ;
        RECT 764.825 217.040 764.995 217.210 ;
        RECT 765.285 217.040 765.455 217.210 ;
        RECT 765.745 217.040 765.915 217.210 ;
        RECT 766.205 217.040 766.375 217.210 ;
        RECT 766.665 217.040 766.835 217.210 ;
        RECT 767.125 217.040 767.295 217.210 ;
        RECT 767.585 217.040 767.755 217.210 ;
        RECT 768.045 217.040 768.215 217.210 ;
        RECT 768.505 217.040 768.675 217.210 ;
        RECT 768.965 217.040 769.135 217.210 ;
        RECT 769.425 217.040 769.595 217.210 ;
        RECT 769.885 217.040 770.055 217.210 ;
        RECT 770.345 217.040 770.515 217.210 ;
        RECT 770.805 217.040 770.975 217.210 ;
        RECT 771.265 217.040 771.435 217.210 ;
        RECT 771.725 217.040 771.895 217.210 ;
        RECT 772.185 217.040 772.355 217.210 ;
        RECT 772.645 217.040 772.815 217.210 ;
        RECT 773.105 217.040 773.275 217.210 ;
        RECT 773.565 217.040 773.735 217.210 ;
        RECT 774.025 217.040 774.195 217.210 ;
        RECT 774.485 217.040 774.655 217.210 ;
        RECT 774.945 217.040 775.115 217.210 ;
        RECT 775.405 217.040 775.575 217.210 ;
        RECT 775.865 217.040 776.035 217.210 ;
        RECT 776.325 217.040 776.495 217.210 ;
        RECT 776.785 217.040 776.955 217.210 ;
        RECT 777.245 217.040 777.415 217.210 ;
        RECT 777.705 217.040 777.875 217.210 ;
        RECT 778.165 217.040 778.335 217.210 ;
        RECT 778.625 217.040 778.795 217.210 ;
        RECT 779.085 217.040 779.255 217.210 ;
        RECT 779.545 217.040 779.715 217.210 ;
        RECT 780.005 217.040 780.175 217.210 ;
        RECT 780.465 217.040 780.635 217.210 ;
        RECT 780.925 217.040 781.095 217.210 ;
        RECT 781.385 217.040 781.555 217.210 ;
        RECT 781.845 217.040 782.015 217.210 ;
        RECT 782.305 217.040 782.475 217.210 ;
        RECT 782.765 217.040 782.935 217.210 ;
        RECT 783.225 217.040 783.395 217.210 ;
        RECT 783.685 217.040 783.855 217.210 ;
        RECT 784.145 217.040 784.315 217.210 ;
        RECT 784.605 217.040 784.775 217.210 ;
        RECT 785.065 217.040 785.235 217.210 ;
        RECT 785.525 217.040 785.695 217.210 ;
        RECT 785.985 217.040 786.155 217.210 ;
        RECT 786.445 217.040 786.615 217.210 ;
        RECT 786.905 217.040 787.075 217.210 ;
        RECT 787.365 217.040 787.535 217.210 ;
        RECT 787.825 217.040 787.995 217.210 ;
        RECT 788.285 217.040 788.455 217.210 ;
        RECT 788.745 217.040 788.915 217.210 ;
      LAYER li1 ;
        RECT 789.060 217.040 789.205 217.210 ;
        RECT 789.375 217.040 794.580 217.210 ;
      LAYER li1 ;
        RECT 794.725 217.040 794.895 217.210 ;
      LAYER li1 ;
        RECT 723.365 216.495 728.710 217.040 ;
        RECT 724.950 215.665 725.290 216.495 ;
        RECT 671.130 212.315 671.470 213.145 ;
        RECT 760.830 212.315 761.170 213.145 ;
        RECT 669.545 211.770 674.890 212.315 ;
        RECT 759.245 211.770 764.590 212.315 ;
      LAYER li1 ;
        RECT 669.145 211.600 669.315 211.770 ;
      LAYER li1 ;
        RECT 669.460 211.600 674.980 211.770 ;
      LAYER li1 ;
        RECT 675.125 211.600 675.295 211.770 ;
        RECT 675.585 211.600 675.755 211.770 ;
        RECT 676.045 211.600 676.215 211.770 ;
        RECT 676.505 211.600 676.675 211.770 ;
        RECT 676.965 211.600 677.135 211.770 ;
        RECT 677.425 211.600 677.595 211.770 ;
        RECT 677.885 211.600 678.055 211.770 ;
        RECT 678.345 211.600 678.515 211.770 ;
        RECT 678.805 211.600 678.975 211.770 ;
        RECT 679.265 211.600 679.435 211.770 ;
        RECT 679.725 211.600 679.895 211.770 ;
        RECT 680.185 211.600 680.355 211.770 ;
        RECT 680.645 211.600 680.815 211.770 ;
        RECT 681.105 211.600 681.275 211.770 ;
        RECT 681.565 211.600 681.735 211.770 ;
        RECT 682.025 211.600 682.195 211.770 ;
        RECT 682.485 211.600 682.655 211.770 ;
        RECT 682.945 211.600 683.115 211.770 ;
        RECT 683.405 211.600 683.575 211.770 ;
        RECT 683.865 211.600 684.035 211.770 ;
        RECT 684.325 211.600 684.495 211.770 ;
        RECT 684.785 211.600 684.955 211.770 ;
        RECT 685.245 211.600 685.415 211.770 ;
        RECT 685.705 211.600 685.875 211.770 ;
        RECT 686.165 211.600 686.335 211.770 ;
        RECT 686.625 211.600 686.795 211.770 ;
        RECT 687.085 211.600 687.255 211.770 ;
        RECT 687.545 211.600 687.715 211.770 ;
        RECT 688.005 211.600 688.175 211.770 ;
        RECT 688.465 211.600 688.635 211.770 ;
        RECT 688.925 211.600 689.095 211.770 ;
        RECT 689.385 211.600 689.555 211.770 ;
        RECT 689.845 211.600 690.015 211.770 ;
        RECT 690.305 211.600 690.475 211.770 ;
        RECT 690.765 211.600 690.935 211.770 ;
        RECT 691.225 211.600 691.395 211.770 ;
        RECT 691.685 211.600 691.855 211.770 ;
        RECT 692.145 211.600 692.315 211.770 ;
        RECT 692.605 211.600 692.775 211.770 ;
        RECT 693.065 211.600 693.235 211.770 ;
        RECT 693.525 211.600 693.695 211.770 ;
        RECT 693.985 211.600 694.155 211.770 ;
        RECT 694.445 211.600 694.615 211.770 ;
        RECT 694.905 211.600 695.075 211.770 ;
        RECT 695.365 211.600 695.535 211.770 ;
        RECT 695.825 211.600 695.995 211.770 ;
        RECT 696.285 211.600 696.455 211.770 ;
        RECT 696.745 211.600 696.915 211.770 ;
        RECT 697.205 211.600 697.375 211.770 ;
        RECT 697.665 211.600 697.835 211.770 ;
        RECT 698.125 211.600 698.295 211.770 ;
        RECT 698.585 211.600 698.755 211.770 ;
        RECT 699.045 211.600 699.215 211.770 ;
        RECT 699.505 211.600 699.675 211.770 ;
        RECT 699.965 211.600 700.135 211.770 ;
        RECT 700.425 211.600 700.595 211.770 ;
        RECT 700.885 211.600 701.055 211.770 ;
        RECT 701.345 211.600 701.515 211.770 ;
        RECT 701.805 211.600 701.975 211.770 ;
        RECT 702.265 211.600 702.435 211.770 ;
        RECT 702.725 211.600 702.895 211.770 ;
        RECT 703.185 211.600 703.355 211.770 ;
        RECT 703.645 211.600 703.815 211.770 ;
        RECT 704.105 211.600 704.275 211.770 ;
        RECT 704.565 211.600 704.735 211.770 ;
        RECT 705.025 211.600 705.195 211.770 ;
        RECT 705.485 211.600 705.655 211.770 ;
        RECT 705.945 211.600 706.115 211.770 ;
        RECT 706.405 211.600 706.575 211.770 ;
        RECT 706.865 211.600 707.035 211.770 ;
        RECT 707.325 211.600 707.495 211.770 ;
        RECT 707.785 211.600 707.955 211.770 ;
        RECT 708.245 211.600 708.415 211.770 ;
        RECT 708.705 211.600 708.875 211.770 ;
        RECT 709.165 211.600 709.335 211.770 ;
        RECT 709.625 211.600 709.795 211.770 ;
        RECT 710.085 211.600 710.255 211.770 ;
        RECT 710.545 211.600 710.715 211.770 ;
        RECT 711.005 211.600 711.175 211.770 ;
        RECT 711.465 211.600 711.635 211.770 ;
        RECT 711.925 211.600 712.095 211.770 ;
        RECT 712.385 211.600 712.555 211.770 ;
        RECT 712.845 211.600 713.015 211.770 ;
        RECT 713.305 211.600 713.475 211.770 ;
        RECT 713.765 211.600 713.935 211.770 ;
        RECT 714.225 211.600 714.395 211.770 ;
        RECT 714.685 211.600 714.855 211.770 ;
        RECT 715.145 211.600 715.315 211.770 ;
        RECT 715.605 211.600 715.775 211.770 ;
        RECT 716.065 211.600 716.235 211.770 ;
        RECT 716.525 211.600 716.695 211.770 ;
        RECT 716.985 211.600 717.155 211.770 ;
        RECT 717.445 211.600 717.615 211.770 ;
        RECT 717.905 211.600 718.075 211.770 ;
        RECT 718.365 211.600 718.535 211.770 ;
        RECT 718.825 211.600 718.995 211.770 ;
        RECT 719.285 211.600 719.455 211.770 ;
        RECT 719.745 211.600 719.915 211.770 ;
        RECT 720.205 211.600 720.375 211.770 ;
        RECT 720.665 211.600 720.835 211.770 ;
        RECT 721.125 211.600 721.295 211.770 ;
        RECT 721.585 211.600 721.755 211.770 ;
        RECT 722.045 211.600 722.215 211.770 ;
        RECT 722.505 211.600 722.675 211.770 ;
        RECT 722.965 211.600 723.135 211.770 ;
        RECT 723.425 211.600 723.595 211.770 ;
        RECT 723.885 211.600 724.055 211.770 ;
        RECT 724.345 211.600 724.515 211.770 ;
        RECT 724.805 211.600 724.975 211.770 ;
        RECT 725.265 211.600 725.435 211.770 ;
        RECT 725.725 211.600 725.895 211.770 ;
        RECT 726.185 211.600 726.355 211.770 ;
        RECT 726.645 211.600 726.815 211.770 ;
        RECT 727.105 211.600 727.275 211.770 ;
        RECT 727.565 211.600 727.735 211.770 ;
        RECT 728.025 211.600 728.195 211.770 ;
        RECT 728.485 211.600 728.655 211.770 ;
        RECT 728.945 211.600 729.115 211.770 ;
        RECT 758.845 211.600 759.015 211.770 ;
      LAYER li1 ;
        RECT 759.160 211.600 764.680 211.770 ;
      LAYER li1 ;
        RECT 764.825 211.600 764.995 211.770 ;
        RECT 765.285 211.600 765.455 211.770 ;
        RECT 765.745 211.600 765.915 211.770 ;
        RECT 766.205 211.600 766.375 211.770 ;
        RECT 766.665 211.600 766.835 211.770 ;
        RECT 767.125 211.600 767.295 211.770 ;
        RECT 767.585 211.600 767.755 211.770 ;
        RECT 768.045 211.600 768.215 211.770 ;
        RECT 768.505 211.600 768.675 211.770 ;
        RECT 768.965 211.600 769.135 211.770 ;
        RECT 769.425 211.600 769.595 211.770 ;
        RECT 769.885 211.600 770.055 211.770 ;
        RECT 770.345 211.600 770.515 211.770 ;
        RECT 770.805 211.600 770.975 211.770 ;
        RECT 771.265 211.600 771.435 211.770 ;
        RECT 771.725 211.600 771.895 211.770 ;
        RECT 772.185 211.600 772.355 211.770 ;
        RECT 772.645 211.600 772.815 211.770 ;
        RECT 773.105 211.600 773.275 211.770 ;
        RECT 773.565 211.600 773.735 211.770 ;
        RECT 774.025 211.600 774.195 211.770 ;
        RECT 774.485 211.600 774.655 211.770 ;
        RECT 774.945 211.600 775.115 211.770 ;
        RECT 775.405 211.600 775.575 211.770 ;
        RECT 775.865 211.600 776.035 211.770 ;
        RECT 776.325 211.600 776.495 211.770 ;
        RECT 776.785 211.600 776.955 211.770 ;
        RECT 777.245 211.600 777.415 211.770 ;
        RECT 777.705 211.600 777.875 211.770 ;
        RECT 778.165 211.600 778.335 211.770 ;
        RECT 778.625 211.600 778.795 211.770 ;
        RECT 779.085 211.600 779.255 211.770 ;
        RECT 779.545 211.600 779.715 211.770 ;
        RECT 780.005 211.600 780.175 211.770 ;
        RECT 780.465 211.600 780.635 211.770 ;
        RECT 780.925 211.600 781.095 211.770 ;
        RECT 781.385 211.600 781.555 211.770 ;
        RECT 781.845 211.600 782.015 211.770 ;
        RECT 782.305 211.600 782.475 211.770 ;
        RECT 782.765 211.600 782.935 211.770 ;
        RECT 783.225 211.600 783.395 211.770 ;
        RECT 783.685 211.600 783.855 211.770 ;
        RECT 784.145 211.600 784.315 211.770 ;
        RECT 784.605 211.600 784.775 211.770 ;
        RECT 785.065 211.600 785.235 211.770 ;
        RECT 785.525 211.600 785.695 211.770 ;
        RECT 785.985 211.600 786.155 211.770 ;
        RECT 786.445 211.600 786.615 211.770 ;
        RECT 786.905 211.600 787.075 211.770 ;
        RECT 787.365 211.600 787.535 211.770 ;
        RECT 787.825 211.600 787.995 211.770 ;
        RECT 788.285 211.600 788.455 211.770 ;
        RECT 788.745 211.600 788.915 211.770 ;
        RECT 789.205 211.600 789.375 211.770 ;
        RECT 789.665 211.600 789.835 211.770 ;
        RECT 790.125 211.600 790.295 211.770 ;
        RECT 790.585 211.600 790.755 211.770 ;
        RECT 791.045 211.600 791.215 211.770 ;
        RECT 791.505 211.600 791.675 211.770 ;
        RECT 791.965 211.600 792.135 211.770 ;
        RECT 792.425 211.600 792.595 211.770 ;
        RECT 792.885 211.600 793.055 211.770 ;
        RECT 793.345 211.600 793.515 211.770 ;
        RECT 793.805 211.600 793.975 211.770 ;
        RECT 794.265 211.600 794.435 211.770 ;
        RECT 794.725 211.600 794.895 211.770 ;
      LAYER mcon ;
        RECT 670.065 217.040 670.235 217.210 ;
        RECT 670.525 217.040 670.695 217.210 ;
        RECT 670.985 217.040 671.155 217.210 ;
        RECT 671.445 217.040 671.615 217.210 ;
        RECT 671.905 217.040 672.075 217.210 ;
        RECT 672.365 217.040 672.535 217.210 ;
        RECT 672.825 217.040 672.995 217.210 ;
        RECT 673.285 217.040 673.455 217.210 ;
        RECT 673.745 217.040 673.915 217.210 ;
        RECT 674.205 217.040 674.375 217.210 ;
        RECT 674.665 217.040 674.835 217.210 ;
        RECT 676.045 217.040 676.215 217.210 ;
        RECT 676.505 217.040 676.675 217.210 ;
        RECT 676.965 217.040 677.135 217.210 ;
        RECT 677.425 217.040 677.595 217.210 ;
        RECT 677.885 217.040 678.055 217.210 ;
        RECT 678.345 217.040 678.515 217.210 ;
        RECT 678.805 217.040 678.975 217.210 ;
        RECT 679.265 217.040 679.435 217.210 ;
        RECT 679.725 217.040 679.895 217.210 ;
        RECT 680.185 217.040 680.355 217.210 ;
        RECT 680.645 217.040 680.815 217.210 ;
        RECT 682.025 217.040 682.195 217.210 ;
        RECT 682.485 217.040 682.655 217.210 ;
        RECT 682.945 217.040 683.115 217.210 ;
        RECT 683.405 217.040 683.575 217.210 ;
        RECT 683.865 217.040 684.035 217.210 ;
        RECT 684.325 217.040 684.495 217.210 ;
        RECT 684.785 217.040 684.955 217.210 ;
        RECT 685.245 217.040 685.415 217.210 ;
        RECT 685.705 217.040 685.875 217.210 ;
        RECT 686.165 217.040 686.335 217.210 ;
        RECT 686.625 217.040 686.795 217.210 ;
        RECT 688.005 217.040 688.175 217.210 ;
        RECT 688.465 217.040 688.635 217.210 ;
        RECT 688.925 217.040 689.095 217.210 ;
        RECT 689.385 217.040 689.555 217.210 ;
        RECT 689.845 217.040 690.015 217.210 ;
        RECT 690.305 217.040 690.475 217.210 ;
        RECT 690.765 217.040 690.935 217.210 ;
        RECT 691.225 217.040 691.395 217.210 ;
        RECT 691.685 217.040 691.855 217.210 ;
        RECT 692.145 217.040 692.315 217.210 ;
        RECT 692.605 217.040 692.775 217.210 ;
        RECT 711.925 217.040 712.095 217.210 ;
        RECT 712.385 217.040 712.555 217.210 ;
        RECT 712.845 217.040 713.015 217.210 ;
        RECT 713.305 217.040 713.475 217.210 ;
        RECT 713.765 217.040 713.935 217.210 ;
        RECT 714.225 217.040 714.395 217.210 ;
        RECT 714.685 217.040 714.855 217.210 ;
        RECT 715.145 217.040 715.315 217.210 ;
        RECT 715.605 217.040 715.775 217.210 ;
        RECT 716.065 217.040 716.235 217.210 ;
        RECT 716.525 217.040 716.695 217.210 ;
        RECT 717.905 217.040 718.075 217.210 ;
        RECT 718.365 217.040 718.535 217.210 ;
        RECT 718.825 217.040 718.995 217.210 ;
        RECT 719.285 217.040 719.455 217.210 ;
        RECT 719.745 217.040 719.915 217.210 ;
        RECT 720.205 217.040 720.375 217.210 ;
        RECT 720.665 217.040 720.835 217.210 ;
        RECT 721.125 217.040 721.295 217.210 ;
        RECT 721.585 217.040 721.755 217.210 ;
        RECT 722.045 217.040 722.215 217.210 ;
        RECT 722.505 217.040 722.675 217.210 ;
        RECT 723.885 217.040 724.055 217.210 ;
        RECT 724.345 217.040 724.515 217.210 ;
        RECT 724.805 217.040 724.975 217.210 ;
        RECT 725.265 217.040 725.435 217.210 ;
        RECT 725.725 217.040 725.895 217.210 ;
        RECT 726.185 217.040 726.355 217.210 ;
        RECT 726.645 217.040 726.815 217.210 ;
        RECT 727.105 217.040 727.275 217.210 ;
        RECT 727.565 217.040 727.735 217.210 ;
        RECT 728.025 217.040 728.195 217.210 ;
        RECT 728.485 217.040 728.655 217.210 ;
        RECT 789.665 217.040 789.835 217.210 ;
        RECT 790.125 217.040 790.295 217.210 ;
        RECT 790.585 217.040 790.755 217.210 ;
        RECT 791.045 217.040 791.215 217.210 ;
        RECT 791.505 217.040 791.675 217.210 ;
        RECT 791.965 217.040 792.135 217.210 ;
        RECT 792.425 217.040 792.595 217.210 ;
        RECT 792.885 217.040 793.055 217.210 ;
        RECT 793.345 217.040 793.515 217.210 ;
        RECT 793.805 217.040 793.975 217.210 ;
        RECT 794.265 217.040 794.435 217.210 ;
        RECT 670.065 211.600 670.235 211.770 ;
        RECT 670.525 211.600 670.695 211.770 ;
        RECT 670.985 211.600 671.155 211.770 ;
        RECT 671.445 211.600 671.615 211.770 ;
        RECT 671.905 211.600 672.075 211.770 ;
        RECT 672.365 211.600 672.535 211.770 ;
        RECT 672.825 211.600 672.995 211.770 ;
        RECT 673.285 211.600 673.455 211.770 ;
        RECT 673.745 211.600 673.915 211.770 ;
        RECT 674.205 211.600 674.375 211.770 ;
        RECT 674.665 211.600 674.835 211.770 ;
        RECT 759.765 211.600 759.935 211.770 ;
        RECT 760.225 211.600 760.395 211.770 ;
        RECT 760.685 211.600 760.855 211.770 ;
        RECT 761.145 211.600 761.315 211.770 ;
        RECT 761.605 211.600 761.775 211.770 ;
        RECT 762.065 211.600 762.235 211.770 ;
        RECT 762.525 211.600 762.695 211.770 ;
        RECT 762.985 211.600 763.155 211.770 ;
        RECT 763.445 211.600 763.615 211.770 ;
        RECT 763.905 211.600 764.075 211.770 ;
        RECT 764.365 211.600 764.535 211.770 ;
      LAYER met1 ;
        RECT 669.000 216.885 795.040 217.365 ;
        RECT 669.000 211.445 795.040 211.925 ;
      LAYER via ;
        RECT 736.975 216.985 738.760 217.285 ;
        RECT 736.975 211.575 738.760 211.875 ;
      LAYER met2 ;
        RECT 736.935 216.915 738.800 217.345 ;
        RECT 736.935 211.490 738.800 211.920 ;
      LAYER via2 ;
        RECT 736.975 216.985 738.760 217.285 ;
        RECT 736.975 211.575 738.760 211.875 ;
      LAYER met3 ;
        RECT 736.940 209.835 738.805 217.360 ;
    END
    PORT
      LAYER li1 ;
        RECT 2148.130 217.755 2148.470 218.585 ;
        RECT 2154.110 217.755 2154.450 218.585 ;
        RECT 2160.090 217.755 2160.430 218.585 ;
        RECT 2166.070 217.755 2166.410 218.585 ;
        RECT 2172.050 217.755 2172.390 218.585 ;
        RECT 2178.030 217.755 2178.370 218.585 ;
        RECT 2184.010 217.755 2184.350 218.585 ;
        RECT 2189.990 217.755 2190.330 218.585 ;
        RECT 2195.970 217.755 2196.310 218.585 ;
        RECT 2201.950 217.755 2202.290 218.585 ;
        RECT 2237.830 217.755 2238.170 218.585 ;
        RECT 2243.810 217.755 2244.150 218.585 ;
        RECT 2249.790 217.755 2250.130 218.585 ;
        RECT 2255.770 217.755 2256.110 218.585 ;
        RECT 2261.750 217.755 2262.090 218.585 ;
        RECT 2267.730 217.755 2268.070 218.585 ;
        RECT 2146.545 217.210 2151.890 217.755 ;
        RECT 2152.525 217.210 2157.870 217.755 ;
        RECT 2158.505 217.210 2163.850 217.755 ;
        RECT 2164.485 217.210 2169.830 217.755 ;
        RECT 2170.465 217.210 2175.810 217.755 ;
        RECT 2176.445 217.210 2181.790 217.755 ;
        RECT 2182.425 217.210 2187.770 217.755 ;
        RECT 2188.405 217.210 2193.750 217.755 ;
        RECT 2194.385 217.210 2199.730 217.755 ;
        RECT 2200.365 217.210 2205.710 217.755 ;
        RECT 2236.245 217.210 2241.590 217.755 ;
        RECT 2242.225 217.210 2247.570 217.755 ;
        RECT 2248.205 217.210 2253.550 217.755 ;
        RECT 2254.185 217.210 2259.530 217.755 ;
        RECT 2260.165 217.210 2265.510 217.755 ;
        RECT 2266.145 217.210 2271.490 217.755 ;
      LAYER li1 ;
        RECT 2146.145 217.040 2146.315 217.210 ;
      LAYER li1 ;
        RECT 2146.460 217.040 2146.605 217.210 ;
        RECT 2146.775 217.040 2151.980 217.210 ;
      LAYER li1 ;
        RECT 2152.125 217.040 2152.295 217.210 ;
      LAYER li1 ;
        RECT 2152.440 217.040 2152.585 217.210 ;
        RECT 2152.755 217.040 2157.960 217.210 ;
      LAYER li1 ;
        RECT 2158.105 217.040 2158.275 217.210 ;
      LAYER li1 ;
        RECT 2158.420 217.040 2158.565 217.210 ;
        RECT 2158.735 217.040 2163.940 217.210 ;
      LAYER li1 ;
        RECT 2164.085 217.040 2164.255 217.210 ;
      LAYER li1 ;
        RECT 2164.400 217.040 2164.545 217.210 ;
        RECT 2164.715 217.040 2169.920 217.210 ;
      LAYER li1 ;
        RECT 2170.065 217.040 2170.235 217.210 ;
      LAYER li1 ;
        RECT 2170.380 217.040 2170.525 217.210 ;
        RECT 2170.695 217.040 2175.900 217.210 ;
      LAYER li1 ;
        RECT 2176.045 217.040 2176.215 217.210 ;
      LAYER li1 ;
        RECT 2176.360 217.040 2176.505 217.210 ;
        RECT 2176.675 217.040 2181.880 217.210 ;
      LAYER li1 ;
        RECT 2182.025 217.040 2182.195 217.210 ;
      LAYER li1 ;
        RECT 2182.340 217.040 2182.485 217.210 ;
        RECT 2182.655 217.040 2187.860 217.210 ;
      LAYER li1 ;
        RECT 2188.005 217.040 2188.175 217.210 ;
      LAYER li1 ;
        RECT 2188.320 217.040 2188.465 217.210 ;
        RECT 2188.635 217.040 2193.840 217.210 ;
      LAYER li1 ;
        RECT 2193.985 217.040 2194.155 217.210 ;
      LAYER li1 ;
        RECT 2194.300 217.040 2194.445 217.210 ;
        RECT 2194.615 217.040 2199.820 217.210 ;
      LAYER li1 ;
        RECT 2199.965 217.040 2200.135 217.210 ;
      LAYER li1 ;
        RECT 2200.280 217.040 2205.800 217.210 ;
      LAYER li1 ;
        RECT 2205.945 217.040 2206.115 217.210 ;
        RECT 2235.845 217.040 2236.015 217.210 ;
      LAYER li1 ;
        RECT 2236.160 217.040 2236.305 217.210 ;
        RECT 2236.475 217.040 2241.680 217.210 ;
      LAYER li1 ;
        RECT 2241.825 217.040 2241.995 217.210 ;
      LAYER li1 ;
        RECT 2242.140 217.040 2242.285 217.210 ;
        RECT 2242.455 217.040 2247.660 217.210 ;
      LAYER li1 ;
        RECT 2247.805 217.040 2247.975 217.210 ;
      LAYER li1 ;
        RECT 2248.120 217.040 2248.265 217.210 ;
        RECT 2248.435 217.040 2253.640 217.210 ;
      LAYER li1 ;
        RECT 2253.785 217.040 2253.955 217.210 ;
      LAYER li1 ;
        RECT 2254.100 217.040 2254.245 217.210 ;
        RECT 2254.415 217.040 2259.620 217.210 ;
      LAYER li1 ;
        RECT 2259.765 217.040 2259.935 217.210 ;
      LAYER li1 ;
        RECT 2260.080 217.040 2260.225 217.210 ;
        RECT 2260.395 217.040 2265.600 217.210 ;
      LAYER li1 ;
        RECT 2265.745 217.040 2265.915 217.210 ;
      LAYER li1 ;
        RECT 2266.060 217.040 2266.205 217.210 ;
        RECT 2266.375 217.040 2271.580 217.210 ;
      LAYER li1 ;
        RECT 2271.725 217.040 2271.895 217.210 ;
      LAYER li1 ;
        RECT 2200.365 216.495 2205.710 217.040 ;
        RECT 2201.950 215.665 2202.290 216.495 ;
        RECT 2148.130 212.315 2148.470 213.145 ;
        RECT 2237.830 212.315 2238.170 213.145 ;
        RECT 2146.545 211.770 2151.890 212.315 ;
        RECT 2236.245 211.770 2241.590 212.315 ;
      LAYER li1 ;
        RECT 2146.145 211.600 2146.315 211.770 ;
      LAYER li1 ;
        RECT 2146.460 211.600 2151.980 211.770 ;
      LAYER li1 ;
        RECT 2152.125 211.600 2152.295 211.770 ;
        RECT 2152.585 211.600 2152.755 211.770 ;
        RECT 2153.045 211.600 2153.215 211.770 ;
        RECT 2153.505 211.600 2153.675 211.770 ;
        RECT 2153.965 211.600 2154.135 211.770 ;
        RECT 2154.425 211.600 2154.595 211.770 ;
        RECT 2154.885 211.600 2155.055 211.770 ;
        RECT 2155.345 211.600 2155.515 211.770 ;
        RECT 2155.805 211.600 2155.975 211.770 ;
        RECT 2156.265 211.600 2156.435 211.770 ;
        RECT 2156.725 211.600 2156.895 211.770 ;
        RECT 2157.185 211.600 2157.355 211.770 ;
        RECT 2157.645 211.600 2157.815 211.770 ;
        RECT 2158.105 211.600 2158.275 211.770 ;
        RECT 2158.565 211.600 2158.735 211.770 ;
        RECT 2159.025 211.600 2159.195 211.770 ;
        RECT 2159.485 211.600 2159.655 211.770 ;
        RECT 2159.945 211.600 2160.115 211.770 ;
        RECT 2160.405 211.600 2160.575 211.770 ;
        RECT 2160.865 211.600 2161.035 211.770 ;
        RECT 2161.325 211.600 2161.495 211.770 ;
        RECT 2161.785 211.600 2161.955 211.770 ;
        RECT 2162.245 211.600 2162.415 211.770 ;
        RECT 2162.705 211.600 2162.875 211.770 ;
        RECT 2163.165 211.600 2163.335 211.770 ;
        RECT 2163.625 211.600 2163.795 211.770 ;
        RECT 2164.085 211.600 2164.255 211.770 ;
        RECT 2164.545 211.600 2164.715 211.770 ;
        RECT 2165.005 211.600 2165.175 211.770 ;
        RECT 2165.465 211.600 2165.635 211.770 ;
        RECT 2165.925 211.600 2166.095 211.770 ;
        RECT 2166.385 211.600 2166.555 211.770 ;
        RECT 2166.845 211.600 2167.015 211.770 ;
        RECT 2167.305 211.600 2167.475 211.770 ;
        RECT 2167.765 211.600 2167.935 211.770 ;
        RECT 2168.225 211.600 2168.395 211.770 ;
        RECT 2168.685 211.600 2168.855 211.770 ;
        RECT 2169.145 211.600 2169.315 211.770 ;
        RECT 2169.605 211.600 2169.775 211.770 ;
        RECT 2170.065 211.600 2170.235 211.770 ;
        RECT 2170.525 211.600 2170.695 211.770 ;
        RECT 2170.985 211.600 2171.155 211.770 ;
        RECT 2171.445 211.600 2171.615 211.770 ;
        RECT 2171.905 211.600 2172.075 211.770 ;
        RECT 2172.365 211.600 2172.535 211.770 ;
        RECT 2172.825 211.600 2172.995 211.770 ;
        RECT 2173.285 211.600 2173.455 211.770 ;
        RECT 2173.745 211.600 2173.915 211.770 ;
        RECT 2174.205 211.600 2174.375 211.770 ;
        RECT 2174.665 211.600 2174.835 211.770 ;
        RECT 2175.125 211.600 2175.295 211.770 ;
        RECT 2175.585 211.600 2175.755 211.770 ;
        RECT 2176.045 211.600 2176.215 211.770 ;
        RECT 2176.505 211.600 2176.675 211.770 ;
        RECT 2176.965 211.600 2177.135 211.770 ;
        RECT 2177.425 211.600 2177.595 211.770 ;
        RECT 2177.885 211.600 2178.055 211.770 ;
        RECT 2178.345 211.600 2178.515 211.770 ;
        RECT 2178.805 211.600 2178.975 211.770 ;
        RECT 2179.265 211.600 2179.435 211.770 ;
        RECT 2179.725 211.600 2179.895 211.770 ;
        RECT 2180.185 211.600 2180.355 211.770 ;
        RECT 2180.645 211.600 2180.815 211.770 ;
        RECT 2181.105 211.600 2181.275 211.770 ;
        RECT 2181.565 211.600 2181.735 211.770 ;
        RECT 2182.025 211.600 2182.195 211.770 ;
        RECT 2182.485 211.600 2182.655 211.770 ;
        RECT 2182.945 211.600 2183.115 211.770 ;
        RECT 2183.405 211.600 2183.575 211.770 ;
        RECT 2183.865 211.600 2184.035 211.770 ;
        RECT 2184.325 211.600 2184.495 211.770 ;
        RECT 2184.785 211.600 2184.955 211.770 ;
        RECT 2185.245 211.600 2185.415 211.770 ;
        RECT 2185.705 211.600 2185.875 211.770 ;
        RECT 2186.165 211.600 2186.335 211.770 ;
        RECT 2186.625 211.600 2186.795 211.770 ;
        RECT 2187.085 211.600 2187.255 211.770 ;
        RECT 2187.545 211.600 2187.715 211.770 ;
        RECT 2188.005 211.600 2188.175 211.770 ;
        RECT 2188.465 211.600 2188.635 211.770 ;
        RECT 2188.925 211.600 2189.095 211.770 ;
        RECT 2189.385 211.600 2189.555 211.770 ;
        RECT 2189.845 211.600 2190.015 211.770 ;
        RECT 2190.305 211.600 2190.475 211.770 ;
        RECT 2190.765 211.600 2190.935 211.770 ;
        RECT 2191.225 211.600 2191.395 211.770 ;
        RECT 2191.685 211.600 2191.855 211.770 ;
        RECT 2192.145 211.600 2192.315 211.770 ;
        RECT 2192.605 211.600 2192.775 211.770 ;
        RECT 2193.065 211.600 2193.235 211.770 ;
        RECT 2193.525 211.600 2193.695 211.770 ;
        RECT 2193.985 211.600 2194.155 211.770 ;
        RECT 2194.445 211.600 2194.615 211.770 ;
        RECT 2194.905 211.600 2195.075 211.770 ;
        RECT 2195.365 211.600 2195.535 211.770 ;
        RECT 2195.825 211.600 2195.995 211.770 ;
        RECT 2196.285 211.600 2196.455 211.770 ;
        RECT 2196.745 211.600 2196.915 211.770 ;
        RECT 2197.205 211.600 2197.375 211.770 ;
        RECT 2197.665 211.600 2197.835 211.770 ;
        RECT 2198.125 211.600 2198.295 211.770 ;
        RECT 2198.585 211.600 2198.755 211.770 ;
        RECT 2199.045 211.600 2199.215 211.770 ;
        RECT 2199.505 211.600 2199.675 211.770 ;
        RECT 2199.965 211.600 2200.135 211.770 ;
        RECT 2200.425 211.600 2200.595 211.770 ;
        RECT 2200.885 211.600 2201.055 211.770 ;
        RECT 2201.345 211.600 2201.515 211.770 ;
        RECT 2201.805 211.600 2201.975 211.770 ;
        RECT 2202.265 211.600 2202.435 211.770 ;
        RECT 2202.725 211.600 2202.895 211.770 ;
        RECT 2203.185 211.600 2203.355 211.770 ;
        RECT 2203.645 211.600 2203.815 211.770 ;
        RECT 2204.105 211.600 2204.275 211.770 ;
        RECT 2204.565 211.600 2204.735 211.770 ;
        RECT 2205.025 211.600 2205.195 211.770 ;
        RECT 2205.485 211.600 2205.655 211.770 ;
        RECT 2205.945 211.600 2206.115 211.770 ;
        RECT 2235.845 211.600 2236.015 211.770 ;
      LAYER li1 ;
        RECT 2236.160 211.600 2241.680 211.770 ;
      LAYER li1 ;
        RECT 2241.825 211.600 2241.995 211.770 ;
        RECT 2242.285 211.600 2242.455 211.770 ;
        RECT 2242.745 211.600 2242.915 211.770 ;
        RECT 2243.205 211.600 2243.375 211.770 ;
        RECT 2243.665 211.600 2243.835 211.770 ;
        RECT 2244.125 211.600 2244.295 211.770 ;
        RECT 2244.585 211.600 2244.755 211.770 ;
        RECT 2245.045 211.600 2245.215 211.770 ;
        RECT 2245.505 211.600 2245.675 211.770 ;
        RECT 2245.965 211.600 2246.135 211.770 ;
        RECT 2246.425 211.600 2246.595 211.770 ;
        RECT 2246.885 211.600 2247.055 211.770 ;
        RECT 2247.345 211.600 2247.515 211.770 ;
        RECT 2247.805 211.600 2247.975 211.770 ;
        RECT 2248.265 211.600 2248.435 211.770 ;
        RECT 2248.725 211.600 2248.895 211.770 ;
        RECT 2249.185 211.600 2249.355 211.770 ;
        RECT 2249.645 211.600 2249.815 211.770 ;
        RECT 2250.105 211.600 2250.275 211.770 ;
        RECT 2250.565 211.600 2250.735 211.770 ;
        RECT 2251.025 211.600 2251.195 211.770 ;
        RECT 2251.485 211.600 2251.655 211.770 ;
        RECT 2251.945 211.600 2252.115 211.770 ;
        RECT 2252.405 211.600 2252.575 211.770 ;
        RECT 2252.865 211.600 2253.035 211.770 ;
        RECT 2253.325 211.600 2253.495 211.770 ;
        RECT 2253.785 211.600 2253.955 211.770 ;
        RECT 2254.245 211.600 2254.415 211.770 ;
        RECT 2254.705 211.600 2254.875 211.770 ;
        RECT 2255.165 211.600 2255.335 211.770 ;
        RECT 2255.625 211.600 2255.795 211.770 ;
        RECT 2256.085 211.600 2256.255 211.770 ;
        RECT 2256.545 211.600 2256.715 211.770 ;
        RECT 2257.005 211.600 2257.175 211.770 ;
        RECT 2257.465 211.600 2257.635 211.770 ;
        RECT 2257.925 211.600 2258.095 211.770 ;
        RECT 2258.385 211.600 2258.555 211.770 ;
        RECT 2258.845 211.600 2259.015 211.770 ;
        RECT 2259.305 211.600 2259.475 211.770 ;
        RECT 2259.765 211.600 2259.935 211.770 ;
        RECT 2260.225 211.600 2260.395 211.770 ;
        RECT 2260.685 211.600 2260.855 211.770 ;
        RECT 2261.145 211.600 2261.315 211.770 ;
        RECT 2261.605 211.600 2261.775 211.770 ;
        RECT 2262.065 211.600 2262.235 211.770 ;
        RECT 2262.525 211.600 2262.695 211.770 ;
        RECT 2262.985 211.600 2263.155 211.770 ;
        RECT 2263.445 211.600 2263.615 211.770 ;
        RECT 2263.905 211.600 2264.075 211.770 ;
        RECT 2264.365 211.600 2264.535 211.770 ;
        RECT 2264.825 211.600 2264.995 211.770 ;
        RECT 2265.285 211.600 2265.455 211.770 ;
        RECT 2265.745 211.600 2265.915 211.770 ;
        RECT 2266.205 211.600 2266.375 211.770 ;
        RECT 2266.665 211.600 2266.835 211.770 ;
        RECT 2267.125 211.600 2267.295 211.770 ;
        RECT 2267.585 211.600 2267.755 211.770 ;
        RECT 2268.045 211.600 2268.215 211.770 ;
        RECT 2268.505 211.600 2268.675 211.770 ;
        RECT 2268.965 211.600 2269.135 211.770 ;
        RECT 2269.425 211.600 2269.595 211.770 ;
        RECT 2269.885 211.600 2270.055 211.770 ;
        RECT 2270.345 211.600 2270.515 211.770 ;
        RECT 2270.805 211.600 2270.975 211.770 ;
        RECT 2271.265 211.600 2271.435 211.770 ;
        RECT 2271.725 211.600 2271.895 211.770 ;
      LAYER mcon ;
        RECT 2147.065 217.040 2147.235 217.210 ;
        RECT 2147.525 217.040 2147.695 217.210 ;
        RECT 2147.985 217.040 2148.155 217.210 ;
        RECT 2148.445 217.040 2148.615 217.210 ;
        RECT 2148.905 217.040 2149.075 217.210 ;
        RECT 2149.365 217.040 2149.535 217.210 ;
        RECT 2149.825 217.040 2149.995 217.210 ;
        RECT 2150.285 217.040 2150.455 217.210 ;
        RECT 2150.745 217.040 2150.915 217.210 ;
        RECT 2151.205 217.040 2151.375 217.210 ;
        RECT 2151.665 217.040 2151.835 217.210 ;
        RECT 2153.045 217.040 2153.215 217.210 ;
        RECT 2153.505 217.040 2153.675 217.210 ;
        RECT 2153.965 217.040 2154.135 217.210 ;
        RECT 2154.425 217.040 2154.595 217.210 ;
        RECT 2154.885 217.040 2155.055 217.210 ;
        RECT 2155.345 217.040 2155.515 217.210 ;
        RECT 2155.805 217.040 2155.975 217.210 ;
        RECT 2156.265 217.040 2156.435 217.210 ;
        RECT 2156.725 217.040 2156.895 217.210 ;
        RECT 2157.185 217.040 2157.355 217.210 ;
        RECT 2157.645 217.040 2157.815 217.210 ;
        RECT 2159.025 217.040 2159.195 217.210 ;
        RECT 2159.485 217.040 2159.655 217.210 ;
        RECT 2159.945 217.040 2160.115 217.210 ;
        RECT 2160.405 217.040 2160.575 217.210 ;
        RECT 2160.865 217.040 2161.035 217.210 ;
        RECT 2161.325 217.040 2161.495 217.210 ;
        RECT 2161.785 217.040 2161.955 217.210 ;
        RECT 2162.245 217.040 2162.415 217.210 ;
        RECT 2162.705 217.040 2162.875 217.210 ;
        RECT 2163.165 217.040 2163.335 217.210 ;
        RECT 2163.625 217.040 2163.795 217.210 ;
        RECT 2165.005 217.040 2165.175 217.210 ;
        RECT 2165.465 217.040 2165.635 217.210 ;
        RECT 2165.925 217.040 2166.095 217.210 ;
        RECT 2166.385 217.040 2166.555 217.210 ;
        RECT 2166.845 217.040 2167.015 217.210 ;
        RECT 2167.305 217.040 2167.475 217.210 ;
        RECT 2167.765 217.040 2167.935 217.210 ;
        RECT 2168.225 217.040 2168.395 217.210 ;
        RECT 2168.685 217.040 2168.855 217.210 ;
        RECT 2169.145 217.040 2169.315 217.210 ;
        RECT 2169.605 217.040 2169.775 217.210 ;
        RECT 2170.985 217.040 2171.155 217.210 ;
        RECT 2171.445 217.040 2171.615 217.210 ;
        RECT 2171.905 217.040 2172.075 217.210 ;
        RECT 2172.365 217.040 2172.535 217.210 ;
        RECT 2172.825 217.040 2172.995 217.210 ;
        RECT 2173.285 217.040 2173.455 217.210 ;
        RECT 2173.745 217.040 2173.915 217.210 ;
        RECT 2174.205 217.040 2174.375 217.210 ;
        RECT 2174.665 217.040 2174.835 217.210 ;
        RECT 2175.125 217.040 2175.295 217.210 ;
        RECT 2175.585 217.040 2175.755 217.210 ;
        RECT 2176.965 217.040 2177.135 217.210 ;
        RECT 2177.425 217.040 2177.595 217.210 ;
        RECT 2177.885 217.040 2178.055 217.210 ;
        RECT 2178.345 217.040 2178.515 217.210 ;
        RECT 2178.805 217.040 2178.975 217.210 ;
        RECT 2179.265 217.040 2179.435 217.210 ;
        RECT 2179.725 217.040 2179.895 217.210 ;
        RECT 2180.185 217.040 2180.355 217.210 ;
        RECT 2180.645 217.040 2180.815 217.210 ;
        RECT 2181.105 217.040 2181.275 217.210 ;
        RECT 2181.565 217.040 2181.735 217.210 ;
        RECT 2182.945 217.040 2183.115 217.210 ;
        RECT 2183.405 217.040 2183.575 217.210 ;
        RECT 2183.865 217.040 2184.035 217.210 ;
        RECT 2184.325 217.040 2184.495 217.210 ;
        RECT 2184.785 217.040 2184.955 217.210 ;
        RECT 2185.245 217.040 2185.415 217.210 ;
        RECT 2185.705 217.040 2185.875 217.210 ;
        RECT 2186.165 217.040 2186.335 217.210 ;
        RECT 2186.625 217.040 2186.795 217.210 ;
        RECT 2187.085 217.040 2187.255 217.210 ;
        RECT 2187.545 217.040 2187.715 217.210 ;
        RECT 2188.925 217.040 2189.095 217.210 ;
        RECT 2189.385 217.040 2189.555 217.210 ;
        RECT 2189.845 217.040 2190.015 217.210 ;
        RECT 2190.305 217.040 2190.475 217.210 ;
        RECT 2190.765 217.040 2190.935 217.210 ;
        RECT 2191.225 217.040 2191.395 217.210 ;
        RECT 2191.685 217.040 2191.855 217.210 ;
        RECT 2192.145 217.040 2192.315 217.210 ;
        RECT 2192.605 217.040 2192.775 217.210 ;
        RECT 2193.065 217.040 2193.235 217.210 ;
        RECT 2193.525 217.040 2193.695 217.210 ;
        RECT 2194.905 217.040 2195.075 217.210 ;
        RECT 2195.365 217.040 2195.535 217.210 ;
        RECT 2195.825 217.040 2195.995 217.210 ;
        RECT 2196.285 217.040 2196.455 217.210 ;
        RECT 2196.745 217.040 2196.915 217.210 ;
        RECT 2197.205 217.040 2197.375 217.210 ;
        RECT 2197.665 217.040 2197.835 217.210 ;
        RECT 2198.125 217.040 2198.295 217.210 ;
        RECT 2198.585 217.040 2198.755 217.210 ;
        RECT 2199.045 217.040 2199.215 217.210 ;
        RECT 2199.505 217.040 2199.675 217.210 ;
        RECT 2200.885 217.040 2201.055 217.210 ;
        RECT 2201.345 217.040 2201.515 217.210 ;
        RECT 2201.805 217.040 2201.975 217.210 ;
        RECT 2202.265 217.040 2202.435 217.210 ;
        RECT 2202.725 217.040 2202.895 217.210 ;
        RECT 2203.185 217.040 2203.355 217.210 ;
        RECT 2203.645 217.040 2203.815 217.210 ;
        RECT 2204.105 217.040 2204.275 217.210 ;
        RECT 2204.565 217.040 2204.735 217.210 ;
        RECT 2205.025 217.040 2205.195 217.210 ;
        RECT 2205.485 217.040 2205.655 217.210 ;
        RECT 2236.765 217.040 2236.935 217.210 ;
        RECT 2237.225 217.040 2237.395 217.210 ;
        RECT 2237.685 217.040 2237.855 217.210 ;
        RECT 2238.145 217.040 2238.315 217.210 ;
        RECT 2238.605 217.040 2238.775 217.210 ;
        RECT 2239.065 217.040 2239.235 217.210 ;
        RECT 2239.525 217.040 2239.695 217.210 ;
        RECT 2239.985 217.040 2240.155 217.210 ;
        RECT 2240.445 217.040 2240.615 217.210 ;
        RECT 2240.905 217.040 2241.075 217.210 ;
        RECT 2241.365 217.040 2241.535 217.210 ;
        RECT 2242.745 217.040 2242.915 217.210 ;
        RECT 2243.205 217.040 2243.375 217.210 ;
        RECT 2243.665 217.040 2243.835 217.210 ;
        RECT 2244.125 217.040 2244.295 217.210 ;
        RECT 2244.585 217.040 2244.755 217.210 ;
        RECT 2245.045 217.040 2245.215 217.210 ;
        RECT 2245.505 217.040 2245.675 217.210 ;
        RECT 2245.965 217.040 2246.135 217.210 ;
        RECT 2246.425 217.040 2246.595 217.210 ;
        RECT 2246.885 217.040 2247.055 217.210 ;
        RECT 2247.345 217.040 2247.515 217.210 ;
        RECT 2248.725 217.040 2248.895 217.210 ;
        RECT 2249.185 217.040 2249.355 217.210 ;
        RECT 2249.645 217.040 2249.815 217.210 ;
        RECT 2250.105 217.040 2250.275 217.210 ;
        RECT 2250.565 217.040 2250.735 217.210 ;
        RECT 2251.025 217.040 2251.195 217.210 ;
        RECT 2251.485 217.040 2251.655 217.210 ;
        RECT 2251.945 217.040 2252.115 217.210 ;
        RECT 2252.405 217.040 2252.575 217.210 ;
        RECT 2252.865 217.040 2253.035 217.210 ;
        RECT 2253.325 217.040 2253.495 217.210 ;
        RECT 2254.705 217.040 2254.875 217.210 ;
        RECT 2255.165 217.040 2255.335 217.210 ;
        RECT 2255.625 217.040 2255.795 217.210 ;
        RECT 2256.085 217.040 2256.255 217.210 ;
        RECT 2256.545 217.040 2256.715 217.210 ;
        RECT 2257.005 217.040 2257.175 217.210 ;
        RECT 2257.465 217.040 2257.635 217.210 ;
        RECT 2257.925 217.040 2258.095 217.210 ;
        RECT 2258.385 217.040 2258.555 217.210 ;
        RECT 2258.845 217.040 2259.015 217.210 ;
        RECT 2259.305 217.040 2259.475 217.210 ;
        RECT 2260.685 217.040 2260.855 217.210 ;
        RECT 2261.145 217.040 2261.315 217.210 ;
        RECT 2261.605 217.040 2261.775 217.210 ;
        RECT 2262.065 217.040 2262.235 217.210 ;
        RECT 2262.525 217.040 2262.695 217.210 ;
        RECT 2262.985 217.040 2263.155 217.210 ;
        RECT 2263.445 217.040 2263.615 217.210 ;
        RECT 2263.905 217.040 2264.075 217.210 ;
        RECT 2264.365 217.040 2264.535 217.210 ;
        RECT 2264.825 217.040 2264.995 217.210 ;
        RECT 2265.285 217.040 2265.455 217.210 ;
        RECT 2266.665 217.040 2266.835 217.210 ;
        RECT 2267.125 217.040 2267.295 217.210 ;
        RECT 2267.585 217.040 2267.755 217.210 ;
        RECT 2268.045 217.040 2268.215 217.210 ;
        RECT 2268.505 217.040 2268.675 217.210 ;
        RECT 2268.965 217.040 2269.135 217.210 ;
        RECT 2269.425 217.040 2269.595 217.210 ;
        RECT 2269.885 217.040 2270.055 217.210 ;
        RECT 2270.345 217.040 2270.515 217.210 ;
        RECT 2270.805 217.040 2270.975 217.210 ;
        RECT 2271.265 217.040 2271.435 217.210 ;
        RECT 2147.065 211.600 2147.235 211.770 ;
        RECT 2147.525 211.600 2147.695 211.770 ;
        RECT 2147.985 211.600 2148.155 211.770 ;
        RECT 2148.445 211.600 2148.615 211.770 ;
        RECT 2148.905 211.600 2149.075 211.770 ;
        RECT 2149.365 211.600 2149.535 211.770 ;
        RECT 2149.825 211.600 2149.995 211.770 ;
        RECT 2150.285 211.600 2150.455 211.770 ;
        RECT 2150.745 211.600 2150.915 211.770 ;
        RECT 2151.205 211.600 2151.375 211.770 ;
        RECT 2151.665 211.600 2151.835 211.770 ;
        RECT 2236.765 211.600 2236.935 211.770 ;
        RECT 2237.225 211.600 2237.395 211.770 ;
        RECT 2237.685 211.600 2237.855 211.770 ;
        RECT 2238.145 211.600 2238.315 211.770 ;
        RECT 2238.605 211.600 2238.775 211.770 ;
        RECT 2239.065 211.600 2239.235 211.770 ;
        RECT 2239.525 211.600 2239.695 211.770 ;
        RECT 2239.985 211.600 2240.155 211.770 ;
        RECT 2240.445 211.600 2240.615 211.770 ;
        RECT 2240.905 211.600 2241.075 211.770 ;
        RECT 2241.365 211.600 2241.535 211.770 ;
      LAYER met1 ;
        RECT 2146.000 216.885 2272.040 217.365 ;
        RECT 2146.000 211.445 2272.040 211.925 ;
      LAYER via ;
        RECT 2208.130 216.950 2209.915 217.250 ;
        RECT 2208.130 211.540 2209.915 211.840 ;
      LAYER met2 ;
        RECT 2208.090 216.880 2209.955 217.310 ;
        RECT 2208.090 211.455 2209.955 211.885 ;
      LAYER via2 ;
        RECT 2208.130 216.950 2209.915 217.250 ;
        RECT 2208.130 211.540 2209.915 211.840 ;
      LAYER met3 ;
        RECT 2208.095 209.800 2209.960 217.325 ;
    END
    PORT
      LAYER li1 ;
        RECT 201.995 1726.870 202.165 1727.040 ;
        RECT 207.435 1726.870 207.605 1727.040 ;
      LAYER li1 ;
        RECT 207.435 1726.640 207.605 1726.725 ;
        RECT 207.435 1726.580 208.150 1726.640 ;
      LAYER li1 ;
        RECT 201.995 1726.410 202.165 1726.580 ;
      LAYER li1 ;
        RECT 207.605 1726.410 208.150 1726.580 ;
      LAYER li1 ;
        RECT 201.995 1725.950 202.165 1726.120 ;
        RECT 201.995 1725.490 202.165 1725.660 ;
        RECT 201.995 1725.030 202.165 1725.200 ;
      LAYER li1 ;
        RECT 207.435 1725.055 208.150 1726.410 ;
      LAYER li1 ;
        RECT 201.995 1724.570 202.165 1724.740 ;
      LAYER li1 ;
        RECT 207.435 1724.715 208.980 1725.055 ;
      LAYER li1 ;
        RECT 201.995 1724.110 202.165 1724.280 ;
        RECT 201.995 1723.650 202.165 1723.820 ;
        RECT 201.995 1723.190 202.165 1723.360 ;
        RECT 201.995 1722.730 202.165 1722.900 ;
        RECT 201.995 1722.270 202.165 1722.440 ;
        RECT 201.995 1721.810 202.165 1721.980 ;
        RECT 201.995 1721.350 202.165 1721.520 ;
      LAYER li1 ;
        RECT 207.435 1721.295 208.150 1724.715 ;
        RECT 207.435 1721.205 207.605 1721.295 ;
      LAYER li1 ;
        RECT 201.995 1720.890 202.165 1721.060 ;
        RECT 207.435 1720.890 207.605 1721.060 ;
      LAYER li1 ;
        RECT 207.435 1720.660 207.605 1720.745 ;
        RECT 207.435 1720.600 208.150 1720.660 ;
      LAYER li1 ;
        RECT 201.995 1720.430 202.165 1720.600 ;
      LAYER li1 ;
        RECT 207.605 1720.430 208.150 1720.600 ;
      LAYER li1 ;
        RECT 201.995 1719.970 202.165 1720.140 ;
        RECT 201.995 1719.510 202.165 1719.680 ;
        RECT 201.995 1719.050 202.165 1719.220 ;
      LAYER li1 ;
        RECT 207.435 1719.075 208.150 1720.430 ;
      LAYER li1 ;
        RECT 201.995 1718.590 202.165 1718.760 ;
      LAYER li1 ;
        RECT 207.435 1718.735 208.980 1719.075 ;
      LAYER li1 ;
        RECT 201.995 1718.130 202.165 1718.300 ;
        RECT 201.995 1717.670 202.165 1717.840 ;
        RECT 201.995 1717.210 202.165 1717.380 ;
        RECT 201.995 1716.750 202.165 1716.920 ;
        RECT 201.995 1716.290 202.165 1716.460 ;
        RECT 201.995 1715.830 202.165 1716.000 ;
        RECT 201.995 1715.370 202.165 1715.540 ;
      LAYER li1 ;
        RECT 207.435 1715.315 208.150 1718.735 ;
        RECT 207.435 1715.225 207.605 1715.315 ;
      LAYER li1 ;
        RECT 201.995 1714.910 202.165 1715.080 ;
        RECT 207.435 1714.910 207.605 1715.080 ;
      LAYER li1 ;
        RECT 207.435 1714.680 207.605 1714.765 ;
        RECT 207.435 1714.620 208.150 1714.680 ;
      LAYER li1 ;
        RECT 201.995 1714.450 202.165 1714.620 ;
      LAYER li1 ;
        RECT 207.605 1714.450 208.150 1714.620 ;
      LAYER li1 ;
        RECT 201.995 1713.990 202.165 1714.160 ;
        RECT 201.995 1713.530 202.165 1713.700 ;
        RECT 201.995 1713.070 202.165 1713.240 ;
      LAYER li1 ;
        RECT 207.435 1713.095 208.150 1714.450 ;
      LAYER li1 ;
        RECT 201.995 1712.610 202.165 1712.780 ;
      LAYER li1 ;
        RECT 207.435 1712.755 208.980 1713.095 ;
      LAYER li1 ;
        RECT 201.995 1712.150 202.165 1712.320 ;
        RECT 201.995 1711.690 202.165 1711.860 ;
        RECT 201.995 1711.230 202.165 1711.400 ;
        RECT 201.995 1710.770 202.165 1710.940 ;
        RECT 201.995 1710.310 202.165 1710.480 ;
        RECT 201.995 1709.850 202.165 1710.020 ;
        RECT 201.995 1709.390 202.165 1709.560 ;
      LAYER li1 ;
        RECT 207.435 1709.335 208.150 1712.755 ;
        RECT 207.435 1709.245 207.605 1709.335 ;
      LAYER li1 ;
        RECT 201.995 1708.930 202.165 1709.100 ;
        RECT 207.435 1708.930 207.605 1709.100 ;
      LAYER li1 ;
        RECT 207.435 1708.700 207.605 1708.785 ;
        RECT 207.435 1708.640 208.150 1708.700 ;
      LAYER li1 ;
        RECT 201.995 1708.470 202.165 1708.640 ;
      LAYER li1 ;
        RECT 207.605 1708.470 208.150 1708.640 ;
      LAYER li1 ;
        RECT 201.995 1708.010 202.165 1708.180 ;
        RECT 201.995 1707.550 202.165 1707.720 ;
        RECT 201.995 1707.090 202.165 1707.260 ;
      LAYER li1 ;
        RECT 207.435 1707.115 208.150 1708.470 ;
      LAYER li1 ;
        RECT 201.995 1706.630 202.165 1706.800 ;
      LAYER li1 ;
        RECT 207.435 1706.775 208.980 1707.115 ;
      LAYER li1 ;
        RECT 201.995 1706.170 202.165 1706.340 ;
        RECT 201.995 1705.710 202.165 1705.880 ;
        RECT 201.995 1705.250 202.165 1705.420 ;
        RECT 201.995 1704.790 202.165 1704.960 ;
        RECT 201.995 1704.330 202.165 1704.500 ;
        RECT 201.995 1703.870 202.165 1704.040 ;
        RECT 201.995 1703.410 202.165 1703.580 ;
      LAYER li1 ;
        RECT 207.435 1703.355 208.150 1706.775 ;
        RECT 207.435 1703.265 207.605 1703.355 ;
      LAYER li1 ;
        RECT 201.995 1702.950 202.165 1703.120 ;
        RECT 207.435 1702.950 207.605 1703.120 ;
      LAYER li1 ;
        RECT 207.435 1702.720 207.605 1702.805 ;
        RECT 207.435 1702.660 208.150 1702.720 ;
      LAYER li1 ;
        RECT 201.995 1702.490 202.165 1702.660 ;
      LAYER li1 ;
        RECT 207.605 1702.490 208.150 1702.660 ;
      LAYER li1 ;
        RECT 201.995 1702.030 202.165 1702.200 ;
        RECT 201.995 1701.570 202.165 1701.740 ;
        RECT 201.995 1701.110 202.165 1701.280 ;
      LAYER li1 ;
        RECT 207.435 1701.135 208.150 1702.490 ;
      LAYER li1 ;
        RECT 201.995 1700.650 202.165 1700.820 ;
      LAYER li1 ;
        RECT 207.435 1700.795 208.980 1701.135 ;
      LAYER li1 ;
        RECT 201.995 1700.190 202.165 1700.360 ;
        RECT 201.995 1699.730 202.165 1699.900 ;
        RECT 201.995 1699.270 202.165 1699.440 ;
        RECT 201.995 1698.810 202.165 1698.980 ;
        RECT 201.995 1698.350 202.165 1698.520 ;
        RECT 201.995 1697.890 202.165 1698.060 ;
        RECT 201.995 1697.430 202.165 1697.600 ;
      LAYER li1 ;
        RECT 207.435 1697.375 208.150 1700.795 ;
        RECT 207.435 1697.285 207.605 1697.375 ;
      LAYER li1 ;
        RECT 201.995 1696.970 202.165 1697.140 ;
        RECT 207.435 1696.970 207.605 1697.140 ;
      LAYER li1 ;
        RECT 207.435 1696.740 207.605 1696.825 ;
        RECT 207.435 1696.680 208.150 1696.740 ;
      LAYER li1 ;
        RECT 201.995 1696.510 202.165 1696.680 ;
      LAYER li1 ;
        RECT 207.605 1696.510 208.150 1696.680 ;
      LAYER li1 ;
        RECT 201.995 1696.050 202.165 1696.220 ;
        RECT 201.995 1695.590 202.165 1695.760 ;
        RECT 201.995 1695.130 202.165 1695.300 ;
      LAYER li1 ;
        RECT 207.435 1695.155 208.150 1696.510 ;
      LAYER li1 ;
        RECT 201.995 1694.670 202.165 1694.840 ;
      LAYER li1 ;
        RECT 207.435 1694.815 208.980 1695.155 ;
      LAYER li1 ;
        RECT 201.995 1694.210 202.165 1694.380 ;
        RECT 201.995 1693.750 202.165 1693.920 ;
        RECT 201.995 1693.290 202.165 1693.460 ;
        RECT 201.995 1692.830 202.165 1693.000 ;
        RECT 201.995 1692.370 202.165 1692.540 ;
        RECT 201.995 1691.910 202.165 1692.080 ;
        RECT 201.995 1691.450 202.165 1691.620 ;
      LAYER li1 ;
        RECT 207.435 1691.395 208.150 1694.815 ;
        RECT 207.435 1691.305 207.605 1691.395 ;
      LAYER li1 ;
        RECT 201.995 1690.990 202.165 1691.160 ;
        RECT 207.435 1690.990 207.605 1691.160 ;
      LAYER li1 ;
        RECT 207.435 1690.760 207.605 1690.845 ;
        RECT 207.435 1690.700 208.150 1690.760 ;
      LAYER li1 ;
        RECT 201.995 1690.530 202.165 1690.700 ;
      LAYER li1 ;
        RECT 207.605 1690.530 208.150 1690.700 ;
      LAYER li1 ;
        RECT 201.995 1690.070 202.165 1690.240 ;
        RECT 201.995 1689.610 202.165 1689.780 ;
        RECT 201.995 1689.150 202.165 1689.320 ;
      LAYER li1 ;
        RECT 207.435 1689.175 208.150 1690.530 ;
      LAYER li1 ;
        RECT 201.995 1688.690 202.165 1688.860 ;
      LAYER li1 ;
        RECT 207.435 1688.835 208.980 1689.175 ;
      LAYER li1 ;
        RECT 201.995 1688.230 202.165 1688.400 ;
        RECT 201.995 1687.770 202.165 1687.940 ;
        RECT 201.995 1687.310 202.165 1687.480 ;
        RECT 201.995 1686.850 202.165 1687.020 ;
        RECT 201.995 1686.390 202.165 1686.560 ;
        RECT 201.995 1685.930 202.165 1686.100 ;
        RECT 201.995 1685.470 202.165 1685.640 ;
      LAYER li1 ;
        RECT 207.435 1685.415 208.150 1688.835 ;
        RECT 207.435 1685.325 207.605 1685.415 ;
      LAYER li1 ;
        RECT 201.995 1685.010 202.165 1685.180 ;
        RECT 207.435 1685.010 207.605 1685.180 ;
      LAYER li1 ;
        RECT 207.435 1684.780 207.605 1684.865 ;
        RECT 207.435 1684.720 208.150 1684.780 ;
      LAYER li1 ;
        RECT 201.995 1684.550 202.165 1684.720 ;
      LAYER li1 ;
        RECT 207.605 1684.550 208.150 1684.720 ;
      LAYER li1 ;
        RECT 201.995 1684.090 202.165 1684.260 ;
        RECT 201.995 1683.630 202.165 1683.800 ;
        RECT 201.995 1683.170 202.165 1683.340 ;
      LAYER li1 ;
        RECT 207.435 1683.195 208.150 1684.550 ;
      LAYER li1 ;
        RECT 201.995 1682.710 202.165 1682.880 ;
      LAYER li1 ;
        RECT 207.435 1682.855 208.980 1683.195 ;
      LAYER li1 ;
        RECT 201.995 1682.250 202.165 1682.420 ;
        RECT 201.995 1681.790 202.165 1681.960 ;
        RECT 201.995 1681.330 202.165 1681.500 ;
        RECT 201.995 1680.870 202.165 1681.040 ;
        RECT 201.995 1680.410 202.165 1680.580 ;
        RECT 201.995 1679.950 202.165 1680.120 ;
        RECT 201.995 1679.490 202.165 1679.660 ;
      LAYER li1 ;
        RECT 207.435 1679.435 208.150 1682.855 ;
        RECT 207.435 1679.345 207.605 1679.435 ;
      LAYER li1 ;
        RECT 201.995 1679.030 202.165 1679.200 ;
        RECT 207.435 1679.030 207.605 1679.200 ;
      LAYER li1 ;
        RECT 207.435 1678.800 207.605 1678.885 ;
        RECT 207.435 1678.740 208.150 1678.800 ;
      LAYER li1 ;
        RECT 201.995 1678.570 202.165 1678.740 ;
      LAYER li1 ;
        RECT 207.605 1678.570 208.150 1678.740 ;
      LAYER li1 ;
        RECT 201.995 1678.110 202.165 1678.280 ;
        RECT 201.995 1677.650 202.165 1677.820 ;
        RECT 201.995 1677.190 202.165 1677.360 ;
      LAYER li1 ;
        RECT 207.435 1677.215 208.150 1678.570 ;
      LAYER li1 ;
        RECT 201.995 1676.730 202.165 1676.900 ;
      LAYER li1 ;
        RECT 207.435 1676.875 208.980 1677.215 ;
      LAYER li1 ;
        RECT 201.995 1676.270 202.165 1676.440 ;
        RECT 201.995 1675.810 202.165 1675.980 ;
        RECT 201.995 1675.350 202.165 1675.520 ;
        RECT 201.995 1674.890 202.165 1675.060 ;
        RECT 201.995 1674.430 202.165 1674.600 ;
        RECT 201.995 1673.970 202.165 1674.140 ;
        RECT 201.995 1673.510 202.165 1673.680 ;
      LAYER li1 ;
        RECT 207.435 1673.455 208.150 1676.875 ;
        RECT 207.435 1673.365 207.605 1673.455 ;
      LAYER li1 ;
        RECT 201.995 1673.050 202.165 1673.220 ;
        RECT 207.435 1673.050 207.605 1673.220 ;
      LAYER mcon ;
        RECT 207.435 1725.950 207.605 1726.120 ;
        RECT 207.435 1725.490 207.605 1725.660 ;
        RECT 207.435 1725.030 207.605 1725.200 ;
        RECT 207.435 1724.570 207.605 1724.740 ;
        RECT 207.435 1724.110 207.605 1724.280 ;
        RECT 207.435 1723.650 207.605 1723.820 ;
        RECT 207.435 1723.190 207.605 1723.360 ;
        RECT 207.435 1722.730 207.605 1722.900 ;
        RECT 207.435 1722.270 207.605 1722.440 ;
        RECT 207.435 1721.810 207.605 1721.980 ;
        RECT 207.435 1721.350 207.605 1721.520 ;
        RECT 207.435 1719.970 207.605 1720.140 ;
        RECT 207.435 1719.510 207.605 1719.680 ;
        RECT 207.435 1719.050 207.605 1719.220 ;
        RECT 207.435 1718.590 207.605 1718.760 ;
        RECT 207.435 1718.130 207.605 1718.300 ;
        RECT 207.435 1717.670 207.605 1717.840 ;
        RECT 207.435 1717.210 207.605 1717.380 ;
        RECT 207.435 1716.750 207.605 1716.920 ;
        RECT 207.435 1716.290 207.605 1716.460 ;
        RECT 207.435 1715.830 207.605 1716.000 ;
        RECT 207.435 1715.370 207.605 1715.540 ;
        RECT 207.435 1713.990 207.605 1714.160 ;
        RECT 207.435 1713.530 207.605 1713.700 ;
        RECT 207.435 1713.070 207.605 1713.240 ;
        RECT 207.435 1712.610 207.605 1712.780 ;
        RECT 207.435 1712.150 207.605 1712.320 ;
        RECT 207.435 1711.690 207.605 1711.860 ;
        RECT 207.435 1711.230 207.605 1711.400 ;
        RECT 207.435 1710.770 207.605 1710.940 ;
        RECT 207.435 1710.310 207.605 1710.480 ;
        RECT 207.435 1709.850 207.605 1710.020 ;
        RECT 207.435 1709.390 207.605 1709.560 ;
        RECT 207.435 1708.010 207.605 1708.180 ;
        RECT 207.435 1707.550 207.605 1707.720 ;
        RECT 207.435 1707.090 207.605 1707.260 ;
        RECT 207.435 1706.630 207.605 1706.800 ;
        RECT 207.435 1706.170 207.605 1706.340 ;
        RECT 207.435 1705.710 207.605 1705.880 ;
        RECT 207.435 1705.250 207.605 1705.420 ;
        RECT 207.435 1704.790 207.605 1704.960 ;
        RECT 207.435 1704.330 207.605 1704.500 ;
        RECT 207.435 1703.870 207.605 1704.040 ;
        RECT 207.435 1703.410 207.605 1703.580 ;
        RECT 207.435 1702.030 207.605 1702.200 ;
        RECT 207.435 1701.570 207.605 1701.740 ;
        RECT 207.435 1701.110 207.605 1701.280 ;
        RECT 207.435 1700.650 207.605 1700.820 ;
        RECT 207.435 1700.190 207.605 1700.360 ;
        RECT 207.435 1699.730 207.605 1699.900 ;
        RECT 207.435 1699.270 207.605 1699.440 ;
        RECT 207.435 1698.810 207.605 1698.980 ;
        RECT 207.435 1698.350 207.605 1698.520 ;
        RECT 207.435 1697.890 207.605 1698.060 ;
        RECT 207.435 1697.430 207.605 1697.600 ;
        RECT 207.435 1696.050 207.605 1696.220 ;
        RECT 207.435 1695.590 207.605 1695.760 ;
        RECT 207.435 1695.130 207.605 1695.300 ;
        RECT 207.435 1694.670 207.605 1694.840 ;
        RECT 207.435 1694.210 207.605 1694.380 ;
        RECT 207.435 1693.750 207.605 1693.920 ;
        RECT 207.435 1693.290 207.605 1693.460 ;
        RECT 207.435 1692.830 207.605 1693.000 ;
        RECT 207.435 1692.370 207.605 1692.540 ;
        RECT 207.435 1691.910 207.605 1692.080 ;
        RECT 207.435 1691.450 207.605 1691.620 ;
        RECT 207.435 1690.070 207.605 1690.240 ;
        RECT 207.435 1689.610 207.605 1689.780 ;
        RECT 207.435 1689.150 207.605 1689.320 ;
        RECT 207.435 1688.690 207.605 1688.860 ;
        RECT 207.435 1688.230 207.605 1688.400 ;
        RECT 207.435 1687.770 207.605 1687.940 ;
        RECT 207.435 1687.310 207.605 1687.480 ;
        RECT 207.435 1686.850 207.605 1687.020 ;
        RECT 207.435 1686.390 207.605 1686.560 ;
        RECT 207.435 1685.930 207.605 1686.100 ;
        RECT 207.435 1685.470 207.605 1685.640 ;
        RECT 207.435 1684.090 207.605 1684.260 ;
        RECT 207.435 1683.630 207.605 1683.800 ;
        RECT 207.435 1683.170 207.605 1683.340 ;
        RECT 207.435 1682.710 207.605 1682.880 ;
        RECT 207.435 1682.250 207.605 1682.420 ;
        RECT 207.435 1681.790 207.605 1681.960 ;
        RECT 207.435 1681.330 207.605 1681.500 ;
        RECT 207.435 1680.870 207.605 1681.040 ;
        RECT 207.435 1680.410 207.605 1680.580 ;
        RECT 207.435 1679.950 207.605 1680.120 ;
        RECT 207.435 1679.490 207.605 1679.660 ;
        RECT 207.435 1678.110 207.605 1678.280 ;
        RECT 207.435 1677.650 207.605 1677.820 ;
        RECT 207.435 1677.190 207.605 1677.360 ;
        RECT 207.435 1676.730 207.605 1676.900 ;
        RECT 207.435 1676.270 207.605 1676.440 ;
        RECT 207.435 1675.810 207.605 1675.980 ;
        RECT 207.435 1675.350 207.605 1675.520 ;
        RECT 207.435 1674.890 207.605 1675.060 ;
        RECT 207.435 1674.430 207.605 1674.600 ;
        RECT 207.435 1673.970 207.605 1674.140 ;
        RECT 207.435 1673.510 207.605 1673.680 ;
      LAYER met1 ;
        RECT 201.840 1672.905 202.320 1736.740 ;
        RECT 207.280 1672.905 207.760 1736.700 ;
      LAYER via ;
        RECT 201.950 1734.795 202.250 1736.580 ;
        RECT 207.360 1734.795 207.660 1736.580 ;
      LAYER met2 ;
        RECT 201.865 1734.755 202.295 1736.620 ;
        RECT 207.290 1734.755 207.720 1736.620 ;
      LAYER via2 ;
        RECT 201.950 1734.795 202.250 1736.580 ;
        RECT 207.360 1734.795 207.660 1736.580 ;
      LAYER met3 ;
        RECT 200.210 1734.750 207.735 1736.615 ;
    END
    PORT
      LAYER li1 ;
        RECT 201.885 3014.775 202.055 3014.945 ;
        RECT 207.325 3014.775 207.495 3014.945 ;
        RECT 201.885 3014.315 202.055 3014.485 ;
        RECT 207.325 3014.315 207.495 3014.485 ;
        RECT 201.885 3013.855 202.055 3014.025 ;
        RECT 207.325 3013.855 207.495 3014.025 ;
        RECT 201.885 3013.395 202.055 3013.565 ;
        RECT 207.325 3013.395 207.495 3013.565 ;
        RECT 201.885 3012.935 202.055 3013.105 ;
        RECT 207.325 3012.935 207.495 3013.105 ;
        RECT 201.885 3012.475 202.055 3012.645 ;
        RECT 207.325 3012.475 207.495 3012.645 ;
        RECT 201.885 3012.015 202.055 3012.185 ;
        RECT 207.325 3012.015 207.495 3012.185 ;
        RECT 201.885 3011.555 202.055 3011.725 ;
        RECT 207.325 3011.555 207.495 3011.725 ;
        RECT 201.885 3011.095 202.055 3011.265 ;
        RECT 207.325 3011.095 207.495 3011.265 ;
        RECT 201.885 3010.635 202.055 3010.805 ;
        RECT 207.325 3010.635 207.495 3010.805 ;
        RECT 201.885 3010.175 202.055 3010.345 ;
        RECT 207.325 3010.175 207.495 3010.345 ;
        RECT 201.885 3009.715 202.055 3009.885 ;
        RECT 207.325 3009.715 207.495 3009.885 ;
        RECT 201.885 3009.255 202.055 3009.425 ;
        RECT 207.325 3009.255 207.495 3009.425 ;
        RECT 201.885 3008.795 202.055 3008.965 ;
        RECT 207.325 3008.795 207.495 3008.965 ;
        RECT 201.885 3008.335 202.055 3008.505 ;
        RECT 207.325 3008.335 207.495 3008.505 ;
        RECT 201.885 3007.875 202.055 3008.045 ;
        RECT 207.325 3007.875 207.495 3008.045 ;
        RECT 201.885 3007.415 202.055 3007.585 ;
        RECT 207.325 3007.415 207.495 3007.585 ;
        RECT 201.885 3006.955 202.055 3007.125 ;
        RECT 207.325 3006.955 207.495 3007.125 ;
        RECT 201.885 3006.495 202.055 3006.665 ;
        RECT 207.325 3006.495 207.495 3006.665 ;
        RECT 201.885 3006.035 202.055 3006.205 ;
        RECT 207.325 3006.035 207.495 3006.205 ;
        RECT 201.885 3005.575 202.055 3005.745 ;
        RECT 207.325 3005.575 207.495 3005.745 ;
        RECT 201.885 3005.115 202.055 3005.285 ;
        RECT 207.325 3005.115 207.495 3005.285 ;
        RECT 201.885 3004.655 202.055 3004.825 ;
        RECT 207.325 3004.655 207.495 3004.825 ;
        RECT 201.885 3004.195 202.055 3004.365 ;
        RECT 207.325 3004.195 207.495 3004.365 ;
        RECT 201.885 3003.735 202.055 3003.905 ;
        RECT 207.325 3003.735 207.495 3003.905 ;
        RECT 201.885 3003.275 202.055 3003.445 ;
        RECT 207.325 3003.275 207.495 3003.445 ;
        RECT 201.885 3002.815 202.055 3002.985 ;
        RECT 207.325 3002.815 207.495 3002.985 ;
        RECT 201.885 3002.355 202.055 3002.525 ;
        RECT 207.325 3002.355 207.495 3002.525 ;
        RECT 201.885 3001.895 202.055 3002.065 ;
        RECT 207.325 3001.895 207.495 3002.065 ;
        RECT 201.885 3001.435 202.055 3001.605 ;
        RECT 207.325 3001.435 207.495 3001.605 ;
        RECT 201.885 3000.975 202.055 3001.145 ;
        RECT 207.325 3000.975 207.495 3001.145 ;
        RECT 201.885 3000.515 202.055 3000.685 ;
        RECT 207.325 3000.515 207.495 3000.685 ;
        RECT 201.885 3000.055 202.055 3000.225 ;
        RECT 207.325 3000.055 207.495 3000.225 ;
        RECT 201.885 2999.595 202.055 2999.765 ;
        RECT 207.325 2999.595 207.495 2999.765 ;
        RECT 201.885 2999.135 202.055 2999.305 ;
        RECT 207.325 2999.135 207.495 2999.305 ;
        RECT 201.885 2998.675 202.055 2998.845 ;
        RECT 207.325 2998.675 207.495 2998.845 ;
        RECT 201.885 2998.215 202.055 2998.385 ;
        RECT 207.325 2998.215 207.495 2998.385 ;
        RECT 201.885 2997.755 202.055 2997.925 ;
        RECT 207.325 2997.755 207.495 2997.925 ;
        RECT 201.885 2997.295 202.055 2997.465 ;
        RECT 207.325 2997.295 207.495 2997.465 ;
        RECT 201.885 2996.835 202.055 2997.005 ;
        RECT 207.325 2996.835 207.495 2997.005 ;
        RECT 201.885 2996.375 202.055 2996.545 ;
        RECT 207.325 2996.375 207.495 2996.545 ;
        RECT 201.885 2995.915 202.055 2996.085 ;
        RECT 207.325 2995.915 207.495 2996.085 ;
        RECT 201.885 2995.455 202.055 2995.625 ;
        RECT 207.325 2995.455 207.495 2995.625 ;
        RECT 201.885 2994.995 202.055 2995.165 ;
        RECT 207.325 2994.995 207.495 2995.165 ;
        RECT 201.885 2994.535 202.055 2994.705 ;
        RECT 207.325 2994.535 207.495 2994.705 ;
        RECT 201.885 2994.075 202.055 2994.245 ;
        RECT 207.325 2994.075 207.495 2994.245 ;
        RECT 201.885 2993.615 202.055 2993.785 ;
        RECT 207.325 2993.615 207.495 2993.785 ;
        RECT 201.885 2993.155 202.055 2993.325 ;
        RECT 207.325 2993.155 207.495 2993.325 ;
        RECT 201.885 2992.695 202.055 2992.865 ;
        RECT 207.325 2992.695 207.495 2992.865 ;
        RECT 201.885 2992.235 202.055 2992.405 ;
        RECT 207.325 2992.235 207.495 2992.405 ;
        RECT 201.885 2991.775 202.055 2991.945 ;
        RECT 207.325 2991.775 207.495 2991.945 ;
        RECT 201.885 2991.315 202.055 2991.485 ;
        RECT 207.325 2991.315 207.495 2991.485 ;
        RECT 201.885 2990.855 202.055 2991.025 ;
        RECT 207.325 2990.855 207.495 2991.025 ;
        RECT 201.885 2990.395 202.055 2990.565 ;
        RECT 207.325 2990.395 207.495 2990.565 ;
        RECT 201.885 2989.935 202.055 2990.105 ;
        RECT 207.325 2989.935 207.495 2990.105 ;
        RECT 201.885 2989.475 202.055 2989.645 ;
        RECT 207.325 2989.475 207.495 2989.645 ;
        RECT 201.885 2989.015 202.055 2989.185 ;
        RECT 207.325 2989.015 207.495 2989.185 ;
        RECT 201.885 2988.555 202.055 2988.725 ;
        RECT 207.325 2988.555 207.495 2988.725 ;
        RECT 201.885 2988.095 202.055 2988.265 ;
        RECT 207.325 2988.095 207.495 2988.265 ;
        RECT 201.885 2987.635 202.055 2987.805 ;
        RECT 207.325 2987.635 207.495 2987.805 ;
        RECT 201.885 2987.175 202.055 2987.345 ;
        RECT 207.325 2987.175 207.495 2987.345 ;
        RECT 201.885 2986.715 202.055 2986.885 ;
        RECT 207.325 2986.715 207.495 2986.885 ;
        RECT 201.885 2986.255 202.055 2986.425 ;
        RECT 207.325 2986.255 207.495 2986.425 ;
        RECT 201.885 2985.795 202.055 2985.965 ;
        RECT 207.325 2985.795 207.495 2985.965 ;
        RECT 201.885 2985.335 202.055 2985.505 ;
        RECT 207.325 2985.335 207.495 2985.505 ;
        RECT 201.885 2984.875 202.055 2985.045 ;
        RECT 207.325 2984.875 207.495 2985.045 ;
      LAYER met1 ;
        RECT 201.730 2984.730 202.210 3024.940 ;
        RECT 207.170 2984.730 207.650 3024.940 ;
      LAYER via ;
        RECT 201.855 3023.050 202.155 3024.835 ;
        RECT 207.265 3023.050 207.565 3024.835 ;
      LAYER met2 ;
        RECT 201.770 3023.010 202.200 3024.875 ;
        RECT 207.195 3023.010 207.625 3024.875 ;
      LAYER via2 ;
        RECT 201.855 3023.050 202.155 3024.835 ;
        RECT 207.265 3023.050 207.565 3024.835 ;
      LAYER met3 ;
        RECT 200.115 3023.005 207.640 3024.870 ;
    END
  END vssd
  PIN vccd
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 3377.780 2238.065 3377.950 2238.235 ;
        RECT 3383.220 2238.065 3383.390 2238.235 ;
      LAYER li1 ;
        RECT 3377.780 2237.835 3377.950 2237.920 ;
        RECT 3377.780 2234.430 3378.385 2237.835 ;
      LAYER li1 ;
        RECT 3383.220 2237.605 3383.390 2237.775 ;
        RECT 3383.220 2237.145 3383.390 2237.315 ;
        RECT 3383.220 2236.685 3383.390 2236.855 ;
        RECT 3383.220 2236.225 3383.390 2236.395 ;
        RECT 3383.220 2235.765 3383.390 2235.935 ;
        RECT 3383.220 2235.305 3383.390 2235.475 ;
        RECT 3383.220 2234.845 3383.390 2235.015 ;
      LAYER li1 ;
        RECT 3377.780 2234.080 3379.635 2234.430 ;
      LAYER li1 ;
        RECT 3383.220 2234.385 3383.390 2234.555 ;
      LAYER li1 ;
        RECT 3377.780 2232.490 3378.385 2234.080 ;
      LAYER li1 ;
        RECT 3383.220 2233.925 3383.390 2234.095 ;
        RECT 3383.220 2233.465 3383.390 2233.635 ;
        RECT 3383.220 2233.005 3383.390 2233.175 ;
        RECT 3383.220 2232.545 3383.390 2232.715 ;
      LAYER li1 ;
        RECT 3377.780 2232.400 3377.950 2232.490 ;
      LAYER li1 ;
        RECT 3377.780 2232.085 3377.950 2232.255 ;
        RECT 3383.220 2232.085 3383.390 2232.255 ;
      LAYER li1 ;
        RECT 3377.780 2231.855 3377.950 2231.940 ;
        RECT 3377.780 2228.450 3378.385 2231.855 ;
      LAYER li1 ;
        RECT 3383.220 2231.625 3383.390 2231.795 ;
        RECT 3383.220 2231.165 3383.390 2231.335 ;
        RECT 3383.220 2230.705 3383.390 2230.875 ;
        RECT 3383.220 2230.245 3383.390 2230.415 ;
        RECT 3383.220 2229.785 3383.390 2229.955 ;
        RECT 3383.220 2229.325 3383.390 2229.495 ;
        RECT 3383.220 2228.865 3383.390 2229.035 ;
      LAYER li1 ;
        RECT 3377.780 2228.100 3379.635 2228.450 ;
      LAYER li1 ;
        RECT 3383.220 2228.405 3383.390 2228.575 ;
      LAYER li1 ;
        RECT 3377.780 2226.510 3378.385 2228.100 ;
      LAYER li1 ;
        RECT 3383.220 2227.945 3383.390 2228.115 ;
        RECT 3383.220 2227.485 3383.390 2227.655 ;
        RECT 3383.220 2227.025 3383.390 2227.195 ;
        RECT 3383.220 2226.565 3383.390 2226.735 ;
      LAYER li1 ;
        RECT 3377.780 2226.420 3377.950 2226.510 ;
      LAYER li1 ;
        RECT 3377.780 2226.105 3377.950 2226.275 ;
        RECT 3383.220 2226.105 3383.390 2226.275 ;
      LAYER li1 ;
        RECT 3377.780 2225.875 3377.950 2225.960 ;
        RECT 3377.780 2222.470 3378.385 2225.875 ;
      LAYER li1 ;
        RECT 3383.220 2225.645 3383.390 2225.815 ;
        RECT 3383.220 2225.185 3383.390 2225.355 ;
        RECT 3383.220 2224.725 3383.390 2224.895 ;
        RECT 3383.220 2224.265 3383.390 2224.435 ;
        RECT 3383.220 2223.805 3383.390 2223.975 ;
        RECT 3383.220 2223.345 3383.390 2223.515 ;
        RECT 3383.220 2222.885 3383.390 2223.055 ;
      LAYER li1 ;
        RECT 3377.780 2222.120 3379.635 2222.470 ;
      LAYER li1 ;
        RECT 3383.220 2222.425 3383.390 2222.595 ;
      LAYER li1 ;
        RECT 3377.780 2220.530 3378.385 2222.120 ;
      LAYER li1 ;
        RECT 3383.220 2221.965 3383.390 2222.135 ;
        RECT 3383.220 2221.505 3383.390 2221.675 ;
        RECT 3383.220 2221.045 3383.390 2221.215 ;
        RECT 3383.220 2220.585 3383.390 2220.755 ;
      LAYER li1 ;
        RECT 3377.780 2220.440 3377.950 2220.530 ;
      LAYER li1 ;
        RECT 3377.780 2220.125 3377.950 2220.295 ;
        RECT 3383.220 2220.125 3383.390 2220.295 ;
      LAYER li1 ;
        RECT 3377.780 2219.895 3377.950 2219.980 ;
        RECT 3377.780 2216.490 3378.385 2219.895 ;
      LAYER li1 ;
        RECT 3383.220 2219.665 3383.390 2219.835 ;
        RECT 3383.220 2219.205 3383.390 2219.375 ;
        RECT 3383.220 2218.745 3383.390 2218.915 ;
        RECT 3383.220 2218.285 3383.390 2218.455 ;
        RECT 3383.220 2217.825 3383.390 2217.995 ;
        RECT 3383.220 2217.365 3383.390 2217.535 ;
        RECT 3383.220 2216.905 3383.390 2217.075 ;
      LAYER li1 ;
        RECT 3377.780 2216.140 3379.635 2216.490 ;
      LAYER li1 ;
        RECT 3383.220 2216.445 3383.390 2216.615 ;
      LAYER li1 ;
        RECT 3377.780 2214.550 3378.385 2216.140 ;
      LAYER li1 ;
        RECT 3383.220 2215.985 3383.390 2216.155 ;
        RECT 3383.220 2215.525 3383.390 2215.695 ;
        RECT 3383.220 2215.065 3383.390 2215.235 ;
        RECT 3383.220 2214.605 3383.390 2214.775 ;
      LAYER li1 ;
        RECT 3377.780 2214.460 3377.950 2214.550 ;
      LAYER li1 ;
        RECT 3377.780 2214.145 3377.950 2214.315 ;
        RECT 3383.220 2214.145 3383.390 2214.315 ;
      LAYER li1 ;
        RECT 3377.780 2213.915 3377.950 2214.000 ;
        RECT 3377.780 2210.510 3378.385 2213.915 ;
      LAYER li1 ;
        RECT 3383.220 2213.685 3383.390 2213.855 ;
        RECT 3383.220 2213.225 3383.390 2213.395 ;
        RECT 3383.220 2212.765 3383.390 2212.935 ;
        RECT 3383.220 2212.305 3383.390 2212.475 ;
        RECT 3383.220 2211.845 3383.390 2212.015 ;
        RECT 3383.220 2211.385 3383.390 2211.555 ;
        RECT 3383.220 2210.925 3383.390 2211.095 ;
      LAYER li1 ;
        RECT 3377.780 2210.160 3379.635 2210.510 ;
      LAYER li1 ;
        RECT 3383.220 2210.465 3383.390 2210.635 ;
      LAYER li1 ;
        RECT 3377.780 2208.570 3378.385 2210.160 ;
      LAYER li1 ;
        RECT 3383.220 2210.005 3383.390 2210.175 ;
        RECT 3383.220 2209.545 3383.390 2209.715 ;
        RECT 3383.220 2209.085 3383.390 2209.255 ;
        RECT 3383.220 2208.625 3383.390 2208.795 ;
      LAYER li1 ;
        RECT 3377.780 2208.480 3377.950 2208.570 ;
      LAYER li1 ;
        RECT 3377.780 2208.165 3377.950 2208.335 ;
        RECT 3383.220 2208.165 3383.390 2208.335 ;
      LAYER li1 ;
        RECT 3377.780 2207.935 3377.950 2208.020 ;
        RECT 3377.780 2204.530 3378.385 2207.935 ;
      LAYER li1 ;
        RECT 3383.220 2207.705 3383.390 2207.875 ;
        RECT 3383.220 2207.245 3383.390 2207.415 ;
        RECT 3383.220 2206.785 3383.390 2206.955 ;
        RECT 3383.220 2206.325 3383.390 2206.495 ;
        RECT 3383.220 2205.865 3383.390 2206.035 ;
        RECT 3383.220 2205.405 3383.390 2205.575 ;
        RECT 3383.220 2204.945 3383.390 2205.115 ;
      LAYER li1 ;
        RECT 3377.780 2204.180 3379.635 2204.530 ;
      LAYER li1 ;
        RECT 3383.220 2204.485 3383.390 2204.655 ;
      LAYER li1 ;
        RECT 3377.780 2202.590 3378.385 2204.180 ;
      LAYER li1 ;
        RECT 3383.220 2204.025 3383.390 2204.195 ;
        RECT 3383.220 2203.565 3383.390 2203.735 ;
        RECT 3383.220 2203.105 3383.390 2203.275 ;
        RECT 3383.220 2202.645 3383.390 2202.815 ;
      LAYER li1 ;
        RECT 3377.780 2202.500 3377.950 2202.590 ;
      LAYER li1 ;
        RECT 3377.780 2202.185 3377.950 2202.355 ;
        RECT 3383.220 2202.185 3383.390 2202.355 ;
      LAYER li1 ;
        RECT 3377.780 2201.955 3377.950 2202.040 ;
        RECT 3377.780 2198.550 3378.385 2201.955 ;
      LAYER li1 ;
        RECT 3383.220 2201.725 3383.390 2201.895 ;
        RECT 3383.220 2201.265 3383.390 2201.435 ;
        RECT 3383.220 2200.805 3383.390 2200.975 ;
        RECT 3383.220 2200.345 3383.390 2200.515 ;
        RECT 3383.220 2199.885 3383.390 2200.055 ;
        RECT 3383.220 2199.425 3383.390 2199.595 ;
        RECT 3383.220 2198.965 3383.390 2199.135 ;
      LAYER li1 ;
        RECT 3377.780 2198.200 3379.635 2198.550 ;
      LAYER li1 ;
        RECT 3383.220 2198.505 3383.390 2198.675 ;
      LAYER li1 ;
        RECT 3377.780 2196.610 3378.385 2198.200 ;
      LAYER li1 ;
        RECT 3383.220 2198.045 3383.390 2198.215 ;
        RECT 3383.220 2197.585 3383.390 2197.755 ;
        RECT 3383.220 2197.125 3383.390 2197.295 ;
        RECT 3383.220 2196.665 3383.390 2196.835 ;
      LAYER li1 ;
        RECT 3377.780 2196.520 3377.950 2196.610 ;
      LAYER li1 ;
        RECT 3377.780 2196.205 3377.950 2196.375 ;
        RECT 3383.220 2196.205 3383.390 2196.375 ;
      LAYER mcon ;
        RECT 3377.780 2237.145 3377.950 2237.315 ;
        RECT 3377.780 2236.685 3377.950 2236.855 ;
        RECT 3377.780 2236.225 3377.950 2236.395 ;
        RECT 3377.780 2235.765 3377.950 2235.935 ;
        RECT 3377.780 2235.305 3377.950 2235.475 ;
        RECT 3377.780 2234.845 3377.950 2235.015 ;
        RECT 3377.780 2234.385 3377.950 2234.555 ;
        RECT 3377.780 2233.925 3377.950 2234.095 ;
        RECT 3377.780 2233.465 3377.950 2233.635 ;
        RECT 3377.780 2233.005 3377.950 2233.175 ;
        RECT 3377.780 2232.545 3377.950 2232.715 ;
        RECT 3377.780 2231.165 3377.950 2231.335 ;
        RECT 3377.780 2230.705 3377.950 2230.875 ;
        RECT 3377.780 2230.245 3377.950 2230.415 ;
        RECT 3377.780 2229.785 3377.950 2229.955 ;
        RECT 3377.780 2229.325 3377.950 2229.495 ;
        RECT 3377.780 2228.865 3377.950 2229.035 ;
        RECT 3377.780 2228.405 3377.950 2228.575 ;
        RECT 3377.780 2227.945 3377.950 2228.115 ;
        RECT 3377.780 2227.485 3377.950 2227.655 ;
        RECT 3377.780 2227.025 3377.950 2227.195 ;
        RECT 3377.780 2226.565 3377.950 2226.735 ;
        RECT 3377.780 2225.185 3377.950 2225.355 ;
        RECT 3377.780 2224.725 3377.950 2224.895 ;
        RECT 3377.780 2224.265 3377.950 2224.435 ;
        RECT 3377.780 2223.805 3377.950 2223.975 ;
        RECT 3377.780 2223.345 3377.950 2223.515 ;
        RECT 3377.780 2222.885 3377.950 2223.055 ;
        RECT 3377.780 2222.425 3377.950 2222.595 ;
        RECT 3377.780 2221.965 3377.950 2222.135 ;
        RECT 3377.780 2221.505 3377.950 2221.675 ;
        RECT 3377.780 2221.045 3377.950 2221.215 ;
        RECT 3377.780 2220.585 3377.950 2220.755 ;
        RECT 3377.780 2219.205 3377.950 2219.375 ;
        RECT 3377.780 2218.745 3377.950 2218.915 ;
        RECT 3377.780 2218.285 3377.950 2218.455 ;
        RECT 3377.780 2217.825 3377.950 2217.995 ;
        RECT 3377.780 2217.365 3377.950 2217.535 ;
        RECT 3377.780 2216.905 3377.950 2217.075 ;
        RECT 3377.780 2216.445 3377.950 2216.615 ;
        RECT 3377.780 2215.985 3377.950 2216.155 ;
        RECT 3377.780 2215.525 3377.950 2215.695 ;
        RECT 3377.780 2215.065 3377.950 2215.235 ;
        RECT 3377.780 2214.605 3377.950 2214.775 ;
        RECT 3377.780 2213.225 3377.950 2213.395 ;
        RECT 3377.780 2212.765 3377.950 2212.935 ;
        RECT 3377.780 2212.305 3377.950 2212.475 ;
        RECT 3377.780 2211.845 3377.950 2212.015 ;
        RECT 3377.780 2211.385 3377.950 2211.555 ;
        RECT 3377.780 2210.925 3377.950 2211.095 ;
        RECT 3377.780 2210.465 3377.950 2210.635 ;
        RECT 3377.780 2210.005 3377.950 2210.175 ;
        RECT 3377.780 2209.545 3377.950 2209.715 ;
        RECT 3377.780 2209.085 3377.950 2209.255 ;
        RECT 3377.780 2208.625 3377.950 2208.795 ;
        RECT 3377.780 2207.245 3377.950 2207.415 ;
        RECT 3377.780 2206.785 3377.950 2206.955 ;
        RECT 3377.780 2206.325 3377.950 2206.495 ;
        RECT 3377.780 2205.865 3377.950 2206.035 ;
        RECT 3377.780 2205.405 3377.950 2205.575 ;
        RECT 3377.780 2204.945 3377.950 2205.115 ;
        RECT 3377.780 2204.485 3377.950 2204.655 ;
        RECT 3377.780 2204.025 3377.950 2204.195 ;
        RECT 3377.780 2203.565 3377.950 2203.735 ;
        RECT 3377.780 2203.105 3377.950 2203.275 ;
        RECT 3377.780 2202.645 3377.950 2202.815 ;
        RECT 3377.780 2201.265 3377.950 2201.435 ;
        RECT 3377.780 2200.805 3377.950 2200.975 ;
        RECT 3377.780 2200.345 3377.950 2200.515 ;
        RECT 3377.780 2199.885 3377.950 2200.055 ;
        RECT 3377.780 2199.425 3377.950 2199.595 ;
        RECT 3377.780 2198.965 3377.950 2199.135 ;
        RECT 3377.780 2198.505 3377.950 2198.675 ;
        RECT 3377.780 2198.045 3377.950 2198.215 ;
        RECT 3377.780 2197.585 3377.950 2197.755 ;
        RECT 3377.780 2197.125 3377.950 2197.295 ;
        RECT 3377.780 2196.665 3377.950 2196.835 ;
      LAYER met1 ;
        RECT 3377.625 2196.060 3378.105 2238.380 ;
        RECT 3383.065 2196.060 3383.545 2238.380 ;
      LAYER via ;
        RECT 3377.690 2234.495 3377.990 2236.280 ;
        RECT 3383.130 2234.495 3383.430 2236.280 ;
      LAYER met2 ;
        RECT 3377.620 2234.455 3378.050 2236.320 ;
        RECT 3383.060 2234.455 3383.490 2236.320 ;
      LAYER via2 ;
        RECT 3377.690 2234.495 3377.990 2236.280 ;
        RECT 3383.130 2234.495 3383.430 2236.280 ;
      LAYER met3 ;
        RECT 3377.620 2234.465 3387.875 2236.315 ;
    END
    PORT
      LAYER li1 ;
        RECT 3377.780 3608.185 3377.950 3608.355 ;
        RECT 3383.220 3608.185 3383.390 3608.355 ;
      LAYER li1 ;
        RECT 3377.780 3607.955 3377.950 3608.040 ;
        RECT 3377.780 3604.550 3378.385 3607.955 ;
      LAYER li1 ;
        RECT 3383.220 3607.725 3383.390 3607.895 ;
        RECT 3383.220 3607.265 3383.390 3607.435 ;
        RECT 3383.220 3606.805 3383.390 3606.975 ;
        RECT 3383.220 3606.345 3383.390 3606.515 ;
        RECT 3383.220 3605.885 3383.390 3606.055 ;
        RECT 3383.220 3605.425 3383.390 3605.595 ;
        RECT 3383.220 3604.965 3383.390 3605.135 ;
      LAYER li1 ;
        RECT 3377.780 3604.200 3379.635 3604.550 ;
      LAYER li1 ;
        RECT 3383.220 3604.505 3383.390 3604.675 ;
      LAYER li1 ;
        RECT 3377.780 3602.610 3378.385 3604.200 ;
      LAYER li1 ;
        RECT 3383.220 3604.045 3383.390 3604.215 ;
        RECT 3383.220 3603.585 3383.390 3603.755 ;
        RECT 3383.220 3603.125 3383.390 3603.295 ;
        RECT 3383.220 3602.665 3383.390 3602.835 ;
      LAYER li1 ;
        RECT 3377.780 3602.520 3377.950 3602.610 ;
      LAYER li1 ;
        RECT 3377.780 3602.205 3377.950 3602.375 ;
        RECT 3383.220 3602.205 3383.390 3602.375 ;
      LAYER mcon ;
        RECT 3377.780 3607.265 3377.950 3607.435 ;
        RECT 3377.780 3606.805 3377.950 3606.975 ;
        RECT 3377.780 3606.345 3377.950 3606.515 ;
        RECT 3377.780 3605.885 3377.950 3606.055 ;
        RECT 3377.780 3605.425 3377.950 3605.595 ;
        RECT 3377.780 3604.965 3377.950 3605.135 ;
        RECT 3377.780 3604.505 3377.950 3604.675 ;
        RECT 3377.780 3604.045 3377.950 3604.215 ;
        RECT 3377.780 3603.585 3377.950 3603.755 ;
        RECT 3377.780 3603.125 3377.950 3603.295 ;
        RECT 3377.780 3602.665 3377.950 3602.835 ;
      LAYER met1 ;
        RECT 3377.625 3602.060 3378.105 3618.470 ;
        RECT 3383.065 3602.060 3383.545 3618.500 ;
      LAYER via ;
        RECT 3377.730 3616.500 3378.030 3618.285 ;
        RECT 3383.170 3616.500 3383.470 3618.285 ;
      LAYER met2 ;
        RECT 3377.660 3616.460 3378.090 3618.325 ;
        RECT 3383.100 3616.460 3383.530 3618.325 ;
      LAYER via2 ;
        RECT 3377.730 3616.500 3378.030 3618.285 ;
        RECT 3383.170 3616.500 3383.470 3618.285 ;
      LAYER met3 ;
        RECT 3377.660 3616.470 3387.915 3618.320 ;
    END
    PORT
      LAYER li1 ;
        RECT 669.145 219.760 669.315 219.930 ;
      LAYER li1 ;
        RECT 669.460 219.760 674.980 219.930 ;
      LAYER li1 ;
        RECT 675.125 219.760 675.295 219.930 ;
      LAYER li1 ;
        RECT 675.440 219.760 680.960 219.930 ;
      LAYER li1 ;
        RECT 681.105 219.760 681.275 219.930 ;
      LAYER li1 ;
        RECT 681.420 219.760 686.940 219.930 ;
      LAYER li1 ;
        RECT 687.085 219.760 687.255 219.930 ;
      LAYER li1 ;
        RECT 687.400 219.760 692.920 219.930 ;
      LAYER li1 ;
        RECT 693.065 219.760 693.235 219.930 ;
      LAYER li1 ;
        RECT 693.380 219.760 698.900 219.930 ;
      LAYER li1 ;
        RECT 699.045 219.760 699.215 219.930 ;
      LAYER li1 ;
        RECT 699.360 219.760 704.880 219.930 ;
      LAYER li1 ;
        RECT 705.025 219.760 705.195 219.930 ;
      LAYER li1 ;
        RECT 705.340 219.760 710.860 219.930 ;
      LAYER li1 ;
        RECT 711.005 219.760 711.175 219.930 ;
      LAYER li1 ;
        RECT 711.320 219.760 716.840 219.930 ;
      LAYER li1 ;
        RECT 716.985 219.760 717.155 219.930 ;
      LAYER li1 ;
        RECT 717.300 219.760 722.820 219.930 ;
      LAYER li1 ;
        RECT 722.965 219.760 723.135 219.930 ;
      LAYER li1 ;
        RECT 723.280 219.760 728.800 219.930 ;
      LAYER li1 ;
        RECT 728.945 219.760 729.115 219.930 ;
        RECT 758.845 219.760 759.015 219.930 ;
      LAYER li1 ;
        RECT 759.160 219.760 764.680 219.930 ;
      LAYER li1 ;
        RECT 764.825 219.760 764.995 219.930 ;
      LAYER li1 ;
        RECT 765.140 219.760 770.660 219.930 ;
      LAYER li1 ;
        RECT 770.805 219.760 770.975 219.930 ;
      LAYER li1 ;
        RECT 771.120 219.760 776.640 219.930 ;
      LAYER li1 ;
        RECT 776.785 219.760 776.955 219.930 ;
      LAYER li1 ;
        RECT 777.100 219.760 782.620 219.930 ;
      LAYER li1 ;
        RECT 782.765 219.760 782.935 219.930 ;
      LAYER li1 ;
        RECT 783.080 219.760 788.600 219.930 ;
      LAYER li1 ;
        RECT 788.745 219.760 788.915 219.930 ;
      LAYER li1 ;
        RECT 789.060 219.760 794.580 219.930 ;
      LAYER li1 ;
        RECT 794.725 219.760 794.895 219.930 ;
      LAYER li1 ;
        RECT 669.545 219.325 674.890 219.760 ;
        RECT 675.525 219.325 680.870 219.760 ;
        RECT 681.505 219.325 686.850 219.760 ;
        RECT 687.485 219.325 692.830 219.760 ;
        RECT 693.465 219.325 698.810 219.760 ;
        RECT 699.445 219.325 704.790 219.760 ;
        RECT 705.425 219.325 710.770 219.760 ;
        RECT 711.405 219.325 716.750 219.760 ;
        RECT 717.385 219.325 722.730 219.760 ;
        RECT 723.365 219.325 728.710 219.760 ;
        RECT 759.245 219.325 764.590 219.760 ;
        RECT 765.225 219.325 770.570 219.760 ;
        RECT 771.205 219.325 776.550 219.760 ;
        RECT 777.185 219.325 782.530 219.760 ;
        RECT 783.165 219.325 788.510 219.760 ;
        RECT 789.145 219.325 794.490 219.760 ;
        RECT 672.950 218.075 673.300 219.325 ;
        RECT 678.930 218.075 679.280 219.325 ;
        RECT 684.910 218.075 685.260 219.325 ;
        RECT 690.890 218.075 691.240 219.325 ;
        RECT 696.870 218.075 697.220 219.325 ;
        RECT 702.850 218.075 703.200 219.325 ;
        RECT 708.830 218.075 709.180 219.325 ;
        RECT 714.810 218.075 715.160 219.325 ;
        RECT 720.790 218.075 721.140 219.325 ;
        RECT 726.770 218.075 727.120 219.325 ;
        RECT 762.650 218.075 763.000 219.325 ;
        RECT 768.630 218.075 768.980 219.325 ;
        RECT 774.610 218.075 774.960 219.325 ;
        RECT 780.590 218.075 780.940 219.325 ;
        RECT 786.570 218.075 786.920 219.325 ;
        RECT 792.550 218.075 792.900 219.325 ;
      LAYER li1 ;
        RECT 669.145 214.320 669.315 214.490 ;
        RECT 669.605 214.320 669.775 214.490 ;
        RECT 670.065 214.320 670.235 214.490 ;
        RECT 670.525 214.320 670.695 214.490 ;
        RECT 670.985 214.320 671.155 214.490 ;
        RECT 671.445 214.320 671.615 214.490 ;
        RECT 671.905 214.320 672.075 214.490 ;
        RECT 672.365 214.320 672.535 214.490 ;
        RECT 672.825 214.320 672.995 214.490 ;
        RECT 673.285 214.320 673.455 214.490 ;
        RECT 673.745 214.320 673.915 214.490 ;
        RECT 674.205 214.320 674.375 214.490 ;
        RECT 674.665 214.320 674.835 214.490 ;
        RECT 675.125 214.320 675.295 214.490 ;
        RECT 675.585 214.320 675.755 214.490 ;
        RECT 676.045 214.320 676.215 214.490 ;
        RECT 676.505 214.320 676.675 214.490 ;
        RECT 676.965 214.320 677.135 214.490 ;
        RECT 677.425 214.320 677.595 214.490 ;
        RECT 677.885 214.320 678.055 214.490 ;
        RECT 678.345 214.320 678.515 214.490 ;
        RECT 678.805 214.320 678.975 214.490 ;
        RECT 679.265 214.320 679.435 214.490 ;
        RECT 679.725 214.320 679.895 214.490 ;
        RECT 680.185 214.320 680.355 214.490 ;
        RECT 680.645 214.320 680.815 214.490 ;
        RECT 681.105 214.320 681.275 214.490 ;
        RECT 681.565 214.320 681.735 214.490 ;
        RECT 682.025 214.320 682.195 214.490 ;
        RECT 682.485 214.320 682.655 214.490 ;
        RECT 682.945 214.320 683.115 214.490 ;
        RECT 683.405 214.320 683.575 214.490 ;
        RECT 683.865 214.320 684.035 214.490 ;
        RECT 684.325 214.320 684.495 214.490 ;
        RECT 684.785 214.320 684.955 214.490 ;
        RECT 685.245 214.320 685.415 214.490 ;
        RECT 685.705 214.320 685.875 214.490 ;
        RECT 686.165 214.320 686.335 214.490 ;
        RECT 686.625 214.320 686.795 214.490 ;
        RECT 687.085 214.320 687.255 214.490 ;
        RECT 687.545 214.320 687.715 214.490 ;
        RECT 688.005 214.320 688.175 214.490 ;
        RECT 688.465 214.320 688.635 214.490 ;
        RECT 688.925 214.320 689.095 214.490 ;
        RECT 689.385 214.320 689.555 214.490 ;
        RECT 689.845 214.320 690.015 214.490 ;
        RECT 690.305 214.320 690.475 214.490 ;
        RECT 690.765 214.320 690.935 214.490 ;
        RECT 691.225 214.320 691.395 214.490 ;
        RECT 691.685 214.320 691.855 214.490 ;
        RECT 692.145 214.320 692.315 214.490 ;
        RECT 692.605 214.320 692.775 214.490 ;
        RECT 693.065 214.320 693.235 214.490 ;
        RECT 693.525 214.320 693.695 214.490 ;
        RECT 693.985 214.320 694.155 214.490 ;
        RECT 694.445 214.320 694.615 214.490 ;
        RECT 694.905 214.320 695.075 214.490 ;
        RECT 695.365 214.320 695.535 214.490 ;
        RECT 695.825 214.320 695.995 214.490 ;
        RECT 696.285 214.320 696.455 214.490 ;
        RECT 696.745 214.320 696.915 214.490 ;
        RECT 697.205 214.320 697.375 214.490 ;
        RECT 697.665 214.320 697.835 214.490 ;
        RECT 698.125 214.320 698.295 214.490 ;
        RECT 698.585 214.320 698.755 214.490 ;
        RECT 699.045 214.320 699.215 214.490 ;
        RECT 699.505 214.320 699.675 214.490 ;
        RECT 699.965 214.320 700.135 214.490 ;
        RECT 700.425 214.320 700.595 214.490 ;
        RECT 700.885 214.320 701.055 214.490 ;
        RECT 701.345 214.320 701.515 214.490 ;
        RECT 701.805 214.320 701.975 214.490 ;
        RECT 702.265 214.320 702.435 214.490 ;
        RECT 702.725 214.320 702.895 214.490 ;
        RECT 703.185 214.320 703.355 214.490 ;
        RECT 703.645 214.320 703.815 214.490 ;
        RECT 704.105 214.320 704.275 214.490 ;
        RECT 704.565 214.320 704.735 214.490 ;
        RECT 705.025 214.320 705.195 214.490 ;
        RECT 705.485 214.320 705.655 214.490 ;
        RECT 705.945 214.320 706.115 214.490 ;
        RECT 706.405 214.320 706.575 214.490 ;
        RECT 706.865 214.320 707.035 214.490 ;
        RECT 707.325 214.320 707.495 214.490 ;
        RECT 707.785 214.320 707.955 214.490 ;
        RECT 708.245 214.320 708.415 214.490 ;
        RECT 708.705 214.320 708.875 214.490 ;
        RECT 709.165 214.320 709.335 214.490 ;
        RECT 709.625 214.320 709.795 214.490 ;
        RECT 710.085 214.320 710.255 214.490 ;
        RECT 710.545 214.320 710.715 214.490 ;
        RECT 711.005 214.320 711.175 214.490 ;
        RECT 711.465 214.320 711.635 214.490 ;
        RECT 711.925 214.320 712.095 214.490 ;
        RECT 712.385 214.320 712.555 214.490 ;
        RECT 712.845 214.320 713.015 214.490 ;
        RECT 713.305 214.320 713.475 214.490 ;
        RECT 713.765 214.320 713.935 214.490 ;
        RECT 714.225 214.320 714.395 214.490 ;
        RECT 714.685 214.320 714.855 214.490 ;
        RECT 715.145 214.320 715.315 214.490 ;
        RECT 715.605 214.320 715.775 214.490 ;
        RECT 716.065 214.320 716.235 214.490 ;
        RECT 716.525 214.320 716.695 214.490 ;
        RECT 716.985 214.320 717.155 214.490 ;
        RECT 717.445 214.320 717.615 214.490 ;
        RECT 717.905 214.320 718.075 214.490 ;
        RECT 718.365 214.320 718.535 214.490 ;
        RECT 718.825 214.320 718.995 214.490 ;
        RECT 719.285 214.320 719.455 214.490 ;
        RECT 719.745 214.320 719.915 214.490 ;
        RECT 720.205 214.320 720.375 214.490 ;
        RECT 720.665 214.320 720.835 214.490 ;
        RECT 721.125 214.320 721.295 214.490 ;
        RECT 721.585 214.320 721.755 214.490 ;
        RECT 722.045 214.320 722.215 214.490 ;
        RECT 722.505 214.320 722.675 214.490 ;
        RECT 722.965 214.320 723.135 214.490 ;
        RECT 723.425 214.320 723.595 214.490 ;
        RECT 723.885 214.320 724.055 214.490 ;
        RECT 724.345 214.320 724.515 214.490 ;
        RECT 724.805 214.320 724.975 214.490 ;
        RECT 725.265 214.320 725.435 214.490 ;
        RECT 725.725 214.320 725.895 214.490 ;
        RECT 726.185 214.320 726.355 214.490 ;
        RECT 726.645 214.320 726.815 214.490 ;
        RECT 727.105 214.320 727.275 214.490 ;
        RECT 727.565 214.320 727.735 214.490 ;
        RECT 728.025 214.320 728.195 214.490 ;
        RECT 728.485 214.320 728.655 214.490 ;
        RECT 728.945 214.320 729.115 214.490 ;
        RECT 758.845 214.320 759.015 214.490 ;
        RECT 759.305 214.320 759.475 214.490 ;
        RECT 759.765 214.320 759.935 214.490 ;
        RECT 760.225 214.320 760.395 214.490 ;
        RECT 760.685 214.320 760.855 214.490 ;
        RECT 761.145 214.320 761.315 214.490 ;
        RECT 761.605 214.320 761.775 214.490 ;
        RECT 762.065 214.320 762.235 214.490 ;
        RECT 762.525 214.320 762.695 214.490 ;
        RECT 762.985 214.320 763.155 214.490 ;
        RECT 763.445 214.320 763.615 214.490 ;
        RECT 763.905 214.320 764.075 214.490 ;
        RECT 764.365 214.320 764.535 214.490 ;
        RECT 764.825 214.320 764.995 214.490 ;
        RECT 765.285 214.320 765.455 214.490 ;
        RECT 765.745 214.320 765.915 214.490 ;
        RECT 766.205 214.320 766.375 214.490 ;
        RECT 766.665 214.320 766.835 214.490 ;
        RECT 767.125 214.320 767.295 214.490 ;
        RECT 767.585 214.320 767.755 214.490 ;
        RECT 768.045 214.320 768.215 214.490 ;
        RECT 768.505 214.320 768.675 214.490 ;
        RECT 768.965 214.320 769.135 214.490 ;
        RECT 769.425 214.320 769.595 214.490 ;
        RECT 769.885 214.320 770.055 214.490 ;
        RECT 770.345 214.320 770.515 214.490 ;
        RECT 770.805 214.320 770.975 214.490 ;
        RECT 771.265 214.320 771.435 214.490 ;
        RECT 771.725 214.320 771.895 214.490 ;
        RECT 772.185 214.320 772.355 214.490 ;
        RECT 772.645 214.320 772.815 214.490 ;
        RECT 773.105 214.320 773.275 214.490 ;
        RECT 773.565 214.320 773.735 214.490 ;
        RECT 774.025 214.320 774.195 214.490 ;
        RECT 774.485 214.320 774.655 214.490 ;
        RECT 774.945 214.320 775.115 214.490 ;
        RECT 775.405 214.320 775.575 214.490 ;
        RECT 775.865 214.320 776.035 214.490 ;
        RECT 776.325 214.320 776.495 214.490 ;
        RECT 776.785 214.320 776.955 214.490 ;
        RECT 777.245 214.320 777.415 214.490 ;
        RECT 777.705 214.320 777.875 214.490 ;
        RECT 778.165 214.320 778.335 214.490 ;
        RECT 778.625 214.320 778.795 214.490 ;
        RECT 779.085 214.320 779.255 214.490 ;
        RECT 779.545 214.320 779.715 214.490 ;
        RECT 780.005 214.320 780.175 214.490 ;
        RECT 780.465 214.320 780.635 214.490 ;
        RECT 780.925 214.320 781.095 214.490 ;
        RECT 781.385 214.320 781.555 214.490 ;
        RECT 781.845 214.320 782.015 214.490 ;
        RECT 782.305 214.320 782.475 214.490 ;
        RECT 782.765 214.320 782.935 214.490 ;
        RECT 783.225 214.320 783.395 214.490 ;
        RECT 783.685 214.320 783.855 214.490 ;
        RECT 784.145 214.320 784.315 214.490 ;
        RECT 784.605 214.320 784.775 214.490 ;
        RECT 785.065 214.320 785.235 214.490 ;
        RECT 785.525 214.320 785.695 214.490 ;
        RECT 785.985 214.320 786.155 214.490 ;
        RECT 786.445 214.320 786.615 214.490 ;
        RECT 786.905 214.320 787.075 214.490 ;
        RECT 787.365 214.320 787.535 214.490 ;
        RECT 787.825 214.320 787.995 214.490 ;
        RECT 788.285 214.320 788.455 214.490 ;
        RECT 788.745 214.320 788.915 214.490 ;
        RECT 789.205 214.320 789.375 214.490 ;
        RECT 789.665 214.320 789.835 214.490 ;
        RECT 790.125 214.320 790.295 214.490 ;
        RECT 790.585 214.320 790.755 214.490 ;
        RECT 791.045 214.320 791.215 214.490 ;
        RECT 791.505 214.320 791.675 214.490 ;
        RECT 791.965 214.320 792.135 214.490 ;
        RECT 792.425 214.320 792.595 214.490 ;
        RECT 792.885 214.320 793.055 214.490 ;
        RECT 793.345 214.320 793.515 214.490 ;
        RECT 793.805 214.320 793.975 214.490 ;
        RECT 794.265 214.320 794.435 214.490 ;
        RECT 794.725 214.320 794.895 214.490 ;
      LAYER mcon ;
        RECT 670.065 219.760 670.235 219.930 ;
        RECT 670.525 219.760 670.695 219.930 ;
        RECT 670.985 219.760 671.155 219.930 ;
        RECT 671.445 219.760 671.615 219.930 ;
        RECT 671.905 219.760 672.075 219.930 ;
        RECT 672.365 219.760 672.535 219.930 ;
        RECT 672.825 219.760 672.995 219.930 ;
        RECT 673.285 219.760 673.455 219.930 ;
        RECT 673.745 219.760 673.915 219.930 ;
        RECT 674.205 219.760 674.375 219.930 ;
        RECT 674.665 219.760 674.835 219.930 ;
        RECT 676.045 219.760 676.215 219.930 ;
        RECT 676.505 219.760 676.675 219.930 ;
        RECT 676.965 219.760 677.135 219.930 ;
        RECT 677.425 219.760 677.595 219.930 ;
        RECT 677.885 219.760 678.055 219.930 ;
        RECT 678.345 219.760 678.515 219.930 ;
        RECT 678.805 219.760 678.975 219.930 ;
        RECT 679.265 219.760 679.435 219.930 ;
        RECT 679.725 219.760 679.895 219.930 ;
        RECT 680.185 219.760 680.355 219.930 ;
        RECT 680.645 219.760 680.815 219.930 ;
        RECT 682.025 219.760 682.195 219.930 ;
        RECT 682.485 219.760 682.655 219.930 ;
        RECT 682.945 219.760 683.115 219.930 ;
        RECT 683.405 219.760 683.575 219.930 ;
        RECT 683.865 219.760 684.035 219.930 ;
        RECT 684.325 219.760 684.495 219.930 ;
        RECT 684.785 219.760 684.955 219.930 ;
        RECT 685.245 219.760 685.415 219.930 ;
        RECT 685.705 219.760 685.875 219.930 ;
        RECT 686.165 219.760 686.335 219.930 ;
        RECT 686.625 219.760 686.795 219.930 ;
        RECT 688.005 219.760 688.175 219.930 ;
        RECT 688.465 219.760 688.635 219.930 ;
        RECT 688.925 219.760 689.095 219.930 ;
        RECT 689.385 219.760 689.555 219.930 ;
        RECT 689.845 219.760 690.015 219.930 ;
        RECT 690.305 219.760 690.475 219.930 ;
        RECT 690.765 219.760 690.935 219.930 ;
        RECT 691.225 219.760 691.395 219.930 ;
        RECT 691.685 219.760 691.855 219.930 ;
        RECT 692.145 219.760 692.315 219.930 ;
        RECT 692.605 219.760 692.775 219.930 ;
        RECT 693.985 219.760 694.155 219.930 ;
        RECT 694.445 219.760 694.615 219.930 ;
        RECT 694.905 219.760 695.075 219.930 ;
        RECT 695.365 219.760 695.535 219.930 ;
        RECT 695.825 219.760 695.995 219.930 ;
        RECT 696.285 219.760 696.455 219.930 ;
        RECT 696.745 219.760 696.915 219.930 ;
        RECT 697.205 219.760 697.375 219.930 ;
        RECT 697.665 219.760 697.835 219.930 ;
        RECT 698.125 219.760 698.295 219.930 ;
        RECT 698.585 219.760 698.755 219.930 ;
        RECT 699.965 219.760 700.135 219.930 ;
        RECT 700.425 219.760 700.595 219.930 ;
        RECT 700.885 219.760 701.055 219.930 ;
        RECT 701.345 219.760 701.515 219.930 ;
        RECT 701.805 219.760 701.975 219.930 ;
        RECT 702.265 219.760 702.435 219.930 ;
        RECT 702.725 219.760 702.895 219.930 ;
        RECT 703.185 219.760 703.355 219.930 ;
        RECT 703.645 219.760 703.815 219.930 ;
        RECT 704.105 219.760 704.275 219.930 ;
        RECT 704.565 219.760 704.735 219.930 ;
        RECT 705.945 219.760 706.115 219.930 ;
        RECT 706.405 219.760 706.575 219.930 ;
        RECT 706.865 219.760 707.035 219.930 ;
        RECT 707.325 219.760 707.495 219.930 ;
        RECT 707.785 219.760 707.955 219.930 ;
        RECT 708.245 219.760 708.415 219.930 ;
        RECT 708.705 219.760 708.875 219.930 ;
        RECT 709.165 219.760 709.335 219.930 ;
        RECT 709.625 219.760 709.795 219.930 ;
        RECT 710.085 219.760 710.255 219.930 ;
        RECT 710.545 219.760 710.715 219.930 ;
        RECT 711.925 219.760 712.095 219.930 ;
        RECT 712.385 219.760 712.555 219.930 ;
        RECT 712.845 219.760 713.015 219.930 ;
        RECT 713.305 219.760 713.475 219.930 ;
        RECT 713.765 219.760 713.935 219.930 ;
        RECT 714.225 219.760 714.395 219.930 ;
        RECT 714.685 219.760 714.855 219.930 ;
        RECT 715.145 219.760 715.315 219.930 ;
        RECT 715.605 219.760 715.775 219.930 ;
        RECT 716.065 219.760 716.235 219.930 ;
        RECT 716.525 219.760 716.695 219.930 ;
        RECT 717.905 219.760 718.075 219.930 ;
        RECT 718.365 219.760 718.535 219.930 ;
        RECT 718.825 219.760 718.995 219.930 ;
        RECT 719.285 219.760 719.455 219.930 ;
        RECT 719.745 219.760 719.915 219.930 ;
        RECT 720.205 219.760 720.375 219.930 ;
        RECT 720.665 219.760 720.835 219.930 ;
        RECT 721.125 219.760 721.295 219.930 ;
        RECT 721.585 219.760 721.755 219.930 ;
        RECT 722.045 219.760 722.215 219.930 ;
        RECT 722.505 219.760 722.675 219.930 ;
        RECT 723.885 219.760 724.055 219.930 ;
        RECT 724.345 219.760 724.515 219.930 ;
        RECT 724.805 219.760 724.975 219.930 ;
        RECT 725.265 219.760 725.435 219.930 ;
        RECT 725.725 219.760 725.895 219.930 ;
        RECT 726.185 219.760 726.355 219.930 ;
        RECT 726.645 219.760 726.815 219.930 ;
        RECT 727.105 219.760 727.275 219.930 ;
        RECT 727.565 219.760 727.735 219.930 ;
        RECT 728.025 219.760 728.195 219.930 ;
        RECT 728.485 219.760 728.655 219.930 ;
        RECT 759.765 219.760 759.935 219.930 ;
        RECT 760.225 219.760 760.395 219.930 ;
        RECT 760.685 219.760 760.855 219.930 ;
        RECT 761.145 219.760 761.315 219.930 ;
        RECT 761.605 219.760 761.775 219.930 ;
        RECT 762.065 219.760 762.235 219.930 ;
        RECT 762.525 219.760 762.695 219.930 ;
        RECT 762.985 219.760 763.155 219.930 ;
        RECT 763.445 219.760 763.615 219.930 ;
        RECT 763.905 219.760 764.075 219.930 ;
        RECT 764.365 219.760 764.535 219.930 ;
        RECT 765.745 219.760 765.915 219.930 ;
        RECT 766.205 219.760 766.375 219.930 ;
        RECT 766.665 219.760 766.835 219.930 ;
        RECT 767.125 219.760 767.295 219.930 ;
        RECT 767.585 219.760 767.755 219.930 ;
        RECT 768.045 219.760 768.215 219.930 ;
        RECT 768.505 219.760 768.675 219.930 ;
        RECT 768.965 219.760 769.135 219.930 ;
        RECT 769.425 219.760 769.595 219.930 ;
        RECT 769.885 219.760 770.055 219.930 ;
        RECT 770.345 219.760 770.515 219.930 ;
        RECT 771.725 219.760 771.895 219.930 ;
        RECT 772.185 219.760 772.355 219.930 ;
        RECT 772.645 219.760 772.815 219.930 ;
        RECT 773.105 219.760 773.275 219.930 ;
        RECT 773.565 219.760 773.735 219.930 ;
        RECT 774.025 219.760 774.195 219.930 ;
        RECT 774.485 219.760 774.655 219.930 ;
        RECT 774.945 219.760 775.115 219.930 ;
        RECT 775.405 219.760 775.575 219.930 ;
        RECT 775.865 219.760 776.035 219.930 ;
        RECT 776.325 219.760 776.495 219.930 ;
        RECT 777.705 219.760 777.875 219.930 ;
        RECT 778.165 219.760 778.335 219.930 ;
        RECT 778.625 219.760 778.795 219.930 ;
        RECT 779.085 219.760 779.255 219.930 ;
        RECT 779.545 219.760 779.715 219.930 ;
        RECT 780.005 219.760 780.175 219.930 ;
        RECT 780.465 219.760 780.635 219.930 ;
        RECT 780.925 219.760 781.095 219.930 ;
        RECT 781.385 219.760 781.555 219.930 ;
        RECT 781.845 219.760 782.015 219.930 ;
        RECT 782.305 219.760 782.475 219.930 ;
        RECT 783.685 219.760 783.855 219.930 ;
        RECT 784.145 219.760 784.315 219.930 ;
        RECT 784.605 219.760 784.775 219.930 ;
        RECT 785.065 219.760 785.235 219.930 ;
        RECT 785.525 219.760 785.695 219.930 ;
        RECT 785.985 219.760 786.155 219.930 ;
        RECT 786.445 219.760 786.615 219.930 ;
        RECT 786.905 219.760 787.075 219.930 ;
        RECT 787.365 219.760 787.535 219.930 ;
        RECT 787.825 219.760 787.995 219.930 ;
        RECT 788.285 219.760 788.455 219.930 ;
        RECT 789.665 219.760 789.835 219.930 ;
        RECT 790.125 219.760 790.295 219.930 ;
        RECT 790.585 219.760 790.755 219.930 ;
        RECT 791.045 219.760 791.215 219.930 ;
        RECT 791.505 219.760 791.675 219.930 ;
        RECT 791.965 219.760 792.135 219.930 ;
        RECT 792.425 219.760 792.595 219.930 ;
        RECT 792.885 219.760 793.055 219.930 ;
        RECT 793.345 219.760 793.515 219.930 ;
        RECT 793.805 219.760 793.975 219.930 ;
        RECT 794.265 219.760 794.435 219.930 ;
      LAYER met1 ;
        RECT 669.000 219.605 795.040 220.085 ;
        RECT 669.000 214.165 795.040 214.645 ;
      LAYER via ;
        RECT 730.995 219.720 732.780 220.020 ;
        RECT 730.995 214.280 732.780 214.580 ;
      LAYER met2 ;
        RECT 730.955 219.660 732.820 220.090 ;
        RECT 730.955 214.220 732.820 214.650 ;
      LAYER via2 ;
        RECT 730.995 219.720 732.780 220.020 ;
        RECT 730.995 214.280 732.780 214.580 ;
      LAYER met3 ;
        RECT 730.965 209.835 732.815 220.090 ;
    END
    PORT
      LAYER li1 ;
        RECT 2146.145 219.760 2146.315 219.930 ;
      LAYER li1 ;
        RECT 2146.460 219.760 2151.980 219.930 ;
      LAYER li1 ;
        RECT 2152.125 219.760 2152.295 219.930 ;
      LAYER li1 ;
        RECT 2152.440 219.760 2157.960 219.930 ;
      LAYER li1 ;
        RECT 2158.105 219.760 2158.275 219.930 ;
      LAYER li1 ;
        RECT 2158.420 219.760 2163.940 219.930 ;
      LAYER li1 ;
        RECT 2164.085 219.760 2164.255 219.930 ;
      LAYER li1 ;
        RECT 2164.400 219.760 2169.920 219.930 ;
      LAYER li1 ;
        RECT 2170.065 219.760 2170.235 219.930 ;
      LAYER li1 ;
        RECT 2170.380 219.760 2175.900 219.930 ;
      LAYER li1 ;
        RECT 2176.045 219.760 2176.215 219.930 ;
      LAYER li1 ;
        RECT 2176.360 219.760 2181.880 219.930 ;
      LAYER li1 ;
        RECT 2182.025 219.760 2182.195 219.930 ;
      LAYER li1 ;
        RECT 2182.340 219.760 2187.860 219.930 ;
      LAYER li1 ;
        RECT 2188.005 219.760 2188.175 219.930 ;
      LAYER li1 ;
        RECT 2188.320 219.760 2193.840 219.930 ;
      LAYER li1 ;
        RECT 2193.985 219.760 2194.155 219.930 ;
      LAYER li1 ;
        RECT 2194.300 219.760 2199.820 219.930 ;
      LAYER li1 ;
        RECT 2199.965 219.760 2200.135 219.930 ;
      LAYER li1 ;
        RECT 2200.280 219.760 2205.800 219.930 ;
      LAYER li1 ;
        RECT 2205.945 219.760 2206.115 219.930 ;
        RECT 2235.845 219.760 2236.015 219.930 ;
      LAYER li1 ;
        RECT 2236.160 219.760 2241.680 219.930 ;
      LAYER li1 ;
        RECT 2241.825 219.760 2241.995 219.930 ;
      LAYER li1 ;
        RECT 2242.140 219.760 2247.660 219.930 ;
      LAYER li1 ;
        RECT 2247.805 219.760 2247.975 219.930 ;
      LAYER li1 ;
        RECT 2248.120 219.760 2253.640 219.930 ;
      LAYER li1 ;
        RECT 2253.785 219.760 2253.955 219.930 ;
      LAYER li1 ;
        RECT 2254.100 219.760 2259.620 219.930 ;
      LAYER li1 ;
        RECT 2259.765 219.760 2259.935 219.930 ;
      LAYER li1 ;
        RECT 2260.080 219.760 2265.600 219.930 ;
      LAYER li1 ;
        RECT 2265.745 219.760 2265.915 219.930 ;
      LAYER li1 ;
        RECT 2266.060 219.760 2271.580 219.930 ;
      LAYER li1 ;
        RECT 2271.725 219.760 2271.895 219.930 ;
      LAYER li1 ;
        RECT 2146.545 219.325 2151.890 219.760 ;
        RECT 2152.525 219.325 2157.870 219.760 ;
        RECT 2158.505 219.325 2163.850 219.760 ;
        RECT 2164.485 219.325 2169.830 219.760 ;
        RECT 2170.465 219.325 2175.810 219.760 ;
        RECT 2176.445 219.325 2181.790 219.760 ;
        RECT 2182.425 219.325 2187.770 219.760 ;
        RECT 2188.405 219.325 2193.750 219.760 ;
        RECT 2194.385 219.325 2199.730 219.760 ;
        RECT 2200.365 219.325 2205.710 219.760 ;
        RECT 2236.245 219.325 2241.590 219.760 ;
        RECT 2242.225 219.325 2247.570 219.760 ;
        RECT 2248.205 219.325 2253.550 219.760 ;
        RECT 2254.185 219.325 2259.530 219.760 ;
        RECT 2260.165 219.325 2265.510 219.760 ;
        RECT 2266.145 219.325 2271.490 219.760 ;
        RECT 2149.950 218.075 2150.300 219.325 ;
        RECT 2155.930 218.075 2156.280 219.325 ;
        RECT 2161.910 218.075 2162.260 219.325 ;
        RECT 2167.890 218.075 2168.240 219.325 ;
        RECT 2173.870 218.075 2174.220 219.325 ;
        RECT 2179.850 218.075 2180.200 219.325 ;
        RECT 2185.830 218.075 2186.180 219.325 ;
        RECT 2191.810 218.075 2192.160 219.325 ;
        RECT 2197.790 218.075 2198.140 219.325 ;
        RECT 2203.770 218.075 2204.120 219.325 ;
        RECT 2239.650 218.075 2240.000 219.325 ;
        RECT 2245.630 218.075 2245.980 219.325 ;
        RECT 2251.610 218.075 2251.960 219.325 ;
        RECT 2257.590 218.075 2257.940 219.325 ;
        RECT 2263.570 218.075 2263.920 219.325 ;
        RECT 2269.550 218.075 2269.900 219.325 ;
      LAYER li1 ;
        RECT 2146.145 214.320 2146.315 214.490 ;
        RECT 2146.605 214.320 2146.775 214.490 ;
        RECT 2147.065 214.320 2147.235 214.490 ;
        RECT 2147.525 214.320 2147.695 214.490 ;
        RECT 2147.985 214.320 2148.155 214.490 ;
        RECT 2148.445 214.320 2148.615 214.490 ;
        RECT 2148.905 214.320 2149.075 214.490 ;
        RECT 2149.365 214.320 2149.535 214.490 ;
        RECT 2149.825 214.320 2149.995 214.490 ;
        RECT 2150.285 214.320 2150.455 214.490 ;
        RECT 2150.745 214.320 2150.915 214.490 ;
        RECT 2151.205 214.320 2151.375 214.490 ;
        RECT 2151.665 214.320 2151.835 214.490 ;
        RECT 2152.125 214.320 2152.295 214.490 ;
        RECT 2152.585 214.320 2152.755 214.490 ;
        RECT 2153.045 214.320 2153.215 214.490 ;
        RECT 2153.505 214.320 2153.675 214.490 ;
        RECT 2153.965 214.320 2154.135 214.490 ;
        RECT 2154.425 214.320 2154.595 214.490 ;
        RECT 2154.885 214.320 2155.055 214.490 ;
        RECT 2155.345 214.320 2155.515 214.490 ;
        RECT 2155.805 214.320 2155.975 214.490 ;
        RECT 2156.265 214.320 2156.435 214.490 ;
        RECT 2156.725 214.320 2156.895 214.490 ;
        RECT 2157.185 214.320 2157.355 214.490 ;
        RECT 2157.645 214.320 2157.815 214.490 ;
        RECT 2158.105 214.320 2158.275 214.490 ;
        RECT 2158.565 214.320 2158.735 214.490 ;
        RECT 2159.025 214.320 2159.195 214.490 ;
        RECT 2159.485 214.320 2159.655 214.490 ;
        RECT 2159.945 214.320 2160.115 214.490 ;
        RECT 2160.405 214.320 2160.575 214.490 ;
        RECT 2160.865 214.320 2161.035 214.490 ;
        RECT 2161.325 214.320 2161.495 214.490 ;
        RECT 2161.785 214.320 2161.955 214.490 ;
        RECT 2162.245 214.320 2162.415 214.490 ;
        RECT 2162.705 214.320 2162.875 214.490 ;
        RECT 2163.165 214.320 2163.335 214.490 ;
        RECT 2163.625 214.320 2163.795 214.490 ;
        RECT 2164.085 214.320 2164.255 214.490 ;
        RECT 2164.545 214.320 2164.715 214.490 ;
        RECT 2165.005 214.320 2165.175 214.490 ;
        RECT 2165.465 214.320 2165.635 214.490 ;
        RECT 2165.925 214.320 2166.095 214.490 ;
        RECT 2166.385 214.320 2166.555 214.490 ;
        RECT 2166.845 214.320 2167.015 214.490 ;
        RECT 2167.305 214.320 2167.475 214.490 ;
        RECT 2167.765 214.320 2167.935 214.490 ;
        RECT 2168.225 214.320 2168.395 214.490 ;
        RECT 2168.685 214.320 2168.855 214.490 ;
        RECT 2169.145 214.320 2169.315 214.490 ;
        RECT 2169.605 214.320 2169.775 214.490 ;
        RECT 2170.065 214.320 2170.235 214.490 ;
        RECT 2170.525 214.320 2170.695 214.490 ;
        RECT 2170.985 214.320 2171.155 214.490 ;
        RECT 2171.445 214.320 2171.615 214.490 ;
        RECT 2171.905 214.320 2172.075 214.490 ;
        RECT 2172.365 214.320 2172.535 214.490 ;
        RECT 2172.825 214.320 2172.995 214.490 ;
        RECT 2173.285 214.320 2173.455 214.490 ;
        RECT 2173.745 214.320 2173.915 214.490 ;
        RECT 2174.205 214.320 2174.375 214.490 ;
        RECT 2174.665 214.320 2174.835 214.490 ;
        RECT 2175.125 214.320 2175.295 214.490 ;
        RECT 2175.585 214.320 2175.755 214.490 ;
        RECT 2176.045 214.320 2176.215 214.490 ;
        RECT 2176.505 214.320 2176.675 214.490 ;
        RECT 2176.965 214.320 2177.135 214.490 ;
        RECT 2177.425 214.320 2177.595 214.490 ;
        RECT 2177.885 214.320 2178.055 214.490 ;
        RECT 2178.345 214.320 2178.515 214.490 ;
        RECT 2178.805 214.320 2178.975 214.490 ;
        RECT 2179.265 214.320 2179.435 214.490 ;
        RECT 2179.725 214.320 2179.895 214.490 ;
        RECT 2180.185 214.320 2180.355 214.490 ;
        RECT 2180.645 214.320 2180.815 214.490 ;
        RECT 2181.105 214.320 2181.275 214.490 ;
        RECT 2181.565 214.320 2181.735 214.490 ;
        RECT 2182.025 214.320 2182.195 214.490 ;
        RECT 2182.485 214.320 2182.655 214.490 ;
        RECT 2182.945 214.320 2183.115 214.490 ;
        RECT 2183.405 214.320 2183.575 214.490 ;
        RECT 2183.865 214.320 2184.035 214.490 ;
        RECT 2184.325 214.320 2184.495 214.490 ;
        RECT 2184.785 214.320 2184.955 214.490 ;
        RECT 2185.245 214.320 2185.415 214.490 ;
        RECT 2185.705 214.320 2185.875 214.490 ;
        RECT 2186.165 214.320 2186.335 214.490 ;
        RECT 2186.625 214.320 2186.795 214.490 ;
        RECT 2187.085 214.320 2187.255 214.490 ;
        RECT 2187.545 214.320 2187.715 214.490 ;
        RECT 2188.005 214.320 2188.175 214.490 ;
        RECT 2188.465 214.320 2188.635 214.490 ;
        RECT 2188.925 214.320 2189.095 214.490 ;
        RECT 2189.385 214.320 2189.555 214.490 ;
        RECT 2189.845 214.320 2190.015 214.490 ;
        RECT 2190.305 214.320 2190.475 214.490 ;
        RECT 2190.765 214.320 2190.935 214.490 ;
        RECT 2191.225 214.320 2191.395 214.490 ;
        RECT 2191.685 214.320 2191.855 214.490 ;
        RECT 2192.145 214.320 2192.315 214.490 ;
        RECT 2192.605 214.320 2192.775 214.490 ;
        RECT 2193.065 214.320 2193.235 214.490 ;
        RECT 2193.525 214.320 2193.695 214.490 ;
        RECT 2193.985 214.320 2194.155 214.490 ;
        RECT 2194.445 214.320 2194.615 214.490 ;
        RECT 2194.905 214.320 2195.075 214.490 ;
        RECT 2195.365 214.320 2195.535 214.490 ;
        RECT 2195.825 214.320 2195.995 214.490 ;
        RECT 2196.285 214.320 2196.455 214.490 ;
        RECT 2196.745 214.320 2196.915 214.490 ;
        RECT 2197.205 214.320 2197.375 214.490 ;
        RECT 2197.665 214.320 2197.835 214.490 ;
        RECT 2198.125 214.320 2198.295 214.490 ;
        RECT 2198.585 214.320 2198.755 214.490 ;
        RECT 2199.045 214.320 2199.215 214.490 ;
        RECT 2199.505 214.320 2199.675 214.490 ;
        RECT 2199.965 214.320 2200.135 214.490 ;
        RECT 2200.425 214.320 2200.595 214.490 ;
        RECT 2200.885 214.320 2201.055 214.490 ;
        RECT 2201.345 214.320 2201.515 214.490 ;
        RECT 2201.805 214.320 2201.975 214.490 ;
        RECT 2202.265 214.320 2202.435 214.490 ;
        RECT 2202.725 214.320 2202.895 214.490 ;
        RECT 2203.185 214.320 2203.355 214.490 ;
        RECT 2203.645 214.320 2203.815 214.490 ;
        RECT 2204.105 214.320 2204.275 214.490 ;
        RECT 2204.565 214.320 2204.735 214.490 ;
        RECT 2205.025 214.320 2205.195 214.490 ;
        RECT 2205.485 214.320 2205.655 214.490 ;
        RECT 2205.945 214.320 2206.115 214.490 ;
        RECT 2235.845 214.320 2236.015 214.490 ;
        RECT 2236.305 214.320 2236.475 214.490 ;
        RECT 2236.765 214.320 2236.935 214.490 ;
        RECT 2237.225 214.320 2237.395 214.490 ;
        RECT 2237.685 214.320 2237.855 214.490 ;
        RECT 2238.145 214.320 2238.315 214.490 ;
        RECT 2238.605 214.320 2238.775 214.490 ;
        RECT 2239.065 214.320 2239.235 214.490 ;
        RECT 2239.525 214.320 2239.695 214.490 ;
        RECT 2239.985 214.320 2240.155 214.490 ;
        RECT 2240.445 214.320 2240.615 214.490 ;
        RECT 2240.905 214.320 2241.075 214.490 ;
        RECT 2241.365 214.320 2241.535 214.490 ;
        RECT 2241.825 214.320 2241.995 214.490 ;
        RECT 2242.285 214.320 2242.455 214.490 ;
        RECT 2242.745 214.320 2242.915 214.490 ;
        RECT 2243.205 214.320 2243.375 214.490 ;
        RECT 2243.665 214.320 2243.835 214.490 ;
        RECT 2244.125 214.320 2244.295 214.490 ;
        RECT 2244.585 214.320 2244.755 214.490 ;
        RECT 2245.045 214.320 2245.215 214.490 ;
        RECT 2245.505 214.320 2245.675 214.490 ;
        RECT 2245.965 214.320 2246.135 214.490 ;
        RECT 2246.425 214.320 2246.595 214.490 ;
        RECT 2246.885 214.320 2247.055 214.490 ;
        RECT 2247.345 214.320 2247.515 214.490 ;
        RECT 2247.805 214.320 2247.975 214.490 ;
        RECT 2248.265 214.320 2248.435 214.490 ;
        RECT 2248.725 214.320 2248.895 214.490 ;
        RECT 2249.185 214.320 2249.355 214.490 ;
        RECT 2249.645 214.320 2249.815 214.490 ;
        RECT 2250.105 214.320 2250.275 214.490 ;
        RECT 2250.565 214.320 2250.735 214.490 ;
        RECT 2251.025 214.320 2251.195 214.490 ;
        RECT 2251.485 214.320 2251.655 214.490 ;
        RECT 2251.945 214.320 2252.115 214.490 ;
        RECT 2252.405 214.320 2252.575 214.490 ;
        RECT 2252.865 214.320 2253.035 214.490 ;
        RECT 2253.325 214.320 2253.495 214.490 ;
        RECT 2253.785 214.320 2253.955 214.490 ;
        RECT 2254.245 214.320 2254.415 214.490 ;
        RECT 2254.705 214.320 2254.875 214.490 ;
        RECT 2255.165 214.320 2255.335 214.490 ;
        RECT 2255.625 214.320 2255.795 214.490 ;
        RECT 2256.085 214.320 2256.255 214.490 ;
        RECT 2256.545 214.320 2256.715 214.490 ;
        RECT 2257.005 214.320 2257.175 214.490 ;
        RECT 2257.465 214.320 2257.635 214.490 ;
        RECT 2257.925 214.320 2258.095 214.490 ;
        RECT 2258.385 214.320 2258.555 214.490 ;
        RECT 2258.845 214.320 2259.015 214.490 ;
        RECT 2259.305 214.320 2259.475 214.490 ;
        RECT 2259.765 214.320 2259.935 214.490 ;
        RECT 2260.225 214.320 2260.395 214.490 ;
        RECT 2260.685 214.320 2260.855 214.490 ;
        RECT 2261.145 214.320 2261.315 214.490 ;
        RECT 2261.605 214.320 2261.775 214.490 ;
        RECT 2262.065 214.320 2262.235 214.490 ;
        RECT 2262.525 214.320 2262.695 214.490 ;
        RECT 2262.985 214.320 2263.155 214.490 ;
        RECT 2263.445 214.320 2263.615 214.490 ;
        RECT 2263.905 214.320 2264.075 214.490 ;
        RECT 2264.365 214.320 2264.535 214.490 ;
        RECT 2264.825 214.320 2264.995 214.490 ;
        RECT 2265.285 214.320 2265.455 214.490 ;
        RECT 2265.745 214.320 2265.915 214.490 ;
        RECT 2266.205 214.320 2266.375 214.490 ;
        RECT 2266.665 214.320 2266.835 214.490 ;
        RECT 2267.125 214.320 2267.295 214.490 ;
        RECT 2267.585 214.320 2267.755 214.490 ;
        RECT 2268.045 214.320 2268.215 214.490 ;
        RECT 2268.505 214.320 2268.675 214.490 ;
        RECT 2268.965 214.320 2269.135 214.490 ;
        RECT 2269.425 214.320 2269.595 214.490 ;
        RECT 2269.885 214.320 2270.055 214.490 ;
        RECT 2270.345 214.320 2270.515 214.490 ;
        RECT 2270.805 214.320 2270.975 214.490 ;
        RECT 2271.265 214.320 2271.435 214.490 ;
        RECT 2271.725 214.320 2271.895 214.490 ;
      LAYER mcon ;
        RECT 2147.065 219.760 2147.235 219.930 ;
        RECT 2147.525 219.760 2147.695 219.930 ;
        RECT 2147.985 219.760 2148.155 219.930 ;
        RECT 2148.445 219.760 2148.615 219.930 ;
        RECT 2148.905 219.760 2149.075 219.930 ;
        RECT 2149.365 219.760 2149.535 219.930 ;
        RECT 2149.825 219.760 2149.995 219.930 ;
        RECT 2150.285 219.760 2150.455 219.930 ;
        RECT 2150.745 219.760 2150.915 219.930 ;
        RECT 2151.205 219.760 2151.375 219.930 ;
        RECT 2151.665 219.760 2151.835 219.930 ;
        RECT 2153.045 219.760 2153.215 219.930 ;
        RECT 2153.505 219.760 2153.675 219.930 ;
        RECT 2153.965 219.760 2154.135 219.930 ;
        RECT 2154.425 219.760 2154.595 219.930 ;
        RECT 2154.885 219.760 2155.055 219.930 ;
        RECT 2155.345 219.760 2155.515 219.930 ;
        RECT 2155.805 219.760 2155.975 219.930 ;
        RECT 2156.265 219.760 2156.435 219.930 ;
        RECT 2156.725 219.760 2156.895 219.930 ;
        RECT 2157.185 219.760 2157.355 219.930 ;
        RECT 2157.645 219.760 2157.815 219.930 ;
        RECT 2159.025 219.760 2159.195 219.930 ;
        RECT 2159.485 219.760 2159.655 219.930 ;
        RECT 2159.945 219.760 2160.115 219.930 ;
        RECT 2160.405 219.760 2160.575 219.930 ;
        RECT 2160.865 219.760 2161.035 219.930 ;
        RECT 2161.325 219.760 2161.495 219.930 ;
        RECT 2161.785 219.760 2161.955 219.930 ;
        RECT 2162.245 219.760 2162.415 219.930 ;
        RECT 2162.705 219.760 2162.875 219.930 ;
        RECT 2163.165 219.760 2163.335 219.930 ;
        RECT 2163.625 219.760 2163.795 219.930 ;
        RECT 2165.005 219.760 2165.175 219.930 ;
        RECT 2165.465 219.760 2165.635 219.930 ;
        RECT 2165.925 219.760 2166.095 219.930 ;
        RECT 2166.385 219.760 2166.555 219.930 ;
        RECT 2166.845 219.760 2167.015 219.930 ;
        RECT 2167.305 219.760 2167.475 219.930 ;
        RECT 2167.765 219.760 2167.935 219.930 ;
        RECT 2168.225 219.760 2168.395 219.930 ;
        RECT 2168.685 219.760 2168.855 219.930 ;
        RECT 2169.145 219.760 2169.315 219.930 ;
        RECT 2169.605 219.760 2169.775 219.930 ;
        RECT 2170.985 219.760 2171.155 219.930 ;
        RECT 2171.445 219.760 2171.615 219.930 ;
        RECT 2171.905 219.760 2172.075 219.930 ;
        RECT 2172.365 219.760 2172.535 219.930 ;
        RECT 2172.825 219.760 2172.995 219.930 ;
        RECT 2173.285 219.760 2173.455 219.930 ;
        RECT 2173.745 219.760 2173.915 219.930 ;
        RECT 2174.205 219.760 2174.375 219.930 ;
        RECT 2174.665 219.760 2174.835 219.930 ;
        RECT 2175.125 219.760 2175.295 219.930 ;
        RECT 2175.585 219.760 2175.755 219.930 ;
        RECT 2176.965 219.760 2177.135 219.930 ;
        RECT 2177.425 219.760 2177.595 219.930 ;
        RECT 2177.885 219.760 2178.055 219.930 ;
        RECT 2178.345 219.760 2178.515 219.930 ;
        RECT 2178.805 219.760 2178.975 219.930 ;
        RECT 2179.265 219.760 2179.435 219.930 ;
        RECT 2179.725 219.760 2179.895 219.930 ;
        RECT 2180.185 219.760 2180.355 219.930 ;
        RECT 2180.645 219.760 2180.815 219.930 ;
        RECT 2181.105 219.760 2181.275 219.930 ;
        RECT 2181.565 219.760 2181.735 219.930 ;
        RECT 2182.945 219.760 2183.115 219.930 ;
        RECT 2183.405 219.760 2183.575 219.930 ;
        RECT 2183.865 219.760 2184.035 219.930 ;
        RECT 2184.325 219.760 2184.495 219.930 ;
        RECT 2184.785 219.760 2184.955 219.930 ;
        RECT 2185.245 219.760 2185.415 219.930 ;
        RECT 2185.705 219.760 2185.875 219.930 ;
        RECT 2186.165 219.760 2186.335 219.930 ;
        RECT 2186.625 219.760 2186.795 219.930 ;
        RECT 2187.085 219.760 2187.255 219.930 ;
        RECT 2187.545 219.760 2187.715 219.930 ;
        RECT 2188.925 219.760 2189.095 219.930 ;
        RECT 2189.385 219.760 2189.555 219.930 ;
        RECT 2189.845 219.760 2190.015 219.930 ;
        RECT 2190.305 219.760 2190.475 219.930 ;
        RECT 2190.765 219.760 2190.935 219.930 ;
        RECT 2191.225 219.760 2191.395 219.930 ;
        RECT 2191.685 219.760 2191.855 219.930 ;
        RECT 2192.145 219.760 2192.315 219.930 ;
        RECT 2192.605 219.760 2192.775 219.930 ;
        RECT 2193.065 219.760 2193.235 219.930 ;
        RECT 2193.525 219.760 2193.695 219.930 ;
        RECT 2194.905 219.760 2195.075 219.930 ;
        RECT 2195.365 219.760 2195.535 219.930 ;
        RECT 2195.825 219.760 2195.995 219.930 ;
        RECT 2196.285 219.760 2196.455 219.930 ;
        RECT 2196.745 219.760 2196.915 219.930 ;
        RECT 2197.205 219.760 2197.375 219.930 ;
        RECT 2197.665 219.760 2197.835 219.930 ;
        RECT 2198.125 219.760 2198.295 219.930 ;
        RECT 2198.585 219.760 2198.755 219.930 ;
        RECT 2199.045 219.760 2199.215 219.930 ;
        RECT 2199.505 219.760 2199.675 219.930 ;
        RECT 2200.885 219.760 2201.055 219.930 ;
        RECT 2201.345 219.760 2201.515 219.930 ;
        RECT 2201.805 219.760 2201.975 219.930 ;
        RECT 2202.265 219.760 2202.435 219.930 ;
        RECT 2202.725 219.760 2202.895 219.930 ;
        RECT 2203.185 219.760 2203.355 219.930 ;
        RECT 2203.645 219.760 2203.815 219.930 ;
        RECT 2204.105 219.760 2204.275 219.930 ;
        RECT 2204.565 219.760 2204.735 219.930 ;
        RECT 2205.025 219.760 2205.195 219.930 ;
        RECT 2205.485 219.760 2205.655 219.930 ;
        RECT 2236.765 219.760 2236.935 219.930 ;
        RECT 2237.225 219.760 2237.395 219.930 ;
        RECT 2237.685 219.760 2237.855 219.930 ;
        RECT 2238.145 219.760 2238.315 219.930 ;
        RECT 2238.605 219.760 2238.775 219.930 ;
        RECT 2239.065 219.760 2239.235 219.930 ;
        RECT 2239.525 219.760 2239.695 219.930 ;
        RECT 2239.985 219.760 2240.155 219.930 ;
        RECT 2240.445 219.760 2240.615 219.930 ;
        RECT 2240.905 219.760 2241.075 219.930 ;
        RECT 2241.365 219.760 2241.535 219.930 ;
        RECT 2242.745 219.760 2242.915 219.930 ;
        RECT 2243.205 219.760 2243.375 219.930 ;
        RECT 2243.665 219.760 2243.835 219.930 ;
        RECT 2244.125 219.760 2244.295 219.930 ;
        RECT 2244.585 219.760 2244.755 219.930 ;
        RECT 2245.045 219.760 2245.215 219.930 ;
        RECT 2245.505 219.760 2245.675 219.930 ;
        RECT 2245.965 219.760 2246.135 219.930 ;
        RECT 2246.425 219.760 2246.595 219.930 ;
        RECT 2246.885 219.760 2247.055 219.930 ;
        RECT 2247.345 219.760 2247.515 219.930 ;
        RECT 2248.725 219.760 2248.895 219.930 ;
        RECT 2249.185 219.760 2249.355 219.930 ;
        RECT 2249.645 219.760 2249.815 219.930 ;
        RECT 2250.105 219.760 2250.275 219.930 ;
        RECT 2250.565 219.760 2250.735 219.930 ;
        RECT 2251.025 219.760 2251.195 219.930 ;
        RECT 2251.485 219.760 2251.655 219.930 ;
        RECT 2251.945 219.760 2252.115 219.930 ;
        RECT 2252.405 219.760 2252.575 219.930 ;
        RECT 2252.865 219.760 2253.035 219.930 ;
        RECT 2253.325 219.760 2253.495 219.930 ;
        RECT 2254.705 219.760 2254.875 219.930 ;
        RECT 2255.165 219.760 2255.335 219.930 ;
        RECT 2255.625 219.760 2255.795 219.930 ;
        RECT 2256.085 219.760 2256.255 219.930 ;
        RECT 2256.545 219.760 2256.715 219.930 ;
        RECT 2257.005 219.760 2257.175 219.930 ;
        RECT 2257.465 219.760 2257.635 219.930 ;
        RECT 2257.925 219.760 2258.095 219.930 ;
        RECT 2258.385 219.760 2258.555 219.930 ;
        RECT 2258.845 219.760 2259.015 219.930 ;
        RECT 2259.305 219.760 2259.475 219.930 ;
        RECT 2260.685 219.760 2260.855 219.930 ;
        RECT 2261.145 219.760 2261.315 219.930 ;
        RECT 2261.605 219.760 2261.775 219.930 ;
        RECT 2262.065 219.760 2262.235 219.930 ;
        RECT 2262.525 219.760 2262.695 219.930 ;
        RECT 2262.985 219.760 2263.155 219.930 ;
        RECT 2263.445 219.760 2263.615 219.930 ;
        RECT 2263.905 219.760 2264.075 219.930 ;
        RECT 2264.365 219.760 2264.535 219.930 ;
        RECT 2264.825 219.760 2264.995 219.930 ;
        RECT 2265.285 219.760 2265.455 219.930 ;
        RECT 2266.665 219.760 2266.835 219.930 ;
        RECT 2267.125 219.760 2267.295 219.930 ;
        RECT 2267.585 219.760 2267.755 219.930 ;
        RECT 2268.045 219.760 2268.215 219.930 ;
        RECT 2268.505 219.760 2268.675 219.930 ;
        RECT 2268.965 219.760 2269.135 219.930 ;
        RECT 2269.425 219.760 2269.595 219.930 ;
        RECT 2269.885 219.760 2270.055 219.930 ;
        RECT 2270.345 219.760 2270.515 219.930 ;
        RECT 2270.805 219.760 2270.975 219.930 ;
        RECT 2271.265 219.760 2271.435 219.930 ;
      LAYER met1 ;
        RECT 2146.000 219.605 2272.040 220.085 ;
        RECT 2146.000 214.165 2272.040 214.645 ;
      LAYER via ;
        RECT 2202.150 219.685 2203.935 219.985 ;
        RECT 2202.150 214.245 2203.935 214.545 ;
      LAYER met2 ;
        RECT 2202.110 219.625 2203.975 220.055 ;
        RECT 2202.110 214.185 2203.975 214.615 ;
      LAYER via2 ;
        RECT 2202.150 219.685 2203.935 219.985 ;
        RECT 2202.150 214.245 2203.935 214.545 ;
      LAYER met3 ;
        RECT 2202.120 209.800 2203.970 220.055 ;
    END
    PORT
      LAYER li1 ;
        RECT 204.715 1726.870 204.885 1727.040 ;
        RECT 210.155 1726.870 210.325 1727.040 ;
      LAYER li1 ;
        RECT 210.155 1726.640 210.325 1726.725 ;
      LAYER li1 ;
        RECT 204.715 1726.410 204.885 1726.580 ;
        RECT 204.715 1725.950 204.885 1726.120 ;
        RECT 204.715 1725.490 204.885 1725.660 ;
        RECT 204.715 1725.030 204.885 1725.200 ;
        RECT 204.715 1724.570 204.885 1724.740 ;
        RECT 204.715 1724.110 204.885 1724.280 ;
        RECT 204.715 1723.650 204.885 1723.820 ;
        RECT 204.715 1723.190 204.885 1723.360 ;
      LAYER li1 ;
        RECT 209.720 1723.235 210.325 1726.640 ;
      LAYER li1 ;
        RECT 204.715 1722.730 204.885 1722.900 ;
      LAYER li1 ;
        RECT 208.470 1722.885 210.325 1723.235 ;
      LAYER li1 ;
        RECT 204.715 1722.270 204.885 1722.440 ;
        RECT 204.715 1721.810 204.885 1721.980 ;
        RECT 204.715 1721.350 204.885 1721.520 ;
      LAYER li1 ;
        RECT 209.720 1721.295 210.325 1722.885 ;
        RECT 210.155 1721.205 210.325 1721.295 ;
      LAYER li1 ;
        RECT 204.715 1720.890 204.885 1721.060 ;
        RECT 210.155 1720.890 210.325 1721.060 ;
      LAYER li1 ;
        RECT 210.155 1720.660 210.325 1720.745 ;
      LAYER li1 ;
        RECT 204.715 1720.430 204.885 1720.600 ;
        RECT 204.715 1719.970 204.885 1720.140 ;
        RECT 204.715 1719.510 204.885 1719.680 ;
        RECT 204.715 1719.050 204.885 1719.220 ;
        RECT 204.715 1718.590 204.885 1718.760 ;
        RECT 204.715 1718.130 204.885 1718.300 ;
        RECT 204.715 1717.670 204.885 1717.840 ;
        RECT 204.715 1717.210 204.885 1717.380 ;
      LAYER li1 ;
        RECT 209.720 1717.255 210.325 1720.660 ;
      LAYER li1 ;
        RECT 204.715 1716.750 204.885 1716.920 ;
      LAYER li1 ;
        RECT 208.470 1716.905 210.325 1717.255 ;
      LAYER li1 ;
        RECT 204.715 1716.290 204.885 1716.460 ;
        RECT 204.715 1715.830 204.885 1716.000 ;
        RECT 204.715 1715.370 204.885 1715.540 ;
      LAYER li1 ;
        RECT 209.720 1715.315 210.325 1716.905 ;
        RECT 210.155 1715.225 210.325 1715.315 ;
      LAYER li1 ;
        RECT 204.715 1714.910 204.885 1715.080 ;
        RECT 210.155 1714.910 210.325 1715.080 ;
      LAYER li1 ;
        RECT 210.155 1714.680 210.325 1714.765 ;
      LAYER li1 ;
        RECT 204.715 1714.450 204.885 1714.620 ;
        RECT 204.715 1713.990 204.885 1714.160 ;
        RECT 204.715 1713.530 204.885 1713.700 ;
        RECT 204.715 1713.070 204.885 1713.240 ;
        RECT 204.715 1712.610 204.885 1712.780 ;
        RECT 204.715 1712.150 204.885 1712.320 ;
        RECT 204.715 1711.690 204.885 1711.860 ;
        RECT 204.715 1711.230 204.885 1711.400 ;
      LAYER li1 ;
        RECT 209.720 1711.275 210.325 1714.680 ;
      LAYER li1 ;
        RECT 204.715 1710.770 204.885 1710.940 ;
      LAYER li1 ;
        RECT 208.470 1710.925 210.325 1711.275 ;
      LAYER li1 ;
        RECT 204.715 1710.310 204.885 1710.480 ;
        RECT 204.715 1709.850 204.885 1710.020 ;
        RECT 204.715 1709.390 204.885 1709.560 ;
      LAYER li1 ;
        RECT 209.720 1709.335 210.325 1710.925 ;
        RECT 210.155 1709.245 210.325 1709.335 ;
      LAYER li1 ;
        RECT 204.715 1708.930 204.885 1709.100 ;
        RECT 210.155 1708.930 210.325 1709.100 ;
      LAYER li1 ;
        RECT 210.155 1708.700 210.325 1708.785 ;
      LAYER li1 ;
        RECT 204.715 1708.470 204.885 1708.640 ;
        RECT 204.715 1708.010 204.885 1708.180 ;
        RECT 204.715 1707.550 204.885 1707.720 ;
        RECT 204.715 1707.090 204.885 1707.260 ;
        RECT 204.715 1706.630 204.885 1706.800 ;
        RECT 204.715 1706.170 204.885 1706.340 ;
        RECT 204.715 1705.710 204.885 1705.880 ;
        RECT 204.715 1705.250 204.885 1705.420 ;
      LAYER li1 ;
        RECT 209.720 1705.295 210.325 1708.700 ;
      LAYER li1 ;
        RECT 204.715 1704.790 204.885 1704.960 ;
      LAYER li1 ;
        RECT 208.470 1704.945 210.325 1705.295 ;
      LAYER li1 ;
        RECT 204.715 1704.330 204.885 1704.500 ;
        RECT 204.715 1703.870 204.885 1704.040 ;
        RECT 204.715 1703.410 204.885 1703.580 ;
      LAYER li1 ;
        RECT 209.720 1703.355 210.325 1704.945 ;
        RECT 210.155 1703.265 210.325 1703.355 ;
      LAYER li1 ;
        RECT 204.715 1702.950 204.885 1703.120 ;
        RECT 210.155 1702.950 210.325 1703.120 ;
      LAYER li1 ;
        RECT 210.155 1702.720 210.325 1702.805 ;
      LAYER li1 ;
        RECT 204.715 1702.490 204.885 1702.660 ;
        RECT 204.715 1702.030 204.885 1702.200 ;
        RECT 204.715 1701.570 204.885 1701.740 ;
        RECT 204.715 1701.110 204.885 1701.280 ;
        RECT 204.715 1700.650 204.885 1700.820 ;
        RECT 204.715 1700.190 204.885 1700.360 ;
        RECT 204.715 1699.730 204.885 1699.900 ;
        RECT 204.715 1699.270 204.885 1699.440 ;
      LAYER li1 ;
        RECT 209.720 1699.315 210.325 1702.720 ;
      LAYER li1 ;
        RECT 204.715 1698.810 204.885 1698.980 ;
      LAYER li1 ;
        RECT 208.470 1698.965 210.325 1699.315 ;
      LAYER li1 ;
        RECT 204.715 1698.350 204.885 1698.520 ;
        RECT 204.715 1697.890 204.885 1698.060 ;
        RECT 204.715 1697.430 204.885 1697.600 ;
      LAYER li1 ;
        RECT 209.720 1697.375 210.325 1698.965 ;
        RECT 210.155 1697.285 210.325 1697.375 ;
      LAYER li1 ;
        RECT 204.715 1696.970 204.885 1697.140 ;
        RECT 210.155 1696.970 210.325 1697.140 ;
      LAYER li1 ;
        RECT 210.155 1696.740 210.325 1696.825 ;
      LAYER li1 ;
        RECT 204.715 1696.510 204.885 1696.680 ;
        RECT 204.715 1696.050 204.885 1696.220 ;
        RECT 204.715 1695.590 204.885 1695.760 ;
        RECT 204.715 1695.130 204.885 1695.300 ;
        RECT 204.715 1694.670 204.885 1694.840 ;
        RECT 204.715 1694.210 204.885 1694.380 ;
        RECT 204.715 1693.750 204.885 1693.920 ;
        RECT 204.715 1693.290 204.885 1693.460 ;
      LAYER li1 ;
        RECT 209.720 1693.335 210.325 1696.740 ;
      LAYER li1 ;
        RECT 204.715 1692.830 204.885 1693.000 ;
      LAYER li1 ;
        RECT 208.470 1692.985 210.325 1693.335 ;
      LAYER li1 ;
        RECT 204.715 1692.370 204.885 1692.540 ;
        RECT 204.715 1691.910 204.885 1692.080 ;
        RECT 204.715 1691.450 204.885 1691.620 ;
      LAYER li1 ;
        RECT 209.720 1691.395 210.325 1692.985 ;
        RECT 210.155 1691.305 210.325 1691.395 ;
      LAYER li1 ;
        RECT 204.715 1690.990 204.885 1691.160 ;
        RECT 210.155 1690.990 210.325 1691.160 ;
      LAYER li1 ;
        RECT 210.155 1690.760 210.325 1690.845 ;
      LAYER li1 ;
        RECT 204.715 1690.530 204.885 1690.700 ;
        RECT 204.715 1690.070 204.885 1690.240 ;
        RECT 204.715 1689.610 204.885 1689.780 ;
        RECT 204.715 1689.150 204.885 1689.320 ;
        RECT 204.715 1688.690 204.885 1688.860 ;
        RECT 204.715 1688.230 204.885 1688.400 ;
        RECT 204.715 1687.770 204.885 1687.940 ;
        RECT 204.715 1687.310 204.885 1687.480 ;
      LAYER li1 ;
        RECT 209.720 1687.355 210.325 1690.760 ;
      LAYER li1 ;
        RECT 204.715 1686.850 204.885 1687.020 ;
      LAYER li1 ;
        RECT 208.470 1687.005 210.325 1687.355 ;
      LAYER li1 ;
        RECT 204.715 1686.390 204.885 1686.560 ;
        RECT 204.715 1685.930 204.885 1686.100 ;
        RECT 204.715 1685.470 204.885 1685.640 ;
      LAYER li1 ;
        RECT 209.720 1685.415 210.325 1687.005 ;
        RECT 210.155 1685.325 210.325 1685.415 ;
      LAYER li1 ;
        RECT 204.715 1685.010 204.885 1685.180 ;
        RECT 210.155 1685.010 210.325 1685.180 ;
      LAYER li1 ;
        RECT 210.155 1684.780 210.325 1684.865 ;
      LAYER li1 ;
        RECT 204.715 1684.550 204.885 1684.720 ;
        RECT 204.715 1684.090 204.885 1684.260 ;
        RECT 204.715 1683.630 204.885 1683.800 ;
        RECT 204.715 1683.170 204.885 1683.340 ;
        RECT 204.715 1682.710 204.885 1682.880 ;
        RECT 204.715 1682.250 204.885 1682.420 ;
        RECT 204.715 1681.790 204.885 1681.960 ;
        RECT 204.715 1681.330 204.885 1681.500 ;
      LAYER li1 ;
        RECT 209.720 1681.375 210.325 1684.780 ;
      LAYER li1 ;
        RECT 204.715 1680.870 204.885 1681.040 ;
      LAYER li1 ;
        RECT 208.470 1681.025 210.325 1681.375 ;
      LAYER li1 ;
        RECT 204.715 1680.410 204.885 1680.580 ;
        RECT 204.715 1679.950 204.885 1680.120 ;
        RECT 204.715 1679.490 204.885 1679.660 ;
      LAYER li1 ;
        RECT 209.720 1679.435 210.325 1681.025 ;
        RECT 210.155 1679.345 210.325 1679.435 ;
      LAYER li1 ;
        RECT 204.715 1679.030 204.885 1679.200 ;
        RECT 210.155 1679.030 210.325 1679.200 ;
      LAYER li1 ;
        RECT 210.155 1678.800 210.325 1678.885 ;
      LAYER li1 ;
        RECT 204.715 1678.570 204.885 1678.740 ;
        RECT 204.715 1678.110 204.885 1678.280 ;
        RECT 204.715 1677.650 204.885 1677.820 ;
        RECT 204.715 1677.190 204.885 1677.360 ;
        RECT 204.715 1676.730 204.885 1676.900 ;
        RECT 204.715 1676.270 204.885 1676.440 ;
        RECT 204.715 1675.810 204.885 1675.980 ;
        RECT 204.715 1675.350 204.885 1675.520 ;
      LAYER li1 ;
        RECT 209.720 1675.395 210.325 1678.800 ;
      LAYER li1 ;
        RECT 204.715 1674.890 204.885 1675.060 ;
      LAYER li1 ;
        RECT 208.470 1675.045 210.325 1675.395 ;
      LAYER li1 ;
        RECT 204.715 1674.430 204.885 1674.600 ;
        RECT 204.715 1673.970 204.885 1674.140 ;
        RECT 204.715 1673.510 204.885 1673.680 ;
      LAYER li1 ;
        RECT 209.720 1673.455 210.325 1675.045 ;
        RECT 210.155 1673.365 210.325 1673.455 ;
      LAYER li1 ;
        RECT 204.715 1673.050 204.885 1673.220 ;
        RECT 210.155 1673.050 210.325 1673.220 ;
      LAYER mcon ;
        RECT 210.155 1725.950 210.325 1726.120 ;
        RECT 210.155 1725.490 210.325 1725.660 ;
        RECT 210.155 1725.030 210.325 1725.200 ;
        RECT 210.155 1724.570 210.325 1724.740 ;
        RECT 210.155 1724.110 210.325 1724.280 ;
        RECT 210.155 1723.650 210.325 1723.820 ;
        RECT 210.155 1723.190 210.325 1723.360 ;
        RECT 210.155 1722.730 210.325 1722.900 ;
        RECT 210.155 1722.270 210.325 1722.440 ;
        RECT 210.155 1721.810 210.325 1721.980 ;
        RECT 210.155 1721.350 210.325 1721.520 ;
        RECT 210.155 1719.970 210.325 1720.140 ;
        RECT 210.155 1719.510 210.325 1719.680 ;
        RECT 210.155 1719.050 210.325 1719.220 ;
        RECT 210.155 1718.590 210.325 1718.760 ;
        RECT 210.155 1718.130 210.325 1718.300 ;
        RECT 210.155 1717.670 210.325 1717.840 ;
        RECT 210.155 1717.210 210.325 1717.380 ;
        RECT 210.155 1716.750 210.325 1716.920 ;
        RECT 210.155 1716.290 210.325 1716.460 ;
        RECT 210.155 1715.830 210.325 1716.000 ;
        RECT 210.155 1715.370 210.325 1715.540 ;
        RECT 210.155 1713.990 210.325 1714.160 ;
        RECT 210.155 1713.530 210.325 1713.700 ;
        RECT 210.155 1713.070 210.325 1713.240 ;
        RECT 210.155 1712.610 210.325 1712.780 ;
        RECT 210.155 1712.150 210.325 1712.320 ;
        RECT 210.155 1711.690 210.325 1711.860 ;
        RECT 210.155 1711.230 210.325 1711.400 ;
        RECT 210.155 1710.770 210.325 1710.940 ;
        RECT 210.155 1710.310 210.325 1710.480 ;
        RECT 210.155 1709.850 210.325 1710.020 ;
        RECT 210.155 1709.390 210.325 1709.560 ;
        RECT 210.155 1708.010 210.325 1708.180 ;
        RECT 210.155 1707.550 210.325 1707.720 ;
        RECT 210.155 1707.090 210.325 1707.260 ;
        RECT 210.155 1706.630 210.325 1706.800 ;
        RECT 210.155 1706.170 210.325 1706.340 ;
        RECT 210.155 1705.710 210.325 1705.880 ;
        RECT 210.155 1705.250 210.325 1705.420 ;
        RECT 210.155 1704.790 210.325 1704.960 ;
        RECT 210.155 1704.330 210.325 1704.500 ;
        RECT 210.155 1703.870 210.325 1704.040 ;
        RECT 210.155 1703.410 210.325 1703.580 ;
        RECT 210.155 1702.030 210.325 1702.200 ;
        RECT 210.155 1701.570 210.325 1701.740 ;
        RECT 210.155 1701.110 210.325 1701.280 ;
        RECT 210.155 1700.650 210.325 1700.820 ;
        RECT 210.155 1700.190 210.325 1700.360 ;
        RECT 210.155 1699.730 210.325 1699.900 ;
        RECT 210.155 1699.270 210.325 1699.440 ;
        RECT 210.155 1698.810 210.325 1698.980 ;
        RECT 210.155 1698.350 210.325 1698.520 ;
        RECT 210.155 1697.890 210.325 1698.060 ;
        RECT 210.155 1697.430 210.325 1697.600 ;
        RECT 210.155 1696.050 210.325 1696.220 ;
        RECT 210.155 1695.590 210.325 1695.760 ;
        RECT 210.155 1695.130 210.325 1695.300 ;
        RECT 210.155 1694.670 210.325 1694.840 ;
        RECT 210.155 1694.210 210.325 1694.380 ;
        RECT 210.155 1693.750 210.325 1693.920 ;
        RECT 210.155 1693.290 210.325 1693.460 ;
        RECT 210.155 1692.830 210.325 1693.000 ;
        RECT 210.155 1692.370 210.325 1692.540 ;
        RECT 210.155 1691.910 210.325 1692.080 ;
        RECT 210.155 1691.450 210.325 1691.620 ;
        RECT 210.155 1690.070 210.325 1690.240 ;
        RECT 210.155 1689.610 210.325 1689.780 ;
        RECT 210.155 1689.150 210.325 1689.320 ;
        RECT 210.155 1688.690 210.325 1688.860 ;
        RECT 210.155 1688.230 210.325 1688.400 ;
        RECT 210.155 1687.770 210.325 1687.940 ;
        RECT 210.155 1687.310 210.325 1687.480 ;
        RECT 210.155 1686.850 210.325 1687.020 ;
        RECT 210.155 1686.390 210.325 1686.560 ;
        RECT 210.155 1685.930 210.325 1686.100 ;
        RECT 210.155 1685.470 210.325 1685.640 ;
        RECT 210.155 1684.090 210.325 1684.260 ;
        RECT 210.155 1683.630 210.325 1683.800 ;
        RECT 210.155 1683.170 210.325 1683.340 ;
        RECT 210.155 1682.710 210.325 1682.880 ;
        RECT 210.155 1682.250 210.325 1682.420 ;
        RECT 210.155 1681.790 210.325 1681.960 ;
        RECT 210.155 1681.330 210.325 1681.500 ;
        RECT 210.155 1680.870 210.325 1681.040 ;
        RECT 210.155 1680.410 210.325 1680.580 ;
        RECT 210.155 1679.950 210.325 1680.120 ;
        RECT 210.155 1679.490 210.325 1679.660 ;
        RECT 210.155 1678.110 210.325 1678.280 ;
        RECT 210.155 1677.650 210.325 1677.820 ;
        RECT 210.155 1677.190 210.325 1677.360 ;
        RECT 210.155 1676.730 210.325 1676.900 ;
        RECT 210.155 1676.270 210.325 1676.440 ;
        RECT 210.155 1675.810 210.325 1675.980 ;
        RECT 210.155 1675.350 210.325 1675.520 ;
        RECT 210.155 1674.890 210.325 1675.060 ;
        RECT 210.155 1674.430 210.325 1674.600 ;
        RECT 210.155 1673.970 210.325 1674.140 ;
        RECT 210.155 1673.510 210.325 1673.680 ;
      LAYER met1 ;
        RECT 204.560 1672.905 205.040 1730.790 ;
        RECT 210.000 1672.905 210.480 1730.800 ;
      LAYER via ;
        RECT 204.655 1728.815 204.955 1730.600 ;
        RECT 210.095 1728.815 210.395 1730.600 ;
      LAYER met2 ;
        RECT 204.595 1728.775 205.025 1730.640 ;
        RECT 210.035 1728.775 210.465 1730.640 ;
      LAYER via2 ;
        RECT 204.655 1728.815 204.955 1730.600 ;
        RECT 210.095 1728.815 210.395 1730.600 ;
      LAYER met3 ;
        RECT 200.210 1728.780 210.465 1730.630 ;
    END
    PORT
      LAYER li1 ;
        RECT 204.605 3014.775 204.775 3014.945 ;
        RECT 210.045 3014.775 210.215 3014.945 ;
      LAYER li1 ;
        RECT 210.045 3014.545 210.215 3014.630 ;
      LAYER li1 ;
        RECT 204.605 3014.315 204.775 3014.485 ;
        RECT 204.605 3013.855 204.775 3014.025 ;
        RECT 204.605 3013.395 204.775 3013.565 ;
        RECT 204.605 3012.935 204.775 3013.105 ;
        RECT 204.605 3012.475 204.775 3012.645 ;
        RECT 204.605 3012.015 204.775 3012.185 ;
        RECT 204.605 3011.555 204.775 3011.725 ;
        RECT 204.605 3011.095 204.775 3011.265 ;
      LAYER li1 ;
        RECT 209.610 3011.140 210.215 3014.545 ;
      LAYER li1 ;
        RECT 204.605 3010.635 204.775 3010.805 ;
      LAYER li1 ;
        RECT 208.360 3010.790 210.215 3011.140 ;
      LAYER li1 ;
        RECT 204.605 3010.175 204.775 3010.345 ;
        RECT 204.605 3009.715 204.775 3009.885 ;
        RECT 204.605 3009.255 204.775 3009.425 ;
      LAYER li1 ;
        RECT 209.610 3009.200 210.215 3010.790 ;
        RECT 210.045 3009.110 210.215 3009.200 ;
      LAYER li1 ;
        RECT 204.605 3008.795 204.775 3008.965 ;
        RECT 210.045 3008.795 210.215 3008.965 ;
      LAYER li1 ;
        RECT 210.045 3008.565 210.215 3008.650 ;
      LAYER li1 ;
        RECT 204.605 3008.335 204.775 3008.505 ;
        RECT 204.605 3007.875 204.775 3008.045 ;
        RECT 204.605 3007.415 204.775 3007.585 ;
        RECT 204.605 3006.955 204.775 3007.125 ;
        RECT 204.605 3006.495 204.775 3006.665 ;
        RECT 204.605 3006.035 204.775 3006.205 ;
        RECT 204.605 3005.575 204.775 3005.745 ;
        RECT 204.605 3005.115 204.775 3005.285 ;
      LAYER li1 ;
        RECT 209.610 3005.160 210.215 3008.565 ;
      LAYER li1 ;
        RECT 204.605 3004.655 204.775 3004.825 ;
      LAYER li1 ;
        RECT 208.360 3004.810 210.215 3005.160 ;
      LAYER li1 ;
        RECT 204.605 3004.195 204.775 3004.365 ;
        RECT 204.605 3003.735 204.775 3003.905 ;
        RECT 204.605 3003.275 204.775 3003.445 ;
      LAYER li1 ;
        RECT 209.610 3003.220 210.215 3004.810 ;
        RECT 210.045 3003.130 210.215 3003.220 ;
      LAYER li1 ;
        RECT 204.605 3002.815 204.775 3002.985 ;
        RECT 210.045 3002.815 210.215 3002.985 ;
      LAYER li1 ;
        RECT 210.045 3002.585 210.215 3002.670 ;
      LAYER li1 ;
        RECT 204.605 3002.355 204.775 3002.525 ;
        RECT 204.605 3001.895 204.775 3002.065 ;
        RECT 204.605 3001.435 204.775 3001.605 ;
        RECT 204.605 3000.975 204.775 3001.145 ;
        RECT 204.605 3000.515 204.775 3000.685 ;
        RECT 204.605 3000.055 204.775 3000.225 ;
        RECT 204.605 2999.595 204.775 2999.765 ;
        RECT 204.605 2999.135 204.775 2999.305 ;
      LAYER li1 ;
        RECT 209.610 2999.180 210.215 3002.585 ;
      LAYER li1 ;
        RECT 204.605 2998.675 204.775 2998.845 ;
      LAYER li1 ;
        RECT 208.360 2998.830 210.215 2999.180 ;
      LAYER li1 ;
        RECT 204.605 2998.215 204.775 2998.385 ;
        RECT 204.605 2997.755 204.775 2997.925 ;
        RECT 204.605 2997.295 204.775 2997.465 ;
      LAYER li1 ;
        RECT 209.610 2997.240 210.215 2998.830 ;
        RECT 210.045 2997.150 210.215 2997.240 ;
      LAYER li1 ;
        RECT 204.605 2996.835 204.775 2997.005 ;
        RECT 210.045 2996.835 210.215 2997.005 ;
      LAYER li1 ;
        RECT 210.045 2996.605 210.215 2996.690 ;
      LAYER li1 ;
        RECT 204.605 2996.375 204.775 2996.545 ;
        RECT 204.605 2995.915 204.775 2996.085 ;
        RECT 204.605 2995.455 204.775 2995.625 ;
        RECT 204.605 2994.995 204.775 2995.165 ;
        RECT 204.605 2994.535 204.775 2994.705 ;
        RECT 204.605 2994.075 204.775 2994.245 ;
        RECT 204.605 2993.615 204.775 2993.785 ;
        RECT 204.605 2993.155 204.775 2993.325 ;
      LAYER li1 ;
        RECT 209.610 2993.200 210.215 2996.605 ;
      LAYER li1 ;
        RECT 204.605 2992.695 204.775 2992.865 ;
      LAYER li1 ;
        RECT 208.360 2992.850 210.215 2993.200 ;
      LAYER li1 ;
        RECT 204.605 2992.235 204.775 2992.405 ;
        RECT 204.605 2991.775 204.775 2991.945 ;
        RECT 204.605 2991.315 204.775 2991.485 ;
      LAYER li1 ;
        RECT 209.610 2991.260 210.215 2992.850 ;
        RECT 210.045 2991.170 210.215 2991.260 ;
      LAYER li1 ;
        RECT 204.605 2990.855 204.775 2991.025 ;
        RECT 210.045 2990.855 210.215 2991.025 ;
      LAYER li1 ;
        RECT 210.045 2990.625 210.215 2990.710 ;
      LAYER li1 ;
        RECT 204.605 2990.395 204.775 2990.565 ;
        RECT 204.605 2989.935 204.775 2990.105 ;
        RECT 204.605 2989.475 204.775 2989.645 ;
        RECT 204.605 2989.015 204.775 2989.185 ;
        RECT 204.605 2988.555 204.775 2988.725 ;
        RECT 204.605 2988.095 204.775 2988.265 ;
        RECT 204.605 2987.635 204.775 2987.805 ;
        RECT 204.605 2987.175 204.775 2987.345 ;
      LAYER li1 ;
        RECT 209.610 2987.220 210.215 2990.625 ;
      LAYER li1 ;
        RECT 204.605 2986.715 204.775 2986.885 ;
      LAYER li1 ;
        RECT 208.360 2986.870 210.215 2987.220 ;
      LAYER li1 ;
        RECT 204.605 2986.255 204.775 2986.425 ;
        RECT 204.605 2985.795 204.775 2985.965 ;
        RECT 204.605 2985.335 204.775 2985.505 ;
      LAYER li1 ;
        RECT 209.610 2985.280 210.215 2986.870 ;
        RECT 210.045 2985.190 210.215 2985.280 ;
      LAYER li1 ;
        RECT 204.605 2984.875 204.775 2985.045 ;
        RECT 210.045 2984.875 210.215 2985.045 ;
      LAYER mcon ;
        RECT 210.045 3013.855 210.215 3014.025 ;
        RECT 210.045 3013.395 210.215 3013.565 ;
        RECT 210.045 3012.935 210.215 3013.105 ;
        RECT 210.045 3012.475 210.215 3012.645 ;
        RECT 210.045 3012.015 210.215 3012.185 ;
        RECT 210.045 3011.555 210.215 3011.725 ;
        RECT 210.045 3011.095 210.215 3011.265 ;
        RECT 210.045 3010.635 210.215 3010.805 ;
        RECT 210.045 3010.175 210.215 3010.345 ;
        RECT 210.045 3009.715 210.215 3009.885 ;
        RECT 210.045 3009.255 210.215 3009.425 ;
        RECT 210.045 3007.875 210.215 3008.045 ;
        RECT 210.045 3007.415 210.215 3007.585 ;
        RECT 210.045 3006.955 210.215 3007.125 ;
        RECT 210.045 3006.495 210.215 3006.665 ;
        RECT 210.045 3006.035 210.215 3006.205 ;
        RECT 210.045 3005.575 210.215 3005.745 ;
        RECT 210.045 3005.115 210.215 3005.285 ;
        RECT 210.045 3004.655 210.215 3004.825 ;
        RECT 210.045 3004.195 210.215 3004.365 ;
        RECT 210.045 3003.735 210.215 3003.905 ;
        RECT 210.045 3003.275 210.215 3003.445 ;
        RECT 210.045 3001.895 210.215 3002.065 ;
        RECT 210.045 3001.435 210.215 3001.605 ;
        RECT 210.045 3000.975 210.215 3001.145 ;
        RECT 210.045 3000.515 210.215 3000.685 ;
        RECT 210.045 3000.055 210.215 3000.225 ;
        RECT 210.045 2999.595 210.215 2999.765 ;
        RECT 210.045 2999.135 210.215 2999.305 ;
        RECT 210.045 2998.675 210.215 2998.845 ;
        RECT 210.045 2998.215 210.215 2998.385 ;
        RECT 210.045 2997.755 210.215 2997.925 ;
        RECT 210.045 2997.295 210.215 2997.465 ;
        RECT 210.045 2995.915 210.215 2996.085 ;
        RECT 210.045 2995.455 210.215 2995.625 ;
        RECT 210.045 2994.995 210.215 2995.165 ;
        RECT 210.045 2994.535 210.215 2994.705 ;
        RECT 210.045 2994.075 210.215 2994.245 ;
        RECT 210.045 2993.615 210.215 2993.785 ;
        RECT 210.045 2993.155 210.215 2993.325 ;
        RECT 210.045 2992.695 210.215 2992.865 ;
        RECT 210.045 2992.235 210.215 2992.405 ;
        RECT 210.045 2991.775 210.215 2991.945 ;
        RECT 210.045 2991.315 210.215 2991.485 ;
        RECT 210.045 2989.935 210.215 2990.105 ;
        RECT 210.045 2989.475 210.215 2989.645 ;
        RECT 210.045 2989.015 210.215 2989.185 ;
        RECT 210.045 2988.555 210.215 2988.725 ;
        RECT 210.045 2988.095 210.215 2988.265 ;
        RECT 210.045 2987.635 210.215 2987.805 ;
        RECT 210.045 2987.175 210.215 2987.345 ;
        RECT 210.045 2986.715 210.215 2986.885 ;
        RECT 210.045 2986.255 210.215 2986.425 ;
        RECT 210.045 2985.795 210.215 2985.965 ;
        RECT 210.045 2985.335 210.215 2985.505 ;
      LAYER met1 ;
        RECT 204.450 2984.730 204.930 3019.020 ;
        RECT 209.890 2984.730 210.370 3019.030 ;
      LAYER via ;
        RECT 204.560 3017.070 204.860 3018.855 ;
        RECT 210.000 3017.070 210.300 3018.855 ;
      LAYER met2 ;
        RECT 204.500 3017.030 204.930 3018.895 ;
        RECT 209.940 3017.030 210.370 3018.895 ;
      LAYER via2 ;
        RECT 204.560 3017.070 204.860 3018.855 ;
        RECT 210.000 3017.070 210.300 3018.855 ;
      LAYER met3 ;
        RECT 200.115 3017.035 210.370 3018.885 ;
    END
  END vccd
  OBS
      LAYER nwell ;
        RECT 3377.675 3601.870 3379.280 3608.690 ;
      LAYER pwell ;
        RECT 3379.610 3608.055 3380.395 3608.485 ;
        RECT 3380.775 3608.055 3381.560 3608.485 ;
        RECT 3380.690 3607.960 3381.600 3608.035 ;
        RECT 3380.435 3607.680 3381.600 3607.960 ;
        RECT 3380.690 3602.905 3381.600 3607.680 ;
        RECT 3379.610 3602.075 3380.395 3602.505 ;
        RECT 3380.775 3602.075 3381.560 3602.505 ;
      LAYER nwell ;
        RECT 3381.890 3601.870 3384.720 3608.690 ;
      LAYER pwell ;
        RECT 3385.050 3608.055 3385.835 3608.485 ;
        RECT 3385.010 3602.840 3385.920 3607.655 ;
        RECT 3385.010 3602.670 3386.110 3602.840 ;
        RECT 3385.010 3602.525 3385.920 3602.670 ;
        RECT 3385.050 3602.075 3385.835 3602.505 ;
        RECT 202.160 3014.645 202.945 3015.075 ;
        RECT 202.075 3009.430 202.985 3014.245 ;
        RECT 201.885 3009.260 202.985 3009.430 ;
        RECT 202.075 3009.115 202.985 3009.260 ;
        RECT 202.160 3008.665 202.945 3009.095 ;
        RECT 202.075 3003.450 202.985 3008.265 ;
        RECT 201.885 3003.280 202.985 3003.450 ;
        RECT 202.075 3003.135 202.985 3003.280 ;
        RECT 202.160 3002.685 202.945 3003.115 ;
        RECT 202.075 2997.470 202.985 3002.285 ;
        RECT 201.885 2997.300 202.985 2997.470 ;
        RECT 202.075 2997.155 202.985 2997.300 ;
        RECT 202.160 2996.705 202.945 2997.135 ;
        RECT 202.075 2991.490 202.985 2996.305 ;
        RECT 201.885 2991.320 202.985 2991.490 ;
        RECT 202.075 2991.175 202.985 2991.320 ;
        RECT 202.160 2990.725 202.945 2991.155 ;
        RECT 202.075 2985.510 202.985 2990.325 ;
        RECT 201.885 2985.340 202.985 2985.510 ;
        RECT 202.075 2985.195 202.985 2985.340 ;
        RECT 202.160 2984.745 202.945 2985.175 ;
      LAYER nwell ;
        RECT 203.275 2984.540 206.105 3015.280 ;
      LAYER pwell ;
        RECT 206.435 3014.645 207.220 3015.075 ;
        RECT 207.600 3014.645 208.385 3015.075 ;
        RECT 206.395 3014.550 207.305 3014.625 ;
        RECT 206.395 3014.270 207.560 3014.550 ;
        RECT 206.395 3009.495 207.305 3014.270 ;
        RECT 206.435 3008.665 207.220 3009.095 ;
        RECT 207.600 3008.665 208.385 3009.095 ;
        RECT 206.395 3008.570 207.305 3008.645 ;
        RECT 206.395 3008.290 207.560 3008.570 ;
        RECT 206.395 3003.515 207.305 3008.290 ;
        RECT 206.435 3002.685 207.220 3003.115 ;
        RECT 207.600 3002.685 208.385 3003.115 ;
        RECT 206.395 3002.590 207.305 3002.665 ;
        RECT 206.395 3002.310 207.560 3002.590 ;
        RECT 206.395 2997.535 207.305 3002.310 ;
        RECT 206.435 2996.705 207.220 2997.135 ;
        RECT 207.600 2996.705 208.385 2997.135 ;
        RECT 206.395 2996.610 207.305 2996.685 ;
        RECT 206.395 2996.330 207.560 2996.610 ;
        RECT 206.395 2991.555 207.305 2996.330 ;
        RECT 206.435 2990.725 207.220 2991.155 ;
        RECT 207.600 2990.725 208.385 2991.155 ;
        RECT 206.395 2990.630 207.305 2990.705 ;
        RECT 206.395 2990.350 207.560 2990.630 ;
        RECT 206.395 2985.575 207.305 2990.350 ;
        RECT 206.435 2984.745 207.220 2985.175 ;
        RECT 207.600 2984.745 208.385 2985.175 ;
      LAYER nwell ;
        RECT 208.715 2984.540 210.320 3015.280 ;
        RECT 3377.675 2195.870 3379.280 2238.570 ;
      LAYER pwell ;
        RECT 3379.610 2237.935 3380.395 2238.365 ;
        RECT 3380.775 2237.935 3381.560 2238.365 ;
        RECT 3380.690 2237.840 3381.600 2237.915 ;
        RECT 3380.435 2237.560 3381.600 2237.840 ;
        RECT 3380.690 2232.785 3381.600 2237.560 ;
        RECT 3379.610 2231.955 3380.395 2232.385 ;
        RECT 3380.775 2231.955 3381.560 2232.385 ;
        RECT 3380.690 2231.860 3381.600 2231.935 ;
        RECT 3380.435 2231.580 3381.600 2231.860 ;
        RECT 3380.690 2226.805 3381.600 2231.580 ;
        RECT 3379.610 2225.975 3380.395 2226.405 ;
        RECT 3380.775 2225.975 3381.560 2226.405 ;
        RECT 3380.690 2225.880 3381.600 2225.955 ;
        RECT 3380.435 2225.600 3381.600 2225.880 ;
        RECT 3380.690 2220.825 3381.600 2225.600 ;
        RECT 3379.610 2219.995 3380.395 2220.425 ;
        RECT 3380.775 2219.995 3381.560 2220.425 ;
        RECT 3380.690 2219.900 3381.600 2219.975 ;
        RECT 3380.435 2219.620 3381.600 2219.900 ;
        RECT 3380.690 2214.845 3381.600 2219.620 ;
        RECT 3379.610 2214.015 3380.395 2214.445 ;
        RECT 3380.775 2214.015 3381.560 2214.445 ;
        RECT 3380.690 2213.920 3381.600 2213.995 ;
        RECT 3380.435 2213.640 3381.600 2213.920 ;
        RECT 3380.690 2208.865 3381.600 2213.640 ;
        RECT 3379.610 2208.035 3380.395 2208.465 ;
        RECT 3380.775 2208.035 3381.560 2208.465 ;
        RECT 3380.690 2207.940 3381.600 2208.015 ;
        RECT 3380.435 2207.660 3381.600 2207.940 ;
        RECT 3380.690 2202.885 3381.600 2207.660 ;
        RECT 3379.610 2202.055 3380.395 2202.485 ;
        RECT 3380.775 2202.055 3381.560 2202.485 ;
        RECT 3380.690 2201.960 3381.600 2202.035 ;
        RECT 3380.435 2201.680 3381.600 2201.960 ;
        RECT 3380.690 2196.905 3381.600 2201.680 ;
        RECT 3379.610 2196.075 3380.395 2196.505 ;
        RECT 3380.775 2196.075 3381.560 2196.505 ;
      LAYER nwell ;
        RECT 3381.890 2195.870 3384.720 2238.570 ;
      LAYER pwell ;
        RECT 3385.050 2237.935 3385.835 2238.365 ;
        RECT 3385.010 2232.720 3385.920 2237.535 ;
        RECT 3385.010 2232.550 3386.110 2232.720 ;
        RECT 3385.010 2232.405 3385.920 2232.550 ;
        RECT 3385.050 2231.955 3385.835 2232.385 ;
        RECT 3385.010 2226.740 3385.920 2231.555 ;
        RECT 3385.010 2226.570 3386.110 2226.740 ;
        RECT 3385.010 2226.425 3385.920 2226.570 ;
        RECT 3385.050 2225.975 3385.835 2226.405 ;
        RECT 3385.010 2220.760 3385.920 2225.575 ;
        RECT 3385.010 2220.590 3386.110 2220.760 ;
        RECT 3385.010 2220.445 3385.920 2220.590 ;
        RECT 3385.050 2219.995 3385.835 2220.425 ;
        RECT 3385.010 2214.780 3385.920 2219.595 ;
        RECT 3385.010 2214.610 3386.110 2214.780 ;
        RECT 3385.010 2214.465 3385.920 2214.610 ;
        RECT 3385.050 2214.015 3385.835 2214.445 ;
        RECT 3385.010 2208.800 3385.920 2213.615 ;
        RECT 3385.010 2208.630 3386.110 2208.800 ;
        RECT 3385.010 2208.485 3385.920 2208.630 ;
        RECT 3385.050 2208.035 3385.835 2208.465 ;
        RECT 3385.010 2202.820 3385.920 2207.635 ;
        RECT 3385.010 2202.650 3386.110 2202.820 ;
        RECT 3385.010 2202.505 3385.920 2202.650 ;
        RECT 3385.050 2202.055 3385.835 2202.485 ;
        RECT 3385.010 2196.840 3385.920 2201.655 ;
        RECT 3385.010 2196.670 3386.110 2196.840 ;
        RECT 3385.010 2196.525 3385.920 2196.670 ;
        RECT 3385.050 2196.075 3385.835 2196.505 ;
        RECT 202.270 1726.740 203.055 1727.170 ;
        RECT 202.185 1721.525 203.095 1726.340 ;
        RECT 201.995 1721.355 203.095 1721.525 ;
        RECT 202.185 1721.210 203.095 1721.355 ;
        RECT 202.270 1720.760 203.055 1721.190 ;
        RECT 202.185 1715.545 203.095 1720.360 ;
        RECT 201.995 1715.375 203.095 1715.545 ;
        RECT 202.185 1715.230 203.095 1715.375 ;
        RECT 202.270 1714.780 203.055 1715.210 ;
        RECT 202.185 1709.565 203.095 1714.380 ;
        RECT 201.995 1709.395 203.095 1709.565 ;
        RECT 202.185 1709.250 203.095 1709.395 ;
        RECT 202.270 1708.800 203.055 1709.230 ;
        RECT 202.185 1703.585 203.095 1708.400 ;
        RECT 201.995 1703.415 203.095 1703.585 ;
        RECT 202.185 1703.270 203.095 1703.415 ;
        RECT 202.270 1702.820 203.055 1703.250 ;
        RECT 202.185 1697.605 203.095 1702.420 ;
        RECT 201.995 1697.435 203.095 1697.605 ;
        RECT 202.185 1697.290 203.095 1697.435 ;
        RECT 202.270 1696.840 203.055 1697.270 ;
        RECT 202.185 1691.625 203.095 1696.440 ;
        RECT 201.995 1691.455 203.095 1691.625 ;
        RECT 202.185 1691.310 203.095 1691.455 ;
        RECT 202.270 1690.860 203.055 1691.290 ;
        RECT 202.185 1685.645 203.095 1690.460 ;
        RECT 201.995 1685.475 203.095 1685.645 ;
        RECT 202.185 1685.330 203.095 1685.475 ;
        RECT 202.270 1684.880 203.055 1685.310 ;
        RECT 202.185 1679.665 203.095 1684.480 ;
        RECT 201.995 1679.495 203.095 1679.665 ;
        RECT 202.185 1679.350 203.095 1679.495 ;
        RECT 202.270 1678.900 203.055 1679.330 ;
        RECT 202.185 1673.685 203.095 1678.500 ;
        RECT 201.995 1673.515 203.095 1673.685 ;
        RECT 202.185 1673.370 203.095 1673.515 ;
        RECT 202.270 1672.920 203.055 1673.350 ;
      LAYER nwell ;
        RECT 203.385 1672.715 206.215 1727.375 ;
      LAYER pwell ;
        RECT 206.545 1726.740 207.330 1727.170 ;
        RECT 207.710 1726.740 208.495 1727.170 ;
        RECT 206.505 1726.645 207.415 1726.720 ;
        RECT 206.505 1726.365 207.670 1726.645 ;
        RECT 206.505 1721.590 207.415 1726.365 ;
        RECT 206.545 1720.760 207.330 1721.190 ;
        RECT 207.710 1720.760 208.495 1721.190 ;
        RECT 206.505 1720.665 207.415 1720.740 ;
        RECT 206.505 1720.385 207.670 1720.665 ;
        RECT 206.505 1715.610 207.415 1720.385 ;
        RECT 206.545 1714.780 207.330 1715.210 ;
        RECT 207.710 1714.780 208.495 1715.210 ;
        RECT 206.505 1714.685 207.415 1714.760 ;
        RECT 206.505 1714.405 207.670 1714.685 ;
        RECT 206.505 1709.630 207.415 1714.405 ;
        RECT 206.545 1708.800 207.330 1709.230 ;
        RECT 207.710 1708.800 208.495 1709.230 ;
        RECT 206.505 1708.705 207.415 1708.780 ;
        RECT 206.505 1708.425 207.670 1708.705 ;
        RECT 206.505 1703.650 207.415 1708.425 ;
        RECT 206.545 1702.820 207.330 1703.250 ;
        RECT 207.710 1702.820 208.495 1703.250 ;
        RECT 206.505 1702.725 207.415 1702.800 ;
        RECT 206.505 1702.445 207.670 1702.725 ;
        RECT 206.505 1697.670 207.415 1702.445 ;
        RECT 206.545 1696.840 207.330 1697.270 ;
        RECT 207.710 1696.840 208.495 1697.270 ;
        RECT 206.505 1696.745 207.415 1696.820 ;
        RECT 206.505 1696.465 207.670 1696.745 ;
        RECT 206.505 1691.690 207.415 1696.465 ;
        RECT 206.545 1690.860 207.330 1691.290 ;
        RECT 207.710 1690.860 208.495 1691.290 ;
        RECT 206.505 1690.765 207.415 1690.840 ;
        RECT 206.505 1690.485 207.670 1690.765 ;
        RECT 206.505 1685.710 207.415 1690.485 ;
        RECT 206.545 1684.880 207.330 1685.310 ;
        RECT 207.710 1684.880 208.495 1685.310 ;
        RECT 206.505 1684.785 207.415 1684.860 ;
        RECT 206.505 1684.505 207.670 1684.785 ;
        RECT 206.505 1679.730 207.415 1684.505 ;
        RECT 206.545 1678.900 207.330 1679.330 ;
        RECT 207.710 1678.900 208.495 1679.330 ;
        RECT 206.505 1678.805 207.415 1678.880 ;
        RECT 206.505 1678.525 207.670 1678.805 ;
        RECT 206.505 1673.750 207.415 1678.525 ;
        RECT 206.545 1672.920 207.330 1673.350 ;
        RECT 207.710 1672.920 208.495 1673.350 ;
      LAYER nwell ;
        RECT 208.825 1672.715 210.430 1727.375 ;
        RECT 668.810 218.430 729.450 220.035 ;
        RECT 758.510 218.430 795.230 220.035 ;
        RECT 2145.810 218.430 2206.450 220.035 ;
        RECT 2235.510 218.430 2272.230 220.035 ;
      LAYER pwell ;
        RECT 669.015 217.315 669.445 218.100 ;
        RECT 674.995 217.315 675.425 218.100 ;
        RECT 680.975 217.315 681.405 218.100 ;
        RECT 686.955 217.315 687.385 218.100 ;
        RECT 692.935 217.315 693.365 218.100 ;
        RECT 698.915 217.315 699.345 218.100 ;
        RECT 704.895 217.315 705.325 218.100 ;
        RECT 710.875 217.315 711.305 218.100 ;
        RECT 716.855 217.315 717.285 218.100 ;
        RECT 722.835 217.315 723.265 218.100 ;
        RECT 728.815 217.315 729.245 218.100 ;
        RECT 758.715 217.315 759.145 218.100 ;
        RECT 764.695 217.315 765.125 218.100 ;
        RECT 770.675 217.315 771.105 218.100 ;
        RECT 776.655 217.315 777.085 218.100 ;
        RECT 782.635 217.315 783.065 218.100 ;
        RECT 788.615 217.315 789.045 218.100 ;
        RECT 794.595 217.315 795.025 218.100 ;
        RECT 2146.015 217.315 2146.445 218.100 ;
        RECT 2151.995 217.315 2152.425 218.100 ;
        RECT 2157.975 217.315 2158.405 218.100 ;
        RECT 2163.955 217.315 2164.385 218.100 ;
        RECT 2169.935 217.315 2170.365 218.100 ;
        RECT 2175.915 217.315 2176.345 218.100 ;
        RECT 2181.895 217.315 2182.325 218.100 ;
        RECT 2187.875 217.315 2188.305 218.100 ;
        RECT 2193.855 217.315 2194.285 218.100 ;
        RECT 2199.835 217.315 2200.265 218.100 ;
        RECT 2205.815 217.315 2206.245 218.100 ;
        RECT 2235.715 217.315 2236.145 218.100 ;
        RECT 2241.695 217.315 2242.125 218.100 ;
        RECT 2247.675 217.315 2248.105 218.100 ;
        RECT 2253.655 217.315 2254.085 218.100 ;
        RECT 2259.635 217.315 2260.065 218.100 ;
        RECT 2265.615 217.315 2266.045 218.100 ;
        RECT 2271.595 217.315 2272.025 218.100 ;
        RECT 669.540 216.995 669.820 217.275 ;
        RECT 674.660 217.020 674.830 217.210 ;
        RECT 669.015 216.150 669.445 216.935 ;
        RECT 669.845 216.110 674.975 217.020 ;
        RECT 675.520 216.995 675.800 217.275 ;
        RECT 680.640 217.020 680.810 217.210 ;
        RECT 674.995 216.150 675.425 216.935 ;
        RECT 675.825 216.110 680.955 217.020 ;
        RECT 681.500 216.995 681.780 217.275 ;
        RECT 686.620 217.020 686.790 217.210 ;
        RECT 680.975 216.150 681.405 216.935 ;
        RECT 681.805 216.110 686.935 217.020 ;
        RECT 687.480 216.995 687.760 217.275 ;
        RECT 692.600 217.020 692.770 217.210 ;
        RECT 686.955 216.150 687.385 216.935 ;
        RECT 687.785 216.110 692.915 217.020 ;
        RECT 693.460 216.995 693.740 217.275 ;
        RECT 698.580 217.020 698.750 217.210 ;
        RECT 692.935 216.150 693.365 216.935 ;
        RECT 693.765 216.110 698.895 217.020 ;
        RECT 699.440 216.995 699.720 217.275 ;
        RECT 704.560 217.020 704.730 217.210 ;
        RECT 698.915 216.150 699.345 216.935 ;
        RECT 699.745 216.110 704.875 217.020 ;
        RECT 705.420 216.995 705.700 217.275 ;
        RECT 710.540 217.020 710.710 217.210 ;
        RECT 704.895 216.150 705.325 216.935 ;
        RECT 705.725 216.110 710.855 217.020 ;
        RECT 711.400 216.995 711.680 217.275 ;
        RECT 716.520 217.020 716.690 217.210 ;
        RECT 710.875 216.150 711.305 216.935 ;
        RECT 711.705 216.110 716.835 217.020 ;
        RECT 717.380 216.995 717.660 217.275 ;
        RECT 722.500 217.020 722.670 217.210 ;
        RECT 716.855 216.150 717.285 216.935 ;
        RECT 717.685 216.110 722.815 217.020 ;
        RECT 723.360 216.975 723.640 217.275 ;
        RECT 759.240 216.995 759.520 217.275 ;
        RECT 764.360 217.020 764.530 217.210 ;
        RECT 722.835 216.150 723.265 216.935 ;
        RECT 728.815 216.150 729.245 216.935 ;
        RECT 758.715 216.150 759.145 216.935 ;
        RECT 759.545 216.110 764.675 217.020 ;
        RECT 765.220 216.995 765.500 217.275 ;
        RECT 770.340 217.020 770.510 217.210 ;
        RECT 764.695 216.150 765.125 216.935 ;
        RECT 765.525 216.110 770.655 217.020 ;
        RECT 771.200 216.995 771.480 217.275 ;
        RECT 776.320 217.020 776.490 217.210 ;
        RECT 770.675 216.150 771.105 216.935 ;
        RECT 771.505 216.110 776.635 217.020 ;
        RECT 777.180 216.995 777.460 217.275 ;
        RECT 782.300 217.020 782.470 217.210 ;
        RECT 776.655 216.150 777.085 216.935 ;
        RECT 777.485 216.110 782.615 217.020 ;
        RECT 783.160 216.995 783.440 217.275 ;
        RECT 788.280 217.020 788.450 217.210 ;
        RECT 782.635 216.150 783.065 216.935 ;
        RECT 783.465 216.110 788.595 217.020 ;
        RECT 789.140 216.995 789.420 217.275 ;
        RECT 794.260 217.020 794.430 217.210 ;
        RECT 788.615 216.150 789.045 216.935 ;
        RECT 789.445 216.110 794.575 217.020 ;
        RECT 2146.540 216.995 2146.820 217.275 ;
        RECT 2151.660 217.020 2151.830 217.210 ;
        RECT 794.595 216.150 795.025 216.935 ;
        RECT 2146.015 216.150 2146.445 216.935 ;
        RECT 2146.845 216.110 2151.975 217.020 ;
        RECT 2152.520 216.995 2152.800 217.275 ;
        RECT 2157.640 217.020 2157.810 217.210 ;
        RECT 2151.995 216.150 2152.425 216.935 ;
        RECT 2152.825 216.110 2157.955 217.020 ;
        RECT 2158.500 216.995 2158.780 217.275 ;
        RECT 2163.620 217.020 2163.790 217.210 ;
        RECT 2157.975 216.150 2158.405 216.935 ;
        RECT 2158.805 216.110 2163.935 217.020 ;
        RECT 2164.480 216.995 2164.760 217.275 ;
        RECT 2169.600 217.020 2169.770 217.210 ;
        RECT 2163.955 216.150 2164.385 216.935 ;
        RECT 2164.785 216.110 2169.915 217.020 ;
        RECT 2170.460 216.995 2170.740 217.275 ;
        RECT 2175.580 217.020 2175.750 217.210 ;
        RECT 2169.935 216.150 2170.365 216.935 ;
        RECT 2170.765 216.110 2175.895 217.020 ;
        RECT 2176.440 216.995 2176.720 217.275 ;
        RECT 2181.560 217.020 2181.730 217.210 ;
        RECT 2175.915 216.150 2176.345 216.935 ;
        RECT 2176.745 216.110 2181.875 217.020 ;
        RECT 2182.420 216.995 2182.700 217.275 ;
        RECT 2187.540 217.020 2187.710 217.210 ;
        RECT 2181.895 216.150 2182.325 216.935 ;
        RECT 2182.725 216.110 2187.855 217.020 ;
        RECT 2188.400 216.995 2188.680 217.275 ;
        RECT 2193.520 217.020 2193.690 217.210 ;
        RECT 2187.875 216.150 2188.305 216.935 ;
        RECT 2188.705 216.110 2193.835 217.020 ;
        RECT 2194.380 216.995 2194.660 217.275 ;
        RECT 2199.500 217.020 2199.670 217.210 ;
        RECT 2193.855 216.150 2194.285 216.935 ;
        RECT 2194.685 216.110 2199.815 217.020 ;
        RECT 2200.360 216.975 2200.640 217.275 ;
        RECT 2236.240 216.995 2236.520 217.275 ;
        RECT 2241.360 217.020 2241.530 217.210 ;
        RECT 2199.835 216.150 2200.265 216.935 ;
        RECT 2205.815 216.150 2206.245 216.935 ;
        RECT 2235.715 216.150 2236.145 216.935 ;
        RECT 2236.545 216.110 2241.675 217.020 ;
        RECT 2242.220 216.995 2242.500 217.275 ;
        RECT 2247.340 217.020 2247.510 217.210 ;
        RECT 2241.695 216.150 2242.125 216.935 ;
        RECT 2242.525 216.110 2247.655 217.020 ;
        RECT 2248.200 216.995 2248.480 217.275 ;
        RECT 2253.320 217.020 2253.490 217.210 ;
        RECT 2247.675 216.150 2248.105 216.935 ;
        RECT 2248.505 216.110 2253.635 217.020 ;
        RECT 2254.180 216.995 2254.460 217.275 ;
        RECT 2259.300 217.020 2259.470 217.210 ;
        RECT 2253.655 216.150 2254.085 216.935 ;
        RECT 2254.485 216.110 2259.615 217.020 ;
        RECT 2260.160 216.995 2260.440 217.275 ;
        RECT 2265.280 217.020 2265.450 217.210 ;
        RECT 2259.635 216.150 2260.065 216.935 ;
        RECT 2260.465 216.110 2265.595 217.020 ;
        RECT 2266.140 216.995 2266.420 217.275 ;
        RECT 2271.260 217.020 2271.430 217.210 ;
        RECT 2265.615 216.150 2266.045 216.935 ;
        RECT 2266.445 216.110 2271.575 217.020 ;
        RECT 2271.595 216.150 2272.025 216.935 ;
      LAYER nwell ;
        RECT 668.810 212.990 729.450 215.820 ;
        RECT 758.510 212.990 795.230 215.820 ;
        RECT 2145.810 212.990 2206.450 215.820 ;
        RECT 2235.510 212.990 2272.230 215.820 ;
      LAYER pwell ;
        RECT 669.015 211.875 669.445 212.660 ;
        RECT 674.995 211.875 675.425 212.660 ;
        RECT 669.540 211.555 669.820 211.835 ;
        RECT 675.445 211.790 680.575 212.700 ;
        RECT 680.975 211.875 681.405 212.660 ;
        RECT 681.425 211.790 686.555 212.700 ;
        RECT 686.955 211.875 687.385 212.660 ;
        RECT 687.405 211.790 692.535 212.700 ;
        RECT 692.935 211.875 693.365 212.660 ;
        RECT 693.385 211.790 698.515 212.700 ;
        RECT 698.915 211.875 699.345 212.660 ;
        RECT 699.365 211.790 704.495 212.700 ;
        RECT 704.895 211.875 705.325 212.660 ;
        RECT 705.345 211.790 710.475 212.700 ;
        RECT 710.875 211.875 711.305 212.660 ;
        RECT 711.325 211.790 716.455 212.700 ;
        RECT 716.855 211.875 717.285 212.660 ;
        RECT 717.305 211.790 722.435 212.700 ;
        RECT 722.835 211.875 723.265 212.660 ;
        RECT 723.285 211.790 728.415 212.700 ;
        RECT 728.815 211.875 729.245 212.660 ;
        RECT 758.715 211.875 759.145 212.660 ;
        RECT 764.695 211.875 765.125 212.660 ;
        RECT 675.590 211.600 675.760 211.790 ;
        RECT 681.570 211.600 681.740 211.790 ;
        RECT 687.550 211.600 687.720 211.790 ;
        RECT 693.530 211.600 693.700 211.790 ;
        RECT 699.510 211.600 699.680 211.790 ;
        RECT 705.490 211.600 705.660 211.790 ;
        RECT 711.470 211.600 711.640 211.790 ;
        RECT 717.450 211.600 717.620 211.790 ;
        RECT 723.430 211.600 723.600 211.790 ;
        RECT 759.240 211.555 759.520 211.835 ;
        RECT 765.145 211.790 770.275 212.700 ;
        RECT 770.675 211.875 771.105 212.660 ;
        RECT 771.125 211.790 776.255 212.700 ;
        RECT 776.655 211.875 777.085 212.660 ;
        RECT 777.105 211.790 782.235 212.700 ;
        RECT 782.635 211.875 783.065 212.660 ;
        RECT 783.085 211.790 788.215 212.700 ;
        RECT 788.615 211.875 789.045 212.660 ;
        RECT 789.445 211.790 794.575 212.700 ;
        RECT 794.595 211.875 795.025 212.660 ;
        RECT 2146.015 211.875 2146.445 212.660 ;
        RECT 2151.995 211.875 2152.425 212.660 ;
        RECT 765.290 211.600 765.460 211.790 ;
        RECT 771.270 211.600 771.440 211.790 ;
        RECT 777.250 211.600 777.420 211.790 ;
        RECT 783.230 211.600 783.400 211.790 ;
        RECT 794.260 211.600 794.430 211.790 ;
        RECT 2146.540 211.555 2146.820 211.835 ;
        RECT 2152.445 211.790 2157.575 212.700 ;
        RECT 2157.975 211.875 2158.405 212.660 ;
        RECT 2158.425 211.790 2163.555 212.700 ;
        RECT 2163.955 211.875 2164.385 212.660 ;
        RECT 2164.405 211.790 2169.535 212.700 ;
        RECT 2169.935 211.875 2170.365 212.660 ;
        RECT 2170.385 211.790 2175.515 212.700 ;
        RECT 2175.915 211.875 2176.345 212.660 ;
        RECT 2176.365 211.790 2181.495 212.700 ;
        RECT 2181.895 211.875 2182.325 212.660 ;
        RECT 2182.345 211.790 2187.475 212.700 ;
        RECT 2187.875 211.875 2188.305 212.660 ;
        RECT 2188.325 211.790 2193.455 212.700 ;
        RECT 2193.855 211.875 2194.285 212.660 ;
        RECT 2194.305 211.790 2199.435 212.700 ;
        RECT 2199.835 211.875 2200.265 212.660 ;
        RECT 2200.285 211.790 2205.415 212.700 ;
        RECT 2205.815 211.875 2206.245 212.660 ;
        RECT 2235.715 211.875 2236.145 212.660 ;
        RECT 2241.695 211.875 2242.125 212.660 ;
        RECT 2152.590 211.600 2152.760 211.790 ;
        RECT 2158.570 211.600 2158.740 211.790 ;
        RECT 2164.550 211.600 2164.720 211.790 ;
        RECT 2170.530 211.600 2170.700 211.790 ;
        RECT 2176.510 211.600 2176.680 211.790 ;
        RECT 2182.490 211.600 2182.660 211.790 ;
        RECT 2188.470 211.600 2188.640 211.790 ;
        RECT 2194.450 211.600 2194.620 211.790 ;
        RECT 2200.430 211.600 2200.600 211.790 ;
        RECT 2236.240 211.555 2236.520 211.835 ;
        RECT 2242.145 211.790 2247.275 212.700 ;
        RECT 2247.675 211.875 2248.105 212.660 ;
        RECT 2248.125 211.790 2253.255 212.700 ;
        RECT 2253.655 211.875 2254.085 212.660 ;
        RECT 2254.105 211.790 2259.235 212.700 ;
        RECT 2259.635 211.875 2260.065 212.660 ;
        RECT 2260.085 211.790 2265.215 212.700 ;
        RECT 2265.615 211.875 2266.045 212.660 ;
        RECT 2266.445 211.790 2271.575 212.700 ;
        RECT 2271.595 211.875 2272.025 212.660 ;
        RECT 2242.290 211.600 2242.460 211.790 ;
        RECT 2248.270 211.600 2248.440 211.790 ;
        RECT 2254.250 211.600 2254.420 211.790 ;
        RECT 2260.230 211.600 2260.400 211.790 ;
        RECT 2271.260 211.600 2271.430 211.790 ;
      LAYER li1 ;
        RECT 3377.780 3608.415 3377.950 3608.500 ;
        RECT 3380.500 3608.415 3380.670 3608.500 ;
        RECT 3383.220 3608.415 3383.390 3608.500 ;
        RECT 3385.940 3608.415 3386.110 3608.500 ;
        RECT 3377.780 3608.355 3379.115 3608.415 ;
        RECT 3377.950 3608.185 3379.115 3608.355 ;
        RECT 3377.780 3608.125 3379.115 3608.185 ;
        RECT 3379.775 3608.355 3381.395 3608.415 ;
        RECT 3379.775 3608.185 3380.500 3608.355 ;
        RECT 3380.670 3608.185 3381.395 3608.355 ;
        RECT 3379.775 3608.125 3381.395 3608.185 ;
        RECT 3382.055 3608.355 3384.555 3608.415 ;
        RECT 3382.055 3608.185 3383.220 3608.355 ;
        RECT 3383.390 3608.185 3384.555 3608.355 ;
        RECT 3382.055 3608.125 3384.555 3608.185 ;
        RECT 3385.215 3608.355 3386.110 3608.415 ;
        RECT 3385.215 3608.185 3385.940 3608.355 ;
        RECT 3385.215 3608.125 3386.110 3608.185 ;
        RECT 3377.780 3608.040 3377.950 3608.125 ;
      LAYER li1 ;
        RECT 3379.955 3606.370 3380.500 3607.955 ;
      LAYER li1 ;
        RECT 3380.500 3607.895 3380.670 3608.125 ;
        RECT 3380.500 3607.525 3380.670 3607.725 ;
        RECT 3380.840 3607.695 3381.490 3607.865 ;
        RECT 3380.500 3607.435 3381.150 3607.525 ;
        RECT 3380.670 3607.265 3381.150 3607.435 ;
        RECT 3380.500 3607.195 3381.150 3607.265 ;
        RECT 3380.500 3606.975 3380.670 3607.195 ;
        RECT 3381.320 3607.025 3381.490 3607.695 ;
        RECT 3380.845 3606.855 3381.490 3607.025 ;
        RECT 3380.500 3606.685 3380.670 3606.805 ;
        RECT 3380.500 3606.515 3381.150 3606.685 ;
      LAYER li1 ;
        RECT 3379.125 3606.030 3380.500 3606.370 ;
      LAYER li1 ;
        RECT 3380.670 3606.355 3381.150 3606.515 ;
        RECT 3381.320 3606.620 3381.490 3606.855 ;
        RECT 3382.030 3607.615 3383.050 3607.945 ;
        RECT 3383.220 3607.895 3383.390 3608.125 ;
        RECT 3385.940 3607.895 3386.110 3608.125 ;
        RECT 3382.030 3607.105 3382.200 3607.615 ;
        RECT 3383.220 3607.565 3383.390 3607.725 ;
        RECT 3385.940 3607.565 3386.110 3607.725 ;
        RECT 3383.220 3607.445 3384.540 3607.565 ;
        RECT 3382.420 3607.435 3384.540 3607.445 ;
        RECT 3382.420 3607.275 3383.220 3607.435 ;
        RECT 3383.390 3607.265 3384.540 3607.435 ;
        RECT 3383.220 3607.235 3384.540 3607.265 ;
        RECT 3385.140 3607.435 3386.110 3607.565 ;
        RECT 3385.140 3607.265 3385.940 3607.435 ;
        RECT 3385.140 3607.235 3386.110 3607.265 ;
        RECT 3382.030 3606.775 3383.050 3607.105 ;
        RECT 3383.220 3606.975 3383.390 3607.235 ;
        RECT 3385.940 3606.975 3386.110 3607.235 ;
        RECT 3382.030 3606.620 3382.200 3606.775 ;
        RECT 3381.320 3606.445 3382.200 3606.620 ;
        RECT 3383.220 3606.725 3383.390 3606.805 ;
        RECT 3385.940 3606.725 3386.110 3606.805 ;
        RECT 3383.220 3606.605 3384.190 3606.725 ;
        RECT 3382.420 3606.515 3384.190 3606.605 ;
        RECT 3380.500 3606.055 3380.670 3606.345 ;
      LAYER li1 ;
        RECT 3379.955 3602.610 3380.500 3606.030 ;
        RECT 3380.840 3606.015 3381.490 3606.185 ;
      LAYER li1 ;
        RECT 3380.500 3605.845 3380.670 3605.885 ;
        RECT 3380.500 3605.595 3381.150 3605.845 ;
        RECT 3380.670 3605.515 3381.150 3605.595 ;
        RECT 3380.500 3605.135 3380.670 3605.425 ;
      LAYER li1 ;
        RECT 3381.320 3605.345 3381.490 3606.015 ;
        RECT 3380.840 3605.175 3381.490 3605.345 ;
      LAYER li1 ;
        RECT 3380.670 3604.965 3381.150 3605.005 ;
        RECT 3380.500 3604.675 3381.150 3604.965 ;
      LAYER li1 ;
        RECT 3381.320 3604.505 3381.490 3605.175 ;
      LAYER li1 ;
        RECT 3380.500 3604.215 3380.670 3604.505 ;
      LAYER li1 ;
        RECT 3380.840 3604.335 3381.490 3604.505 ;
      LAYER li1 ;
        RECT 3380.670 3604.045 3381.150 3604.165 ;
        RECT 3380.500 3603.835 3381.150 3604.045 ;
        RECT 3380.500 3603.755 3380.670 3603.835 ;
      LAYER li1 ;
        RECT 3381.320 3603.750 3381.490 3604.335 ;
      LAYER li1 ;
        RECT 3381.660 3603.995 3381.830 3606.445 ;
        RECT 3382.420 3606.435 3383.220 3606.515 ;
        RECT 3383.390 3606.395 3384.190 3606.515 ;
      LAYER li1 ;
        RECT 3382.030 3606.015 3383.050 3606.185 ;
      LAYER li1 ;
        RECT 3383.220 3606.055 3383.390 3606.345 ;
      LAYER li1 ;
        RECT 3382.030 3605.345 3382.200 3606.015 ;
      LAYER li1 ;
        RECT 3383.220 3605.845 3384.190 3605.885 ;
        RECT 3382.420 3605.595 3384.190 3605.845 ;
        RECT 3382.420 3605.515 3383.220 3605.595 ;
        RECT 3383.390 3605.555 3384.190 3605.595 ;
      LAYER li1 ;
        RECT 3382.030 3605.175 3383.050 3605.345 ;
        RECT 3382.030 3604.505 3382.200 3605.175 ;
      LAYER li1 ;
        RECT 3383.220 3605.135 3383.390 3605.425 ;
        RECT 3382.420 3604.965 3383.220 3605.005 ;
        RECT 3383.390 3604.965 3384.190 3605.045 ;
        RECT 3382.420 3604.715 3384.190 3604.965 ;
        RECT 3382.420 3604.675 3383.390 3604.715 ;
      LAYER li1 ;
        RECT 3382.030 3604.335 3383.050 3604.505 ;
        RECT 3382.030 3603.750 3382.200 3604.335 ;
      LAYER li1 ;
        RECT 3383.220 3604.215 3383.390 3604.505 ;
        RECT 3382.420 3604.045 3383.220 3604.165 ;
        RECT 3383.390 3604.045 3384.190 3604.125 ;
        RECT 3384.780 3604.115 3384.950 3606.565 ;
        RECT 3385.460 3606.515 3386.110 3606.725 ;
        RECT 3385.460 3606.395 3385.940 3606.515 ;
        RECT 3385.940 3606.055 3386.110 3606.345 ;
        RECT 3385.460 3605.595 3386.110 3605.885 ;
        RECT 3385.460 3605.555 3385.940 3605.595 ;
        RECT 3385.940 3605.135 3386.110 3605.425 ;
        RECT 3385.460 3604.965 3385.940 3605.045 ;
        RECT 3385.460 3604.715 3386.110 3604.965 ;
        RECT 3385.940 3604.675 3386.110 3604.715 ;
        RECT 3385.940 3604.215 3386.110 3604.505 ;
        RECT 3382.420 3603.955 3384.190 3604.045 ;
        RECT 3382.420 3603.835 3383.390 3603.955 ;
        RECT 3383.220 3603.755 3383.390 3603.835 ;
        RECT 3384.410 3603.940 3385.290 3604.115 ;
        RECT 3384.410 3603.785 3384.580 3603.940 ;
      LAYER li1 ;
        RECT 3381.320 3603.665 3382.200 3603.750 ;
      LAYER li1 ;
        RECT 3380.500 3603.325 3380.670 3603.585 ;
      LAYER li1 ;
        RECT 3380.840 3603.495 3383.050 3603.665 ;
      LAYER li1 ;
        RECT 3383.220 3603.325 3383.390 3603.585 ;
        RECT 3383.560 3603.455 3384.580 3603.785 ;
        RECT 3380.500 3603.295 3381.470 3603.325 ;
        RECT 3380.670 3603.125 3381.470 3603.295 ;
        RECT 3380.500 3602.995 3381.470 3603.125 ;
        RECT 3382.070 3603.295 3383.390 3603.325 ;
        RECT 3382.070 3603.125 3383.220 3603.295 ;
        RECT 3383.390 3603.125 3384.190 3603.285 ;
        RECT 3382.070 3603.115 3384.190 3603.125 ;
        RECT 3382.070 3602.995 3383.390 3603.115 ;
        RECT 3380.500 3602.835 3380.670 3602.995 ;
        RECT 3383.220 3602.835 3383.390 3602.995 ;
        RECT 3384.410 3602.945 3384.580 3603.455 ;
        RECT 3377.780 3602.435 3377.950 3602.520 ;
        RECT 3380.500 3602.435 3380.670 3602.665 ;
        RECT 3383.220 3602.435 3383.390 3602.665 ;
        RECT 3383.560 3602.615 3384.580 3602.945 ;
      LAYER li1 ;
        RECT 3384.750 3602.660 3384.950 3603.760 ;
      LAYER li1 ;
        RECT 3385.120 3603.705 3385.290 3603.940 ;
        RECT 3385.460 3604.045 3385.940 3604.205 ;
        RECT 3385.460 3603.875 3386.110 3604.045 ;
        RECT 3385.940 3603.755 3386.110 3603.875 ;
        RECT 3385.120 3603.535 3385.765 3603.705 ;
        RECT 3385.120 3602.865 3385.290 3603.535 ;
        RECT 3385.940 3603.365 3386.110 3603.585 ;
        RECT 3385.460 3603.295 3386.110 3603.365 ;
        RECT 3385.460 3603.125 3385.940 3603.295 ;
        RECT 3385.460 3603.035 3386.110 3603.125 ;
        RECT 3385.120 3602.695 3385.770 3602.865 ;
        RECT 3385.940 3602.835 3386.110 3603.035 ;
        RECT 3385.940 3602.435 3386.110 3602.665 ;
        RECT 3377.780 3602.375 3379.115 3602.435 ;
        RECT 3377.950 3602.205 3379.115 3602.375 ;
        RECT 3377.780 3602.145 3379.115 3602.205 ;
        RECT 3379.775 3602.375 3381.395 3602.435 ;
        RECT 3379.775 3602.205 3380.500 3602.375 ;
        RECT 3380.670 3602.205 3381.395 3602.375 ;
        RECT 3379.775 3602.145 3381.395 3602.205 ;
        RECT 3382.055 3602.375 3384.555 3602.435 ;
        RECT 3382.055 3602.205 3383.220 3602.375 ;
        RECT 3383.390 3602.205 3384.555 3602.375 ;
        RECT 3382.055 3602.145 3384.555 3602.205 ;
        RECT 3385.215 3602.375 3386.110 3602.435 ;
        RECT 3385.215 3602.205 3385.940 3602.375 ;
        RECT 3385.215 3602.145 3386.110 3602.205 ;
        RECT 3377.780 3602.060 3377.950 3602.145 ;
        RECT 3380.500 3602.060 3380.670 3602.145 ;
        RECT 3383.220 3602.060 3383.390 3602.145 ;
        RECT 3385.940 3602.060 3386.110 3602.145 ;
        RECT 201.885 3015.005 202.055 3015.090 ;
        RECT 204.605 3015.005 204.775 3015.090 ;
        RECT 207.325 3015.005 207.495 3015.090 ;
        RECT 210.045 3015.005 210.215 3015.090 ;
        RECT 201.885 3014.945 202.780 3015.005 ;
        RECT 202.055 3014.775 202.780 3014.945 ;
        RECT 201.885 3014.715 202.780 3014.775 ;
        RECT 203.440 3014.945 205.940 3015.005 ;
        RECT 203.440 3014.775 204.605 3014.945 ;
        RECT 204.775 3014.775 205.940 3014.945 ;
        RECT 203.440 3014.715 205.940 3014.775 ;
        RECT 206.600 3014.945 208.220 3015.005 ;
        RECT 206.600 3014.775 207.325 3014.945 ;
        RECT 207.495 3014.775 208.220 3014.945 ;
        RECT 206.600 3014.715 208.220 3014.775 ;
        RECT 208.880 3014.945 210.215 3015.005 ;
        RECT 208.880 3014.775 210.045 3014.945 ;
        RECT 208.880 3014.715 210.215 3014.775 ;
        RECT 201.885 3014.485 202.055 3014.715 ;
        RECT 204.605 3014.485 204.775 3014.715 ;
        RECT 201.885 3014.155 202.055 3014.315 ;
        RECT 204.605 3014.155 204.775 3014.315 ;
        RECT 204.945 3014.205 205.965 3014.535 ;
        RECT 207.325 3014.485 207.495 3014.715 ;
        RECT 210.045 3014.630 210.215 3014.715 ;
        RECT 201.885 3014.025 202.855 3014.155 ;
        RECT 202.055 3013.855 202.855 3014.025 ;
        RECT 201.885 3013.825 202.855 3013.855 ;
        RECT 203.455 3014.035 204.775 3014.155 ;
        RECT 203.455 3014.025 205.575 3014.035 ;
        RECT 203.455 3013.855 204.605 3014.025 ;
        RECT 204.775 3013.865 205.575 3014.025 ;
        RECT 203.455 3013.825 204.775 3013.855 ;
        RECT 201.885 3013.565 202.055 3013.825 ;
        RECT 204.605 3013.565 204.775 3013.825 ;
        RECT 205.795 3013.695 205.965 3014.205 ;
        RECT 201.885 3013.315 202.055 3013.395 ;
        RECT 204.605 3013.315 204.775 3013.395 ;
        RECT 204.945 3013.365 205.965 3013.695 ;
        RECT 201.885 3013.105 202.535 3013.315 ;
        RECT 203.805 3013.195 204.775 3013.315 ;
        RECT 205.795 3013.210 205.965 3013.365 ;
        RECT 206.505 3014.285 207.155 3014.455 ;
        RECT 206.505 3013.615 206.675 3014.285 ;
        RECT 207.325 3014.115 207.495 3014.315 ;
        RECT 206.845 3014.025 207.495 3014.115 ;
        RECT 206.845 3013.855 207.325 3014.025 ;
        RECT 206.845 3013.785 207.495 3013.855 ;
        RECT 206.505 3013.445 207.150 3013.615 ;
        RECT 207.325 3013.565 207.495 3013.785 ;
        RECT 206.505 3013.210 206.675 3013.445 ;
        RECT 207.325 3013.275 207.495 3013.395 ;
        RECT 202.055 3012.985 202.535 3013.105 ;
        RECT 201.885 3012.645 202.055 3012.935 ;
        RECT 201.885 3012.185 202.535 3012.475 ;
        RECT 202.055 3012.145 202.535 3012.185 ;
        RECT 201.885 3011.725 202.055 3012.015 ;
        RECT 202.055 3011.555 202.535 3011.635 ;
        RECT 201.885 3011.305 202.535 3011.555 ;
        RECT 201.885 3011.265 202.055 3011.305 ;
        RECT 201.885 3010.805 202.055 3011.095 ;
        RECT 202.055 3010.635 202.535 3010.795 ;
        RECT 203.045 3010.705 203.215 3013.155 ;
        RECT 203.805 3013.105 205.575 3013.195 ;
        RECT 203.805 3012.985 204.605 3013.105 ;
        RECT 204.775 3013.025 205.575 3013.105 ;
        RECT 205.795 3013.035 206.675 3013.210 ;
        RECT 206.845 3013.105 207.495 3013.275 ;
        RECT 204.605 3012.645 204.775 3012.935 ;
      LAYER li1 ;
        RECT 204.945 3012.605 205.965 3012.775 ;
      LAYER li1 ;
        RECT 203.805 3012.435 204.775 3012.475 ;
        RECT 203.805 3012.185 205.575 3012.435 ;
        RECT 203.805 3012.145 204.605 3012.185 ;
        RECT 204.775 3012.105 205.575 3012.185 ;
        RECT 204.605 3011.725 204.775 3012.015 ;
      LAYER li1 ;
        RECT 205.795 3011.935 205.965 3012.605 ;
        RECT 204.945 3011.765 205.965 3011.935 ;
      LAYER li1 ;
        RECT 203.805 3011.555 204.605 3011.635 ;
        RECT 204.775 3011.555 205.575 3011.595 ;
        RECT 203.805 3011.305 205.575 3011.555 ;
        RECT 204.605 3011.265 205.575 3011.305 ;
      LAYER li1 ;
        RECT 205.795 3011.095 205.965 3011.765 ;
      LAYER li1 ;
        RECT 204.605 3010.805 204.775 3011.095 ;
      LAYER li1 ;
        RECT 204.945 3010.925 205.965 3011.095 ;
      LAYER li1 ;
        RECT 201.885 3010.465 202.535 3010.635 ;
        RECT 202.705 3010.530 203.585 3010.705 ;
        RECT 203.805 3010.635 204.605 3010.715 ;
        RECT 204.775 3010.635 205.575 3010.755 ;
        RECT 203.805 3010.545 205.575 3010.635 ;
        RECT 201.885 3010.345 202.055 3010.465 ;
        RECT 202.705 3010.295 202.875 3010.530 ;
        RECT 203.415 3010.375 203.585 3010.530 ;
        RECT 204.605 3010.425 205.575 3010.545 ;
        RECT 201.885 3009.955 202.055 3010.175 ;
        RECT 202.230 3010.125 202.875 3010.295 ;
        RECT 201.885 3009.885 202.535 3009.955 ;
        RECT 202.055 3009.715 202.535 3009.885 ;
        RECT 201.885 3009.625 202.535 3009.715 ;
        RECT 201.885 3009.425 202.055 3009.625 ;
        RECT 202.705 3009.455 202.875 3010.125 ;
        RECT 202.225 3009.285 202.875 3009.455 ;
        RECT 201.885 3009.025 202.055 3009.255 ;
      LAYER li1 ;
        RECT 203.045 3009.250 203.245 3010.350 ;
      LAYER li1 ;
        RECT 203.415 3010.045 204.435 3010.375 ;
        RECT 204.605 3010.345 204.775 3010.425 ;
      LAYER li1 ;
        RECT 205.795 3010.340 205.965 3010.925 ;
      LAYER li1 ;
        RECT 206.165 3010.585 206.335 3013.035 ;
        RECT 206.845 3012.945 207.325 3013.105 ;
      LAYER li1 ;
        RECT 207.495 3012.960 208.040 3014.545 ;
        RECT 206.505 3012.605 207.155 3012.775 ;
      LAYER li1 ;
        RECT 207.325 3012.645 207.495 3012.935 ;
      LAYER li1 ;
        RECT 207.495 3012.620 208.870 3012.960 ;
        RECT 206.505 3011.935 206.675 3012.605 ;
      LAYER li1 ;
        RECT 207.325 3012.435 207.495 3012.475 ;
        RECT 206.845 3012.185 207.495 3012.435 ;
        RECT 206.845 3012.105 207.325 3012.185 ;
      LAYER li1 ;
        RECT 206.505 3011.765 207.155 3011.935 ;
        RECT 206.505 3011.095 206.675 3011.765 ;
      LAYER li1 ;
        RECT 207.325 3011.725 207.495 3012.015 ;
        RECT 206.845 3011.555 207.325 3011.595 ;
        RECT 206.845 3011.265 207.495 3011.555 ;
      LAYER li1 ;
        RECT 206.505 3010.925 207.155 3011.095 ;
        RECT 206.505 3010.340 206.675 3010.925 ;
      LAYER li1 ;
        RECT 207.325 3010.805 207.495 3011.095 ;
        RECT 206.845 3010.635 207.325 3010.755 ;
        RECT 206.845 3010.425 207.495 3010.635 ;
        RECT 207.325 3010.345 207.495 3010.425 ;
      LAYER li1 ;
        RECT 205.795 3010.255 206.675 3010.340 ;
      LAYER li1 ;
        RECT 203.415 3009.535 203.585 3010.045 ;
        RECT 204.605 3009.915 204.775 3010.175 ;
      LAYER li1 ;
        RECT 204.945 3010.085 207.155 3010.255 ;
      LAYER li1 ;
        RECT 207.325 3009.915 207.495 3010.175 ;
        RECT 204.605 3009.885 205.925 3009.915 ;
        RECT 203.805 3009.715 204.605 3009.875 ;
        RECT 204.775 3009.715 205.925 3009.885 ;
        RECT 203.805 3009.705 205.925 3009.715 ;
        RECT 204.605 3009.585 205.925 3009.705 ;
        RECT 206.525 3009.885 207.495 3009.915 ;
        RECT 206.525 3009.715 207.325 3009.885 ;
        RECT 206.525 3009.585 207.495 3009.715 ;
        RECT 203.415 3009.205 204.435 3009.535 ;
        RECT 204.605 3009.425 204.775 3009.585 ;
        RECT 207.325 3009.425 207.495 3009.585 ;
        RECT 204.605 3009.025 204.775 3009.255 ;
        RECT 207.325 3009.025 207.495 3009.255 ;
      LAYER li1 ;
        RECT 207.495 3009.200 208.040 3012.620 ;
      LAYER li1 ;
        RECT 210.045 3009.025 210.215 3009.110 ;
        RECT 201.885 3008.965 202.780 3009.025 ;
        RECT 202.055 3008.795 202.780 3008.965 ;
        RECT 201.885 3008.735 202.780 3008.795 ;
        RECT 203.440 3008.965 205.940 3009.025 ;
        RECT 203.440 3008.795 204.605 3008.965 ;
        RECT 204.775 3008.795 205.940 3008.965 ;
        RECT 203.440 3008.735 205.940 3008.795 ;
        RECT 206.600 3008.965 208.220 3009.025 ;
        RECT 206.600 3008.795 207.325 3008.965 ;
        RECT 207.495 3008.795 208.220 3008.965 ;
        RECT 206.600 3008.735 208.220 3008.795 ;
        RECT 208.880 3008.965 210.215 3009.025 ;
        RECT 208.880 3008.795 210.045 3008.965 ;
        RECT 208.880 3008.735 210.215 3008.795 ;
        RECT 201.885 3008.505 202.055 3008.735 ;
        RECT 204.605 3008.505 204.775 3008.735 ;
        RECT 201.885 3008.175 202.055 3008.335 ;
        RECT 204.605 3008.175 204.775 3008.335 ;
        RECT 204.945 3008.225 205.965 3008.555 ;
        RECT 207.325 3008.505 207.495 3008.735 ;
        RECT 210.045 3008.650 210.215 3008.735 ;
        RECT 201.885 3008.045 202.855 3008.175 ;
        RECT 202.055 3007.875 202.855 3008.045 ;
        RECT 201.885 3007.845 202.855 3007.875 ;
        RECT 203.455 3008.055 204.775 3008.175 ;
        RECT 203.455 3008.045 205.575 3008.055 ;
        RECT 203.455 3007.875 204.605 3008.045 ;
        RECT 204.775 3007.885 205.575 3008.045 ;
        RECT 203.455 3007.845 204.775 3007.875 ;
        RECT 201.885 3007.585 202.055 3007.845 ;
        RECT 204.605 3007.585 204.775 3007.845 ;
        RECT 205.795 3007.715 205.965 3008.225 ;
        RECT 201.885 3007.335 202.055 3007.415 ;
        RECT 204.605 3007.335 204.775 3007.415 ;
        RECT 204.945 3007.385 205.965 3007.715 ;
        RECT 201.885 3007.125 202.535 3007.335 ;
        RECT 203.805 3007.215 204.775 3007.335 ;
        RECT 205.795 3007.230 205.965 3007.385 ;
        RECT 206.505 3008.305 207.155 3008.475 ;
        RECT 206.505 3007.635 206.675 3008.305 ;
        RECT 207.325 3008.135 207.495 3008.335 ;
        RECT 206.845 3008.045 207.495 3008.135 ;
        RECT 206.845 3007.875 207.325 3008.045 ;
        RECT 206.845 3007.805 207.495 3007.875 ;
        RECT 206.505 3007.465 207.150 3007.635 ;
        RECT 207.325 3007.585 207.495 3007.805 ;
        RECT 206.505 3007.230 206.675 3007.465 ;
        RECT 207.325 3007.295 207.495 3007.415 ;
        RECT 202.055 3007.005 202.535 3007.125 ;
        RECT 201.885 3006.665 202.055 3006.955 ;
        RECT 201.885 3006.205 202.535 3006.495 ;
        RECT 202.055 3006.165 202.535 3006.205 ;
        RECT 201.885 3005.745 202.055 3006.035 ;
        RECT 202.055 3005.575 202.535 3005.655 ;
        RECT 201.885 3005.325 202.535 3005.575 ;
        RECT 201.885 3005.285 202.055 3005.325 ;
        RECT 201.885 3004.825 202.055 3005.115 ;
        RECT 202.055 3004.655 202.535 3004.815 ;
        RECT 203.045 3004.725 203.215 3007.175 ;
        RECT 203.805 3007.125 205.575 3007.215 ;
        RECT 203.805 3007.005 204.605 3007.125 ;
        RECT 204.775 3007.045 205.575 3007.125 ;
        RECT 205.795 3007.055 206.675 3007.230 ;
        RECT 206.845 3007.125 207.495 3007.295 ;
        RECT 204.605 3006.665 204.775 3006.955 ;
      LAYER li1 ;
        RECT 204.945 3006.625 205.965 3006.795 ;
      LAYER li1 ;
        RECT 203.805 3006.455 204.775 3006.495 ;
        RECT 203.805 3006.205 205.575 3006.455 ;
        RECT 203.805 3006.165 204.605 3006.205 ;
        RECT 204.775 3006.125 205.575 3006.205 ;
        RECT 204.605 3005.745 204.775 3006.035 ;
      LAYER li1 ;
        RECT 205.795 3005.955 205.965 3006.625 ;
        RECT 204.945 3005.785 205.965 3005.955 ;
      LAYER li1 ;
        RECT 203.805 3005.575 204.605 3005.655 ;
        RECT 204.775 3005.575 205.575 3005.615 ;
        RECT 203.805 3005.325 205.575 3005.575 ;
        RECT 204.605 3005.285 205.575 3005.325 ;
      LAYER li1 ;
        RECT 205.795 3005.115 205.965 3005.785 ;
      LAYER li1 ;
        RECT 204.605 3004.825 204.775 3005.115 ;
      LAYER li1 ;
        RECT 204.945 3004.945 205.965 3005.115 ;
      LAYER li1 ;
        RECT 201.885 3004.485 202.535 3004.655 ;
        RECT 202.705 3004.550 203.585 3004.725 ;
        RECT 203.805 3004.655 204.605 3004.735 ;
        RECT 204.775 3004.655 205.575 3004.775 ;
        RECT 203.805 3004.565 205.575 3004.655 ;
        RECT 201.885 3004.365 202.055 3004.485 ;
        RECT 202.705 3004.315 202.875 3004.550 ;
        RECT 203.415 3004.395 203.585 3004.550 ;
        RECT 204.605 3004.445 205.575 3004.565 ;
        RECT 201.885 3003.975 202.055 3004.195 ;
        RECT 202.230 3004.145 202.875 3004.315 ;
        RECT 201.885 3003.905 202.535 3003.975 ;
        RECT 202.055 3003.735 202.535 3003.905 ;
        RECT 201.885 3003.645 202.535 3003.735 ;
        RECT 201.885 3003.445 202.055 3003.645 ;
        RECT 202.705 3003.475 202.875 3004.145 ;
        RECT 202.225 3003.305 202.875 3003.475 ;
        RECT 201.885 3003.045 202.055 3003.275 ;
      LAYER li1 ;
        RECT 203.045 3003.270 203.245 3004.370 ;
      LAYER li1 ;
        RECT 203.415 3004.065 204.435 3004.395 ;
        RECT 204.605 3004.365 204.775 3004.445 ;
      LAYER li1 ;
        RECT 205.795 3004.360 205.965 3004.945 ;
      LAYER li1 ;
        RECT 206.165 3004.605 206.335 3007.055 ;
        RECT 206.845 3006.965 207.325 3007.125 ;
      LAYER li1 ;
        RECT 207.495 3006.980 208.040 3008.565 ;
        RECT 206.505 3006.625 207.155 3006.795 ;
      LAYER li1 ;
        RECT 207.325 3006.665 207.495 3006.955 ;
      LAYER li1 ;
        RECT 207.495 3006.640 208.870 3006.980 ;
        RECT 206.505 3005.955 206.675 3006.625 ;
      LAYER li1 ;
        RECT 207.325 3006.455 207.495 3006.495 ;
        RECT 206.845 3006.205 207.495 3006.455 ;
        RECT 206.845 3006.125 207.325 3006.205 ;
      LAYER li1 ;
        RECT 206.505 3005.785 207.155 3005.955 ;
        RECT 206.505 3005.115 206.675 3005.785 ;
      LAYER li1 ;
        RECT 207.325 3005.745 207.495 3006.035 ;
        RECT 206.845 3005.575 207.325 3005.615 ;
        RECT 206.845 3005.285 207.495 3005.575 ;
      LAYER li1 ;
        RECT 206.505 3004.945 207.155 3005.115 ;
        RECT 206.505 3004.360 206.675 3004.945 ;
      LAYER li1 ;
        RECT 207.325 3004.825 207.495 3005.115 ;
        RECT 206.845 3004.655 207.325 3004.775 ;
        RECT 206.845 3004.445 207.495 3004.655 ;
        RECT 207.325 3004.365 207.495 3004.445 ;
      LAYER li1 ;
        RECT 205.795 3004.275 206.675 3004.360 ;
      LAYER li1 ;
        RECT 203.415 3003.555 203.585 3004.065 ;
        RECT 204.605 3003.935 204.775 3004.195 ;
      LAYER li1 ;
        RECT 204.945 3004.105 207.155 3004.275 ;
      LAYER li1 ;
        RECT 207.325 3003.935 207.495 3004.195 ;
        RECT 204.605 3003.905 205.925 3003.935 ;
        RECT 203.805 3003.735 204.605 3003.895 ;
        RECT 204.775 3003.735 205.925 3003.905 ;
        RECT 203.805 3003.725 205.925 3003.735 ;
        RECT 204.605 3003.605 205.925 3003.725 ;
        RECT 206.525 3003.905 207.495 3003.935 ;
        RECT 206.525 3003.735 207.325 3003.905 ;
        RECT 206.525 3003.605 207.495 3003.735 ;
        RECT 203.415 3003.225 204.435 3003.555 ;
        RECT 204.605 3003.445 204.775 3003.605 ;
        RECT 207.325 3003.445 207.495 3003.605 ;
        RECT 204.605 3003.045 204.775 3003.275 ;
        RECT 207.325 3003.045 207.495 3003.275 ;
      LAYER li1 ;
        RECT 207.495 3003.220 208.040 3006.640 ;
      LAYER li1 ;
        RECT 210.045 3003.045 210.215 3003.130 ;
        RECT 201.885 3002.985 202.780 3003.045 ;
        RECT 202.055 3002.815 202.780 3002.985 ;
        RECT 201.885 3002.755 202.780 3002.815 ;
        RECT 203.440 3002.985 205.940 3003.045 ;
        RECT 203.440 3002.815 204.605 3002.985 ;
        RECT 204.775 3002.815 205.940 3002.985 ;
        RECT 203.440 3002.755 205.940 3002.815 ;
        RECT 206.600 3002.985 208.220 3003.045 ;
        RECT 206.600 3002.815 207.325 3002.985 ;
        RECT 207.495 3002.815 208.220 3002.985 ;
        RECT 206.600 3002.755 208.220 3002.815 ;
        RECT 208.880 3002.985 210.215 3003.045 ;
        RECT 208.880 3002.815 210.045 3002.985 ;
        RECT 208.880 3002.755 210.215 3002.815 ;
        RECT 201.885 3002.525 202.055 3002.755 ;
        RECT 204.605 3002.525 204.775 3002.755 ;
        RECT 201.885 3002.195 202.055 3002.355 ;
        RECT 204.605 3002.195 204.775 3002.355 ;
        RECT 204.945 3002.245 205.965 3002.575 ;
        RECT 207.325 3002.525 207.495 3002.755 ;
        RECT 210.045 3002.670 210.215 3002.755 ;
        RECT 201.885 3002.065 202.855 3002.195 ;
        RECT 202.055 3001.895 202.855 3002.065 ;
        RECT 201.885 3001.865 202.855 3001.895 ;
        RECT 203.455 3002.075 204.775 3002.195 ;
        RECT 203.455 3002.065 205.575 3002.075 ;
        RECT 203.455 3001.895 204.605 3002.065 ;
        RECT 204.775 3001.905 205.575 3002.065 ;
        RECT 203.455 3001.865 204.775 3001.895 ;
        RECT 201.885 3001.605 202.055 3001.865 ;
        RECT 204.605 3001.605 204.775 3001.865 ;
        RECT 205.795 3001.735 205.965 3002.245 ;
        RECT 201.885 3001.355 202.055 3001.435 ;
        RECT 204.605 3001.355 204.775 3001.435 ;
        RECT 204.945 3001.405 205.965 3001.735 ;
        RECT 201.885 3001.145 202.535 3001.355 ;
        RECT 203.805 3001.235 204.775 3001.355 ;
        RECT 205.795 3001.250 205.965 3001.405 ;
        RECT 206.505 3002.325 207.155 3002.495 ;
        RECT 206.505 3001.655 206.675 3002.325 ;
        RECT 207.325 3002.155 207.495 3002.355 ;
        RECT 206.845 3002.065 207.495 3002.155 ;
        RECT 206.845 3001.895 207.325 3002.065 ;
        RECT 206.845 3001.825 207.495 3001.895 ;
        RECT 206.505 3001.485 207.150 3001.655 ;
        RECT 207.325 3001.605 207.495 3001.825 ;
        RECT 206.505 3001.250 206.675 3001.485 ;
        RECT 207.325 3001.315 207.495 3001.435 ;
        RECT 202.055 3001.025 202.535 3001.145 ;
        RECT 201.885 3000.685 202.055 3000.975 ;
        RECT 201.885 3000.225 202.535 3000.515 ;
        RECT 202.055 3000.185 202.535 3000.225 ;
        RECT 201.885 2999.765 202.055 3000.055 ;
        RECT 202.055 2999.595 202.535 2999.675 ;
        RECT 201.885 2999.345 202.535 2999.595 ;
        RECT 201.885 2999.305 202.055 2999.345 ;
        RECT 201.885 2998.845 202.055 2999.135 ;
        RECT 202.055 2998.675 202.535 2998.835 ;
        RECT 203.045 2998.745 203.215 3001.195 ;
        RECT 203.805 3001.145 205.575 3001.235 ;
        RECT 203.805 3001.025 204.605 3001.145 ;
        RECT 204.775 3001.065 205.575 3001.145 ;
        RECT 205.795 3001.075 206.675 3001.250 ;
        RECT 206.845 3001.145 207.495 3001.315 ;
        RECT 204.605 3000.685 204.775 3000.975 ;
      LAYER li1 ;
        RECT 204.945 3000.645 205.965 3000.815 ;
      LAYER li1 ;
        RECT 203.805 3000.475 204.775 3000.515 ;
        RECT 203.805 3000.225 205.575 3000.475 ;
        RECT 203.805 3000.185 204.605 3000.225 ;
        RECT 204.775 3000.145 205.575 3000.225 ;
        RECT 204.605 2999.765 204.775 3000.055 ;
      LAYER li1 ;
        RECT 205.795 2999.975 205.965 3000.645 ;
        RECT 204.945 2999.805 205.965 2999.975 ;
      LAYER li1 ;
        RECT 203.805 2999.595 204.605 2999.675 ;
        RECT 204.775 2999.595 205.575 2999.635 ;
        RECT 203.805 2999.345 205.575 2999.595 ;
        RECT 204.605 2999.305 205.575 2999.345 ;
      LAYER li1 ;
        RECT 205.795 2999.135 205.965 2999.805 ;
      LAYER li1 ;
        RECT 204.605 2998.845 204.775 2999.135 ;
      LAYER li1 ;
        RECT 204.945 2998.965 205.965 2999.135 ;
      LAYER li1 ;
        RECT 201.885 2998.505 202.535 2998.675 ;
        RECT 202.705 2998.570 203.585 2998.745 ;
        RECT 203.805 2998.675 204.605 2998.755 ;
        RECT 204.775 2998.675 205.575 2998.795 ;
        RECT 203.805 2998.585 205.575 2998.675 ;
        RECT 201.885 2998.385 202.055 2998.505 ;
        RECT 202.705 2998.335 202.875 2998.570 ;
        RECT 203.415 2998.415 203.585 2998.570 ;
        RECT 204.605 2998.465 205.575 2998.585 ;
        RECT 201.885 2997.995 202.055 2998.215 ;
        RECT 202.230 2998.165 202.875 2998.335 ;
        RECT 201.885 2997.925 202.535 2997.995 ;
        RECT 202.055 2997.755 202.535 2997.925 ;
        RECT 201.885 2997.665 202.535 2997.755 ;
        RECT 201.885 2997.465 202.055 2997.665 ;
        RECT 202.705 2997.495 202.875 2998.165 ;
        RECT 202.225 2997.325 202.875 2997.495 ;
        RECT 201.885 2997.065 202.055 2997.295 ;
      LAYER li1 ;
        RECT 203.045 2997.290 203.245 2998.390 ;
      LAYER li1 ;
        RECT 203.415 2998.085 204.435 2998.415 ;
        RECT 204.605 2998.385 204.775 2998.465 ;
      LAYER li1 ;
        RECT 205.795 2998.380 205.965 2998.965 ;
      LAYER li1 ;
        RECT 206.165 2998.625 206.335 3001.075 ;
        RECT 206.845 3000.985 207.325 3001.145 ;
      LAYER li1 ;
        RECT 207.495 3001.000 208.040 3002.585 ;
        RECT 206.505 3000.645 207.155 3000.815 ;
      LAYER li1 ;
        RECT 207.325 3000.685 207.495 3000.975 ;
      LAYER li1 ;
        RECT 207.495 3000.660 208.870 3001.000 ;
        RECT 206.505 2999.975 206.675 3000.645 ;
      LAYER li1 ;
        RECT 207.325 3000.475 207.495 3000.515 ;
        RECT 206.845 3000.225 207.495 3000.475 ;
        RECT 206.845 3000.145 207.325 3000.225 ;
      LAYER li1 ;
        RECT 206.505 2999.805 207.155 2999.975 ;
        RECT 206.505 2999.135 206.675 2999.805 ;
      LAYER li1 ;
        RECT 207.325 2999.765 207.495 3000.055 ;
        RECT 206.845 2999.595 207.325 2999.635 ;
        RECT 206.845 2999.305 207.495 2999.595 ;
      LAYER li1 ;
        RECT 206.505 2998.965 207.155 2999.135 ;
        RECT 206.505 2998.380 206.675 2998.965 ;
      LAYER li1 ;
        RECT 207.325 2998.845 207.495 2999.135 ;
        RECT 206.845 2998.675 207.325 2998.795 ;
        RECT 206.845 2998.465 207.495 2998.675 ;
        RECT 207.325 2998.385 207.495 2998.465 ;
      LAYER li1 ;
        RECT 205.795 2998.295 206.675 2998.380 ;
      LAYER li1 ;
        RECT 203.415 2997.575 203.585 2998.085 ;
        RECT 204.605 2997.955 204.775 2998.215 ;
      LAYER li1 ;
        RECT 204.945 2998.125 207.155 2998.295 ;
      LAYER li1 ;
        RECT 207.325 2997.955 207.495 2998.215 ;
        RECT 204.605 2997.925 205.925 2997.955 ;
        RECT 203.805 2997.755 204.605 2997.915 ;
        RECT 204.775 2997.755 205.925 2997.925 ;
        RECT 203.805 2997.745 205.925 2997.755 ;
        RECT 204.605 2997.625 205.925 2997.745 ;
        RECT 206.525 2997.925 207.495 2997.955 ;
        RECT 206.525 2997.755 207.325 2997.925 ;
        RECT 206.525 2997.625 207.495 2997.755 ;
        RECT 203.415 2997.245 204.435 2997.575 ;
        RECT 204.605 2997.465 204.775 2997.625 ;
        RECT 207.325 2997.465 207.495 2997.625 ;
        RECT 204.605 2997.065 204.775 2997.295 ;
        RECT 207.325 2997.065 207.495 2997.295 ;
      LAYER li1 ;
        RECT 207.495 2997.240 208.040 3000.660 ;
      LAYER li1 ;
        RECT 210.045 2997.065 210.215 2997.150 ;
        RECT 201.885 2997.005 202.780 2997.065 ;
        RECT 202.055 2996.835 202.780 2997.005 ;
        RECT 201.885 2996.775 202.780 2996.835 ;
        RECT 203.440 2997.005 205.940 2997.065 ;
        RECT 203.440 2996.835 204.605 2997.005 ;
        RECT 204.775 2996.835 205.940 2997.005 ;
        RECT 203.440 2996.775 205.940 2996.835 ;
        RECT 206.600 2997.005 208.220 2997.065 ;
        RECT 206.600 2996.835 207.325 2997.005 ;
        RECT 207.495 2996.835 208.220 2997.005 ;
        RECT 206.600 2996.775 208.220 2996.835 ;
        RECT 208.880 2997.005 210.215 2997.065 ;
        RECT 208.880 2996.835 210.045 2997.005 ;
        RECT 208.880 2996.775 210.215 2996.835 ;
        RECT 201.885 2996.545 202.055 2996.775 ;
        RECT 204.605 2996.545 204.775 2996.775 ;
        RECT 201.885 2996.215 202.055 2996.375 ;
        RECT 204.605 2996.215 204.775 2996.375 ;
        RECT 204.945 2996.265 205.965 2996.595 ;
        RECT 207.325 2996.545 207.495 2996.775 ;
        RECT 210.045 2996.690 210.215 2996.775 ;
        RECT 201.885 2996.085 202.855 2996.215 ;
        RECT 202.055 2995.915 202.855 2996.085 ;
        RECT 201.885 2995.885 202.855 2995.915 ;
        RECT 203.455 2996.095 204.775 2996.215 ;
        RECT 203.455 2996.085 205.575 2996.095 ;
        RECT 203.455 2995.915 204.605 2996.085 ;
        RECT 204.775 2995.925 205.575 2996.085 ;
        RECT 203.455 2995.885 204.775 2995.915 ;
        RECT 201.885 2995.625 202.055 2995.885 ;
        RECT 204.605 2995.625 204.775 2995.885 ;
        RECT 205.795 2995.755 205.965 2996.265 ;
        RECT 201.885 2995.375 202.055 2995.455 ;
        RECT 204.605 2995.375 204.775 2995.455 ;
        RECT 204.945 2995.425 205.965 2995.755 ;
        RECT 201.885 2995.165 202.535 2995.375 ;
        RECT 203.805 2995.255 204.775 2995.375 ;
        RECT 205.795 2995.270 205.965 2995.425 ;
        RECT 206.505 2996.345 207.155 2996.515 ;
        RECT 206.505 2995.675 206.675 2996.345 ;
        RECT 207.325 2996.175 207.495 2996.375 ;
        RECT 206.845 2996.085 207.495 2996.175 ;
        RECT 206.845 2995.915 207.325 2996.085 ;
        RECT 206.845 2995.845 207.495 2995.915 ;
        RECT 206.505 2995.505 207.150 2995.675 ;
        RECT 207.325 2995.625 207.495 2995.845 ;
        RECT 206.505 2995.270 206.675 2995.505 ;
        RECT 207.325 2995.335 207.495 2995.455 ;
        RECT 202.055 2995.045 202.535 2995.165 ;
        RECT 201.885 2994.705 202.055 2994.995 ;
        RECT 201.885 2994.245 202.535 2994.535 ;
        RECT 202.055 2994.205 202.535 2994.245 ;
        RECT 201.885 2993.785 202.055 2994.075 ;
        RECT 202.055 2993.615 202.535 2993.695 ;
        RECT 201.885 2993.365 202.535 2993.615 ;
        RECT 201.885 2993.325 202.055 2993.365 ;
        RECT 201.885 2992.865 202.055 2993.155 ;
        RECT 202.055 2992.695 202.535 2992.855 ;
        RECT 203.045 2992.765 203.215 2995.215 ;
        RECT 203.805 2995.165 205.575 2995.255 ;
        RECT 203.805 2995.045 204.605 2995.165 ;
        RECT 204.775 2995.085 205.575 2995.165 ;
        RECT 205.795 2995.095 206.675 2995.270 ;
        RECT 206.845 2995.165 207.495 2995.335 ;
        RECT 204.605 2994.705 204.775 2994.995 ;
      LAYER li1 ;
        RECT 204.945 2994.665 205.965 2994.835 ;
      LAYER li1 ;
        RECT 203.805 2994.495 204.775 2994.535 ;
        RECT 203.805 2994.245 205.575 2994.495 ;
        RECT 203.805 2994.205 204.605 2994.245 ;
        RECT 204.775 2994.165 205.575 2994.245 ;
        RECT 204.605 2993.785 204.775 2994.075 ;
      LAYER li1 ;
        RECT 205.795 2993.995 205.965 2994.665 ;
        RECT 204.945 2993.825 205.965 2993.995 ;
      LAYER li1 ;
        RECT 203.805 2993.615 204.605 2993.695 ;
        RECT 204.775 2993.615 205.575 2993.655 ;
        RECT 203.805 2993.365 205.575 2993.615 ;
        RECT 204.605 2993.325 205.575 2993.365 ;
      LAYER li1 ;
        RECT 205.795 2993.155 205.965 2993.825 ;
      LAYER li1 ;
        RECT 204.605 2992.865 204.775 2993.155 ;
      LAYER li1 ;
        RECT 204.945 2992.985 205.965 2993.155 ;
      LAYER li1 ;
        RECT 201.885 2992.525 202.535 2992.695 ;
        RECT 202.705 2992.590 203.585 2992.765 ;
        RECT 203.805 2992.695 204.605 2992.775 ;
        RECT 204.775 2992.695 205.575 2992.815 ;
        RECT 203.805 2992.605 205.575 2992.695 ;
        RECT 201.885 2992.405 202.055 2992.525 ;
        RECT 202.705 2992.355 202.875 2992.590 ;
        RECT 203.415 2992.435 203.585 2992.590 ;
        RECT 204.605 2992.485 205.575 2992.605 ;
        RECT 201.885 2992.015 202.055 2992.235 ;
        RECT 202.230 2992.185 202.875 2992.355 ;
        RECT 201.885 2991.945 202.535 2992.015 ;
        RECT 202.055 2991.775 202.535 2991.945 ;
        RECT 201.885 2991.685 202.535 2991.775 ;
        RECT 201.885 2991.485 202.055 2991.685 ;
        RECT 202.705 2991.515 202.875 2992.185 ;
        RECT 202.225 2991.345 202.875 2991.515 ;
        RECT 201.885 2991.085 202.055 2991.315 ;
      LAYER li1 ;
        RECT 203.045 2991.310 203.245 2992.410 ;
      LAYER li1 ;
        RECT 203.415 2992.105 204.435 2992.435 ;
        RECT 204.605 2992.405 204.775 2992.485 ;
      LAYER li1 ;
        RECT 205.795 2992.400 205.965 2992.985 ;
      LAYER li1 ;
        RECT 206.165 2992.645 206.335 2995.095 ;
        RECT 206.845 2995.005 207.325 2995.165 ;
      LAYER li1 ;
        RECT 207.495 2995.020 208.040 2996.605 ;
        RECT 206.505 2994.665 207.155 2994.835 ;
      LAYER li1 ;
        RECT 207.325 2994.705 207.495 2994.995 ;
      LAYER li1 ;
        RECT 207.495 2994.680 208.870 2995.020 ;
        RECT 206.505 2993.995 206.675 2994.665 ;
      LAYER li1 ;
        RECT 207.325 2994.495 207.495 2994.535 ;
        RECT 206.845 2994.245 207.495 2994.495 ;
        RECT 206.845 2994.165 207.325 2994.245 ;
      LAYER li1 ;
        RECT 206.505 2993.825 207.155 2993.995 ;
        RECT 206.505 2993.155 206.675 2993.825 ;
      LAYER li1 ;
        RECT 207.325 2993.785 207.495 2994.075 ;
        RECT 206.845 2993.615 207.325 2993.655 ;
        RECT 206.845 2993.325 207.495 2993.615 ;
      LAYER li1 ;
        RECT 206.505 2992.985 207.155 2993.155 ;
        RECT 206.505 2992.400 206.675 2992.985 ;
      LAYER li1 ;
        RECT 207.325 2992.865 207.495 2993.155 ;
        RECT 206.845 2992.695 207.325 2992.815 ;
        RECT 206.845 2992.485 207.495 2992.695 ;
        RECT 207.325 2992.405 207.495 2992.485 ;
      LAYER li1 ;
        RECT 205.795 2992.315 206.675 2992.400 ;
      LAYER li1 ;
        RECT 203.415 2991.595 203.585 2992.105 ;
        RECT 204.605 2991.975 204.775 2992.235 ;
      LAYER li1 ;
        RECT 204.945 2992.145 207.155 2992.315 ;
      LAYER li1 ;
        RECT 207.325 2991.975 207.495 2992.235 ;
        RECT 204.605 2991.945 205.925 2991.975 ;
        RECT 203.805 2991.775 204.605 2991.935 ;
        RECT 204.775 2991.775 205.925 2991.945 ;
        RECT 203.805 2991.765 205.925 2991.775 ;
        RECT 204.605 2991.645 205.925 2991.765 ;
        RECT 206.525 2991.945 207.495 2991.975 ;
        RECT 206.525 2991.775 207.325 2991.945 ;
        RECT 206.525 2991.645 207.495 2991.775 ;
        RECT 203.415 2991.265 204.435 2991.595 ;
        RECT 204.605 2991.485 204.775 2991.645 ;
        RECT 207.325 2991.485 207.495 2991.645 ;
        RECT 204.605 2991.085 204.775 2991.315 ;
        RECT 207.325 2991.085 207.495 2991.315 ;
      LAYER li1 ;
        RECT 207.495 2991.260 208.040 2994.680 ;
      LAYER li1 ;
        RECT 210.045 2991.085 210.215 2991.170 ;
        RECT 201.885 2991.025 202.780 2991.085 ;
        RECT 202.055 2990.855 202.780 2991.025 ;
        RECT 201.885 2990.795 202.780 2990.855 ;
        RECT 203.440 2991.025 205.940 2991.085 ;
        RECT 203.440 2990.855 204.605 2991.025 ;
        RECT 204.775 2990.855 205.940 2991.025 ;
        RECT 203.440 2990.795 205.940 2990.855 ;
        RECT 206.600 2991.025 208.220 2991.085 ;
        RECT 206.600 2990.855 207.325 2991.025 ;
        RECT 207.495 2990.855 208.220 2991.025 ;
        RECT 206.600 2990.795 208.220 2990.855 ;
        RECT 208.880 2991.025 210.215 2991.085 ;
        RECT 208.880 2990.855 210.045 2991.025 ;
        RECT 208.880 2990.795 210.215 2990.855 ;
        RECT 201.885 2990.565 202.055 2990.795 ;
        RECT 204.605 2990.565 204.775 2990.795 ;
        RECT 201.885 2990.235 202.055 2990.395 ;
        RECT 204.605 2990.235 204.775 2990.395 ;
        RECT 204.945 2990.285 205.965 2990.615 ;
        RECT 207.325 2990.565 207.495 2990.795 ;
        RECT 210.045 2990.710 210.215 2990.795 ;
        RECT 201.885 2990.105 202.855 2990.235 ;
        RECT 202.055 2989.935 202.855 2990.105 ;
        RECT 201.885 2989.905 202.855 2989.935 ;
        RECT 203.455 2990.115 204.775 2990.235 ;
        RECT 203.455 2990.105 205.575 2990.115 ;
        RECT 203.455 2989.935 204.605 2990.105 ;
        RECT 204.775 2989.945 205.575 2990.105 ;
        RECT 203.455 2989.905 204.775 2989.935 ;
        RECT 201.885 2989.645 202.055 2989.905 ;
        RECT 204.605 2989.645 204.775 2989.905 ;
        RECT 205.795 2989.775 205.965 2990.285 ;
        RECT 201.885 2989.395 202.055 2989.475 ;
        RECT 204.605 2989.395 204.775 2989.475 ;
        RECT 204.945 2989.445 205.965 2989.775 ;
        RECT 201.885 2989.185 202.535 2989.395 ;
        RECT 203.805 2989.275 204.775 2989.395 ;
        RECT 205.795 2989.290 205.965 2989.445 ;
        RECT 206.505 2990.365 207.155 2990.535 ;
        RECT 206.505 2989.695 206.675 2990.365 ;
        RECT 207.325 2990.195 207.495 2990.395 ;
        RECT 206.845 2990.105 207.495 2990.195 ;
        RECT 206.845 2989.935 207.325 2990.105 ;
        RECT 206.845 2989.865 207.495 2989.935 ;
        RECT 206.505 2989.525 207.150 2989.695 ;
        RECT 207.325 2989.645 207.495 2989.865 ;
        RECT 206.505 2989.290 206.675 2989.525 ;
        RECT 207.325 2989.355 207.495 2989.475 ;
        RECT 202.055 2989.065 202.535 2989.185 ;
        RECT 201.885 2988.725 202.055 2989.015 ;
        RECT 201.885 2988.265 202.535 2988.555 ;
        RECT 202.055 2988.225 202.535 2988.265 ;
        RECT 201.885 2987.805 202.055 2988.095 ;
        RECT 202.055 2987.635 202.535 2987.715 ;
        RECT 201.885 2987.385 202.535 2987.635 ;
        RECT 201.885 2987.345 202.055 2987.385 ;
        RECT 201.885 2986.885 202.055 2987.175 ;
        RECT 202.055 2986.715 202.535 2986.875 ;
        RECT 203.045 2986.785 203.215 2989.235 ;
        RECT 203.805 2989.185 205.575 2989.275 ;
        RECT 203.805 2989.065 204.605 2989.185 ;
        RECT 204.775 2989.105 205.575 2989.185 ;
        RECT 205.795 2989.115 206.675 2989.290 ;
        RECT 206.845 2989.185 207.495 2989.355 ;
        RECT 204.605 2988.725 204.775 2989.015 ;
      LAYER li1 ;
        RECT 204.945 2988.685 205.965 2988.855 ;
      LAYER li1 ;
        RECT 203.805 2988.515 204.775 2988.555 ;
        RECT 203.805 2988.265 205.575 2988.515 ;
        RECT 203.805 2988.225 204.605 2988.265 ;
        RECT 204.775 2988.185 205.575 2988.265 ;
        RECT 204.605 2987.805 204.775 2988.095 ;
      LAYER li1 ;
        RECT 205.795 2988.015 205.965 2988.685 ;
        RECT 204.945 2987.845 205.965 2988.015 ;
      LAYER li1 ;
        RECT 203.805 2987.635 204.605 2987.715 ;
        RECT 204.775 2987.635 205.575 2987.675 ;
        RECT 203.805 2987.385 205.575 2987.635 ;
        RECT 204.605 2987.345 205.575 2987.385 ;
      LAYER li1 ;
        RECT 205.795 2987.175 205.965 2987.845 ;
      LAYER li1 ;
        RECT 204.605 2986.885 204.775 2987.175 ;
      LAYER li1 ;
        RECT 204.945 2987.005 205.965 2987.175 ;
      LAYER li1 ;
        RECT 201.885 2986.545 202.535 2986.715 ;
        RECT 202.705 2986.610 203.585 2986.785 ;
        RECT 203.805 2986.715 204.605 2986.795 ;
        RECT 204.775 2986.715 205.575 2986.835 ;
        RECT 203.805 2986.625 205.575 2986.715 ;
        RECT 201.885 2986.425 202.055 2986.545 ;
        RECT 202.705 2986.375 202.875 2986.610 ;
        RECT 203.415 2986.455 203.585 2986.610 ;
        RECT 204.605 2986.505 205.575 2986.625 ;
        RECT 201.885 2986.035 202.055 2986.255 ;
        RECT 202.230 2986.205 202.875 2986.375 ;
        RECT 201.885 2985.965 202.535 2986.035 ;
        RECT 202.055 2985.795 202.535 2985.965 ;
        RECT 201.885 2985.705 202.535 2985.795 ;
        RECT 201.885 2985.505 202.055 2985.705 ;
        RECT 202.705 2985.535 202.875 2986.205 ;
        RECT 202.225 2985.365 202.875 2985.535 ;
        RECT 201.885 2985.105 202.055 2985.335 ;
      LAYER li1 ;
        RECT 203.045 2985.330 203.245 2986.430 ;
      LAYER li1 ;
        RECT 203.415 2986.125 204.435 2986.455 ;
        RECT 204.605 2986.425 204.775 2986.505 ;
      LAYER li1 ;
        RECT 205.795 2986.420 205.965 2987.005 ;
      LAYER li1 ;
        RECT 206.165 2986.665 206.335 2989.115 ;
        RECT 206.845 2989.025 207.325 2989.185 ;
      LAYER li1 ;
        RECT 207.495 2989.040 208.040 2990.625 ;
        RECT 206.505 2988.685 207.155 2988.855 ;
      LAYER li1 ;
        RECT 207.325 2988.725 207.495 2989.015 ;
      LAYER li1 ;
        RECT 207.495 2988.700 208.870 2989.040 ;
        RECT 206.505 2988.015 206.675 2988.685 ;
      LAYER li1 ;
        RECT 207.325 2988.515 207.495 2988.555 ;
        RECT 206.845 2988.265 207.495 2988.515 ;
        RECT 206.845 2988.185 207.325 2988.265 ;
      LAYER li1 ;
        RECT 206.505 2987.845 207.155 2988.015 ;
        RECT 206.505 2987.175 206.675 2987.845 ;
      LAYER li1 ;
        RECT 207.325 2987.805 207.495 2988.095 ;
        RECT 206.845 2987.635 207.325 2987.675 ;
        RECT 206.845 2987.345 207.495 2987.635 ;
      LAYER li1 ;
        RECT 206.505 2987.005 207.155 2987.175 ;
        RECT 206.505 2986.420 206.675 2987.005 ;
      LAYER li1 ;
        RECT 207.325 2986.885 207.495 2987.175 ;
        RECT 206.845 2986.715 207.325 2986.835 ;
        RECT 206.845 2986.505 207.495 2986.715 ;
        RECT 207.325 2986.425 207.495 2986.505 ;
      LAYER li1 ;
        RECT 205.795 2986.335 206.675 2986.420 ;
      LAYER li1 ;
        RECT 203.415 2985.615 203.585 2986.125 ;
        RECT 204.605 2985.995 204.775 2986.255 ;
      LAYER li1 ;
        RECT 204.945 2986.165 207.155 2986.335 ;
      LAYER li1 ;
        RECT 207.325 2985.995 207.495 2986.255 ;
        RECT 204.605 2985.965 205.925 2985.995 ;
        RECT 203.805 2985.795 204.605 2985.955 ;
        RECT 204.775 2985.795 205.925 2985.965 ;
        RECT 203.805 2985.785 205.925 2985.795 ;
        RECT 204.605 2985.665 205.925 2985.785 ;
        RECT 206.525 2985.965 207.495 2985.995 ;
        RECT 206.525 2985.795 207.325 2985.965 ;
        RECT 206.525 2985.665 207.495 2985.795 ;
        RECT 203.415 2985.285 204.435 2985.615 ;
        RECT 204.605 2985.505 204.775 2985.665 ;
        RECT 207.325 2985.505 207.495 2985.665 ;
        RECT 204.605 2985.105 204.775 2985.335 ;
        RECT 207.325 2985.105 207.495 2985.335 ;
      LAYER li1 ;
        RECT 207.495 2985.280 208.040 2988.700 ;
      LAYER li1 ;
        RECT 210.045 2985.105 210.215 2985.190 ;
        RECT 201.885 2985.045 202.780 2985.105 ;
        RECT 202.055 2984.875 202.780 2985.045 ;
        RECT 201.885 2984.815 202.780 2984.875 ;
        RECT 203.440 2985.045 205.940 2985.105 ;
        RECT 203.440 2984.875 204.605 2985.045 ;
        RECT 204.775 2984.875 205.940 2985.045 ;
        RECT 203.440 2984.815 205.940 2984.875 ;
        RECT 206.600 2985.045 208.220 2985.105 ;
        RECT 206.600 2984.875 207.325 2985.045 ;
        RECT 207.495 2984.875 208.220 2985.045 ;
        RECT 206.600 2984.815 208.220 2984.875 ;
        RECT 208.880 2985.045 210.215 2985.105 ;
        RECT 208.880 2984.875 210.045 2985.045 ;
        RECT 208.880 2984.815 210.215 2984.875 ;
        RECT 201.885 2984.730 202.055 2984.815 ;
        RECT 204.605 2984.730 204.775 2984.815 ;
        RECT 207.325 2984.730 207.495 2984.815 ;
        RECT 210.045 2984.730 210.215 2984.815 ;
        RECT 3377.780 2238.295 3377.950 2238.380 ;
        RECT 3380.500 2238.295 3380.670 2238.380 ;
        RECT 3383.220 2238.295 3383.390 2238.380 ;
        RECT 3385.940 2238.295 3386.110 2238.380 ;
        RECT 3377.780 2238.235 3379.115 2238.295 ;
        RECT 3377.950 2238.065 3379.115 2238.235 ;
        RECT 3377.780 2238.005 3379.115 2238.065 ;
        RECT 3379.775 2238.235 3381.395 2238.295 ;
        RECT 3379.775 2238.065 3380.500 2238.235 ;
        RECT 3380.670 2238.065 3381.395 2238.235 ;
        RECT 3379.775 2238.005 3381.395 2238.065 ;
        RECT 3377.780 2237.920 3377.950 2238.005 ;
        RECT 3380.500 2237.920 3380.670 2238.005 ;
        RECT 3380.840 2237.575 3381.490 2237.745 ;
        RECT 3380.670 2237.075 3381.150 2237.405 ;
        RECT 3381.320 2236.905 3381.490 2237.575 ;
        RECT 3380.845 2236.735 3381.490 2236.905 ;
        RECT 3380.670 2236.235 3381.150 2236.565 ;
        RECT 3381.320 2236.500 3381.490 2236.735 ;
      LAYER li1 ;
        RECT 3381.660 2236.680 3381.860 2238.270 ;
      LAYER li1 ;
        RECT 3382.055 2238.235 3384.555 2238.295 ;
        RECT 3382.055 2238.065 3383.220 2238.235 ;
        RECT 3383.390 2238.065 3384.555 2238.235 ;
        RECT 3382.055 2238.005 3384.555 2238.065 ;
        RECT 3385.215 2238.235 3386.110 2238.295 ;
        RECT 3385.215 2238.065 3385.940 2238.235 ;
        RECT 3385.215 2238.005 3386.110 2238.065 ;
        RECT 3382.030 2237.495 3383.050 2237.825 ;
        RECT 3383.220 2237.775 3383.390 2238.005 ;
        RECT 3385.940 2237.775 3386.110 2238.005 ;
        RECT 3382.030 2236.985 3382.200 2237.495 ;
        RECT 3383.220 2237.445 3383.390 2237.605 ;
        RECT 3385.940 2237.445 3386.110 2237.605 ;
        RECT 3383.220 2237.325 3384.540 2237.445 ;
        RECT 3382.420 2237.315 3384.540 2237.325 ;
        RECT 3382.420 2237.155 3383.220 2237.315 ;
        RECT 3383.390 2237.145 3384.540 2237.315 ;
        RECT 3383.220 2237.115 3384.540 2237.145 ;
        RECT 3385.140 2237.315 3386.110 2237.445 ;
        RECT 3385.140 2237.145 3385.940 2237.315 ;
        RECT 3385.140 2237.115 3386.110 2237.145 ;
        RECT 3382.030 2236.655 3383.050 2236.985 ;
        RECT 3383.220 2236.855 3383.390 2237.115 ;
      LAYER li1 ;
        RECT 3383.560 2236.775 3385.770 2236.945 ;
      LAYER li1 ;
        RECT 3385.940 2236.855 3386.110 2237.115 ;
      LAYER li1 ;
        RECT 3384.410 2236.690 3385.290 2236.775 ;
      LAYER li1 ;
        RECT 3382.030 2236.500 3382.200 2236.655 ;
        RECT 3381.320 2236.325 3382.200 2236.500 ;
        RECT 3383.220 2236.605 3383.390 2236.685 ;
        RECT 3383.220 2236.485 3384.190 2236.605 ;
        RECT 3382.420 2236.395 3384.190 2236.485 ;
        RECT 3380.670 2235.395 3381.150 2235.725 ;
        RECT 3380.670 2234.555 3381.150 2234.885 ;
        RECT 3380.670 2233.715 3381.150 2234.045 ;
        RECT 3381.660 2233.875 3381.830 2236.325 ;
        RECT 3382.420 2236.315 3383.220 2236.395 ;
        RECT 3383.390 2236.275 3384.190 2236.395 ;
        RECT 3383.220 2235.935 3383.390 2236.225 ;
      LAYER li1 ;
        RECT 3384.410 2236.105 3384.580 2236.690 ;
        RECT 3383.560 2235.935 3384.580 2236.105 ;
      LAYER li1 ;
        RECT 3383.220 2235.725 3384.190 2235.765 ;
        RECT 3382.420 2235.475 3384.190 2235.725 ;
        RECT 3382.420 2235.395 3383.220 2235.475 ;
        RECT 3383.390 2235.435 3384.190 2235.475 ;
        RECT 3383.220 2235.015 3383.390 2235.305 ;
      LAYER li1 ;
        RECT 3384.410 2235.265 3384.580 2235.935 ;
        RECT 3383.560 2235.095 3384.580 2235.265 ;
      LAYER li1 ;
        RECT 3382.420 2234.845 3383.220 2234.885 ;
        RECT 3383.390 2234.845 3384.190 2234.925 ;
        RECT 3382.420 2234.595 3384.190 2234.845 ;
        RECT 3382.420 2234.555 3383.390 2234.595 ;
      LAYER li1 ;
        RECT 3384.410 2234.425 3384.580 2235.095 ;
      LAYER li1 ;
        RECT 3383.220 2234.095 3383.390 2234.385 ;
      LAYER li1 ;
        RECT 3383.560 2234.255 3384.580 2234.425 ;
      LAYER li1 ;
        RECT 3382.420 2233.925 3383.220 2234.045 ;
        RECT 3383.390 2233.925 3384.190 2234.005 ;
        RECT 3384.780 2233.995 3384.950 2236.445 ;
      LAYER li1 ;
        RECT 3385.120 2236.105 3385.290 2236.690 ;
      LAYER li1 ;
        RECT 3385.940 2236.605 3386.110 2236.685 ;
        RECT 3385.460 2236.395 3386.110 2236.605 ;
        RECT 3385.460 2236.275 3385.940 2236.395 ;
      LAYER li1 ;
        RECT 3385.120 2235.935 3385.770 2236.105 ;
      LAYER li1 ;
        RECT 3385.940 2235.935 3386.110 2236.225 ;
      LAYER li1 ;
        RECT 3385.120 2235.265 3385.290 2235.935 ;
      LAYER li1 ;
        RECT 3385.460 2235.475 3386.110 2235.765 ;
        RECT 3385.460 2235.435 3385.940 2235.475 ;
      LAYER li1 ;
        RECT 3385.120 2235.095 3385.770 2235.265 ;
        RECT 3385.120 2234.425 3385.290 2235.095 ;
      LAYER li1 ;
        RECT 3385.940 2235.015 3386.110 2235.305 ;
        RECT 3385.460 2234.845 3385.940 2234.925 ;
        RECT 3385.460 2234.595 3386.110 2234.845 ;
        RECT 3385.940 2234.555 3386.110 2234.595 ;
      LAYER li1 ;
        RECT 3385.120 2234.255 3385.770 2234.425 ;
      LAYER li1 ;
        RECT 3385.940 2234.095 3386.110 2234.385 ;
        RECT 3382.420 2233.835 3384.190 2233.925 ;
        RECT 3382.420 2233.715 3383.390 2233.835 ;
        RECT 3383.220 2233.635 3383.390 2233.715 ;
        RECT 3384.410 2233.820 3385.290 2233.995 ;
        RECT 3384.410 2233.665 3384.580 2233.820 ;
        RECT 3383.220 2233.205 3383.390 2233.465 ;
        RECT 3383.560 2233.335 3384.580 2233.665 ;
        RECT 3380.670 2232.875 3381.470 2233.205 ;
        RECT 3382.070 2233.175 3383.390 2233.205 ;
        RECT 3382.070 2233.005 3383.220 2233.175 ;
        RECT 3383.390 2233.005 3384.190 2233.165 ;
        RECT 3382.070 2232.995 3384.190 2233.005 ;
        RECT 3382.070 2232.875 3383.390 2232.995 ;
        RECT 3383.220 2232.715 3383.390 2232.875 ;
        RECT 3384.410 2232.825 3384.580 2233.335 ;
        RECT 3377.780 2232.315 3377.950 2232.400 ;
        RECT 3380.500 2232.315 3380.670 2232.400 ;
        RECT 3383.220 2232.315 3383.390 2232.545 ;
        RECT 3383.560 2232.495 3384.580 2232.825 ;
        RECT 3385.120 2233.585 3385.290 2233.820 ;
        RECT 3385.460 2233.925 3385.940 2234.085 ;
        RECT 3385.460 2233.755 3386.110 2233.925 ;
        RECT 3385.940 2233.635 3386.110 2233.755 ;
        RECT 3385.120 2233.415 3385.765 2233.585 ;
        RECT 3385.120 2232.745 3385.290 2233.415 ;
        RECT 3385.940 2233.245 3386.110 2233.465 ;
        RECT 3385.460 2233.175 3386.110 2233.245 ;
        RECT 3385.460 2233.005 3385.940 2233.175 ;
        RECT 3385.460 2232.915 3386.110 2233.005 ;
        RECT 3385.120 2232.575 3385.770 2232.745 ;
        RECT 3385.940 2232.715 3386.110 2232.915 ;
        RECT 3385.940 2232.315 3386.110 2232.545 ;
        RECT 3377.780 2232.255 3379.115 2232.315 ;
        RECT 3377.950 2232.085 3379.115 2232.255 ;
        RECT 3377.780 2232.025 3379.115 2232.085 ;
        RECT 3379.775 2232.255 3381.395 2232.315 ;
        RECT 3379.775 2232.085 3380.500 2232.255 ;
        RECT 3380.670 2232.085 3381.395 2232.255 ;
        RECT 3379.775 2232.025 3381.395 2232.085 ;
        RECT 3382.055 2232.255 3384.555 2232.315 ;
        RECT 3382.055 2232.085 3383.220 2232.255 ;
        RECT 3383.390 2232.085 3384.555 2232.255 ;
        RECT 3382.055 2232.025 3384.555 2232.085 ;
        RECT 3385.215 2232.255 3386.110 2232.315 ;
        RECT 3385.215 2232.085 3385.940 2232.255 ;
        RECT 3385.215 2232.025 3386.110 2232.085 ;
        RECT 3377.780 2231.940 3377.950 2232.025 ;
      LAYER li1 ;
        RECT 3379.955 2230.270 3380.500 2231.855 ;
      LAYER li1 ;
        RECT 3380.500 2231.795 3380.670 2232.025 ;
        RECT 3380.500 2231.425 3380.670 2231.625 ;
        RECT 3380.840 2231.595 3381.490 2231.765 ;
        RECT 3380.500 2231.335 3381.150 2231.425 ;
        RECT 3380.670 2231.165 3381.150 2231.335 ;
        RECT 3380.500 2231.095 3381.150 2231.165 ;
        RECT 3380.500 2230.875 3380.670 2231.095 ;
        RECT 3381.320 2230.925 3381.490 2231.595 ;
        RECT 3380.845 2230.755 3381.490 2230.925 ;
        RECT 3380.500 2230.585 3380.670 2230.705 ;
        RECT 3380.500 2230.415 3381.150 2230.585 ;
      LAYER li1 ;
        RECT 3379.125 2229.930 3380.500 2230.270 ;
      LAYER li1 ;
        RECT 3380.670 2230.255 3381.150 2230.415 ;
        RECT 3381.320 2230.520 3381.490 2230.755 ;
        RECT 3382.030 2231.515 3383.050 2231.845 ;
        RECT 3383.220 2231.795 3383.390 2232.025 ;
        RECT 3385.940 2231.795 3386.110 2232.025 ;
        RECT 3382.030 2231.005 3382.200 2231.515 ;
        RECT 3383.220 2231.465 3383.390 2231.625 ;
        RECT 3385.940 2231.465 3386.110 2231.625 ;
        RECT 3383.220 2231.345 3384.540 2231.465 ;
        RECT 3382.420 2231.335 3384.540 2231.345 ;
        RECT 3382.420 2231.175 3383.220 2231.335 ;
        RECT 3383.390 2231.165 3384.540 2231.335 ;
        RECT 3383.220 2231.135 3384.540 2231.165 ;
        RECT 3385.140 2231.335 3386.110 2231.465 ;
        RECT 3385.140 2231.165 3385.940 2231.335 ;
        RECT 3385.140 2231.135 3386.110 2231.165 ;
        RECT 3382.030 2230.675 3383.050 2231.005 ;
        RECT 3383.220 2230.875 3383.390 2231.135 ;
        RECT 3385.940 2230.875 3386.110 2231.135 ;
        RECT 3382.030 2230.520 3382.200 2230.675 ;
        RECT 3381.320 2230.345 3382.200 2230.520 ;
        RECT 3383.220 2230.625 3383.390 2230.705 ;
        RECT 3385.940 2230.625 3386.110 2230.705 ;
        RECT 3383.220 2230.505 3384.190 2230.625 ;
        RECT 3382.420 2230.415 3384.190 2230.505 ;
        RECT 3380.500 2229.955 3380.670 2230.245 ;
      LAYER li1 ;
        RECT 3379.955 2226.510 3380.500 2229.930 ;
      LAYER li1 ;
        RECT 3380.500 2229.745 3380.670 2229.785 ;
        RECT 3380.500 2229.495 3381.150 2229.745 ;
        RECT 3380.670 2229.415 3381.150 2229.495 ;
        RECT 3380.500 2229.035 3380.670 2229.325 ;
        RECT 3380.670 2228.865 3381.150 2228.905 ;
        RECT 3380.500 2228.575 3381.150 2228.865 ;
        RECT 3380.500 2228.115 3380.670 2228.405 ;
        RECT 3380.670 2227.945 3381.150 2228.065 ;
        RECT 3380.500 2227.735 3381.150 2227.945 ;
        RECT 3381.660 2227.895 3381.830 2230.345 ;
        RECT 3382.420 2230.335 3383.220 2230.415 ;
        RECT 3383.390 2230.295 3384.190 2230.415 ;
        RECT 3383.220 2229.955 3383.390 2230.245 ;
        RECT 3383.220 2229.745 3384.190 2229.785 ;
        RECT 3382.420 2229.495 3384.190 2229.745 ;
        RECT 3382.420 2229.415 3383.220 2229.495 ;
        RECT 3383.390 2229.455 3384.190 2229.495 ;
        RECT 3383.220 2229.035 3383.390 2229.325 ;
        RECT 3382.420 2228.865 3383.220 2228.905 ;
        RECT 3383.390 2228.865 3384.190 2228.945 ;
        RECT 3382.420 2228.615 3384.190 2228.865 ;
        RECT 3382.420 2228.575 3383.390 2228.615 ;
        RECT 3383.220 2228.115 3383.390 2228.405 ;
        RECT 3382.420 2227.945 3383.220 2228.065 ;
        RECT 3383.390 2227.945 3384.190 2228.025 ;
        RECT 3384.780 2228.015 3384.950 2230.465 ;
        RECT 3385.460 2230.415 3386.110 2230.625 ;
        RECT 3385.460 2230.295 3385.940 2230.415 ;
        RECT 3385.940 2229.955 3386.110 2230.245 ;
        RECT 3385.460 2229.495 3386.110 2229.785 ;
        RECT 3385.460 2229.455 3385.940 2229.495 ;
        RECT 3385.940 2229.035 3386.110 2229.325 ;
        RECT 3385.460 2228.865 3385.940 2228.945 ;
        RECT 3385.460 2228.615 3386.110 2228.865 ;
        RECT 3385.940 2228.575 3386.110 2228.615 ;
        RECT 3385.940 2228.115 3386.110 2228.405 ;
        RECT 3382.420 2227.855 3384.190 2227.945 ;
        RECT 3382.420 2227.735 3383.390 2227.855 ;
        RECT 3380.500 2227.655 3380.670 2227.735 ;
        RECT 3383.220 2227.655 3383.390 2227.735 ;
        RECT 3384.410 2227.840 3385.290 2228.015 ;
        RECT 3384.410 2227.685 3384.580 2227.840 ;
        RECT 3380.500 2227.225 3380.670 2227.485 ;
        RECT 3383.220 2227.225 3383.390 2227.485 ;
        RECT 3383.560 2227.355 3384.580 2227.685 ;
        RECT 3380.500 2227.195 3381.470 2227.225 ;
        RECT 3380.670 2227.025 3381.470 2227.195 ;
        RECT 3380.500 2226.895 3381.470 2227.025 ;
        RECT 3382.070 2227.195 3383.390 2227.225 ;
        RECT 3382.070 2227.025 3383.220 2227.195 ;
        RECT 3383.390 2227.025 3384.190 2227.185 ;
        RECT 3382.070 2227.015 3384.190 2227.025 ;
        RECT 3382.070 2226.895 3383.390 2227.015 ;
        RECT 3380.500 2226.735 3380.670 2226.895 ;
        RECT 3383.220 2226.735 3383.390 2226.895 ;
        RECT 3384.410 2226.845 3384.580 2227.355 ;
        RECT 3377.780 2226.335 3377.950 2226.420 ;
        RECT 3380.500 2226.335 3380.670 2226.565 ;
        RECT 3383.220 2226.335 3383.390 2226.565 ;
        RECT 3383.560 2226.515 3384.580 2226.845 ;
        RECT 3385.120 2227.605 3385.290 2227.840 ;
        RECT 3385.460 2227.945 3385.940 2228.105 ;
        RECT 3385.460 2227.775 3386.110 2227.945 ;
        RECT 3385.940 2227.655 3386.110 2227.775 ;
        RECT 3385.120 2227.435 3385.765 2227.605 ;
        RECT 3385.120 2226.765 3385.290 2227.435 ;
        RECT 3385.940 2227.265 3386.110 2227.485 ;
        RECT 3385.460 2227.195 3386.110 2227.265 ;
        RECT 3385.460 2227.025 3385.940 2227.195 ;
        RECT 3385.460 2226.935 3386.110 2227.025 ;
        RECT 3385.120 2226.595 3385.770 2226.765 ;
        RECT 3385.940 2226.735 3386.110 2226.935 ;
        RECT 3385.940 2226.335 3386.110 2226.565 ;
        RECT 3377.780 2226.275 3379.115 2226.335 ;
        RECT 3377.950 2226.105 3379.115 2226.275 ;
        RECT 3377.780 2226.045 3379.115 2226.105 ;
        RECT 3379.775 2226.275 3381.395 2226.335 ;
        RECT 3379.775 2226.105 3380.500 2226.275 ;
        RECT 3380.670 2226.105 3381.395 2226.275 ;
        RECT 3379.775 2226.045 3381.395 2226.105 ;
        RECT 3382.055 2226.275 3384.555 2226.335 ;
        RECT 3382.055 2226.105 3383.220 2226.275 ;
        RECT 3383.390 2226.105 3384.555 2226.275 ;
        RECT 3382.055 2226.045 3384.555 2226.105 ;
        RECT 3385.215 2226.275 3386.110 2226.335 ;
        RECT 3385.215 2226.105 3385.940 2226.275 ;
        RECT 3385.215 2226.045 3386.110 2226.105 ;
        RECT 3377.780 2225.960 3377.950 2226.045 ;
      LAYER li1 ;
        RECT 3379.955 2224.290 3380.500 2225.875 ;
      LAYER li1 ;
        RECT 3380.500 2225.815 3380.670 2226.045 ;
        RECT 3380.500 2225.445 3380.670 2225.645 ;
        RECT 3380.840 2225.615 3381.490 2225.785 ;
        RECT 3380.500 2225.355 3381.150 2225.445 ;
        RECT 3380.670 2225.185 3381.150 2225.355 ;
        RECT 3380.500 2225.115 3381.150 2225.185 ;
        RECT 3380.500 2224.895 3380.670 2225.115 ;
        RECT 3381.320 2224.945 3381.490 2225.615 ;
        RECT 3380.845 2224.775 3381.490 2224.945 ;
        RECT 3380.500 2224.605 3380.670 2224.725 ;
        RECT 3380.500 2224.435 3381.150 2224.605 ;
      LAYER li1 ;
        RECT 3379.125 2223.950 3380.500 2224.290 ;
      LAYER li1 ;
        RECT 3380.670 2224.275 3381.150 2224.435 ;
        RECT 3381.320 2224.540 3381.490 2224.775 ;
        RECT 3382.030 2225.535 3383.050 2225.865 ;
        RECT 3383.220 2225.815 3383.390 2226.045 ;
        RECT 3385.940 2225.815 3386.110 2226.045 ;
        RECT 3382.030 2225.025 3382.200 2225.535 ;
        RECT 3383.220 2225.485 3383.390 2225.645 ;
        RECT 3385.940 2225.485 3386.110 2225.645 ;
        RECT 3383.220 2225.365 3384.540 2225.485 ;
        RECT 3382.420 2225.355 3384.540 2225.365 ;
        RECT 3382.420 2225.195 3383.220 2225.355 ;
        RECT 3383.390 2225.185 3384.540 2225.355 ;
        RECT 3383.220 2225.155 3384.540 2225.185 ;
        RECT 3385.140 2225.355 3386.110 2225.485 ;
        RECT 3385.140 2225.185 3385.940 2225.355 ;
        RECT 3385.140 2225.155 3386.110 2225.185 ;
        RECT 3382.030 2224.695 3383.050 2225.025 ;
        RECT 3383.220 2224.895 3383.390 2225.155 ;
        RECT 3385.940 2224.895 3386.110 2225.155 ;
        RECT 3382.030 2224.540 3382.200 2224.695 ;
        RECT 3381.320 2224.365 3382.200 2224.540 ;
        RECT 3383.220 2224.645 3383.390 2224.725 ;
        RECT 3385.940 2224.645 3386.110 2224.725 ;
        RECT 3383.220 2224.525 3384.190 2224.645 ;
        RECT 3382.420 2224.435 3384.190 2224.525 ;
        RECT 3380.500 2223.975 3380.670 2224.265 ;
      LAYER li1 ;
        RECT 3379.955 2220.530 3380.500 2223.950 ;
      LAYER li1 ;
        RECT 3380.500 2223.765 3380.670 2223.805 ;
        RECT 3380.500 2223.515 3381.150 2223.765 ;
        RECT 3380.670 2223.435 3381.150 2223.515 ;
        RECT 3380.500 2223.055 3380.670 2223.345 ;
        RECT 3380.670 2222.885 3381.150 2222.925 ;
        RECT 3380.500 2222.595 3381.150 2222.885 ;
        RECT 3380.500 2222.135 3380.670 2222.425 ;
        RECT 3380.670 2221.965 3381.150 2222.085 ;
        RECT 3380.500 2221.755 3381.150 2221.965 ;
        RECT 3381.660 2221.915 3381.830 2224.365 ;
        RECT 3382.420 2224.355 3383.220 2224.435 ;
        RECT 3383.390 2224.315 3384.190 2224.435 ;
        RECT 3383.220 2223.975 3383.390 2224.265 ;
        RECT 3383.220 2223.765 3384.190 2223.805 ;
        RECT 3382.420 2223.515 3384.190 2223.765 ;
        RECT 3382.420 2223.435 3383.220 2223.515 ;
        RECT 3383.390 2223.475 3384.190 2223.515 ;
        RECT 3383.220 2223.055 3383.390 2223.345 ;
        RECT 3382.420 2222.885 3383.220 2222.925 ;
        RECT 3383.390 2222.885 3384.190 2222.965 ;
        RECT 3382.420 2222.635 3384.190 2222.885 ;
        RECT 3382.420 2222.595 3383.390 2222.635 ;
        RECT 3383.220 2222.135 3383.390 2222.425 ;
        RECT 3382.420 2221.965 3383.220 2222.085 ;
        RECT 3383.390 2221.965 3384.190 2222.045 ;
        RECT 3384.780 2222.035 3384.950 2224.485 ;
        RECT 3385.460 2224.435 3386.110 2224.645 ;
        RECT 3385.460 2224.315 3385.940 2224.435 ;
        RECT 3385.940 2223.975 3386.110 2224.265 ;
        RECT 3385.460 2223.515 3386.110 2223.805 ;
        RECT 3385.460 2223.475 3385.940 2223.515 ;
        RECT 3385.940 2223.055 3386.110 2223.345 ;
        RECT 3385.460 2222.885 3385.940 2222.965 ;
        RECT 3385.460 2222.635 3386.110 2222.885 ;
        RECT 3385.940 2222.595 3386.110 2222.635 ;
        RECT 3385.940 2222.135 3386.110 2222.425 ;
        RECT 3382.420 2221.875 3384.190 2221.965 ;
        RECT 3382.420 2221.755 3383.390 2221.875 ;
        RECT 3380.500 2221.675 3380.670 2221.755 ;
        RECT 3383.220 2221.675 3383.390 2221.755 ;
        RECT 3384.410 2221.860 3385.290 2222.035 ;
        RECT 3384.410 2221.705 3384.580 2221.860 ;
        RECT 3380.500 2221.245 3380.670 2221.505 ;
        RECT 3383.220 2221.245 3383.390 2221.505 ;
        RECT 3383.560 2221.375 3384.580 2221.705 ;
        RECT 3380.500 2221.215 3381.470 2221.245 ;
        RECT 3380.670 2221.045 3381.470 2221.215 ;
        RECT 3380.500 2220.915 3381.470 2221.045 ;
        RECT 3382.070 2221.215 3383.390 2221.245 ;
        RECT 3382.070 2221.045 3383.220 2221.215 ;
        RECT 3383.390 2221.045 3384.190 2221.205 ;
        RECT 3382.070 2221.035 3384.190 2221.045 ;
        RECT 3382.070 2220.915 3383.390 2221.035 ;
        RECT 3380.500 2220.755 3380.670 2220.915 ;
        RECT 3383.220 2220.755 3383.390 2220.915 ;
        RECT 3384.410 2220.865 3384.580 2221.375 ;
        RECT 3377.780 2220.355 3377.950 2220.440 ;
        RECT 3380.500 2220.355 3380.670 2220.585 ;
        RECT 3383.220 2220.355 3383.390 2220.585 ;
        RECT 3383.560 2220.535 3384.580 2220.865 ;
        RECT 3385.120 2221.625 3385.290 2221.860 ;
        RECT 3385.460 2221.965 3385.940 2222.125 ;
        RECT 3385.460 2221.795 3386.110 2221.965 ;
        RECT 3385.940 2221.675 3386.110 2221.795 ;
        RECT 3385.120 2221.455 3385.765 2221.625 ;
        RECT 3385.120 2220.785 3385.290 2221.455 ;
        RECT 3385.940 2221.285 3386.110 2221.505 ;
        RECT 3385.460 2221.215 3386.110 2221.285 ;
        RECT 3385.460 2221.045 3385.940 2221.215 ;
        RECT 3385.460 2220.955 3386.110 2221.045 ;
        RECT 3385.120 2220.615 3385.770 2220.785 ;
        RECT 3385.940 2220.755 3386.110 2220.955 ;
        RECT 3385.940 2220.355 3386.110 2220.585 ;
        RECT 3377.780 2220.295 3379.115 2220.355 ;
        RECT 3377.950 2220.125 3379.115 2220.295 ;
        RECT 3377.780 2220.065 3379.115 2220.125 ;
        RECT 3379.775 2220.295 3381.395 2220.355 ;
        RECT 3379.775 2220.125 3380.500 2220.295 ;
        RECT 3380.670 2220.125 3381.395 2220.295 ;
        RECT 3379.775 2220.065 3381.395 2220.125 ;
        RECT 3382.055 2220.295 3384.555 2220.355 ;
        RECT 3382.055 2220.125 3383.220 2220.295 ;
        RECT 3383.390 2220.125 3384.555 2220.295 ;
        RECT 3382.055 2220.065 3384.555 2220.125 ;
        RECT 3385.215 2220.295 3386.110 2220.355 ;
        RECT 3385.215 2220.125 3385.940 2220.295 ;
        RECT 3385.215 2220.065 3386.110 2220.125 ;
        RECT 3377.780 2219.980 3377.950 2220.065 ;
      LAYER li1 ;
        RECT 3379.955 2218.310 3380.500 2219.895 ;
      LAYER li1 ;
        RECT 3380.500 2219.835 3380.670 2220.065 ;
        RECT 3380.500 2219.465 3380.670 2219.665 ;
        RECT 3380.840 2219.635 3381.490 2219.805 ;
        RECT 3380.500 2219.375 3381.150 2219.465 ;
        RECT 3380.670 2219.205 3381.150 2219.375 ;
        RECT 3380.500 2219.135 3381.150 2219.205 ;
        RECT 3380.500 2218.915 3380.670 2219.135 ;
        RECT 3381.320 2218.965 3381.490 2219.635 ;
        RECT 3380.845 2218.795 3381.490 2218.965 ;
        RECT 3380.500 2218.625 3380.670 2218.745 ;
        RECT 3380.500 2218.455 3381.150 2218.625 ;
      LAYER li1 ;
        RECT 3379.125 2217.970 3380.500 2218.310 ;
      LAYER li1 ;
        RECT 3380.670 2218.295 3381.150 2218.455 ;
        RECT 3381.320 2218.560 3381.490 2218.795 ;
        RECT 3382.030 2219.555 3383.050 2219.885 ;
        RECT 3383.220 2219.835 3383.390 2220.065 ;
        RECT 3385.940 2219.835 3386.110 2220.065 ;
        RECT 3382.030 2219.045 3382.200 2219.555 ;
        RECT 3383.220 2219.505 3383.390 2219.665 ;
        RECT 3385.940 2219.505 3386.110 2219.665 ;
        RECT 3383.220 2219.385 3384.540 2219.505 ;
        RECT 3382.420 2219.375 3384.540 2219.385 ;
        RECT 3382.420 2219.215 3383.220 2219.375 ;
        RECT 3383.390 2219.205 3384.540 2219.375 ;
        RECT 3383.220 2219.175 3384.540 2219.205 ;
        RECT 3385.140 2219.375 3386.110 2219.505 ;
        RECT 3385.140 2219.205 3385.940 2219.375 ;
        RECT 3385.140 2219.175 3386.110 2219.205 ;
        RECT 3382.030 2218.715 3383.050 2219.045 ;
        RECT 3383.220 2218.915 3383.390 2219.175 ;
        RECT 3385.940 2218.915 3386.110 2219.175 ;
        RECT 3382.030 2218.560 3382.200 2218.715 ;
        RECT 3381.320 2218.385 3382.200 2218.560 ;
        RECT 3383.220 2218.665 3383.390 2218.745 ;
        RECT 3385.940 2218.665 3386.110 2218.745 ;
        RECT 3383.220 2218.545 3384.190 2218.665 ;
        RECT 3382.420 2218.455 3384.190 2218.545 ;
        RECT 3380.500 2217.995 3380.670 2218.285 ;
      LAYER li1 ;
        RECT 3379.955 2214.550 3380.500 2217.970 ;
      LAYER li1 ;
        RECT 3380.500 2217.785 3380.670 2217.825 ;
        RECT 3380.500 2217.535 3381.150 2217.785 ;
        RECT 3380.670 2217.455 3381.150 2217.535 ;
        RECT 3380.500 2217.075 3380.670 2217.365 ;
        RECT 3380.670 2216.905 3381.150 2216.945 ;
        RECT 3380.500 2216.615 3381.150 2216.905 ;
        RECT 3380.500 2216.155 3380.670 2216.445 ;
        RECT 3380.670 2215.985 3381.150 2216.105 ;
        RECT 3380.500 2215.775 3381.150 2215.985 ;
        RECT 3381.660 2215.935 3381.830 2218.385 ;
        RECT 3382.420 2218.375 3383.220 2218.455 ;
        RECT 3383.390 2218.335 3384.190 2218.455 ;
        RECT 3383.220 2217.995 3383.390 2218.285 ;
        RECT 3383.220 2217.785 3384.190 2217.825 ;
        RECT 3382.420 2217.535 3384.190 2217.785 ;
        RECT 3382.420 2217.455 3383.220 2217.535 ;
        RECT 3383.390 2217.495 3384.190 2217.535 ;
        RECT 3383.220 2217.075 3383.390 2217.365 ;
        RECT 3382.420 2216.905 3383.220 2216.945 ;
        RECT 3383.390 2216.905 3384.190 2216.985 ;
        RECT 3382.420 2216.655 3384.190 2216.905 ;
        RECT 3382.420 2216.615 3383.390 2216.655 ;
        RECT 3383.220 2216.155 3383.390 2216.445 ;
        RECT 3382.420 2215.985 3383.220 2216.105 ;
        RECT 3383.390 2215.985 3384.190 2216.065 ;
        RECT 3384.780 2216.055 3384.950 2218.505 ;
        RECT 3385.460 2218.455 3386.110 2218.665 ;
        RECT 3385.460 2218.335 3385.940 2218.455 ;
        RECT 3385.940 2217.995 3386.110 2218.285 ;
        RECT 3385.460 2217.535 3386.110 2217.825 ;
        RECT 3385.460 2217.495 3385.940 2217.535 ;
        RECT 3385.940 2217.075 3386.110 2217.365 ;
        RECT 3385.460 2216.905 3385.940 2216.985 ;
        RECT 3385.460 2216.655 3386.110 2216.905 ;
        RECT 3385.940 2216.615 3386.110 2216.655 ;
        RECT 3385.940 2216.155 3386.110 2216.445 ;
        RECT 3382.420 2215.895 3384.190 2215.985 ;
        RECT 3382.420 2215.775 3383.390 2215.895 ;
        RECT 3380.500 2215.695 3380.670 2215.775 ;
        RECT 3383.220 2215.695 3383.390 2215.775 ;
        RECT 3384.410 2215.880 3385.290 2216.055 ;
        RECT 3384.410 2215.725 3384.580 2215.880 ;
        RECT 3380.500 2215.265 3380.670 2215.525 ;
        RECT 3383.220 2215.265 3383.390 2215.525 ;
        RECT 3383.560 2215.395 3384.580 2215.725 ;
        RECT 3380.500 2215.235 3381.470 2215.265 ;
        RECT 3380.670 2215.065 3381.470 2215.235 ;
        RECT 3380.500 2214.935 3381.470 2215.065 ;
        RECT 3382.070 2215.235 3383.390 2215.265 ;
        RECT 3382.070 2215.065 3383.220 2215.235 ;
        RECT 3383.390 2215.065 3384.190 2215.225 ;
        RECT 3382.070 2215.055 3384.190 2215.065 ;
        RECT 3382.070 2214.935 3383.390 2215.055 ;
        RECT 3380.500 2214.775 3380.670 2214.935 ;
        RECT 3383.220 2214.775 3383.390 2214.935 ;
        RECT 3384.410 2214.885 3384.580 2215.395 ;
        RECT 3377.780 2214.375 3377.950 2214.460 ;
        RECT 3380.500 2214.375 3380.670 2214.605 ;
        RECT 3383.220 2214.375 3383.390 2214.605 ;
        RECT 3383.560 2214.555 3384.580 2214.885 ;
        RECT 3385.120 2215.645 3385.290 2215.880 ;
        RECT 3385.460 2215.985 3385.940 2216.145 ;
        RECT 3385.460 2215.815 3386.110 2215.985 ;
        RECT 3385.940 2215.695 3386.110 2215.815 ;
        RECT 3385.120 2215.475 3385.765 2215.645 ;
        RECT 3385.120 2214.805 3385.290 2215.475 ;
        RECT 3385.940 2215.305 3386.110 2215.525 ;
        RECT 3385.460 2215.235 3386.110 2215.305 ;
        RECT 3385.460 2215.065 3385.940 2215.235 ;
        RECT 3385.460 2214.975 3386.110 2215.065 ;
        RECT 3385.120 2214.635 3385.770 2214.805 ;
        RECT 3385.940 2214.775 3386.110 2214.975 ;
        RECT 3385.940 2214.375 3386.110 2214.605 ;
        RECT 3377.780 2214.315 3379.115 2214.375 ;
        RECT 3377.950 2214.145 3379.115 2214.315 ;
        RECT 3377.780 2214.085 3379.115 2214.145 ;
        RECT 3379.775 2214.315 3381.395 2214.375 ;
        RECT 3379.775 2214.145 3380.500 2214.315 ;
        RECT 3380.670 2214.145 3381.395 2214.315 ;
        RECT 3379.775 2214.085 3381.395 2214.145 ;
        RECT 3382.055 2214.315 3384.555 2214.375 ;
        RECT 3382.055 2214.145 3383.220 2214.315 ;
        RECT 3383.390 2214.145 3384.555 2214.315 ;
        RECT 3382.055 2214.085 3384.555 2214.145 ;
        RECT 3385.215 2214.315 3386.110 2214.375 ;
        RECT 3385.215 2214.145 3385.940 2214.315 ;
        RECT 3385.215 2214.085 3386.110 2214.145 ;
        RECT 3377.780 2214.000 3377.950 2214.085 ;
      LAYER li1 ;
        RECT 3379.955 2212.330 3380.500 2213.915 ;
      LAYER li1 ;
        RECT 3380.500 2213.855 3380.670 2214.085 ;
        RECT 3380.500 2213.485 3380.670 2213.685 ;
        RECT 3380.840 2213.655 3381.490 2213.825 ;
        RECT 3380.500 2213.395 3381.150 2213.485 ;
        RECT 3380.670 2213.225 3381.150 2213.395 ;
        RECT 3380.500 2213.155 3381.150 2213.225 ;
        RECT 3380.500 2212.935 3380.670 2213.155 ;
        RECT 3381.320 2212.985 3381.490 2213.655 ;
        RECT 3380.845 2212.815 3381.490 2212.985 ;
        RECT 3380.500 2212.645 3380.670 2212.765 ;
        RECT 3380.500 2212.475 3381.150 2212.645 ;
      LAYER li1 ;
        RECT 3379.125 2211.990 3380.500 2212.330 ;
      LAYER li1 ;
        RECT 3380.670 2212.315 3381.150 2212.475 ;
        RECT 3381.320 2212.580 3381.490 2212.815 ;
        RECT 3382.030 2213.575 3383.050 2213.905 ;
        RECT 3383.220 2213.855 3383.390 2214.085 ;
        RECT 3385.940 2213.855 3386.110 2214.085 ;
        RECT 3382.030 2213.065 3382.200 2213.575 ;
        RECT 3383.220 2213.525 3383.390 2213.685 ;
        RECT 3385.940 2213.525 3386.110 2213.685 ;
        RECT 3383.220 2213.405 3384.540 2213.525 ;
        RECT 3382.420 2213.395 3384.540 2213.405 ;
        RECT 3382.420 2213.235 3383.220 2213.395 ;
        RECT 3383.390 2213.225 3384.540 2213.395 ;
        RECT 3383.220 2213.195 3384.540 2213.225 ;
        RECT 3385.140 2213.395 3386.110 2213.525 ;
        RECT 3385.140 2213.225 3385.940 2213.395 ;
        RECT 3385.140 2213.195 3386.110 2213.225 ;
        RECT 3382.030 2212.735 3383.050 2213.065 ;
        RECT 3383.220 2212.935 3383.390 2213.195 ;
        RECT 3385.940 2212.935 3386.110 2213.195 ;
        RECT 3382.030 2212.580 3382.200 2212.735 ;
        RECT 3381.320 2212.405 3382.200 2212.580 ;
        RECT 3383.220 2212.685 3383.390 2212.765 ;
        RECT 3385.940 2212.685 3386.110 2212.765 ;
        RECT 3383.220 2212.565 3384.190 2212.685 ;
        RECT 3382.420 2212.475 3384.190 2212.565 ;
        RECT 3380.500 2212.015 3380.670 2212.305 ;
      LAYER li1 ;
        RECT 3379.955 2208.570 3380.500 2211.990 ;
      LAYER li1 ;
        RECT 3380.500 2211.805 3380.670 2211.845 ;
        RECT 3380.500 2211.555 3381.150 2211.805 ;
        RECT 3380.670 2211.475 3381.150 2211.555 ;
        RECT 3380.500 2211.095 3380.670 2211.385 ;
        RECT 3380.670 2210.925 3381.150 2210.965 ;
        RECT 3380.500 2210.635 3381.150 2210.925 ;
        RECT 3380.500 2210.175 3380.670 2210.465 ;
        RECT 3380.670 2210.005 3381.150 2210.125 ;
        RECT 3380.500 2209.795 3381.150 2210.005 ;
        RECT 3381.660 2209.955 3381.830 2212.405 ;
        RECT 3382.420 2212.395 3383.220 2212.475 ;
        RECT 3383.390 2212.355 3384.190 2212.475 ;
        RECT 3383.220 2212.015 3383.390 2212.305 ;
        RECT 3383.220 2211.805 3384.190 2211.845 ;
        RECT 3382.420 2211.555 3384.190 2211.805 ;
        RECT 3382.420 2211.475 3383.220 2211.555 ;
        RECT 3383.390 2211.515 3384.190 2211.555 ;
        RECT 3383.220 2211.095 3383.390 2211.385 ;
        RECT 3382.420 2210.925 3383.220 2210.965 ;
        RECT 3383.390 2210.925 3384.190 2211.005 ;
        RECT 3382.420 2210.675 3384.190 2210.925 ;
        RECT 3382.420 2210.635 3383.390 2210.675 ;
        RECT 3383.220 2210.175 3383.390 2210.465 ;
        RECT 3382.420 2210.005 3383.220 2210.125 ;
        RECT 3383.390 2210.005 3384.190 2210.085 ;
        RECT 3384.780 2210.075 3384.950 2212.525 ;
        RECT 3385.460 2212.475 3386.110 2212.685 ;
        RECT 3385.460 2212.355 3385.940 2212.475 ;
        RECT 3385.940 2212.015 3386.110 2212.305 ;
        RECT 3385.460 2211.555 3386.110 2211.845 ;
        RECT 3385.460 2211.515 3385.940 2211.555 ;
        RECT 3385.940 2211.095 3386.110 2211.385 ;
        RECT 3385.460 2210.925 3385.940 2211.005 ;
        RECT 3385.460 2210.675 3386.110 2210.925 ;
        RECT 3385.940 2210.635 3386.110 2210.675 ;
        RECT 3385.940 2210.175 3386.110 2210.465 ;
        RECT 3382.420 2209.915 3384.190 2210.005 ;
        RECT 3382.420 2209.795 3383.390 2209.915 ;
        RECT 3380.500 2209.715 3380.670 2209.795 ;
        RECT 3383.220 2209.715 3383.390 2209.795 ;
        RECT 3384.410 2209.900 3385.290 2210.075 ;
        RECT 3384.410 2209.745 3384.580 2209.900 ;
        RECT 3380.500 2209.285 3380.670 2209.545 ;
        RECT 3383.220 2209.285 3383.390 2209.545 ;
        RECT 3383.560 2209.415 3384.580 2209.745 ;
        RECT 3380.500 2209.255 3381.470 2209.285 ;
        RECT 3380.670 2209.085 3381.470 2209.255 ;
        RECT 3380.500 2208.955 3381.470 2209.085 ;
        RECT 3382.070 2209.255 3383.390 2209.285 ;
        RECT 3382.070 2209.085 3383.220 2209.255 ;
        RECT 3383.390 2209.085 3384.190 2209.245 ;
        RECT 3382.070 2209.075 3384.190 2209.085 ;
        RECT 3382.070 2208.955 3383.390 2209.075 ;
        RECT 3380.500 2208.795 3380.670 2208.955 ;
        RECT 3383.220 2208.795 3383.390 2208.955 ;
        RECT 3384.410 2208.905 3384.580 2209.415 ;
        RECT 3377.780 2208.395 3377.950 2208.480 ;
        RECT 3380.500 2208.395 3380.670 2208.625 ;
        RECT 3383.220 2208.395 3383.390 2208.625 ;
        RECT 3383.560 2208.575 3384.580 2208.905 ;
        RECT 3385.120 2209.665 3385.290 2209.900 ;
        RECT 3385.460 2210.005 3385.940 2210.165 ;
        RECT 3385.460 2209.835 3386.110 2210.005 ;
        RECT 3385.940 2209.715 3386.110 2209.835 ;
        RECT 3385.120 2209.495 3385.765 2209.665 ;
        RECT 3385.120 2208.825 3385.290 2209.495 ;
        RECT 3385.940 2209.325 3386.110 2209.545 ;
        RECT 3385.460 2209.255 3386.110 2209.325 ;
        RECT 3385.460 2209.085 3385.940 2209.255 ;
        RECT 3385.460 2208.995 3386.110 2209.085 ;
        RECT 3385.120 2208.655 3385.770 2208.825 ;
        RECT 3385.940 2208.795 3386.110 2208.995 ;
        RECT 3385.940 2208.395 3386.110 2208.625 ;
        RECT 3377.780 2208.335 3379.115 2208.395 ;
        RECT 3377.950 2208.165 3379.115 2208.335 ;
        RECT 3377.780 2208.105 3379.115 2208.165 ;
        RECT 3379.775 2208.335 3381.395 2208.395 ;
        RECT 3379.775 2208.165 3380.500 2208.335 ;
        RECT 3380.670 2208.165 3381.395 2208.335 ;
        RECT 3379.775 2208.105 3381.395 2208.165 ;
        RECT 3382.055 2208.335 3384.555 2208.395 ;
        RECT 3382.055 2208.165 3383.220 2208.335 ;
        RECT 3383.390 2208.165 3384.555 2208.335 ;
        RECT 3382.055 2208.105 3384.555 2208.165 ;
        RECT 3385.215 2208.335 3386.110 2208.395 ;
        RECT 3385.215 2208.165 3385.940 2208.335 ;
        RECT 3385.215 2208.105 3386.110 2208.165 ;
        RECT 3377.780 2208.020 3377.950 2208.105 ;
      LAYER li1 ;
        RECT 3379.955 2206.350 3380.500 2207.935 ;
      LAYER li1 ;
        RECT 3380.500 2207.875 3380.670 2208.105 ;
        RECT 3380.500 2207.505 3380.670 2207.705 ;
        RECT 3380.840 2207.675 3381.490 2207.845 ;
        RECT 3380.500 2207.415 3381.150 2207.505 ;
        RECT 3380.670 2207.245 3381.150 2207.415 ;
        RECT 3380.500 2207.175 3381.150 2207.245 ;
        RECT 3380.500 2206.955 3380.670 2207.175 ;
        RECT 3381.320 2207.005 3381.490 2207.675 ;
        RECT 3380.845 2206.835 3381.490 2207.005 ;
        RECT 3380.500 2206.665 3380.670 2206.785 ;
        RECT 3380.500 2206.495 3381.150 2206.665 ;
      LAYER li1 ;
        RECT 3379.125 2206.010 3380.500 2206.350 ;
      LAYER li1 ;
        RECT 3380.670 2206.335 3381.150 2206.495 ;
        RECT 3381.320 2206.600 3381.490 2206.835 ;
        RECT 3382.030 2207.595 3383.050 2207.925 ;
        RECT 3383.220 2207.875 3383.390 2208.105 ;
        RECT 3385.940 2207.875 3386.110 2208.105 ;
        RECT 3382.030 2207.085 3382.200 2207.595 ;
        RECT 3383.220 2207.545 3383.390 2207.705 ;
        RECT 3385.940 2207.545 3386.110 2207.705 ;
        RECT 3383.220 2207.425 3384.540 2207.545 ;
        RECT 3382.420 2207.415 3384.540 2207.425 ;
        RECT 3382.420 2207.255 3383.220 2207.415 ;
        RECT 3383.390 2207.245 3384.540 2207.415 ;
        RECT 3383.220 2207.215 3384.540 2207.245 ;
        RECT 3385.140 2207.415 3386.110 2207.545 ;
        RECT 3385.140 2207.245 3385.940 2207.415 ;
        RECT 3385.140 2207.215 3386.110 2207.245 ;
        RECT 3382.030 2206.755 3383.050 2207.085 ;
        RECT 3383.220 2206.955 3383.390 2207.215 ;
        RECT 3385.940 2206.955 3386.110 2207.215 ;
        RECT 3382.030 2206.600 3382.200 2206.755 ;
        RECT 3381.320 2206.425 3382.200 2206.600 ;
        RECT 3383.220 2206.705 3383.390 2206.785 ;
        RECT 3385.940 2206.705 3386.110 2206.785 ;
        RECT 3383.220 2206.585 3384.190 2206.705 ;
        RECT 3382.420 2206.495 3384.190 2206.585 ;
        RECT 3380.500 2206.035 3380.670 2206.325 ;
      LAYER li1 ;
        RECT 3379.955 2202.590 3380.500 2206.010 ;
      LAYER li1 ;
        RECT 3380.500 2205.825 3380.670 2205.865 ;
        RECT 3380.500 2205.575 3381.150 2205.825 ;
        RECT 3380.670 2205.495 3381.150 2205.575 ;
        RECT 3380.500 2205.115 3380.670 2205.405 ;
        RECT 3380.670 2204.945 3381.150 2204.985 ;
        RECT 3380.500 2204.655 3381.150 2204.945 ;
        RECT 3380.500 2204.195 3380.670 2204.485 ;
        RECT 3380.670 2204.025 3381.150 2204.145 ;
        RECT 3380.500 2203.815 3381.150 2204.025 ;
        RECT 3381.660 2203.975 3381.830 2206.425 ;
        RECT 3382.420 2206.415 3383.220 2206.495 ;
        RECT 3383.390 2206.375 3384.190 2206.495 ;
        RECT 3383.220 2206.035 3383.390 2206.325 ;
        RECT 3383.220 2205.825 3384.190 2205.865 ;
        RECT 3382.420 2205.575 3384.190 2205.825 ;
        RECT 3382.420 2205.495 3383.220 2205.575 ;
        RECT 3383.390 2205.535 3384.190 2205.575 ;
        RECT 3383.220 2205.115 3383.390 2205.405 ;
        RECT 3382.420 2204.945 3383.220 2204.985 ;
        RECT 3383.390 2204.945 3384.190 2205.025 ;
        RECT 3382.420 2204.695 3384.190 2204.945 ;
        RECT 3382.420 2204.655 3383.390 2204.695 ;
        RECT 3383.220 2204.195 3383.390 2204.485 ;
        RECT 3382.420 2204.025 3383.220 2204.145 ;
        RECT 3383.390 2204.025 3384.190 2204.105 ;
        RECT 3384.780 2204.095 3384.950 2206.545 ;
        RECT 3385.460 2206.495 3386.110 2206.705 ;
        RECT 3385.460 2206.375 3385.940 2206.495 ;
        RECT 3385.940 2206.035 3386.110 2206.325 ;
        RECT 3385.460 2205.575 3386.110 2205.865 ;
        RECT 3385.460 2205.535 3385.940 2205.575 ;
        RECT 3385.940 2205.115 3386.110 2205.405 ;
        RECT 3385.460 2204.945 3385.940 2205.025 ;
        RECT 3385.460 2204.695 3386.110 2204.945 ;
        RECT 3385.940 2204.655 3386.110 2204.695 ;
        RECT 3385.940 2204.195 3386.110 2204.485 ;
        RECT 3382.420 2203.935 3384.190 2204.025 ;
        RECT 3382.420 2203.815 3383.390 2203.935 ;
        RECT 3380.500 2203.735 3380.670 2203.815 ;
        RECT 3383.220 2203.735 3383.390 2203.815 ;
        RECT 3384.410 2203.920 3385.290 2204.095 ;
        RECT 3384.410 2203.765 3384.580 2203.920 ;
        RECT 3380.500 2203.305 3380.670 2203.565 ;
        RECT 3383.220 2203.305 3383.390 2203.565 ;
        RECT 3383.560 2203.435 3384.580 2203.765 ;
        RECT 3380.500 2203.275 3381.470 2203.305 ;
        RECT 3380.670 2203.105 3381.470 2203.275 ;
        RECT 3380.500 2202.975 3381.470 2203.105 ;
        RECT 3382.070 2203.275 3383.390 2203.305 ;
        RECT 3382.070 2203.105 3383.220 2203.275 ;
        RECT 3383.390 2203.105 3384.190 2203.265 ;
        RECT 3382.070 2203.095 3384.190 2203.105 ;
        RECT 3382.070 2202.975 3383.390 2203.095 ;
        RECT 3380.500 2202.815 3380.670 2202.975 ;
        RECT 3383.220 2202.815 3383.390 2202.975 ;
        RECT 3384.410 2202.925 3384.580 2203.435 ;
        RECT 3377.780 2202.415 3377.950 2202.500 ;
        RECT 3380.500 2202.415 3380.670 2202.645 ;
        RECT 3383.220 2202.415 3383.390 2202.645 ;
        RECT 3383.560 2202.595 3384.580 2202.925 ;
        RECT 3385.120 2203.685 3385.290 2203.920 ;
        RECT 3385.460 2204.025 3385.940 2204.185 ;
        RECT 3385.460 2203.855 3386.110 2204.025 ;
        RECT 3385.940 2203.735 3386.110 2203.855 ;
        RECT 3385.120 2203.515 3385.765 2203.685 ;
        RECT 3385.120 2202.845 3385.290 2203.515 ;
        RECT 3385.940 2203.345 3386.110 2203.565 ;
        RECT 3385.460 2203.275 3386.110 2203.345 ;
        RECT 3385.460 2203.105 3385.940 2203.275 ;
        RECT 3385.460 2203.015 3386.110 2203.105 ;
        RECT 3385.120 2202.675 3385.770 2202.845 ;
        RECT 3385.940 2202.815 3386.110 2203.015 ;
        RECT 3385.940 2202.415 3386.110 2202.645 ;
        RECT 3377.780 2202.355 3379.115 2202.415 ;
        RECT 3377.950 2202.185 3379.115 2202.355 ;
        RECT 3377.780 2202.125 3379.115 2202.185 ;
        RECT 3379.775 2202.355 3381.395 2202.415 ;
        RECT 3379.775 2202.185 3380.500 2202.355 ;
        RECT 3380.670 2202.185 3381.395 2202.355 ;
        RECT 3379.775 2202.125 3381.395 2202.185 ;
        RECT 3382.055 2202.355 3384.555 2202.415 ;
        RECT 3382.055 2202.185 3383.220 2202.355 ;
        RECT 3383.390 2202.185 3384.555 2202.355 ;
        RECT 3382.055 2202.125 3384.555 2202.185 ;
        RECT 3385.215 2202.355 3386.110 2202.415 ;
        RECT 3385.215 2202.185 3385.940 2202.355 ;
        RECT 3385.215 2202.125 3386.110 2202.185 ;
        RECT 3377.780 2202.040 3377.950 2202.125 ;
      LAYER li1 ;
        RECT 3379.955 2200.370 3380.500 2201.955 ;
      LAYER li1 ;
        RECT 3380.500 2201.895 3380.670 2202.125 ;
        RECT 3380.500 2201.525 3380.670 2201.725 ;
        RECT 3380.840 2201.695 3381.490 2201.865 ;
        RECT 3380.500 2201.435 3381.150 2201.525 ;
        RECT 3380.670 2201.265 3381.150 2201.435 ;
        RECT 3380.500 2201.195 3381.150 2201.265 ;
        RECT 3380.500 2200.975 3380.670 2201.195 ;
        RECT 3381.320 2201.025 3381.490 2201.695 ;
        RECT 3380.845 2200.855 3381.490 2201.025 ;
        RECT 3380.500 2200.685 3380.670 2200.805 ;
        RECT 3380.500 2200.515 3381.150 2200.685 ;
      LAYER li1 ;
        RECT 3379.125 2200.030 3380.500 2200.370 ;
      LAYER li1 ;
        RECT 3380.670 2200.355 3381.150 2200.515 ;
        RECT 3381.320 2200.620 3381.490 2200.855 ;
        RECT 3382.030 2201.615 3383.050 2201.945 ;
        RECT 3383.220 2201.895 3383.390 2202.125 ;
        RECT 3385.940 2201.895 3386.110 2202.125 ;
        RECT 3382.030 2201.105 3382.200 2201.615 ;
        RECT 3383.220 2201.565 3383.390 2201.725 ;
        RECT 3385.940 2201.565 3386.110 2201.725 ;
        RECT 3383.220 2201.445 3384.540 2201.565 ;
        RECT 3382.420 2201.435 3384.540 2201.445 ;
        RECT 3382.420 2201.275 3383.220 2201.435 ;
        RECT 3383.390 2201.265 3384.540 2201.435 ;
        RECT 3383.220 2201.235 3384.540 2201.265 ;
        RECT 3385.140 2201.435 3386.110 2201.565 ;
        RECT 3385.140 2201.265 3385.940 2201.435 ;
        RECT 3385.140 2201.235 3386.110 2201.265 ;
        RECT 3382.030 2200.775 3383.050 2201.105 ;
        RECT 3383.220 2200.975 3383.390 2201.235 ;
        RECT 3385.940 2200.975 3386.110 2201.235 ;
        RECT 3382.030 2200.620 3382.200 2200.775 ;
        RECT 3381.320 2200.445 3382.200 2200.620 ;
        RECT 3383.220 2200.725 3383.390 2200.805 ;
        RECT 3385.940 2200.725 3386.110 2200.805 ;
        RECT 3383.220 2200.605 3384.190 2200.725 ;
        RECT 3382.420 2200.515 3384.190 2200.605 ;
        RECT 3380.500 2200.055 3380.670 2200.345 ;
      LAYER li1 ;
        RECT 3379.955 2196.610 3380.500 2200.030 ;
      LAYER li1 ;
        RECT 3380.500 2199.845 3380.670 2199.885 ;
        RECT 3380.500 2199.595 3381.150 2199.845 ;
        RECT 3380.670 2199.515 3381.150 2199.595 ;
        RECT 3380.500 2199.135 3380.670 2199.425 ;
        RECT 3380.670 2198.965 3381.150 2199.005 ;
        RECT 3380.500 2198.675 3381.150 2198.965 ;
        RECT 3380.500 2198.215 3380.670 2198.505 ;
        RECT 3380.670 2198.045 3381.150 2198.165 ;
        RECT 3380.500 2197.835 3381.150 2198.045 ;
        RECT 3381.660 2197.995 3381.830 2200.445 ;
        RECT 3382.420 2200.435 3383.220 2200.515 ;
        RECT 3383.390 2200.395 3384.190 2200.515 ;
        RECT 3383.220 2200.055 3383.390 2200.345 ;
        RECT 3383.220 2199.845 3384.190 2199.885 ;
        RECT 3382.420 2199.595 3384.190 2199.845 ;
        RECT 3382.420 2199.515 3383.220 2199.595 ;
        RECT 3383.390 2199.555 3384.190 2199.595 ;
        RECT 3383.220 2199.135 3383.390 2199.425 ;
        RECT 3382.420 2198.965 3383.220 2199.005 ;
        RECT 3383.390 2198.965 3384.190 2199.045 ;
        RECT 3382.420 2198.715 3384.190 2198.965 ;
        RECT 3382.420 2198.675 3383.390 2198.715 ;
        RECT 3383.220 2198.215 3383.390 2198.505 ;
        RECT 3382.420 2198.045 3383.220 2198.165 ;
        RECT 3383.390 2198.045 3384.190 2198.125 ;
        RECT 3384.780 2198.115 3384.950 2200.565 ;
        RECT 3385.460 2200.515 3386.110 2200.725 ;
        RECT 3385.460 2200.395 3385.940 2200.515 ;
        RECT 3385.940 2200.055 3386.110 2200.345 ;
        RECT 3385.460 2199.595 3386.110 2199.885 ;
        RECT 3385.460 2199.555 3385.940 2199.595 ;
        RECT 3385.940 2199.135 3386.110 2199.425 ;
        RECT 3385.460 2198.965 3385.940 2199.045 ;
        RECT 3385.460 2198.715 3386.110 2198.965 ;
        RECT 3385.940 2198.675 3386.110 2198.715 ;
        RECT 3385.940 2198.215 3386.110 2198.505 ;
        RECT 3382.420 2197.955 3384.190 2198.045 ;
        RECT 3382.420 2197.835 3383.390 2197.955 ;
        RECT 3380.500 2197.755 3380.670 2197.835 ;
        RECT 3383.220 2197.755 3383.390 2197.835 ;
        RECT 3384.410 2197.940 3385.290 2198.115 ;
        RECT 3384.410 2197.785 3384.580 2197.940 ;
        RECT 3380.500 2197.325 3380.670 2197.585 ;
        RECT 3383.220 2197.325 3383.390 2197.585 ;
        RECT 3383.560 2197.455 3384.580 2197.785 ;
        RECT 3380.500 2197.295 3381.470 2197.325 ;
        RECT 3380.670 2197.125 3381.470 2197.295 ;
        RECT 3380.500 2196.995 3381.470 2197.125 ;
        RECT 3382.070 2197.295 3383.390 2197.325 ;
        RECT 3382.070 2197.125 3383.220 2197.295 ;
        RECT 3383.390 2197.125 3384.190 2197.285 ;
        RECT 3382.070 2197.115 3384.190 2197.125 ;
        RECT 3382.070 2196.995 3383.390 2197.115 ;
        RECT 3380.500 2196.835 3380.670 2196.995 ;
        RECT 3383.220 2196.835 3383.390 2196.995 ;
        RECT 3384.410 2196.945 3384.580 2197.455 ;
        RECT 3377.780 2196.435 3377.950 2196.520 ;
        RECT 3380.500 2196.435 3380.670 2196.665 ;
        RECT 3383.220 2196.435 3383.390 2196.665 ;
        RECT 3383.560 2196.615 3384.580 2196.945 ;
        RECT 3385.120 2197.705 3385.290 2197.940 ;
        RECT 3385.460 2198.045 3385.940 2198.205 ;
        RECT 3385.460 2197.875 3386.110 2198.045 ;
        RECT 3385.940 2197.755 3386.110 2197.875 ;
        RECT 3385.120 2197.535 3385.765 2197.705 ;
        RECT 3385.120 2196.865 3385.290 2197.535 ;
        RECT 3385.940 2197.365 3386.110 2197.585 ;
        RECT 3385.460 2197.295 3386.110 2197.365 ;
        RECT 3385.460 2197.125 3385.940 2197.295 ;
        RECT 3385.460 2197.035 3386.110 2197.125 ;
        RECT 3385.120 2196.695 3385.770 2196.865 ;
        RECT 3385.940 2196.835 3386.110 2197.035 ;
        RECT 3385.940 2196.435 3386.110 2196.665 ;
        RECT 3377.780 2196.375 3379.115 2196.435 ;
        RECT 3377.950 2196.205 3379.115 2196.375 ;
        RECT 3377.780 2196.145 3379.115 2196.205 ;
        RECT 3379.775 2196.375 3381.395 2196.435 ;
        RECT 3379.775 2196.205 3380.500 2196.375 ;
        RECT 3380.670 2196.205 3381.395 2196.375 ;
        RECT 3379.775 2196.145 3381.395 2196.205 ;
        RECT 3382.055 2196.375 3384.555 2196.435 ;
        RECT 3382.055 2196.205 3383.220 2196.375 ;
        RECT 3383.390 2196.205 3384.555 2196.375 ;
        RECT 3382.055 2196.145 3384.555 2196.205 ;
        RECT 3385.215 2196.375 3386.110 2196.435 ;
        RECT 3385.215 2196.205 3385.940 2196.375 ;
        RECT 3385.215 2196.145 3386.110 2196.205 ;
        RECT 3377.780 2196.060 3377.950 2196.145 ;
        RECT 3380.500 2196.060 3380.670 2196.145 ;
        RECT 3383.220 2196.060 3383.390 2196.145 ;
        RECT 3385.940 2196.060 3386.110 2196.145 ;
        RECT 201.995 1727.100 202.165 1727.185 ;
        RECT 204.715 1727.100 204.885 1727.185 ;
        RECT 207.435 1727.100 207.605 1727.185 ;
        RECT 210.155 1727.100 210.325 1727.185 ;
        RECT 201.995 1727.040 202.890 1727.100 ;
        RECT 202.165 1726.870 202.890 1727.040 ;
        RECT 201.995 1726.810 202.890 1726.870 ;
        RECT 203.550 1727.040 206.050 1727.100 ;
        RECT 203.550 1726.870 204.715 1727.040 ;
        RECT 204.885 1726.870 206.050 1727.040 ;
        RECT 203.550 1726.810 206.050 1726.870 ;
        RECT 201.995 1726.580 202.165 1726.810 ;
        RECT 204.715 1726.580 204.885 1726.810 ;
        RECT 201.995 1726.250 202.165 1726.410 ;
        RECT 204.715 1726.250 204.885 1726.410 ;
        RECT 205.055 1726.300 206.075 1726.630 ;
        RECT 201.995 1726.120 202.965 1726.250 ;
        RECT 202.165 1725.950 202.965 1726.120 ;
        RECT 201.995 1725.920 202.965 1725.950 ;
        RECT 203.565 1726.130 204.885 1726.250 ;
        RECT 203.565 1726.120 205.685 1726.130 ;
        RECT 203.565 1725.950 204.715 1726.120 ;
        RECT 204.885 1725.960 205.685 1726.120 ;
        RECT 203.565 1725.920 204.885 1725.950 ;
        RECT 201.995 1725.660 202.165 1725.920 ;
      LAYER li1 ;
        RECT 202.335 1725.580 204.545 1725.750 ;
      LAYER li1 ;
        RECT 204.715 1725.660 204.885 1725.920 ;
        RECT 205.905 1725.790 206.075 1726.300 ;
      LAYER li1 ;
        RECT 202.815 1725.495 203.695 1725.580 ;
      LAYER li1 ;
        RECT 201.995 1725.410 202.165 1725.490 ;
        RECT 201.995 1725.200 202.645 1725.410 ;
        RECT 202.165 1725.080 202.645 1725.200 ;
        RECT 201.995 1724.740 202.165 1725.030 ;
      LAYER li1 ;
        RECT 202.815 1724.910 202.985 1725.495 ;
        RECT 202.335 1724.740 202.985 1724.910 ;
      LAYER li1 ;
        RECT 201.995 1724.280 202.645 1724.570 ;
        RECT 202.165 1724.240 202.645 1724.280 ;
        RECT 201.995 1723.820 202.165 1724.110 ;
      LAYER li1 ;
        RECT 202.815 1724.070 202.985 1724.740 ;
        RECT 202.335 1723.900 202.985 1724.070 ;
      LAYER li1 ;
        RECT 202.165 1723.650 202.645 1723.730 ;
        RECT 201.995 1723.400 202.645 1723.650 ;
        RECT 201.995 1723.360 202.165 1723.400 ;
      LAYER li1 ;
        RECT 202.815 1723.230 202.985 1723.900 ;
      LAYER li1 ;
        RECT 201.995 1722.900 202.165 1723.190 ;
      LAYER li1 ;
        RECT 202.335 1723.060 202.985 1723.230 ;
      LAYER li1 ;
        RECT 202.165 1722.730 202.645 1722.890 ;
        RECT 203.155 1722.800 203.325 1725.250 ;
      LAYER li1 ;
        RECT 203.525 1724.910 203.695 1725.495 ;
      LAYER li1 ;
        RECT 204.715 1725.410 204.885 1725.490 ;
        RECT 205.055 1725.460 206.075 1725.790 ;
      LAYER li1 ;
        RECT 206.245 1725.485 206.445 1727.075 ;
      LAYER li1 ;
        RECT 206.710 1727.040 208.330 1727.100 ;
        RECT 206.710 1726.870 207.435 1727.040 ;
        RECT 207.605 1726.870 208.330 1727.040 ;
        RECT 206.710 1726.810 208.330 1726.870 ;
        RECT 208.990 1727.040 210.325 1727.100 ;
        RECT 208.990 1726.870 210.155 1727.040 ;
        RECT 208.990 1726.810 210.325 1726.870 ;
        RECT 207.435 1726.725 207.605 1726.810 ;
        RECT 210.155 1726.725 210.325 1726.810 ;
        RECT 206.615 1726.380 207.265 1726.550 ;
        RECT 206.615 1725.710 206.785 1726.380 ;
        RECT 206.955 1725.880 207.435 1726.210 ;
        RECT 206.615 1725.540 207.260 1725.710 ;
        RECT 203.915 1725.290 204.885 1725.410 ;
        RECT 205.905 1725.305 206.075 1725.460 ;
        RECT 206.615 1725.305 206.785 1725.540 ;
        RECT 203.915 1725.200 205.685 1725.290 ;
        RECT 203.915 1725.080 204.715 1725.200 ;
        RECT 204.885 1725.120 205.685 1725.200 ;
        RECT 205.905 1725.130 206.785 1725.305 ;
      LAYER li1 ;
        RECT 203.525 1724.740 204.545 1724.910 ;
      LAYER li1 ;
        RECT 204.715 1724.740 204.885 1725.030 ;
      LAYER li1 ;
        RECT 203.525 1724.070 203.695 1724.740 ;
        RECT 205.055 1724.700 206.075 1724.870 ;
      LAYER li1 ;
        RECT 203.915 1724.530 204.885 1724.570 ;
        RECT 203.915 1724.280 205.685 1724.530 ;
        RECT 203.915 1724.240 204.715 1724.280 ;
        RECT 204.885 1724.200 205.685 1724.280 ;
      LAYER li1 ;
        RECT 203.525 1723.900 204.545 1724.070 ;
        RECT 203.525 1723.230 203.695 1723.900 ;
      LAYER li1 ;
        RECT 204.715 1723.820 204.885 1724.110 ;
      LAYER li1 ;
        RECT 205.905 1724.030 206.075 1724.700 ;
        RECT 205.055 1723.860 206.075 1724.030 ;
      LAYER li1 ;
        RECT 203.915 1723.650 204.715 1723.730 ;
        RECT 204.885 1723.650 205.685 1723.690 ;
        RECT 203.915 1723.400 205.685 1723.650 ;
        RECT 204.715 1723.360 205.685 1723.400 ;
      LAYER li1 ;
        RECT 203.525 1723.060 204.545 1723.230 ;
        RECT 205.905 1723.190 206.075 1723.860 ;
      LAYER li1 ;
        RECT 204.715 1722.900 204.885 1723.190 ;
      LAYER li1 ;
        RECT 205.055 1723.020 206.075 1723.190 ;
      LAYER li1 ;
        RECT 201.995 1722.560 202.645 1722.730 ;
        RECT 202.815 1722.625 203.695 1722.800 ;
        RECT 203.915 1722.730 204.715 1722.810 ;
        RECT 204.885 1722.730 205.685 1722.850 ;
        RECT 203.915 1722.640 205.685 1722.730 ;
        RECT 201.995 1722.440 202.165 1722.560 ;
        RECT 202.815 1722.390 202.985 1722.625 ;
        RECT 203.525 1722.470 203.695 1722.625 ;
        RECT 204.715 1722.520 205.685 1722.640 ;
        RECT 201.995 1722.050 202.165 1722.270 ;
        RECT 202.340 1722.220 202.985 1722.390 ;
        RECT 201.995 1721.980 202.645 1722.050 ;
        RECT 202.165 1721.810 202.645 1721.980 ;
        RECT 201.995 1721.720 202.645 1721.810 ;
        RECT 201.995 1721.520 202.165 1721.720 ;
        RECT 202.815 1721.550 202.985 1722.220 ;
        RECT 202.335 1721.380 202.985 1721.550 ;
        RECT 201.995 1721.120 202.165 1721.350 ;
      LAYER li1 ;
        RECT 203.155 1721.345 203.355 1722.445 ;
      LAYER li1 ;
        RECT 203.525 1722.140 204.545 1722.470 ;
        RECT 204.715 1722.440 204.885 1722.520 ;
      LAYER li1 ;
        RECT 205.905 1722.435 206.075 1723.020 ;
      LAYER li1 ;
        RECT 206.275 1722.680 206.445 1725.130 ;
        RECT 206.955 1725.040 207.435 1725.370 ;
      LAYER li1 ;
        RECT 206.615 1724.700 207.265 1724.870 ;
        RECT 206.615 1724.030 206.785 1724.700 ;
      LAYER li1 ;
        RECT 206.955 1724.200 207.435 1724.530 ;
      LAYER li1 ;
        RECT 206.615 1723.860 207.265 1724.030 ;
        RECT 206.615 1723.190 206.785 1723.860 ;
      LAYER li1 ;
        RECT 206.955 1723.360 207.435 1723.690 ;
      LAYER li1 ;
        RECT 206.615 1723.020 207.265 1723.190 ;
        RECT 206.615 1722.435 206.785 1723.020 ;
      LAYER li1 ;
        RECT 206.955 1722.520 207.435 1722.850 ;
      LAYER li1 ;
        RECT 205.905 1722.350 206.785 1722.435 ;
      LAYER li1 ;
        RECT 203.525 1721.630 203.695 1722.140 ;
        RECT 204.715 1722.010 204.885 1722.270 ;
      LAYER li1 ;
        RECT 205.055 1722.180 207.265 1722.350 ;
      LAYER li1 ;
        RECT 204.715 1721.980 206.035 1722.010 ;
        RECT 203.915 1721.810 204.715 1721.970 ;
        RECT 204.885 1721.810 206.035 1721.980 ;
        RECT 203.915 1721.800 206.035 1721.810 ;
        RECT 204.715 1721.680 206.035 1721.800 ;
        RECT 206.635 1721.680 207.435 1722.010 ;
        RECT 203.525 1721.300 204.545 1721.630 ;
        RECT 204.715 1721.520 204.885 1721.680 ;
        RECT 204.715 1721.120 204.885 1721.350 ;
        RECT 207.435 1721.120 207.605 1721.205 ;
        RECT 210.155 1721.120 210.325 1721.205 ;
        RECT 201.995 1721.060 202.890 1721.120 ;
        RECT 202.165 1720.890 202.890 1721.060 ;
        RECT 201.995 1720.830 202.890 1720.890 ;
        RECT 203.550 1721.060 206.050 1721.120 ;
        RECT 203.550 1720.890 204.715 1721.060 ;
        RECT 204.885 1720.890 206.050 1721.060 ;
        RECT 203.550 1720.830 206.050 1720.890 ;
        RECT 201.995 1720.600 202.165 1720.830 ;
        RECT 204.715 1720.600 204.885 1720.830 ;
        RECT 201.995 1720.270 202.165 1720.430 ;
        RECT 204.715 1720.270 204.885 1720.430 ;
        RECT 205.055 1720.320 206.075 1720.650 ;
        RECT 201.995 1720.140 202.965 1720.270 ;
        RECT 202.165 1719.970 202.965 1720.140 ;
        RECT 201.995 1719.940 202.965 1719.970 ;
        RECT 203.565 1720.150 204.885 1720.270 ;
        RECT 203.565 1720.140 205.685 1720.150 ;
        RECT 203.565 1719.970 204.715 1720.140 ;
        RECT 204.885 1719.980 205.685 1720.140 ;
        RECT 203.565 1719.940 204.885 1719.970 ;
        RECT 201.995 1719.680 202.165 1719.940 ;
      LAYER li1 ;
        RECT 202.335 1719.600 204.545 1719.770 ;
      LAYER li1 ;
        RECT 204.715 1719.680 204.885 1719.940 ;
        RECT 205.905 1719.810 206.075 1720.320 ;
      LAYER li1 ;
        RECT 202.815 1719.515 203.695 1719.600 ;
      LAYER li1 ;
        RECT 201.995 1719.430 202.165 1719.510 ;
        RECT 201.995 1719.220 202.645 1719.430 ;
        RECT 202.165 1719.100 202.645 1719.220 ;
        RECT 201.995 1718.760 202.165 1719.050 ;
      LAYER li1 ;
        RECT 202.815 1718.930 202.985 1719.515 ;
        RECT 202.335 1718.760 202.985 1718.930 ;
      LAYER li1 ;
        RECT 201.995 1718.300 202.645 1718.590 ;
        RECT 202.165 1718.260 202.645 1718.300 ;
        RECT 201.995 1717.840 202.165 1718.130 ;
      LAYER li1 ;
        RECT 202.815 1718.090 202.985 1718.760 ;
        RECT 202.335 1717.920 202.985 1718.090 ;
      LAYER li1 ;
        RECT 202.165 1717.670 202.645 1717.750 ;
        RECT 201.995 1717.420 202.645 1717.670 ;
        RECT 201.995 1717.380 202.165 1717.420 ;
      LAYER li1 ;
        RECT 202.815 1717.250 202.985 1717.920 ;
      LAYER li1 ;
        RECT 201.995 1716.920 202.165 1717.210 ;
      LAYER li1 ;
        RECT 202.335 1717.080 202.985 1717.250 ;
      LAYER li1 ;
        RECT 202.165 1716.750 202.645 1716.910 ;
        RECT 203.155 1716.820 203.325 1719.270 ;
      LAYER li1 ;
        RECT 203.525 1718.930 203.695 1719.515 ;
      LAYER li1 ;
        RECT 204.715 1719.430 204.885 1719.510 ;
        RECT 205.055 1719.480 206.075 1719.810 ;
      LAYER li1 ;
        RECT 206.245 1719.505 206.445 1721.095 ;
      LAYER li1 ;
        RECT 206.710 1721.060 208.330 1721.120 ;
        RECT 206.710 1720.890 207.435 1721.060 ;
        RECT 207.605 1720.890 208.330 1721.060 ;
        RECT 206.710 1720.830 208.330 1720.890 ;
        RECT 208.990 1721.060 210.325 1721.120 ;
        RECT 208.990 1720.890 210.155 1721.060 ;
        RECT 208.990 1720.830 210.325 1720.890 ;
        RECT 207.435 1720.745 207.605 1720.830 ;
        RECT 210.155 1720.745 210.325 1720.830 ;
        RECT 206.615 1720.400 207.265 1720.570 ;
        RECT 206.615 1719.730 206.785 1720.400 ;
        RECT 206.955 1719.900 207.435 1720.230 ;
        RECT 206.615 1719.560 207.260 1719.730 ;
        RECT 203.915 1719.310 204.885 1719.430 ;
        RECT 205.905 1719.325 206.075 1719.480 ;
        RECT 206.615 1719.325 206.785 1719.560 ;
        RECT 203.915 1719.220 205.685 1719.310 ;
        RECT 203.915 1719.100 204.715 1719.220 ;
        RECT 204.885 1719.140 205.685 1719.220 ;
        RECT 205.905 1719.150 206.785 1719.325 ;
      LAYER li1 ;
        RECT 203.525 1718.760 204.545 1718.930 ;
      LAYER li1 ;
        RECT 204.715 1718.760 204.885 1719.050 ;
      LAYER li1 ;
        RECT 203.525 1718.090 203.695 1718.760 ;
        RECT 205.055 1718.720 206.075 1718.890 ;
      LAYER li1 ;
        RECT 203.915 1718.550 204.885 1718.590 ;
        RECT 203.915 1718.300 205.685 1718.550 ;
        RECT 203.915 1718.260 204.715 1718.300 ;
        RECT 204.885 1718.220 205.685 1718.300 ;
      LAYER li1 ;
        RECT 203.525 1717.920 204.545 1718.090 ;
        RECT 203.525 1717.250 203.695 1717.920 ;
      LAYER li1 ;
        RECT 204.715 1717.840 204.885 1718.130 ;
      LAYER li1 ;
        RECT 205.905 1718.050 206.075 1718.720 ;
        RECT 205.055 1717.880 206.075 1718.050 ;
      LAYER li1 ;
        RECT 203.915 1717.670 204.715 1717.750 ;
        RECT 204.885 1717.670 205.685 1717.710 ;
        RECT 203.915 1717.420 205.685 1717.670 ;
        RECT 204.715 1717.380 205.685 1717.420 ;
      LAYER li1 ;
        RECT 203.525 1717.080 204.545 1717.250 ;
        RECT 205.905 1717.210 206.075 1717.880 ;
      LAYER li1 ;
        RECT 204.715 1716.920 204.885 1717.210 ;
      LAYER li1 ;
        RECT 205.055 1717.040 206.075 1717.210 ;
      LAYER li1 ;
        RECT 201.995 1716.580 202.645 1716.750 ;
        RECT 202.815 1716.645 203.695 1716.820 ;
        RECT 203.915 1716.750 204.715 1716.830 ;
        RECT 204.885 1716.750 205.685 1716.870 ;
        RECT 203.915 1716.660 205.685 1716.750 ;
        RECT 201.995 1716.460 202.165 1716.580 ;
        RECT 202.815 1716.410 202.985 1716.645 ;
        RECT 203.525 1716.490 203.695 1716.645 ;
        RECT 204.715 1716.540 205.685 1716.660 ;
        RECT 201.995 1716.070 202.165 1716.290 ;
        RECT 202.340 1716.240 202.985 1716.410 ;
        RECT 201.995 1716.000 202.645 1716.070 ;
        RECT 202.165 1715.830 202.645 1716.000 ;
        RECT 201.995 1715.740 202.645 1715.830 ;
        RECT 201.995 1715.540 202.165 1715.740 ;
        RECT 202.815 1715.570 202.985 1716.240 ;
        RECT 202.335 1715.400 202.985 1715.570 ;
        RECT 201.995 1715.140 202.165 1715.370 ;
      LAYER li1 ;
        RECT 203.155 1715.365 203.355 1716.465 ;
      LAYER li1 ;
        RECT 203.525 1716.160 204.545 1716.490 ;
        RECT 204.715 1716.460 204.885 1716.540 ;
      LAYER li1 ;
        RECT 205.905 1716.455 206.075 1717.040 ;
      LAYER li1 ;
        RECT 206.275 1716.700 206.445 1719.150 ;
        RECT 206.955 1719.060 207.435 1719.390 ;
      LAYER li1 ;
        RECT 206.615 1718.720 207.265 1718.890 ;
        RECT 206.615 1718.050 206.785 1718.720 ;
      LAYER li1 ;
        RECT 206.955 1718.220 207.435 1718.550 ;
      LAYER li1 ;
        RECT 206.615 1717.880 207.265 1718.050 ;
        RECT 206.615 1717.210 206.785 1717.880 ;
      LAYER li1 ;
        RECT 206.955 1717.380 207.435 1717.710 ;
      LAYER li1 ;
        RECT 206.615 1717.040 207.265 1717.210 ;
        RECT 206.615 1716.455 206.785 1717.040 ;
      LAYER li1 ;
        RECT 206.955 1716.540 207.435 1716.870 ;
      LAYER li1 ;
        RECT 205.905 1716.370 206.785 1716.455 ;
      LAYER li1 ;
        RECT 203.525 1715.650 203.695 1716.160 ;
        RECT 204.715 1716.030 204.885 1716.290 ;
      LAYER li1 ;
        RECT 205.055 1716.200 207.265 1716.370 ;
      LAYER li1 ;
        RECT 204.715 1716.000 206.035 1716.030 ;
        RECT 203.915 1715.830 204.715 1715.990 ;
        RECT 204.885 1715.830 206.035 1716.000 ;
        RECT 203.915 1715.820 206.035 1715.830 ;
        RECT 204.715 1715.700 206.035 1715.820 ;
        RECT 206.635 1715.700 207.435 1716.030 ;
        RECT 203.525 1715.320 204.545 1715.650 ;
        RECT 204.715 1715.540 204.885 1715.700 ;
        RECT 204.715 1715.140 204.885 1715.370 ;
        RECT 207.435 1715.140 207.605 1715.225 ;
        RECT 210.155 1715.140 210.325 1715.225 ;
        RECT 201.995 1715.080 202.890 1715.140 ;
        RECT 202.165 1714.910 202.890 1715.080 ;
        RECT 201.995 1714.850 202.890 1714.910 ;
        RECT 203.550 1715.080 206.050 1715.140 ;
        RECT 203.550 1714.910 204.715 1715.080 ;
        RECT 204.885 1714.910 206.050 1715.080 ;
        RECT 203.550 1714.850 206.050 1714.910 ;
        RECT 201.995 1714.620 202.165 1714.850 ;
        RECT 204.715 1714.620 204.885 1714.850 ;
        RECT 201.995 1714.290 202.165 1714.450 ;
        RECT 204.715 1714.290 204.885 1714.450 ;
        RECT 205.055 1714.340 206.075 1714.670 ;
        RECT 201.995 1714.160 202.965 1714.290 ;
        RECT 202.165 1713.990 202.965 1714.160 ;
        RECT 201.995 1713.960 202.965 1713.990 ;
        RECT 203.565 1714.170 204.885 1714.290 ;
        RECT 203.565 1714.160 205.685 1714.170 ;
        RECT 203.565 1713.990 204.715 1714.160 ;
        RECT 204.885 1714.000 205.685 1714.160 ;
        RECT 203.565 1713.960 204.885 1713.990 ;
        RECT 201.995 1713.700 202.165 1713.960 ;
      LAYER li1 ;
        RECT 202.335 1713.620 204.545 1713.790 ;
      LAYER li1 ;
        RECT 204.715 1713.700 204.885 1713.960 ;
        RECT 205.905 1713.830 206.075 1714.340 ;
      LAYER li1 ;
        RECT 202.815 1713.535 203.695 1713.620 ;
      LAYER li1 ;
        RECT 201.995 1713.450 202.165 1713.530 ;
        RECT 201.995 1713.240 202.645 1713.450 ;
        RECT 202.165 1713.120 202.645 1713.240 ;
        RECT 201.995 1712.780 202.165 1713.070 ;
      LAYER li1 ;
        RECT 202.815 1712.950 202.985 1713.535 ;
        RECT 202.335 1712.780 202.985 1712.950 ;
      LAYER li1 ;
        RECT 201.995 1712.320 202.645 1712.610 ;
        RECT 202.165 1712.280 202.645 1712.320 ;
        RECT 201.995 1711.860 202.165 1712.150 ;
      LAYER li1 ;
        RECT 202.815 1712.110 202.985 1712.780 ;
        RECT 202.335 1711.940 202.985 1712.110 ;
      LAYER li1 ;
        RECT 202.165 1711.690 202.645 1711.770 ;
        RECT 201.995 1711.440 202.645 1711.690 ;
        RECT 201.995 1711.400 202.165 1711.440 ;
      LAYER li1 ;
        RECT 202.815 1711.270 202.985 1711.940 ;
      LAYER li1 ;
        RECT 201.995 1710.940 202.165 1711.230 ;
      LAYER li1 ;
        RECT 202.335 1711.100 202.985 1711.270 ;
      LAYER li1 ;
        RECT 202.165 1710.770 202.645 1710.930 ;
        RECT 203.155 1710.840 203.325 1713.290 ;
      LAYER li1 ;
        RECT 203.525 1712.950 203.695 1713.535 ;
      LAYER li1 ;
        RECT 204.715 1713.450 204.885 1713.530 ;
        RECT 205.055 1713.500 206.075 1713.830 ;
      LAYER li1 ;
        RECT 206.245 1713.525 206.445 1715.115 ;
      LAYER li1 ;
        RECT 206.710 1715.080 208.330 1715.140 ;
        RECT 206.710 1714.910 207.435 1715.080 ;
        RECT 207.605 1714.910 208.330 1715.080 ;
        RECT 206.710 1714.850 208.330 1714.910 ;
        RECT 208.990 1715.080 210.325 1715.140 ;
        RECT 208.990 1714.910 210.155 1715.080 ;
        RECT 208.990 1714.850 210.325 1714.910 ;
        RECT 207.435 1714.765 207.605 1714.850 ;
        RECT 210.155 1714.765 210.325 1714.850 ;
        RECT 206.615 1714.420 207.265 1714.590 ;
        RECT 206.615 1713.750 206.785 1714.420 ;
        RECT 206.955 1713.920 207.435 1714.250 ;
        RECT 206.615 1713.580 207.260 1713.750 ;
        RECT 203.915 1713.330 204.885 1713.450 ;
        RECT 205.905 1713.345 206.075 1713.500 ;
        RECT 206.615 1713.345 206.785 1713.580 ;
        RECT 203.915 1713.240 205.685 1713.330 ;
        RECT 203.915 1713.120 204.715 1713.240 ;
        RECT 204.885 1713.160 205.685 1713.240 ;
        RECT 205.905 1713.170 206.785 1713.345 ;
      LAYER li1 ;
        RECT 203.525 1712.780 204.545 1712.950 ;
      LAYER li1 ;
        RECT 204.715 1712.780 204.885 1713.070 ;
      LAYER li1 ;
        RECT 203.525 1712.110 203.695 1712.780 ;
        RECT 205.055 1712.740 206.075 1712.910 ;
      LAYER li1 ;
        RECT 203.915 1712.570 204.885 1712.610 ;
        RECT 203.915 1712.320 205.685 1712.570 ;
        RECT 203.915 1712.280 204.715 1712.320 ;
        RECT 204.885 1712.240 205.685 1712.320 ;
      LAYER li1 ;
        RECT 203.525 1711.940 204.545 1712.110 ;
        RECT 203.525 1711.270 203.695 1711.940 ;
      LAYER li1 ;
        RECT 204.715 1711.860 204.885 1712.150 ;
      LAYER li1 ;
        RECT 205.905 1712.070 206.075 1712.740 ;
        RECT 205.055 1711.900 206.075 1712.070 ;
      LAYER li1 ;
        RECT 203.915 1711.690 204.715 1711.770 ;
        RECT 204.885 1711.690 205.685 1711.730 ;
        RECT 203.915 1711.440 205.685 1711.690 ;
        RECT 204.715 1711.400 205.685 1711.440 ;
      LAYER li1 ;
        RECT 203.525 1711.100 204.545 1711.270 ;
        RECT 205.905 1711.230 206.075 1711.900 ;
      LAYER li1 ;
        RECT 204.715 1710.940 204.885 1711.230 ;
      LAYER li1 ;
        RECT 205.055 1711.060 206.075 1711.230 ;
      LAYER li1 ;
        RECT 201.995 1710.600 202.645 1710.770 ;
        RECT 202.815 1710.665 203.695 1710.840 ;
        RECT 203.915 1710.770 204.715 1710.850 ;
        RECT 204.885 1710.770 205.685 1710.890 ;
        RECT 203.915 1710.680 205.685 1710.770 ;
        RECT 201.995 1710.480 202.165 1710.600 ;
        RECT 202.815 1710.430 202.985 1710.665 ;
        RECT 203.525 1710.510 203.695 1710.665 ;
        RECT 204.715 1710.560 205.685 1710.680 ;
        RECT 201.995 1710.090 202.165 1710.310 ;
        RECT 202.340 1710.260 202.985 1710.430 ;
        RECT 201.995 1710.020 202.645 1710.090 ;
        RECT 202.165 1709.850 202.645 1710.020 ;
        RECT 201.995 1709.760 202.645 1709.850 ;
        RECT 201.995 1709.560 202.165 1709.760 ;
        RECT 202.815 1709.590 202.985 1710.260 ;
        RECT 202.335 1709.420 202.985 1709.590 ;
        RECT 201.995 1709.160 202.165 1709.390 ;
      LAYER li1 ;
        RECT 203.155 1709.385 203.355 1710.485 ;
      LAYER li1 ;
        RECT 203.525 1710.180 204.545 1710.510 ;
        RECT 204.715 1710.480 204.885 1710.560 ;
      LAYER li1 ;
        RECT 205.905 1710.475 206.075 1711.060 ;
      LAYER li1 ;
        RECT 206.275 1710.720 206.445 1713.170 ;
        RECT 206.955 1713.080 207.435 1713.410 ;
      LAYER li1 ;
        RECT 206.615 1712.740 207.265 1712.910 ;
        RECT 206.615 1712.070 206.785 1712.740 ;
      LAYER li1 ;
        RECT 206.955 1712.240 207.435 1712.570 ;
      LAYER li1 ;
        RECT 206.615 1711.900 207.265 1712.070 ;
        RECT 206.615 1711.230 206.785 1711.900 ;
      LAYER li1 ;
        RECT 206.955 1711.400 207.435 1711.730 ;
      LAYER li1 ;
        RECT 206.615 1711.060 207.265 1711.230 ;
        RECT 206.615 1710.475 206.785 1711.060 ;
      LAYER li1 ;
        RECT 206.955 1710.560 207.435 1710.890 ;
      LAYER li1 ;
        RECT 205.905 1710.390 206.785 1710.475 ;
      LAYER li1 ;
        RECT 203.525 1709.670 203.695 1710.180 ;
        RECT 204.715 1710.050 204.885 1710.310 ;
      LAYER li1 ;
        RECT 205.055 1710.220 207.265 1710.390 ;
      LAYER li1 ;
        RECT 204.715 1710.020 206.035 1710.050 ;
        RECT 203.915 1709.850 204.715 1710.010 ;
        RECT 204.885 1709.850 206.035 1710.020 ;
        RECT 203.915 1709.840 206.035 1709.850 ;
        RECT 204.715 1709.720 206.035 1709.840 ;
        RECT 206.635 1709.720 207.435 1710.050 ;
        RECT 203.525 1709.340 204.545 1709.670 ;
        RECT 204.715 1709.560 204.885 1709.720 ;
        RECT 204.715 1709.160 204.885 1709.390 ;
        RECT 207.435 1709.160 207.605 1709.245 ;
        RECT 210.155 1709.160 210.325 1709.245 ;
        RECT 201.995 1709.100 202.890 1709.160 ;
        RECT 202.165 1708.930 202.890 1709.100 ;
        RECT 201.995 1708.870 202.890 1708.930 ;
        RECT 203.550 1709.100 206.050 1709.160 ;
        RECT 203.550 1708.930 204.715 1709.100 ;
        RECT 204.885 1708.930 206.050 1709.100 ;
        RECT 203.550 1708.870 206.050 1708.930 ;
        RECT 201.995 1708.640 202.165 1708.870 ;
        RECT 204.715 1708.640 204.885 1708.870 ;
        RECT 201.995 1708.310 202.165 1708.470 ;
        RECT 204.715 1708.310 204.885 1708.470 ;
        RECT 205.055 1708.360 206.075 1708.690 ;
        RECT 201.995 1708.180 202.965 1708.310 ;
        RECT 202.165 1708.010 202.965 1708.180 ;
        RECT 201.995 1707.980 202.965 1708.010 ;
        RECT 203.565 1708.190 204.885 1708.310 ;
        RECT 203.565 1708.180 205.685 1708.190 ;
        RECT 203.565 1708.010 204.715 1708.180 ;
        RECT 204.885 1708.020 205.685 1708.180 ;
        RECT 203.565 1707.980 204.885 1708.010 ;
        RECT 201.995 1707.720 202.165 1707.980 ;
      LAYER li1 ;
        RECT 202.335 1707.640 204.545 1707.810 ;
      LAYER li1 ;
        RECT 204.715 1707.720 204.885 1707.980 ;
        RECT 205.905 1707.850 206.075 1708.360 ;
      LAYER li1 ;
        RECT 202.815 1707.555 203.695 1707.640 ;
      LAYER li1 ;
        RECT 201.995 1707.470 202.165 1707.550 ;
        RECT 201.995 1707.260 202.645 1707.470 ;
        RECT 202.165 1707.140 202.645 1707.260 ;
        RECT 201.995 1706.800 202.165 1707.090 ;
      LAYER li1 ;
        RECT 202.815 1706.970 202.985 1707.555 ;
        RECT 202.335 1706.800 202.985 1706.970 ;
      LAYER li1 ;
        RECT 201.995 1706.340 202.645 1706.630 ;
        RECT 202.165 1706.300 202.645 1706.340 ;
        RECT 201.995 1705.880 202.165 1706.170 ;
      LAYER li1 ;
        RECT 202.815 1706.130 202.985 1706.800 ;
        RECT 202.335 1705.960 202.985 1706.130 ;
      LAYER li1 ;
        RECT 202.165 1705.710 202.645 1705.790 ;
        RECT 201.995 1705.460 202.645 1705.710 ;
        RECT 201.995 1705.420 202.165 1705.460 ;
      LAYER li1 ;
        RECT 202.815 1705.290 202.985 1705.960 ;
      LAYER li1 ;
        RECT 201.995 1704.960 202.165 1705.250 ;
      LAYER li1 ;
        RECT 202.335 1705.120 202.985 1705.290 ;
      LAYER li1 ;
        RECT 202.165 1704.790 202.645 1704.950 ;
        RECT 203.155 1704.860 203.325 1707.310 ;
      LAYER li1 ;
        RECT 203.525 1706.970 203.695 1707.555 ;
      LAYER li1 ;
        RECT 204.715 1707.470 204.885 1707.550 ;
        RECT 205.055 1707.520 206.075 1707.850 ;
      LAYER li1 ;
        RECT 206.245 1707.545 206.445 1709.135 ;
      LAYER li1 ;
        RECT 206.710 1709.100 208.330 1709.160 ;
        RECT 206.710 1708.930 207.435 1709.100 ;
        RECT 207.605 1708.930 208.330 1709.100 ;
        RECT 206.710 1708.870 208.330 1708.930 ;
        RECT 208.990 1709.100 210.325 1709.160 ;
        RECT 208.990 1708.930 210.155 1709.100 ;
        RECT 208.990 1708.870 210.325 1708.930 ;
        RECT 207.435 1708.785 207.605 1708.870 ;
        RECT 210.155 1708.785 210.325 1708.870 ;
        RECT 206.615 1708.440 207.265 1708.610 ;
        RECT 206.615 1707.770 206.785 1708.440 ;
        RECT 206.955 1707.940 207.435 1708.270 ;
        RECT 206.615 1707.600 207.260 1707.770 ;
        RECT 203.915 1707.350 204.885 1707.470 ;
        RECT 205.905 1707.365 206.075 1707.520 ;
        RECT 206.615 1707.365 206.785 1707.600 ;
        RECT 203.915 1707.260 205.685 1707.350 ;
        RECT 203.915 1707.140 204.715 1707.260 ;
        RECT 204.885 1707.180 205.685 1707.260 ;
        RECT 205.905 1707.190 206.785 1707.365 ;
      LAYER li1 ;
        RECT 203.525 1706.800 204.545 1706.970 ;
      LAYER li1 ;
        RECT 204.715 1706.800 204.885 1707.090 ;
      LAYER li1 ;
        RECT 203.525 1706.130 203.695 1706.800 ;
        RECT 205.055 1706.760 206.075 1706.930 ;
      LAYER li1 ;
        RECT 203.915 1706.590 204.885 1706.630 ;
        RECT 203.915 1706.340 205.685 1706.590 ;
        RECT 203.915 1706.300 204.715 1706.340 ;
        RECT 204.885 1706.260 205.685 1706.340 ;
      LAYER li1 ;
        RECT 203.525 1705.960 204.545 1706.130 ;
        RECT 203.525 1705.290 203.695 1705.960 ;
      LAYER li1 ;
        RECT 204.715 1705.880 204.885 1706.170 ;
      LAYER li1 ;
        RECT 205.905 1706.090 206.075 1706.760 ;
        RECT 205.055 1705.920 206.075 1706.090 ;
      LAYER li1 ;
        RECT 203.915 1705.710 204.715 1705.790 ;
        RECT 204.885 1705.710 205.685 1705.750 ;
        RECT 203.915 1705.460 205.685 1705.710 ;
        RECT 204.715 1705.420 205.685 1705.460 ;
      LAYER li1 ;
        RECT 203.525 1705.120 204.545 1705.290 ;
        RECT 205.905 1705.250 206.075 1705.920 ;
      LAYER li1 ;
        RECT 204.715 1704.960 204.885 1705.250 ;
      LAYER li1 ;
        RECT 205.055 1705.080 206.075 1705.250 ;
      LAYER li1 ;
        RECT 201.995 1704.620 202.645 1704.790 ;
        RECT 202.815 1704.685 203.695 1704.860 ;
        RECT 203.915 1704.790 204.715 1704.870 ;
        RECT 204.885 1704.790 205.685 1704.910 ;
        RECT 203.915 1704.700 205.685 1704.790 ;
        RECT 201.995 1704.500 202.165 1704.620 ;
        RECT 202.815 1704.450 202.985 1704.685 ;
        RECT 203.525 1704.530 203.695 1704.685 ;
        RECT 204.715 1704.580 205.685 1704.700 ;
        RECT 201.995 1704.110 202.165 1704.330 ;
        RECT 202.340 1704.280 202.985 1704.450 ;
        RECT 201.995 1704.040 202.645 1704.110 ;
        RECT 202.165 1703.870 202.645 1704.040 ;
        RECT 201.995 1703.780 202.645 1703.870 ;
        RECT 201.995 1703.580 202.165 1703.780 ;
        RECT 202.815 1703.610 202.985 1704.280 ;
        RECT 202.335 1703.440 202.985 1703.610 ;
        RECT 201.995 1703.180 202.165 1703.410 ;
      LAYER li1 ;
        RECT 203.155 1703.405 203.355 1704.505 ;
      LAYER li1 ;
        RECT 203.525 1704.200 204.545 1704.530 ;
        RECT 204.715 1704.500 204.885 1704.580 ;
      LAYER li1 ;
        RECT 205.905 1704.495 206.075 1705.080 ;
      LAYER li1 ;
        RECT 206.275 1704.740 206.445 1707.190 ;
        RECT 206.955 1707.100 207.435 1707.430 ;
      LAYER li1 ;
        RECT 206.615 1706.760 207.265 1706.930 ;
        RECT 206.615 1706.090 206.785 1706.760 ;
      LAYER li1 ;
        RECT 206.955 1706.260 207.435 1706.590 ;
      LAYER li1 ;
        RECT 206.615 1705.920 207.265 1706.090 ;
        RECT 206.615 1705.250 206.785 1705.920 ;
      LAYER li1 ;
        RECT 206.955 1705.420 207.435 1705.750 ;
      LAYER li1 ;
        RECT 206.615 1705.080 207.265 1705.250 ;
        RECT 206.615 1704.495 206.785 1705.080 ;
      LAYER li1 ;
        RECT 206.955 1704.580 207.435 1704.910 ;
      LAYER li1 ;
        RECT 205.905 1704.410 206.785 1704.495 ;
      LAYER li1 ;
        RECT 203.525 1703.690 203.695 1704.200 ;
        RECT 204.715 1704.070 204.885 1704.330 ;
      LAYER li1 ;
        RECT 205.055 1704.240 207.265 1704.410 ;
      LAYER li1 ;
        RECT 204.715 1704.040 206.035 1704.070 ;
        RECT 203.915 1703.870 204.715 1704.030 ;
        RECT 204.885 1703.870 206.035 1704.040 ;
        RECT 203.915 1703.860 206.035 1703.870 ;
        RECT 204.715 1703.740 206.035 1703.860 ;
        RECT 206.635 1703.740 207.435 1704.070 ;
        RECT 203.525 1703.360 204.545 1703.690 ;
        RECT 204.715 1703.580 204.885 1703.740 ;
        RECT 204.715 1703.180 204.885 1703.410 ;
        RECT 207.435 1703.180 207.605 1703.265 ;
        RECT 210.155 1703.180 210.325 1703.265 ;
        RECT 201.995 1703.120 202.890 1703.180 ;
        RECT 202.165 1702.950 202.890 1703.120 ;
        RECT 201.995 1702.890 202.890 1702.950 ;
        RECT 203.550 1703.120 206.050 1703.180 ;
        RECT 203.550 1702.950 204.715 1703.120 ;
        RECT 204.885 1702.950 206.050 1703.120 ;
        RECT 203.550 1702.890 206.050 1702.950 ;
        RECT 201.995 1702.660 202.165 1702.890 ;
        RECT 204.715 1702.660 204.885 1702.890 ;
        RECT 201.995 1702.330 202.165 1702.490 ;
        RECT 204.715 1702.330 204.885 1702.490 ;
        RECT 205.055 1702.380 206.075 1702.710 ;
        RECT 201.995 1702.200 202.965 1702.330 ;
        RECT 202.165 1702.030 202.965 1702.200 ;
        RECT 201.995 1702.000 202.965 1702.030 ;
        RECT 203.565 1702.210 204.885 1702.330 ;
        RECT 203.565 1702.200 205.685 1702.210 ;
        RECT 203.565 1702.030 204.715 1702.200 ;
        RECT 204.885 1702.040 205.685 1702.200 ;
        RECT 203.565 1702.000 204.885 1702.030 ;
        RECT 201.995 1701.740 202.165 1702.000 ;
      LAYER li1 ;
        RECT 202.335 1701.660 204.545 1701.830 ;
      LAYER li1 ;
        RECT 204.715 1701.740 204.885 1702.000 ;
        RECT 205.905 1701.870 206.075 1702.380 ;
      LAYER li1 ;
        RECT 202.815 1701.575 203.695 1701.660 ;
      LAYER li1 ;
        RECT 201.995 1701.490 202.165 1701.570 ;
        RECT 201.995 1701.280 202.645 1701.490 ;
        RECT 202.165 1701.160 202.645 1701.280 ;
        RECT 201.995 1700.820 202.165 1701.110 ;
      LAYER li1 ;
        RECT 202.815 1700.990 202.985 1701.575 ;
        RECT 202.335 1700.820 202.985 1700.990 ;
      LAYER li1 ;
        RECT 201.995 1700.360 202.645 1700.650 ;
        RECT 202.165 1700.320 202.645 1700.360 ;
        RECT 201.995 1699.900 202.165 1700.190 ;
      LAYER li1 ;
        RECT 202.815 1700.150 202.985 1700.820 ;
        RECT 202.335 1699.980 202.985 1700.150 ;
      LAYER li1 ;
        RECT 202.165 1699.730 202.645 1699.810 ;
        RECT 201.995 1699.480 202.645 1699.730 ;
        RECT 201.995 1699.440 202.165 1699.480 ;
      LAYER li1 ;
        RECT 202.815 1699.310 202.985 1699.980 ;
      LAYER li1 ;
        RECT 201.995 1698.980 202.165 1699.270 ;
      LAYER li1 ;
        RECT 202.335 1699.140 202.985 1699.310 ;
      LAYER li1 ;
        RECT 202.165 1698.810 202.645 1698.970 ;
        RECT 203.155 1698.880 203.325 1701.330 ;
      LAYER li1 ;
        RECT 203.525 1700.990 203.695 1701.575 ;
      LAYER li1 ;
        RECT 204.715 1701.490 204.885 1701.570 ;
        RECT 205.055 1701.540 206.075 1701.870 ;
      LAYER li1 ;
        RECT 206.245 1701.565 206.445 1703.155 ;
      LAYER li1 ;
        RECT 206.710 1703.120 208.330 1703.180 ;
        RECT 206.710 1702.950 207.435 1703.120 ;
        RECT 207.605 1702.950 208.330 1703.120 ;
        RECT 206.710 1702.890 208.330 1702.950 ;
        RECT 208.990 1703.120 210.325 1703.180 ;
        RECT 208.990 1702.950 210.155 1703.120 ;
        RECT 208.990 1702.890 210.325 1702.950 ;
        RECT 207.435 1702.805 207.605 1702.890 ;
        RECT 210.155 1702.805 210.325 1702.890 ;
        RECT 206.615 1702.460 207.265 1702.630 ;
        RECT 206.615 1701.790 206.785 1702.460 ;
        RECT 206.955 1701.960 207.435 1702.290 ;
        RECT 206.615 1701.620 207.260 1701.790 ;
        RECT 203.915 1701.370 204.885 1701.490 ;
        RECT 205.905 1701.385 206.075 1701.540 ;
        RECT 206.615 1701.385 206.785 1701.620 ;
        RECT 203.915 1701.280 205.685 1701.370 ;
        RECT 203.915 1701.160 204.715 1701.280 ;
        RECT 204.885 1701.200 205.685 1701.280 ;
        RECT 205.905 1701.210 206.785 1701.385 ;
      LAYER li1 ;
        RECT 203.525 1700.820 204.545 1700.990 ;
      LAYER li1 ;
        RECT 204.715 1700.820 204.885 1701.110 ;
      LAYER li1 ;
        RECT 203.525 1700.150 203.695 1700.820 ;
        RECT 205.055 1700.780 206.075 1700.950 ;
      LAYER li1 ;
        RECT 203.915 1700.610 204.885 1700.650 ;
        RECT 203.915 1700.360 205.685 1700.610 ;
        RECT 203.915 1700.320 204.715 1700.360 ;
        RECT 204.885 1700.280 205.685 1700.360 ;
      LAYER li1 ;
        RECT 203.525 1699.980 204.545 1700.150 ;
        RECT 203.525 1699.310 203.695 1699.980 ;
      LAYER li1 ;
        RECT 204.715 1699.900 204.885 1700.190 ;
      LAYER li1 ;
        RECT 205.905 1700.110 206.075 1700.780 ;
        RECT 205.055 1699.940 206.075 1700.110 ;
      LAYER li1 ;
        RECT 203.915 1699.730 204.715 1699.810 ;
        RECT 204.885 1699.730 205.685 1699.770 ;
        RECT 203.915 1699.480 205.685 1699.730 ;
        RECT 204.715 1699.440 205.685 1699.480 ;
      LAYER li1 ;
        RECT 203.525 1699.140 204.545 1699.310 ;
        RECT 205.905 1699.270 206.075 1699.940 ;
      LAYER li1 ;
        RECT 204.715 1698.980 204.885 1699.270 ;
      LAYER li1 ;
        RECT 205.055 1699.100 206.075 1699.270 ;
      LAYER li1 ;
        RECT 201.995 1698.640 202.645 1698.810 ;
        RECT 202.815 1698.705 203.695 1698.880 ;
        RECT 203.915 1698.810 204.715 1698.890 ;
        RECT 204.885 1698.810 205.685 1698.930 ;
        RECT 203.915 1698.720 205.685 1698.810 ;
        RECT 201.995 1698.520 202.165 1698.640 ;
        RECT 202.815 1698.470 202.985 1698.705 ;
        RECT 203.525 1698.550 203.695 1698.705 ;
        RECT 204.715 1698.600 205.685 1698.720 ;
        RECT 201.995 1698.130 202.165 1698.350 ;
        RECT 202.340 1698.300 202.985 1698.470 ;
        RECT 201.995 1698.060 202.645 1698.130 ;
        RECT 202.165 1697.890 202.645 1698.060 ;
        RECT 201.995 1697.800 202.645 1697.890 ;
        RECT 201.995 1697.600 202.165 1697.800 ;
        RECT 202.815 1697.630 202.985 1698.300 ;
        RECT 202.335 1697.460 202.985 1697.630 ;
        RECT 201.995 1697.200 202.165 1697.430 ;
      LAYER li1 ;
        RECT 203.155 1697.425 203.355 1698.525 ;
      LAYER li1 ;
        RECT 203.525 1698.220 204.545 1698.550 ;
        RECT 204.715 1698.520 204.885 1698.600 ;
      LAYER li1 ;
        RECT 205.905 1698.515 206.075 1699.100 ;
      LAYER li1 ;
        RECT 206.275 1698.760 206.445 1701.210 ;
        RECT 206.955 1701.120 207.435 1701.450 ;
      LAYER li1 ;
        RECT 206.615 1700.780 207.265 1700.950 ;
        RECT 206.615 1700.110 206.785 1700.780 ;
      LAYER li1 ;
        RECT 206.955 1700.280 207.435 1700.610 ;
      LAYER li1 ;
        RECT 206.615 1699.940 207.265 1700.110 ;
        RECT 206.615 1699.270 206.785 1699.940 ;
      LAYER li1 ;
        RECT 206.955 1699.440 207.435 1699.770 ;
      LAYER li1 ;
        RECT 206.615 1699.100 207.265 1699.270 ;
        RECT 206.615 1698.515 206.785 1699.100 ;
      LAYER li1 ;
        RECT 206.955 1698.600 207.435 1698.930 ;
      LAYER li1 ;
        RECT 205.905 1698.430 206.785 1698.515 ;
      LAYER li1 ;
        RECT 203.525 1697.710 203.695 1698.220 ;
        RECT 204.715 1698.090 204.885 1698.350 ;
      LAYER li1 ;
        RECT 205.055 1698.260 207.265 1698.430 ;
      LAYER li1 ;
        RECT 204.715 1698.060 206.035 1698.090 ;
        RECT 203.915 1697.890 204.715 1698.050 ;
        RECT 204.885 1697.890 206.035 1698.060 ;
        RECT 203.915 1697.880 206.035 1697.890 ;
        RECT 204.715 1697.760 206.035 1697.880 ;
        RECT 206.635 1697.760 207.435 1698.090 ;
        RECT 203.525 1697.380 204.545 1697.710 ;
        RECT 204.715 1697.600 204.885 1697.760 ;
        RECT 204.715 1697.200 204.885 1697.430 ;
        RECT 207.435 1697.200 207.605 1697.285 ;
        RECT 210.155 1697.200 210.325 1697.285 ;
        RECT 201.995 1697.140 202.890 1697.200 ;
        RECT 202.165 1696.970 202.890 1697.140 ;
        RECT 201.995 1696.910 202.890 1696.970 ;
        RECT 203.550 1697.140 206.050 1697.200 ;
        RECT 203.550 1696.970 204.715 1697.140 ;
        RECT 204.885 1696.970 206.050 1697.140 ;
        RECT 203.550 1696.910 206.050 1696.970 ;
        RECT 206.710 1697.140 208.330 1697.200 ;
        RECT 206.710 1696.970 207.435 1697.140 ;
        RECT 207.605 1696.970 208.330 1697.140 ;
        RECT 206.710 1696.910 208.330 1696.970 ;
        RECT 208.990 1697.140 210.325 1697.200 ;
        RECT 208.990 1696.970 210.155 1697.140 ;
        RECT 208.990 1696.910 210.325 1696.970 ;
        RECT 201.995 1696.680 202.165 1696.910 ;
        RECT 204.715 1696.680 204.885 1696.910 ;
        RECT 207.435 1696.825 207.605 1696.910 ;
        RECT 210.155 1696.825 210.325 1696.910 ;
        RECT 201.995 1696.350 202.165 1696.510 ;
        RECT 204.715 1696.350 204.885 1696.510 ;
        RECT 205.055 1696.400 206.075 1696.730 ;
        RECT 201.995 1696.220 202.965 1696.350 ;
        RECT 202.165 1696.050 202.965 1696.220 ;
        RECT 201.995 1696.020 202.965 1696.050 ;
        RECT 203.565 1696.230 204.885 1696.350 ;
        RECT 203.565 1696.220 205.685 1696.230 ;
        RECT 203.565 1696.050 204.715 1696.220 ;
        RECT 204.885 1696.060 205.685 1696.220 ;
        RECT 203.565 1696.020 204.885 1696.050 ;
        RECT 201.995 1695.760 202.165 1696.020 ;
        RECT 204.715 1695.760 204.885 1696.020 ;
        RECT 205.905 1695.890 206.075 1696.400 ;
        RECT 201.995 1695.510 202.165 1695.590 ;
        RECT 204.715 1695.510 204.885 1695.590 ;
        RECT 205.055 1695.560 206.075 1695.890 ;
        RECT 201.995 1695.300 202.645 1695.510 ;
        RECT 203.915 1695.390 204.885 1695.510 ;
        RECT 205.905 1695.405 206.075 1695.560 ;
        RECT 206.615 1696.480 207.265 1696.650 ;
        RECT 206.615 1695.810 206.785 1696.480 ;
        RECT 206.955 1695.980 207.435 1696.310 ;
        RECT 206.615 1695.640 207.260 1695.810 ;
        RECT 206.615 1695.405 206.785 1695.640 ;
        RECT 202.165 1695.180 202.645 1695.300 ;
        RECT 201.995 1694.840 202.165 1695.130 ;
        RECT 201.995 1694.380 202.645 1694.670 ;
        RECT 202.165 1694.340 202.645 1694.380 ;
        RECT 201.995 1693.920 202.165 1694.210 ;
        RECT 202.165 1693.750 202.645 1693.830 ;
        RECT 201.995 1693.500 202.645 1693.750 ;
        RECT 201.995 1693.460 202.165 1693.500 ;
        RECT 201.995 1693.000 202.165 1693.290 ;
        RECT 202.165 1692.830 202.645 1692.990 ;
        RECT 203.155 1692.900 203.325 1695.350 ;
        RECT 203.915 1695.300 205.685 1695.390 ;
        RECT 203.915 1695.180 204.715 1695.300 ;
        RECT 204.885 1695.220 205.685 1695.300 ;
        RECT 205.905 1695.230 206.785 1695.405 ;
        RECT 204.715 1694.840 204.885 1695.130 ;
      LAYER li1 ;
        RECT 205.055 1694.800 206.075 1694.970 ;
      LAYER li1 ;
        RECT 203.915 1694.630 204.885 1694.670 ;
        RECT 203.915 1694.380 205.685 1694.630 ;
        RECT 203.915 1694.340 204.715 1694.380 ;
        RECT 204.885 1694.300 205.685 1694.380 ;
        RECT 204.715 1693.920 204.885 1694.210 ;
      LAYER li1 ;
        RECT 205.905 1694.130 206.075 1694.800 ;
        RECT 205.055 1693.960 206.075 1694.130 ;
      LAYER li1 ;
        RECT 203.915 1693.750 204.715 1693.830 ;
        RECT 204.885 1693.750 205.685 1693.790 ;
        RECT 203.915 1693.500 205.685 1693.750 ;
        RECT 204.715 1693.460 205.685 1693.500 ;
      LAYER li1 ;
        RECT 205.905 1693.290 206.075 1693.960 ;
      LAYER li1 ;
        RECT 204.715 1693.000 204.885 1693.290 ;
      LAYER li1 ;
        RECT 205.055 1693.120 206.075 1693.290 ;
      LAYER li1 ;
        RECT 201.995 1692.660 202.645 1692.830 ;
        RECT 202.815 1692.725 203.695 1692.900 ;
        RECT 203.915 1692.830 204.715 1692.910 ;
        RECT 204.885 1692.830 205.685 1692.950 ;
        RECT 203.915 1692.740 205.685 1692.830 ;
        RECT 201.995 1692.540 202.165 1692.660 ;
        RECT 202.815 1692.490 202.985 1692.725 ;
        RECT 203.525 1692.570 203.695 1692.725 ;
        RECT 204.715 1692.620 205.685 1692.740 ;
        RECT 201.995 1692.150 202.165 1692.370 ;
        RECT 202.340 1692.320 202.985 1692.490 ;
        RECT 201.995 1692.080 202.645 1692.150 ;
        RECT 202.165 1691.910 202.645 1692.080 ;
        RECT 201.995 1691.820 202.645 1691.910 ;
        RECT 201.995 1691.620 202.165 1691.820 ;
        RECT 202.815 1691.650 202.985 1692.320 ;
        RECT 202.335 1691.480 202.985 1691.650 ;
        RECT 201.995 1691.220 202.165 1691.450 ;
      LAYER li1 ;
        RECT 203.155 1691.445 203.355 1692.545 ;
      LAYER li1 ;
        RECT 203.525 1692.240 204.545 1692.570 ;
        RECT 204.715 1692.540 204.885 1692.620 ;
      LAYER li1 ;
        RECT 205.905 1692.535 206.075 1693.120 ;
      LAYER li1 ;
        RECT 206.275 1692.780 206.445 1695.230 ;
        RECT 206.955 1695.140 207.435 1695.470 ;
      LAYER li1 ;
        RECT 206.615 1694.800 207.265 1694.970 ;
        RECT 206.615 1694.130 206.785 1694.800 ;
      LAYER li1 ;
        RECT 206.955 1694.300 207.435 1694.630 ;
      LAYER li1 ;
        RECT 206.615 1693.960 207.265 1694.130 ;
        RECT 206.615 1693.290 206.785 1693.960 ;
      LAYER li1 ;
        RECT 206.955 1693.460 207.435 1693.790 ;
      LAYER li1 ;
        RECT 206.615 1693.120 207.265 1693.290 ;
        RECT 206.615 1692.535 206.785 1693.120 ;
      LAYER li1 ;
        RECT 206.955 1692.620 207.435 1692.950 ;
      LAYER li1 ;
        RECT 205.905 1692.450 206.785 1692.535 ;
      LAYER li1 ;
        RECT 203.525 1691.730 203.695 1692.240 ;
        RECT 204.715 1692.110 204.885 1692.370 ;
      LAYER li1 ;
        RECT 205.055 1692.280 207.265 1692.450 ;
      LAYER li1 ;
        RECT 204.715 1692.080 206.035 1692.110 ;
        RECT 203.915 1691.910 204.715 1692.070 ;
        RECT 204.885 1691.910 206.035 1692.080 ;
        RECT 203.915 1691.900 206.035 1691.910 ;
        RECT 204.715 1691.780 206.035 1691.900 ;
        RECT 206.635 1691.780 207.435 1692.110 ;
        RECT 203.525 1691.400 204.545 1691.730 ;
        RECT 204.715 1691.620 204.885 1691.780 ;
        RECT 204.715 1691.220 204.885 1691.450 ;
        RECT 207.435 1691.220 207.605 1691.305 ;
        RECT 210.155 1691.220 210.325 1691.305 ;
        RECT 201.995 1691.160 202.890 1691.220 ;
        RECT 202.165 1690.990 202.890 1691.160 ;
        RECT 201.995 1690.930 202.890 1690.990 ;
        RECT 203.550 1691.160 206.050 1691.220 ;
        RECT 203.550 1690.990 204.715 1691.160 ;
        RECT 204.885 1690.990 206.050 1691.160 ;
        RECT 203.550 1690.930 206.050 1690.990 ;
        RECT 206.710 1691.160 208.330 1691.220 ;
        RECT 206.710 1690.990 207.435 1691.160 ;
        RECT 207.605 1690.990 208.330 1691.160 ;
        RECT 206.710 1690.930 208.330 1690.990 ;
        RECT 208.990 1691.160 210.325 1691.220 ;
        RECT 208.990 1690.990 210.155 1691.160 ;
        RECT 208.990 1690.930 210.325 1690.990 ;
        RECT 201.995 1690.700 202.165 1690.930 ;
        RECT 204.715 1690.700 204.885 1690.930 ;
        RECT 207.435 1690.845 207.605 1690.930 ;
        RECT 210.155 1690.845 210.325 1690.930 ;
        RECT 201.995 1690.370 202.165 1690.530 ;
        RECT 204.715 1690.370 204.885 1690.530 ;
        RECT 205.055 1690.420 206.075 1690.750 ;
        RECT 201.995 1690.240 202.965 1690.370 ;
        RECT 202.165 1690.070 202.965 1690.240 ;
        RECT 201.995 1690.040 202.965 1690.070 ;
        RECT 203.565 1690.250 204.885 1690.370 ;
        RECT 203.565 1690.240 205.685 1690.250 ;
        RECT 203.565 1690.070 204.715 1690.240 ;
        RECT 204.885 1690.080 205.685 1690.240 ;
        RECT 203.565 1690.040 204.885 1690.070 ;
        RECT 201.995 1689.780 202.165 1690.040 ;
        RECT 204.715 1689.780 204.885 1690.040 ;
        RECT 205.905 1689.910 206.075 1690.420 ;
        RECT 201.995 1689.530 202.165 1689.610 ;
        RECT 204.715 1689.530 204.885 1689.610 ;
        RECT 205.055 1689.580 206.075 1689.910 ;
        RECT 201.995 1689.320 202.645 1689.530 ;
        RECT 203.915 1689.410 204.885 1689.530 ;
        RECT 205.905 1689.425 206.075 1689.580 ;
        RECT 206.615 1690.500 207.265 1690.670 ;
        RECT 206.615 1689.830 206.785 1690.500 ;
        RECT 206.955 1690.000 207.435 1690.330 ;
        RECT 206.615 1689.660 207.260 1689.830 ;
        RECT 206.615 1689.425 206.785 1689.660 ;
        RECT 202.165 1689.200 202.645 1689.320 ;
        RECT 201.995 1688.860 202.165 1689.150 ;
        RECT 201.995 1688.400 202.645 1688.690 ;
        RECT 202.165 1688.360 202.645 1688.400 ;
        RECT 201.995 1687.940 202.165 1688.230 ;
        RECT 202.165 1687.770 202.645 1687.850 ;
        RECT 201.995 1687.520 202.645 1687.770 ;
        RECT 201.995 1687.480 202.165 1687.520 ;
        RECT 201.995 1687.020 202.165 1687.310 ;
        RECT 202.165 1686.850 202.645 1687.010 ;
        RECT 203.155 1686.920 203.325 1689.370 ;
        RECT 203.915 1689.320 205.685 1689.410 ;
        RECT 203.915 1689.200 204.715 1689.320 ;
        RECT 204.885 1689.240 205.685 1689.320 ;
        RECT 205.905 1689.250 206.785 1689.425 ;
        RECT 204.715 1688.860 204.885 1689.150 ;
      LAYER li1 ;
        RECT 205.055 1688.820 206.075 1688.990 ;
      LAYER li1 ;
        RECT 203.915 1688.650 204.885 1688.690 ;
        RECT 203.915 1688.400 205.685 1688.650 ;
        RECT 203.915 1688.360 204.715 1688.400 ;
        RECT 204.885 1688.320 205.685 1688.400 ;
        RECT 204.715 1687.940 204.885 1688.230 ;
      LAYER li1 ;
        RECT 205.905 1688.150 206.075 1688.820 ;
        RECT 205.055 1687.980 206.075 1688.150 ;
      LAYER li1 ;
        RECT 203.915 1687.770 204.715 1687.850 ;
        RECT 204.885 1687.770 205.685 1687.810 ;
        RECT 203.915 1687.520 205.685 1687.770 ;
        RECT 204.715 1687.480 205.685 1687.520 ;
      LAYER li1 ;
        RECT 205.905 1687.310 206.075 1687.980 ;
      LAYER li1 ;
        RECT 204.715 1687.020 204.885 1687.310 ;
      LAYER li1 ;
        RECT 205.055 1687.140 206.075 1687.310 ;
      LAYER li1 ;
        RECT 201.995 1686.680 202.645 1686.850 ;
        RECT 202.815 1686.745 203.695 1686.920 ;
        RECT 203.915 1686.850 204.715 1686.930 ;
        RECT 204.885 1686.850 205.685 1686.970 ;
        RECT 203.915 1686.760 205.685 1686.850 ;
        RECT 201.995 1686.560 202.165 1686.680 ;
        RECT 202.815 1686.510 202.985 1686.745 ;
        RECT 203.525 1686.590 203.695 1686.745 ;
        RECT 204.715 1686.640 205.685 1686.760 ;
        RECT 201.995 1686.170 202.165 1686.390 ;
        RECT 202.340 1686.340 202.985 1686.510 ;
        RECT 201.995 1686.100 202.645 1686.170 ;
        RECT 202.165 1685.930 202.645 1686.100 ;
        RECT 201.995 1685.840 202.645 1685.930 ;
        RECT 201.995 1685.640 202.165 1685.840 ;
        RECT 202.815 1685.670 202.985 1686.340 ;
        RECT 202.335 1685.500 202.985 1685.670 ;
        RECT 201.995 1685.240 202.165 1685.470 ;
      LAYER li1 ;
        RECT 203.155 1685.465 203.355 1686.565 ;
      LAYER li1 ;
        RECT 203.525 1686.260 204.545 1686.590 ;
        RECT 204.715 1686.560 204.885 1686.640 ;
      LAYER li1 ;
        RECT 205.905 1686.555 206.075 1687.140 ;
      LAYER li1 ;
        RECT 206.275 1686.800 206.445 1689.250 ;
        RECT 206.955 1689.160 207.435 1689.490 ;
      LAYER li1 ;
        RECT 206.615 1688.820 207.265 1688.990 ;
        RECT 206.615 1688.150 206.785 1688.820 ;
      LAYER li1 ;
        RECT 206.955 1688.320 207.435 1688.650 ;
      LAYER li1 ;
        RECT 206.615 1687.980 207.265 1688.150 ;
        RECT 206.615 1687.310 206.785 1687.980 ;
      LAYER li1 ;
        RECT 206.955 1687.480 207.435 1687.810 ;
      LAYER li1 ;
        RECT 206.615 1687.140 207.265 1687.310 ;
        RECT 206.615 1686.555 206.785 1687.140 ;
      LAYER li1 ;
        RECT 206.955 1686.640 207.435 1686.970 ;
      LAYER li1 ;
        RECT 205.905 1686.470 206.785 1686.555 ;
      LAYER li1 ;
        RECT 203.525 1685.750 203.695 1686.260 ;
        RECT 204.715 1686.130 204.885 1686.390 ;
      LAYER li1 ;
        RECT 205.055 1686.300 207.265 1686.470 ;
      LAYER li1 ;
        RECT 204.715 1686.100 206.035 1686.130 ;
        RECT 203.915 1685.930 204.715 1686.090 ;
        RECT 204.885 1685.930 206.035 1686.100 ;
        RECT 203.915 1685.920 206.035 1685.930 ;
        RECT 204.715 1685.800 206.035 1685.920 ;
        RECT 206.635 1685.800 207.435 1686.130 ;
        RECT 203.525 1685.420 204.545 1685.750 ;
        RECT 204.715 1685.640 204.885 1685.800 ;
        RECT 204.715 1685.240 204.885 1685.470 ;
        RECT 207.435 1685.240 207.605 1685.325 ;
        RECT 210.155 1685.240 210.325 1685.325 ;
        RECT 201.995 1685.180 202.890 1685.240 ;
        RECT 202.165 1685.010 202.890 1685.180 ;
        RECT 201.995 1684.950 202.890 1685.010 ;
        RECT 203.550 1685.180 206.050 1685.240 ;
        RECT 203.550 1685.010 204.715 1685.180 ;
        RECT 204.885 1685.010 206.050 1685.180 ;
        RECT 203.550 1684.950 206.050 1685.010 ;
        RECT 206.710 1685.180 208.330 1685.240 ;
        RECT 206.710 1685.010 207.435 1685.180 ;
        RECT 207.605 1685.010 208.330 1685.180 ;
        RECT 206.710 1684.950 208.330 1685.010 ;
        RECT 208.990 1685.180 210.325 1685.240 ;
        RECT 208.990 1685.010 210.155 1685.180 ;
        RECT 208.990 1684.950 210.325 1685.010 ;
        RECT 201.995 1684.720 202.165 1684.950 ;
        RECT 204.715 1684.720 204.885 1684.950 ;
        RECT 207.435 1684.865 207.605 1684.950 ;
        RECT 210.155 1684.865 210.325 1684.950 ;
        RECT 201.995 1684.390 202.165 1684.550 ;
        RECT 204.715 1684.390 204.885 1684.550 ;
        RECT 205.055 1684.440 206.075 1684.770 ;
        RECT 201.995 1684.260 202.965 1684.390 ;
        RECT 202.165 1684.090 202.965 1684.260 ;
        RECT 201.995 1684.060 202.965 1684.090 ;
        RECT 203.565 1684.270 204.885 1684.390 ;
        RECT 203.565 1684.260 205.685 1684.270 ;
        RECT 203.565 1684.090 204.715 1684.260 ;
        RECT 204.885 1684.100 205.685 1684.260 ;
        RECT 203.565 1684.060 204.885 1684.090 ;
        RECT 201.995 1683.800 202.165 1684.060 ;
        RECT 204.715 1683.800 204.885 1684.060 ;
        RECT 205.905 1683.930 206.075 1684.440 ;
        RECT 201.995 1683.550 202.165 1683.630 ;
        RECT 204.715 1683.550 204.885 1683.630 ;
        RECT 205.055 1683.600 206.075 1683.930 ;
        RECT 201.995 1683.340 202.645 1683.550 ;
        RECT 203.915 1683.430 204.885 1683.550 ;
        RECT 205.905 1683.445 206.075 1683.600 ;
        RECT 206.615 1684.520 207.265 1684.690 ;
        RECT 206.615 1683.850 206.785 1684.520 ;
        RECT 206.955 1684.020 207.435 1684.350 ;
        RECT 206.615 1683.680 207.260 1683.850 ;
        RECT 206.615 1683.445 206.785 1683.680 ;
        RECT 202.165 1683.220 202.645 1683.340 ;
        RECT 201.995 1682.880 202.165 1683.170 ;
        RECT 201.995 1682.420 202.645 1682.710 ;
        RECT 202.165 1682.380 202.645 1682.420 ;
        RECT 201.995 1681.960 202.165 1682.250 ;
        RECT 202.165 1681.790 202.645 1681.870 ;
        RECT 201.995 1681.540 202.645 1681.790 ;
        RECT 201.995 1681.500 202.165 1681.540 ;
        RECT 201.995 1681.040 202.165 1681.330 ;
        RECT 202.165 1680.870 202.645 1681.030 ;
        RECT 203.155 1680.940 203.325 1683.390 ;
        RECT 203.915 1683.340 205.685 1683.430 ;
        RECT 203.915 1683.220 204.715 1683.340 ;
        RECT 204.885 1683.260 205.685 1683.340 ;
        RECT 205.905 1683.270 206.785 1683.445 ;
        RECT 204.715 1682.880 204.885 1683.170 ;
      LAYER li1 ;
        RECT 205.055 1682.840 206.075 1683.010 ;
      LAYER li1 ;
        RECT 203.915 1682.670 204.885 1682.710 ;
        RECT 203.915 1682.420 205.685 1682.670 ;
        RECT 203.915 1682.380 204.715 1682.420 ;
        RECT 204.885 1682.340 205.685 1682.420 ;
        RECT 204.715 1681.960 204.885 1682.250 ;
      LAYER li1 ;
        RECT 205.905 1682.170 206.075 1682.840 ;
        RECT 205.055 1682.000 206.075 1682.170 ;
      LAYER li1 ;
        RECT 203.915 1681.790 204.715 1681.870 ;
        RECT 204.885 1681.790 205.685 1681.830 ;
        RECT 203.915 1681.540 205.685 1681.790 ;
        RECT 204.715 1681.500 205.685 1681.540 ;
      LAYER li1 ;
        RECT 205.905 1681.330 206.075 1682.000 ;
      LAYER li1 ;
        RECT 204.715 1681.040 204.885 1681.330 ;
      LAYER li1 ;
        RECT 205.055 1681.160 206.075 1681.330 ;
      LAYER li1 ;
        RECT 201.995 1680.700 202.645 1680.870 ;
        RECT 202.815 1680.765 203.695 1680.940 ;
        RECT 203.915 1680.870 204.715 1680.950 ;
        RECT 204.885 1680.870 205.685 1680.990 ;
        RECT 203.915 1680.780 205.685 1680.870 ;
        RECT 201.995 1680.580 202.165 1680.700 ;
        RECT 202.815 1680.530 202.985 1680.765 ;
        RECT 203.525 1680.610 203.695 1680.765 ;
        RECT 204.715 1680.660 205.685 1680.780 ;
        RECT 201.995 1680.190 202.165 1680.410 ;
        RECT 202.340 1680.360 202.985 1680.530 ;
        RECT 201.995 1680.120 202.645 1680.190 ;
        RECT 202.165 1679.950 202.645 1680.120 ;
        RECT 201.995 1679.860 202.645 1679.950 ;
        RECT 201.995 1679.660 202.165 1679.860 ;
        RECT 202.815 1679.690 202.985 1680.360 ;
        RECT 202.335 1679.520 202.985 1679.690 ;
        RECT 201.995 1679.260 202.165 1679.490 ;
      LAYER li1 ;
        RECT 203.155 1679.485 203.355 1680.585 ;
      LAYER li1 ;
        RECT 203.525 1680.280 204.545 1680.610 ;
        RECT 204.715 1680.580 204.885 1680.660 ;
      LAYER li1 ;
        RECT 205.905 1680.575 206.075 1681.160 ;
      LAYER li1 ;
        RECT 206.275 1680.820 206.445 1683.270 ;
        RECT 206.955 1683.180 207.435 1683.510 ;
      LAYER li1 ;
        RECT 206.615 1682.840 207.265 1683.010 ;
        RECT 206.615 1682.170 206.785 1682.840 ;
      LAYER li1 ;
        RECT 206.955 1682.340 207.435 1682.670 ;
      LAYER li1 ;
        RECT 206.615 1682.000 207.265 1682.170 ;
        RECT 206.615 1681.330 206.785 1682.000 ;
      LAYER li1 ;
        RECT 206.955 1681.500 207.435 1681.830 ;
      LAYER li1 ;
        RECT 206.615 1681.160 207.265 1681.330 ;
        RECT 206.615 1680.575 206.785 1681.160 ;
      LAYER li1 ;
        RECT 206.955 1680.660 207.435 1680.990 ;
      LAYER li1 ;
        RECT 205.905 1680.490 206.785 1680.575 ;
      LAYER li1 ;
        RECT 203.525 1679.770 203.695 1680.280 ;
        RECT 204.715 1680.150 204.885 1680.410 ;
      LAYER li1 ;
        RECT 205.055 1680.320 207.265 1680.490 ;
      LAYER li1 ;
        RECT 204.715 1680.120 206.035 1680.150 ;
        RECT 203.915 1679.950 204.715 1680.110 ;
        RECT 204.885 1679.950 206.035 1680.120 ;
        RECT 203.915 1679.940 206.035 1679.950 ;
        RECT 204.715 1679.820 206.035 1679.940 ;
        RECT 206.635 1679.820 207.435 1680.150 ;
        RECT 203.525 1679.440 204.545 1679.770 ;
        RECT 204.715 1679.660 204.885 1679.820 ;
        RECT 204.715 1679.260 204.885 1679.490 ;
        RECT 207.435 1679.260 207.605 1679.345 ;
        RECT 210.155 1679.260 210.325 1679.345 ;
        RECT 201.995 1679.200 202.890 1679.260 ;
        RECT 202.165 1679.030 202.890 1679.200 ;
        RECT 201.995 1678.970 202.890 1679.030 ;
        RECT 203.550 1679.200 206.050 1679.260 ;
        RECT 203.550 1679.030 204.715 1679.200 ;
        RECT 204.885 1679.030 206.050 1679.200 ;
        RECT 203.550 1678.970 206.050 1679.030 ;
        RECT 206.710 1679.200 208.330 1679.260 ;
        RECT 206.710 1679.030 207.435 1679.200 ;
        RECT 207.605 1679.030 208.330 1679.200 ;
        RECT 206.710 1678.970 208.330 1679.030 ;
        RECT 208.990 1679.200 210.325 1679.260 ;
        RECT 208.990 1679.030 210.155 1679.200 ;
        RECT 208.990 1678.970 210.325 1679.030 ;
        RECT 201.995 1678.740 202.165 1678.970 ;
        RECT 204.715 1678.740 204.885 1678.970 ;
        RECT 207.435 1678.885 207.605 1678.970 ;
        RECT 210.155 1678.885 210.325 1678.970 ;
        RECT 201.995 1678.410 202.165 1678.570 ;
        RECT 204.715 1678.410 204.885 1678.570 ;
        RECT 205.055 1678.460 206.075 1678.790 ;
        RECT 201.995 1678.280 202.965 1678.410 ;
        RECT 202.165 1678.110 202.965 1678.280 ;
        RECT 201.995 1678.080 202.965 1678.110 ;
        RECT 203.565 1678.290 204.885 1678.410 ;
        RECT 203.565 1678.280 205.685 1678.290 ;
        RECT 203.565 1678.110 204.715 1678.280 ;
        RECT 204.885 1678.120 205.685 1678.280 ;
        RECT 203.565 1678.080 204.885 1678.110 ;
        RECT 201.995 1677.820 202.165 1678.080 ;
        RECT 204.715 1677.820 204.885 1678.080 ;
        RECT 205.905 1677.950 206.075 1678.460 ;
        RECT 201.995 1677.570 202.165 1677.650 ;
        RECT 204.715 1677.570 204.885 1677.650 ;
        RECT 205.055 1677.620 206.075 1677.950 ;
        RECT 201.995 1677.360 202.645 1677.570 ;
        RECT 203.915 1677.450 204.885 1677.570 ;
        RECT 205.905 1677.465 206.075 1677.620 ;
        RECT 206.615 1678.540 207.265 1678.710 ;
        RECT 206.615 1677.870 206.785 1678.540 ;
        RECT 206.955 1678.040 207.435 1678.370 ;
        RECT 206.615 1677.700 207.260 1677.870 ;
        RECT 206.615 1677.465 206.785 1677.700 ;
        RECT 202.165 1677.240 202.645 1677.360 ;
        RECT 201.995 1676.900 202.165 1677.190 ;
        RECT 201.995 1676.440 202.645 1676.730 ;
        RECT 202.165 1676.400 202.645 1676.440 ;
        RECT 201.995 1675.980 202.165 1676.270 ;
        RECT 202.165 1675.810 202.645 1675.890 ;
        RECT 201.995 1675.560 202.645 1675.810 ;
        RECT 201.995 1675.520 202.165 1675.560 ;
        RECT 201.995 1675.060 202.165 1675.350 ;
        RECT 202.165 1674.890 202.645 1675.050 ;
        RECT 203.155 1674.960 203.325 1677.410 ;
        RECT 203.915 1677.360 205.685 1677.450 ;
        RECT 203.915 1677.240 204.715 1677.360 ;
        RECT 204.885 1677.280 205.685 1677.360 ;
        RECT 205.905 1677.290 206.785 1677.465 ;
        RECT 204.715 1676.900 204.885 1677.190 ;
      LAYER li1 ;
        RECT 205.055 1676.860 206.075 1677.030 ;
      LAYER li1 ;
        RECT 203.915 1676.690 204.885 1676.730 ;
        RECT 203.915 1676.440 205.685 1676.690 ;
        RECT 203.915 1676.400 204.715 1676.440 ;
        RECT 204.885 1676.360 205.685 1676.440 ;
        RECT 204.715 1675.980 204.885 1676.270 ;
      LAYER li1 ;
        RECT 205.905 1676.190 206.075 1676.860 ;
        RECT 205.055 1676.020 206.075 1676.190 ;
      LAYER li1 ;
        RECT 203.915 1675.810 204.715 1675.890 ;
        RECT 204.885 1675.810 205.685 1675.850 ;
        RECT 203.915 1675.560 205.685 1675.810 ;
        RECT 204.715 1675.520 205.685 1675.560 ;
      LAYER li1 ;
        RECT 205.905 1675.350 206.075 1676.020 ;
      LAYER li1 ;
        RECT 204.715 1675.060 204.885 1675.350 ;
      LAYER li1 ;
        RECT 205.055 1675.180 206.075 1675.350 ;
      LAYER li1 ;
        RECT 201.995 1674.720 202.645 1674.890 ;
        RECT 202.815 1674.785 203.695 1674.960 ;
        RECT 203.915 1674.890 204.715 1674.970 ;
        RECT 204.885 1674.890 205.685 1675.010 ;
        RECT 203.915 1674.800 205.685 1674.890 ;
        RECT 201.995 1674.600 202.165 1674.720 ;
        RECT 202.815 1674.550 202.985 1674.785 ;
        RECT 203.525 1674.630 203.695 1674.785 ;
        RECT 204.715 1674.680 205.685 1674.800 ;
        RECT 201.995 1674.210 202.165 1674.430 ;
        RECT 202.340 1674.380 202.985 1674.550 ;
        RECT 201.995 1674.140 202.645 1674.210 ;
        RECT 202.165 1673.970 202.645 1674.140 ;
        RECT 201.995 1673.880 202.645 1673.970 ;
        RECT 201.995 1673.680 202.165 1673.880 ;
        RECT 202.815 1673.710 202.985 1674.380 ;
        RECT 202.335 1673.540 202.985 1673.710 ;
        RECT 201.995 1673.280 202.165 1673.510 ;
      LAYER li1 ;
        RECT 203.155 1673.505 203.355 1674.605 ;
      LAYER li1 ;
        RECT 203.525 1674.300 204.545 1674.630 ;
        RECT 204.715 1674.600 204.885 1674.680 ;
      LAYER li1 ;
        RECT 205.905 1674.595 206.075 1675.180 ;
      LAYER li1 ;
        RECT 206.275 1674.840 206.445 1677.290 ;
        RECT 206.955 1677.200 207.435 1677.530 ;
      LAYER li1 ;
        RECT 206.615 1676.860 207.265 1677.030 ;
        RECT 206.615 1676.190 206.785 1676.860 ;
      LAYER li1 ;
        RECT 206.955 1676.360 207.435 1676.690 ;
      LAYER li1 ;
        RECT 206.615 1676.020 207.265 1676.190 ;
        RECT 206.615 1675.350 206.785 1676.020 ;
      LAYER li1 ;
        RECT 206.955 1675.520 207.435 1675.850 ;
      LAYER li1 ;
        RECT 206.615 1675.180 207.265 1675.350 ;
        RECT 206.615 1674.595 206.785 1675.180 ;
      LAYER li1 ;
        RECT 206.955 1674.680 207.435 1675.010 ;
      LAYER li1 ;
        RECT 205.905 1674.510 206.785 1674.595 ;
      LAYER li1 ;
        RECT 203.525 1673.790 203.695 1674.300 ;
        RECT 204.715 1674.170 204.885 1674.430 ;
      LAYER li1 ;
        RECT 205.055 1674.340 207.265 1674.510 ;
      LAYER li1 ;
        RECT 204.715 1674.140 206.035 1674.170 ;
        RECT 203.915 1673.970 204.715 1674.130 ;
        RECT 204.885 1673.970 206.035 1674.140 ;
        RECT 203.915 1673.960 206.035 1673.970 ;
        RECT 204.715 1673.840 206.035 1673.960 ;
        RECT 206.635 1673.840 207.435 1674.170 ;
        RECT 203.525 1673.460 204.545 1673.790 ;
        RECT 204.715 1673.680 204.885 1673.840 ;
        RECT 204.715 1673.280 204.885 1673.510 ;
        RECT 207.435 1673.280 207.605 1673.365 ;
        RECT 210.155 1673.280 210.325 1673.365 ;
        RECT 201.995 1673.220 202.890 1673.280 ;
        RECT 202.165 1673.050 202.890 1673.220 ;
        RECT 201.995 1672.990 202.890 1673.050 ;
        RECT 203.550 1673.220 206.050 1673.280 ;
        RECT 203.550 1673.050 204.715 1673.220 ;
        RECT 204.885 1673.050 206.050 1673.220 ;
        RECT 203.550 1672.990 206.050 1673.050 ;
        RECT 206.710 1673.220 208.330 1673.280 ;
        RECT 206.710 1673.050 207.435 1673.220 ;
        RECT 207.605 1673.050 208.330 1673.220 ;
        RECT 206.710 1672.990 208.330 1673.050 ;
        RECT 208.990 1673.220 210.325 1673.280 ;
        RECT 208.990 1673.050 210.155 1673.220 ;
        RECT 208.990 1672.990 210.325 1673.050 ;
        RECT 201.995 1672.905 202.165 1672.990 ;
        RECT 204.715 1672.905 204.885 1672.990 ;
        RECT 207.435 1672.905 207.605 1672.990 ;
        RECT 210.155 1672.905 210.325 1672.990 ;
        RECT 669.000 219.760 669.145 219.930 ;
        RECT 669.315 219.760 669.460 219.930 ;
        RECT 674.980 219.760 675.125 219.930 ;
        RECT 675.295 219.760 675.440 219.930 ;
        RECT 680.960 219.760 681.105 219.930 ;
        RECT 681.275 219.760 681.420 219.930 ;
        RECT 686.940 219.760 687.085 219.930 ;
        RECT 687.255 219.760 687.400 219.930 ;
        RECT 692.920 219.760 693.065 219.930 ;
        RECT 693.235 219.760 693.380 219.930 ;
        RECT 698.900 219.760 699.045 219.930 ;
        RECT 699.215 219.760 699.360 219.930 ;
        RECT 704.880 219.760 705.025 219.930 ;
        RECT 705.195 219.760 705.340 219.930 ;
        RECT 710.860 219.760 711.005 219.930 ;
        RECT 711.175 219.760 711.320 219.930 ;
        RECT 716.840 219.760 716.985 219.930 ;
        RECT 717.155 219.760 717.300 219.930 ;
        RECT 722.820 219.760 722.965 219.930 ;
        RECT 723.135 219.760 723.280 219.930 ;
        RECT 728.800 219.760 728.945 219.930 ;
        RECT 729.115 219.760 729.260 219.930 ;
        RECT 758.700 219.760 758.845 219.930 ;
        RECT 759.015 219.760 759.160 219.930 ;
        RECT 764.680 219.760 764.825 219.930 ;
        RECT 764.995 219.760 765.140 219.930 ;
        RECT 770.660 219.760 770.805 219.930 ;
        RECT 770.975 219.760 771.120 219.930 ;
        RECT 776.640 219.760 776.785 219.930 ;
        RECT 776.955 219.760 777.100 219.930 ;
        RECT 782.620 219.760 782.765 219.930 ;
        RECT 782.935 219.760 783.080 219.930 ;
        RECT 788.600 219.760 788.745 219.930 ;
        RECT 788.915 219.760 789.060 219.930 ;
        RECT 794.580 219.760 794.725 219.930 ;
        RECT 794.895 219.760 795.040 219.930 ;
        RECT 2146.000 219.760 2146.145 219.930 ;
        RECT 2146.315 219.760 2146.460 219.930 ;
        RECT 2151.980 219.760 2152.125 219.930 ;
        RECT 2152.295 219.760 2152.440 219.930 ;
        RECT 2157.960 219.760 2158.105 219.930 ;
        RECT 2158.275 219.760 2158.420 219.930 ;
        RECT 2163.940 219.760 2164.085 219.930 ;
        RECT 2164.255 219.760 2164.400 219.930 ;
        RECT 2169.920 219.760 2170.065 219.930 ;
        RECT 2170.235 219.760 2170.380 219.930 ;
        RECT 2175.900 219.760 2176.045 219.930 ;
        RECT 2176.215 219.760 2176.360 219.930 ;
        RECT 2181.880 219.760 2182.025 219.930 ;
        RECT 2182.195 219.760 2182.340 219.930 ;
        RECT 2187.860 219.760 2188.005 219.930 ;
        RECT 2188.175 219.760 2188.320 219.930 ;
        RECT 2193.840 219.760 2193.985 219.930 ;
        RECT 2194.155 219.760 2194.300 219.930 ;
        RECT 2199.820 219.760 2199.965 219.930 ;
        RECT 2200.135 219.760 2200.280 219.930 ;
        RECT 2205.800 219.760 2205.945 219.930 ;
        RECT 2206.115 219.760 2206.260 219.930 ;
        RECT 2235.700 219.760 2235.845 219.930 ;
        RECT 2236.015 219.760 2236.160 219.930 ;
        RECT 2241.680 219.760 2241.825 219.930 ;
        RECT 2241.995 219.760 2242.140 219.930 ;
        RECT 2247.660 219.760 2247.805 219.930 ;
        RECT 2247.975 219.760 2248.120 219.930 ;
        RECT 2253.640 219.760 2253.785 219.930 ;
        RECT 2253.955 219.760 2254.100 219.930 ;
        RECT 2259.620 219.760 2259.765 219.930 ;
        RECT 2259.935 219.760 2260.080 219.930 ;
        RECT 2265.600 219.760 2265.745 219.930 ;
        RECT 2265.915 219.760 2266.060 219.930 ;
        RECT 2271.580 219.760 2271.725 219.930 ;
        RECT 2271.895 219.760 2272.040 219.930 ;
        RECT 669.085 218.595 669.375 219.760 ;
        RECT 675.065 218.595 675.355 219.760 ;
        RECT 681.045 218.595 681.335 219.760 ;
        RECT 687.025 218.595 687.315 219.760 ;
        RECT 693.005 218.595 693.295 219.760 ;
        RECT 698.985 218.595 699.275 219.760 ;
        RECT 704.965 218.595 705.255 219.760 ;
        RECT 710.945 218.595 711.235 219.760 ;
        RECT 716.925 218.595 717.215 219.760 ;
        RECT 722.905 218.595 723.195 219.760 ;
        RECT 728.885 218.595 729.175 219.760 ;
        RECT 758.785 218.595 759.075 219.760 ;
        RECT 764.765 218.595 765.055 219.760 ;
        RECT 770.745 218.595 771.035 219.760 ;
        RECT 776.725 218.595 777.015 219.760 ;
        RECT 782.705 218.595 782.995 219.760 ;
        RECT 788.685 218.595 788.975 219.760 ;
        RECT 794.665 218.595 794.955 219.760 ;
        RECT 2146.085 218.595 2146.375 219.760 ;
        RECT 2152.065 218.595 2152.355 219.760 ;
        RECT 2158.045 218.595 2158.335 219.760 ;
        RECT 2164.025 218.595 2164.315 219.760 ;
        RECT 2170.005 218.595 2170.295 219.760 ;
        RECT 2175.985 218.595 2176.275 219.760 ;
        RECT 2181.965 218.595 2182.255 219.760 ;
        RECT 2187.945 218.595 2188.235 219.760 ;
        RECT 2193.925 218.595 2194.215 219.760 ;
        RECT 2199.905 218.595 2200.195 219.760 ;
        RECT 2205.885 218.595 2206.175 219.760 ;
        RECT 2235.785 218.595 2236.075 219.760 ;
        RECT 2241.765 218.595 2242.055 219.760 ;
        RECT 2247.745 218.595 2248.035 219.760 ;
        RECT 2253.725 218.595 2254.015 219.760 ;
        RECT 2259.705 218.595 2259.995 219.760 ;
        RECT 2265.685 218.595 2265.975 219.760 ;
        RECT 2271.665 218.595 2271.955 219.760 ;
        RECT 669.085 217.210 669.375 217.935 ;
        RECT 675.065 217.210 675.355 217.935 ;
        RECT 681.045 217.210 681.335 217.935 ;
        RECT 687.025 217.210 687.315 217.935 ;
        RECT 693.005 217.210 693.295 217.935 ;
      LAYER li1 ;
        RECT 695.050 217.755 695.390 218.585 ;
        RECT 693.465 217.210 698.810 217.755 ;
      LAYER li1 ;
        RECT 698.985 217.210 699.275 217.935 ;
      LAYER li1 ;
        RECT 701.030 217.755 701.370 218.585 ;
        RECT 699.445 217.210 704.790 217.755 ;
      LAYER li1 ;
        RECT 704.965 217.210 705.255 217.935 ;
      LAYER li1 ;
        RECT 707.010 217.755 707.350 218.585 ;
        RECT 705.425 217.210 710.770 217.755 ;
      LAYER li1 ;
        RECT 710.945 217.210 711.235 217.935 ;
        RECT 716.925 217.210 717.215 217.935 ;
        RECT 722.905 217.210 723.195 217.935 ;
        RECT 728.885 217.210 729.175 217.935 ;
        RECT 758.785 217.210 759.075 217.935 ;
      LAYER li1 ;
        RECT 760.830 217.755 761.170 218.585 ;
        RECT 759.245 217.210 764.590 217.755 ;
      LAYER li1 ;
        RECT 764.765 217.210 765.055 217.935 ;
      LAYER li1 ;
        RECT 766.810 217.755 767.150 218.585 ;
        RECT 765.225 217.210 770.570 217.755 ;
      LAYER li1 ;
        RECT 770.745 217.210 771.035 217.935 ;
      LAYER li1 ;
        RECT 772.790 217.755 773.130 218.585 ;
        RECT 771.205 217.210 776.550 217.755 ;
      LAYER li1 ;
        RECT 776.725 217.210 777.015 217.935 ;
      LAYER li1 ;
        RECT 778.770 217.755 779.110 218.585 ;
        RECT 777.185 217.210 782.530 217.755 ;
      LAYER li1 ;
        RECT 782.705 217.210 782.995 217.935 ;
      LAYER li1 ;
        RECT 784.750 217.755 785.090 218.585 ;
        RECT 783.165 217.210 788.510 217.755 ;
      LAYER li1 ;
        RECT 788.685 217.210 788.975 217.935 ;
        RECT 794.665 217.210 794.955 217.935 ;
        RECT 2146.085 217.210 2146.375 217.935 ;
        RECT 2152.065 217.210 2152.355 217.935 ;
        RECT 2158.045 217.210 2158.335 217.935 ;
        RECT 2164.025 217.210 2164.315 217.935 ;
        RECT 2170.005 217.210 2170.295 217.935 ;
        RECT 2175.985 217.210 2176.275 217.935 ;
        RECT 2181.965 217.210 2182.255 217.935 ;
        RECT 2187.945 217.210 2188.235 217.935 ;
        RECT 2193.925 217.210 2194.215 217.935 ;
        RECT 2199.905 217.210 2200.195 217.935 ;
        RECT 2205.885 217.210 2206.175 217.935 ;
        RECT 2235.785 217.210 2236.075 217.935 ;
        RECT 2241.765 217.210 2242.055 217.935 ;
        RECT 2247.745 217.210 2248.035 217.935 ;
        RECT 2253.725 217.210 2254.015 217.935 ;
        RECT 2259.705 217.210 2259.995 217.935 ;
        RECT 2265.685 217.210 2265.975 217.935 ;
        RECT 2271.665 217.210 2271.955 217.935 ;
        RECT 669.000 217.040 669.145 217.210 ;
        RECT 669.315 217.040 669.460 217.210 ;
        RECT 674.980 217.040 675.125 217.210 ;
        RECT 675.295 217.040 675.440 217.210 ;
        RECT 680.960 217.040 681.105 217.210 ;
        RECT 681.275 217.040 681.420 217.210 ;
        RECT 686.940 217.040 687.085 217.210 ;
        RECT 687.255 217.040 687.400 217.210 ;
        RECT 692.920 217.040 693.065 217.210 ;
        RECT 693.235 217.040 693.525 217.210 ;
        RECT 693.695 217.040 693.985 217.210 ;
        RECT 694.155 217.040 694.445 217.210 ;
        RECT 694.615 217.040 694.905 217.210 ;
        RECT 695.075 217.040 695.365 217.210 ;
        RECT 695.535 217.040 695.825 217.210 ;
        RECT 695.995 217.040 696.285 217.210 ;
        RECT 696.455 217.040 696.745 217.210 ;
        RECT 696.915 217.040 697.205 217.210 ;
        RECT 697.375 217.040 697.665 217.210 ;
        RECT 697.835 217.040 698.125 217.210 ;
        RECT 698.295 217.040 698.585 217.210 ;
        RECT 698.755 217.040 699.045 217.210 ;
        RECT 699.215 217.040 699.505 217.210 ;
        RECT 699.675 217.040 699.965 217.210 ;
        RECT 700.135 217.040 700.425 217.210 ;
        RECT 700.595 217.040 700.885 217.210 ;
        RECT 701.055 217.040 701.345 217.210 ;
        RECT 701.515 217.040 701.805 217.210 ;
        RECT 701.975 217.040 702.265 217.210 ;
        RECT 702.435 217.040 702.725 217.210 ;
        RECT 702.895 217.040 703.185 217.210 ;
        RECT 703.355 217.040 703.645 217.210 ;
        RECT 703.815 217.040 704.105 217.210 ;
        RECT 704.275 217.040 704.565 217.210 ;
        RECT 704.735 217.040 705.025 217.210 ;
        RECT 705.195 217.040 705.485 217.210 ;
        RECT 705.655 217.040 705.945 217.210 ;
        RECT 706.115 217.040 706.405 217.210 ;
        RECT 706.575 217.040 706.865 217.210 ;
        RECT 707.035 217.040 707.325 217.210 ;
        RECT 707.495 217.040 707.785 217.210 ;
        RECT 707.955 217.040 708.245 217.210 ;
        RECT 708.415 217.040 708.705 217.210 ;
        RECT 708.875 217.040 709.165 217.210 ;
        RECT 709.335 217.040 709.625 217.210 ;
        RECT 709.795 217.040 710.085 217.210 ;
        RECT 710.255 217.040 710.545 217.210 ;
        RECT 710.715 217.040 711.005 217.210 ;
        RECT 711.175 217.040 711.320 217.210 ;
        RECT 716.840 217.040 716.985 217.210 ;
        RECT 717.155 217.040 717.300 217.210 ;
        RECT 722.820 217.040 722.965 217.210 ;
        RECT 723.135 217.040 723.280 217.210 ;
        RECT 728.800 217.040 728.945 217.210 ;
        RECT 729.115 217.040 729.260 217.210 ;
        RECT 758.700 217.040 758.845 217.210 ;
        RECT 759.015 217.040 759.305 217.210 ;
        RECT 759.475 217.040 759.765 217.210 ;
        RECT 759.935 217.040 760.225 217.210 ;
        RECT 760.395 217.040 760.685 217.210 ;
        RECT 760.855 217.040 761.145 217.210 ;
        RECT 761.315 217.040 761.605 217.210 ;
        RECT 761.775 217.040 762.065 217.210 ;
        RECT 762.235 217.040 762.525 217.210 ;
        RECT 762.695 217.040 762.985 217.210 ;
        RECT 763.155 217.040 763.445 217.210 ;
        RECT 763.615 217.040 763.905 217.210 ;
        RECT 764.075 217.040 764.365 217.210 ;
        RECT 764.535 217.040 764.825 217.210 ;
        RECT 764.995 217.040 765.285 217.210 ;
        RECT 765.455 217.040 765.745 217.210 ;
        RECT 765.915 217.040 766.205 217.210 ;
        RECT 766.375 217.040 766.665 217.210 ;
        RECT 766.835 217.040 767.125 217.210 ;
        RECT 767.295 217.040 767.585 217.210 ;
        RECT 767.755 217.040 768.045 217.210 ;
        RECT 768.215 217.040 768.505 217.210 ;
        RECT 768.675 217.040 768.965 217.210 ;
        RECT 769.135 217.040 769.425 217.210 ;
        RECT 769.595 217.040 769.885 217.210 ;
        RECT 770.055 217.040 770.345 217.210 ;
        RECT 770.515 217.040 770.805 217.210 ;
        RECT 770.975 217.040 771.265 217.210 ;
        RECT 771.435 217.040 771.725 217.210 ;
        RECT 771.895 217.040 772.185 217.210 ;
        RECT 772.355 217.040 772.645 217.210 ;
        RECT 772.815 217.040 773.105 217.210 ;
        RECT 773.275 217.040 773.565 217.210 ;
        RECT 773.735 217.040 774.025 217.210 ;
        RECT 774.195 217.040 774.485 217.210 ;
        RECT 774.655 217.040 774.945 217.210 ;
        RECT 775.115 217.040 775.405 217.210 ;
        RECT 775.575 217.040 775.865 217.210 ;
        RECT 776.035 217.040 776.325 217.210 ;
        RECT 776.495 217.040 776.785 217.210 ;
        RECT 776.955 217.040 777.245 217.210 ;
        RECT 777.415 217.040 777.705 217.210 ;
        RECT 777.875 217.040 778.165 217.210 ;
        RECT 778.335 217.040 778.625 217.210 ;
        RECT 778.795 217.040 779.085 217.210 ;
        RECT 779.255 217.040 779.545 217.210 ;
        RECT 779.715 217.040 780.005 217.210 ;
        RECT 780.175 217.040 780.465 217.210 ;
        RECT 780.635 217.040 780.925 217.210 ;
        RECT 781.095 217.040 781.385 217.210 ;
        RECT 781.555 217.040 781.845 217.210 ;
        RECT 782.015 217.040 782.305 217.210 ;
        RECT 782.475 217.040 782.765 217.210 ;
        RECT 782.935 217.040 783.225 217.210 ;
        RECT 783.395 217.040 783.685 217.210 ;
        RECT 783.855 217.040 784.145 217.210 ;
        RECT 784.315 217.040 784.605 217.210 ;
        RECT 784.775 217.040 785.065 217.210 ;
        RECT 785.235 217.040 785.525 217.210 ;
        RECT 785.695 217.040 785.985 217.210 ;
        RECT 786.155 217.040 786.445 217.210 ;
        RECT 786.615 217.040 786.905 217.210 ;
        RECT 787.075 217.040 787.365 217.210 ;
        RECT 787.535 217.040 787.825 217.210 ;
        RECT 787.995 217.040 788.285 217.210 ;
        RECT 788.455 217.040 788.745 217.210 ;
        RECT 788.915 217.040 789.060 217.210 ;
        RECT 794.580 217.040 794.725 217.210 ;
        RECT 794.895 217.040 795.040 217.210 ;
        RECT 2146.000 217.040 2146.145 217.210 ;
        RECT 2146.315 217.040 2146.460 217.210 ;
        RECT 2151.980 217.040 2152.125 217.210 ;
        RECT 2152.295 217.040 2152.440 217.210 ;
        RECT 2157.960 217.040 2158.105 217.210 ;
        RECT 2158.275 217.040 2158.420 217.210 ;
        RECT 2163.940 217.040 2164.085 217.210 ;
        RECT 2164.255 217.040 2164.400 217.210 ;
        RECT 2169.920 217.040 2170.065 217.210 ;
        RECT 2170.235 217.040 2170.380 217.210 ;
        RECT 2175.900 217.040 2176.045 217.210 ;
        RECT 2176.215 217.040 2176.360 217.210 ;
        RECT 2181.880 217.040 2182.025 217.210 ;
        RECT 2182.195 217.040 2182.340 217.210 ;
        RECT 2187.860 217.040 2188.005 217.210 ;
        RECT 2188.175 217.040 2188.320 217.210 ;
        RECT 2193.840 217.040 2193.985 217.210 ;
        RECT 2194.155 217.040 2194.300 217.210 ;
        RECT 2199.820 217.040 2199.965 217.210 ;
        RECT 2200.135 217.040 2200.280 217.210 ;
        RECT 2205.800 217.040 2205.945 217.210 ;
        RECT 2206.115 217.040 2206.260 217.210 ;
        RECT 2235.700 217.040 2235.845 217.210 ;
        RECT 2236.015 217.040 2236.160 217.210 ;
        RECT 2241.680 217.040 2241.825 217.210 ;
        RECT 2241.995 217.040 2242.140 217.210 ;
        RECT 2247.660 217.040 2247.805 217.210 ;
        RECT 2247.975 217.040 2248.120 217.210 ;
        RECT 2253.640 217.040 2253.785 217.210 ;
        RECT 2253.955 217.040 2254.100 217.210 ;
        RECT 2259.620 217.040 2259.765 217.210 ;
        RECT 2259.935 217.040 2260.080 217.210 ;
        RECT 2265.600 217.040 2265.745 217.210 ;
        RECT 2265.915 217.040 2266.060 217.210 ;
        RECT 2271.580 217.040 2271.725 217.210 ;
        RECT 2271.895 217.040 2272.040 217.210 ;
        RECT 669.085 216.315 669.375 217.040 ;
        RECT 669.935 216.240 670.265 217.040 ;
      LAYER li1 ;
        RECT 670.435 216.390 670.605 216.870 ;
      LAYER li1 ;
        RECT 670.775 216.560 671.105 217.040 ;
      LAYER li1 ;
        RECT 671.275 216.390 671.445 216.870 ;
      LAYER li1 ;
        RECT 671.615 216.560 671.945 217.040 ;
      LAYER li1 ;
        RECT 672.115 216.390 672.285 216.870 ;
      LAYER li1 ;
        RECT 672.455 216.560 672.785 217.040 ;
      LAYER li1 ;
        RECT 672.955 216.390 673.125 216.870 ;
      LAYER li1 ;
        RECT 673.295 216.560 673.625 217.040 ;
        RECT 673.795 216.390 673.965 216.865 ;
        RECT 674.135 216.560 674.465 217.040 ;
        RECT 674.635 216.390 674.805 216.870 ;
      LAYER li1 ;
        RECT 670.435 216.220 673.125 216.390 ;
      LAYER li1 ;
        RECT 673.385 216.220 674.805 216.390 ;
        RECT 675.065 216.315 675.355 217.040 ;
        RECT 675.915 216.240 676.245 217.040 ;
      LAYER li1 ;
        RECT 676.415 216.390 676.585 216.870 ;
      LAYER li1 ;
        RECT 676.755 216.560 677.085 217.040 ;
      LAYER li1 ;
        RECT 677.255 216.390 677.425 216.870 ;
      LAYER li1 ;
        RECT 677.595 216.560 677.925 217.040 ;
      LAYER li1 ;
        RECT 678.095 216.390 678.265 216.870 ;
      LAYER li1 ;
        RECT 678.435 216.560 678.765 217.040 ;
      LAYER li1 ;
        RECT 678.935 216.390 679.105 216.870 ;
      LAYER li1 ;
        RECT 679.275 216.560 679.605 217.040 ;
        RECT 679.775 216.390 679.945 216.865 ;
        RECT 680.115 216.560 680.445 217.040 ;
        RECT 680.615 216.390 680.785 216.870 ;
      LAYER li1 ;
        RECT 676.415 216.220 679.105 216.390 ;
      LAYER li1 ;
        RECT 679.365 216.220 680.785 216.390 ;
        RECT 681.045 216.315 681.335 217.040 ;
        RECT 681.895 216.240 682.225 217.040 ;
      LAYER li1 ;
        RECT 682.395 216.390 682.565 216.870 ;
      LAYER li1 ;
        RECT 682.735 216.560 683.065 217.040 ;
      LAYER li1 ;
        RECT 683.235 216.390 683.405 216.870 ;
      LAYER li1 ;
        RECT 683.575 216.560 683.905 217.040 ;
      LAYER li1 ;
        RECT 684.075 216.390 684.245 216.870 ;
      LAYER li1 ;
        RECT 684.415 216.560 684.745 217.040 ;
      LAYER li1 ;
        RECT 684.915 216.390 685.085 216.870 ;
      LAYER li1 ;
        RECT 685.255 216.560 685.585 217.040 ;
        RECT 685.755 216.390 685.925 216.865 ;
        RECT 686.095 216.560 686.425 217.040 ;
        RECT 686.595 216.390 686.765 216.870 ;
      LAYER li1 ;
        RECT 682.395 216.220 685.085 216.390 ;
      LAYER li1 ;
        RECT 685.345 216.220 686.765 216.390 ;
        RECT 687.025 216.315 687.315 217.040 ;
        RECT 687.875 216.240 688.205 217.040 ;
      LAYER li1 ;
        RECT 688.375 216.390 688.545 216.870 ;
      LAYER li1 ;
        RECT 688.715 216.560 689.045 217.040 ;
      LAYER li1 ;
        RECT 689.215 216.390 689.385 216.870 ;
      LAYER li1 ;
        RECT 689.555 216.560 689.885 217.040 ;
      LAYER li1 ;
        RECT 690.055 216.390 690.225 216.870 ;
      LAYER li1 ;
        RECT 690.395 216.560 690.725 217.040 ;
      LAYER li1 ;
        RECT 690.895 216.390 691.065 216.870 ;
      LAYER li1 ;
        RECT 691.235 216.560 691.565 217.040 ;
        RECT 691.735 216.390 691.905 216.865 ;
        RECT 692.075 216.560 692.405 217.040 ;
        RECT 692.575 216.390 692.745 216.870 ;
      LAYER li1 ;
        RECT 688.375 216.220 691.065 216.390 ;
      LAYER li1 ;
        RECT 691.325 216.220 692.745 216.390 ;
        RECT 693.005 216.315 693.295 217.040 ;
        RECT 693.855 216.240 694.185 217.040 ;
      LAYER li1 ;
        RECT 694.355 216.390 694.525 216.870 ;
      LAYER li1 ;
        RECT 694.695 216.560 695.025 217.040 ;
      LAYER li1 ;
        RECT 695.195 216.390 695.365 216.870 ;
      LAYER li1 ;
        RECT 695.535 216.560 695.865 217.040 ;
      LAYER li1 ;
        RECT 696.035 216.390 696.205 216.870 ;
      LAYER li1 ;
        RECT 696.375 216.560 696.705 217.040 ;
      LAYER li1 ;
        RECT 696.875 216.390 697.045 216.870 ;
      LAYER li1 ;
        RECT 697.215 216.560 697.545 217.040 ;
        RECT 697.715 216.390 697.885 216.865 ;
        RECT 698.055 216.560 698.385 217.040 ;
        RECT 698.555 216.390 698.725 216.870 ;
      LAYER li1 ;
        RECT 694.355 216.220 697.045 216.390 ;
      LAYER li1 ;
        RECT 697.305 216.220 698.725 216.390 ;
        RECT 698.985 216.315 699.275 217.040 ;
        RECT 699.835 216.240 700.165 217.040 ;
      LAYER li1 ;
        RECT 700.335 216.390 700.505 216.870 ;
      LAYER li1 ;
        RECT 700.675 216.560 701.005 217.040 ;
      LAYER li1 ;
        RECT 701.175 216.390 701.345 216.870 ;
      LAYER li1 ;
        RECT 701.515 216.560 701.845 217.040 ;
      LAYER li1 ;
        RECT 702.015 216.390 702.185 216.870 ;
      LAYER li1 ;
        RECT 702.355 216.560 702.685 217.040 ;
      LAYER li1 ;
        RECT 702.855 216.390 703.025 216.870 ;
      LAYER li1 ;
        RECT 703.195 216.560 703.525 217.040 ;
        RECT 703.695 216.390 703.865 216.865 ;
        RECT 704.035 216.560 704.365 217.040 ;
        RECT 704.535 216.390 704.705 216.870 ;
      LAYER li1 ;
        RECT 700.335 216.220 703.025 216.390 ;
      LAYER li1 ;
        RECT 703.285 216.220 704.705 216.390 ;
        RECT 704.965 216.315 705.255 217.040 ;
        RECT 705.815 216.240 706.145 217.040 ;
      LAYER li1 ;
        RECT 706.315 216.390 706.485 216.870 ;
      LAYER li1 ;
        RECT 706.655 216.560 706.985 217.040 ;
      LAYER li1 ;
        RECT 707.155 216.390 707.325 216.870 ;
      LAYER li1 ;
        RECT 707.495 216.560 707.825 217.040 ;
      LAYER li1 ;
        RECT 707.995 216.390 708.165 216.870 ;
      LAYER li1 ;
        RECT 708.335 216.560 708.665 217.040 ;
      LAYER li1 ;
        RECT 708.835 216.390 709.005 216.870 ;
      LAYER li1 ;
        RECT 709.175 216.560 709.505 217.040 ;
        RECT 709.675 216.390 709.845 216.865 ;
        RECT 710.015 216.560 710.345 217.040 ;
        RECT 710.515 216.390 710.685 216.870 ;
      LAYER li1 ;
        RECT 706.315 216.220 709.005 216.390 ;
      LAYER li1 ;
        RECT 709.265 216.220 710.685 216.390 ;
        RECT 710.945 216.315 711.235 217.040 ;
        RECT 711.795 216.240 712.125 217.040 ;
      LAYER li1 ;
        RECT 712.295 216.390 712.465 216.870 ;
      LAYER li1 ;
        RECT 712.635 216.560 712.965 217.040 ;
      LAYER li1 ;
        RECT 713.135 216.390 713.305 216.870 ;
      LAYER li1 ;
        RECT 713.475 216.560 713.805 217.040 ;
      LAYER li1 ;
        RECT 713.975 216.390 714.145 216.870 ;
      LAYER li1 ;
        RECT 714.315 216.560 714.645 217.040 ;
      LAYER li1 ;
        RECT 714.815 216.390 714.985 216.870 ;
      LAYER li1 ;
        RECT 715.155 216.560 715.485 217.040 ;
        RECT 715.655 216.390 715.825 216.865 ;
        RECT 715.995 216.560 716.325 217.040 ;
        RECT 716.495 216.390 716.665 216.870 ;
      LAYER li1 ;
        RECT 712.295 216.220 714.985 216.390 ;
      LAYER li1 ;
        RECT 715.245 216.220 716.665 216.390 ;
        RECT 716.925 216.315 717.215 217.040 ;
        RECT 717.775 216.240 718.105 217.040 ;
      LAYER li1 ;
        RECT 718.275 216.390 718.445 216.870 ;
      LAYER li1 ;
        RECT 718.615 216.560 718.945 217.040 ;
      LAYER li1 ;
        RECT 719.115 216.390 719.285 216.870 ;
      LAYER li1 ;
        RECT 719.455 216.560 719.785 217.040 ;
      LAYER li1 ;
        RECT 719.955 216.390 720.125 216.870 ;
      LAYER li1 ;
        RECT 720.295 216.560 720.625 217.040 ;
      LAYER li1 ;
        RECT 720.795 216.390 720.965 216.870 ;
      LAYER li1 ;
        RECT 721.135 216.560 721.465 217.040 ;
        RECT 721.635 216.390 721.805 216.865 ;
        RECT 721.975 216.560 722.305 217.040 ;
        RECT 722.475 216.390 722.645 216.870 ;
      LAYER li1 ;
        RECT 718.275 216.220 720.965 216.390 ;
      LAYER li1 ;
        RECT 721.225 216.220 722.645 216.390 ;
        RECT 722.905 216.315 723.195 217.040 ;
        RECT 728.885 216.315 729.175 217.040 ;
        RECT 758.785 216.315 759.075 217.040 ;
        RECT 759.635 216.240 759.965 217.040 ;
        RECT 760.475 216.560 760.805 217.040 ;
        RECT 761.315 216.560 761.645 217.040 ;
        RECT 762.155 216.560 762.485 217.040 ;
        RECT 762.995 216.560 763.325 217.040 ;
        RECT 763.495 216.390 763.665 216.865 ;
        RECT 763.835 216.560 764.165 217.040 ;
        RECT 764.335 216.390 764.505 216.870 ;
        RECT 763.085 216.220 764.505 216.390 ;
        RECT 764.765 216.315 765.055 217.040 ;
        RECT 765.615 216.240 765.945 217.040 ;
        RECT 766.455 216.560 766.785 217.040 ;
        RECT 767.295 216.560 767.625 217.040 ;
        RECT 768.135 216.560 768.465 217.040 ;
        RECT 768.975 216.560 769.305 217.040 ;
        RECT 769.475 216.390 769.645 216.865 ;
        RECT 769.815 216.560 770.145 217.040 ;
        RECT 770.315 216.390 770.485 216.870 ;
        RECT 769.065 216.220 770.485 216.390 ;
        RECT 770.745 216.315 771.035 217.040 ;
        RECT 771.595 216.240 771.925 217.040 ;
        RECT 772.435 216.560 772.765 217.040 ;
        RECT 773.275 216.560 773.605 217.040 ;
        RECT 774.115 216.560 774.445 217.040 ;
        RECT 774.955 216.560 775.285 217.040 ;
        RECT 775.455 216.390 775.625 216.865 ;
        RECT 775.795 216.560 776.125 217.040 ;
        RECT 776.295 216.390 776.465 216.870 ;
        RECT 775.045 216.220 776.465 216.390 ;
        RECT 776.725 216.315 777.015 217.040 ;
        RECT 777.575 216.240 777.905 217.040 ;
        RECT 778.415 216.560 778.745 217.040 ;
        RECT 779.255 216.560 779.585 217.040 ;
        RECT 780.095 216.560 780.425 217.040 ;
        RECT 780.935 216.560 781.265 217.040 ;
        RECT 781.435 216.390 781.605 216.865 ;
        RECT 781.775 216.560 782.105 217.040 ;
        RECT 782.275 216.390 782.445 216.870 ;
        RECT 781.025 216.220 782.445 216.390 ;
        RECT 782.705 216.315 782.995 217.040 ;
        RECT 783.555 216.240 783.885 217.040 ;
        RECT 784.395 216.560 784.725 217.040 ;
        RECT 785.235 216.560 785.565 217.040 ;
        RECT 786.075 216.560 786.405 217.040 ;
        RECT 786.915 216.560 787.245 217.040 ;
        RECT 787.415 216.390 787.585 216.865 ;
        RECT 787.755 216.560 788.085 217.040 ;
        RECT 788.255 216.390 788.425 216.870 ;
        RECT 787.005 216.220 788.425 216.390 ;
        RECT 788.685 216.315 788.975 217.040 ;
        RECT 789.535 216.240 789.865 217.040 ;
        RECT 790.375 216.560 790.705 217.040 ;
        RECT 791.215 216.560 791.545 217.040 ;
        RECT 792.055 216.560 792.385 217.040 ;
        RECT 792.895 216.560 793.225 217.040 ;
        RECT 793.395 216.390 793.565 216.865 ;
        RECT 793.735 216.560 794.065 217.040 ;
        RECT 794.235 216.390 794.405 216.870 ;
        RECT 792.985 216.220 794.405 216.390 ;
        RECT 794.665 216.315 794.955 217.040 ;
        RECT 2146.085 216.315 2146.375 217.040 ;
        RECT 2146.935 216.240 2147.265 217.040 ;
      LAYER li1 ;
        RECT 2147.435 216.390 2147.605 216.870 ;
      LAYER li1 ;
        RECT 2147.775 216.560 2148.105 217.040 ;
      LAYER li1 ;
        RECT 2148.275 216.390 2148.445 216.870 ;
      LAYER li1 ;
        RECT 2148.615 216.560 2148.945 217.040 ;
      LAYER li1 ;
        RECT 2149.115 216.390 2149.285 216.870 ;
      LAYER li1 ;
        RECT 2149.455 216.560 2149.785 217.040 ;
      LAYER li1 ;
        RECT 2149.955 216.390 2150.125 216.870 ;
      LAYER li1 ;
        RECT 2150.295 216.560 2150.625 217.040 ;
        RECT 2150.795 216.390 2150.965 216.865 ;
        RECT 2151.135 216.560 2151.465 217.040 ;
        RECT 2151.635 216.390 2151.805 216.870 ;
      LAYER li1 ;
        RECT 2147.435 216.220 2150.125 216.390 ;
      LAYER li1 ;
        RECT 2150.385 216.220 2151.805 216.390 ;
        RECT 2152.065 216.315 2152.355 217.040 ;
        RECT 2152.915 216.240 2153.245 217.040 ;
      LAYER li1 ;
        RECT 2153.415 216.390 2153.585 216.870 ;
      LAYER li1 ;
        RECT 2153.755 216.560 2154.085 217.040 ;
      LAYER li1 ;
        RECT 2154.255 216.390 2154.425 216.870 ;
      LAYER li1 ;
        RECT 2154.595 216.560 2154.925 217.040 ;
      LAYER li1 ;
        RECT 2155.095 216.390 2155.265 216.870 ;
      LAYER li1 ;
        RECT 2155.435 216.560 2155.765 217.040 ;
      LAYER li1 ;
        RECT 2155.935 216.390 2156.105 216.870 ;
      LAYER li1 ;
        RECT 2156.275 216.560 2156.605 217.040 ;
        RECT 2156.775 216.390 2156.945 216.865 ;
        RECT 2157.115 216.560 2157.445 217.040 ;
        RECT 2157.615 216.390 2157.785 216.870 ;
      LAYER li1 ;
        RECT 2153.415 216.220 2156.105 216.390 ;
      LAYER li1 ;
        RECT 2156.365 216.220 2157.785 216.390 ;
        RECT 2158.045 216.315 2158.335 217.040 ;
        RECT 2158.895 216.240 2159.225 217.040 ;
      LAYER li1 ;
        RECT 2159.395 216.390 2159.565 216.870 ;
      LAYER li1 ;
        RECT 2159.735 216.560 2160.065 217.040 ;
      LAYER li1 ;
        RECT 2160.235 216.390 2160.405 216.870 ;
      LAYER li1 ;
        RECT 2160.575 216.560 2160.905 217.040 ;
      LAYER li1 ;
        RECT 2161.075 216.390 2161.245 216.870 ;
      LAYER li1 ;
        RECT 2161.415 216.560 2161.745 217.040 ;
      LAYER li1 ;
        RECT 2161.915 216.390 2162.085 216.870 ;
      LAYER li1 ;
        RECT 2162.255 216.560 2162.585 217.040 ;
        RECT 2162.755 216.390 2162.925 216.865 ;
        RECT 2163.095 216.560 2163.425 217.040 ;
        RECT 2163.595 216.390 2163.765 216.870 ;
      LAYER li1 ;
        RECT 2159.395 216.220 2162.085 216.390 ;
      LAYER li1 ;
        RECT 2162.345 216.220 2163.765 216.390 ;
        RECT 2164.025 216.315 2164.315 217.040 ;
        RECT 2164.875 216.240 2165.205 217.040 ;
      LAYER li1 ;
        RECT 2165.375 216.390 2165.545 216.870 ;
      LAYER li1 ;
        RECT 2165.715 216.560 2166.045 217.040 ;
      LAYER li1 ;
        RECT 2166.215 216.390 2166.385 216.870 ;
      LAYER li1 ;
        RECT 2166.555 216.560 2166.885 217.040 ;
      LAYER li1 ;
        RECT 2167.055 216.390 2167.225 216.870 ;
      LAYER li1 ;
        RECT 2167.395 216.560 2167.725 217.040 ;
      LAYER li1 ;
        RECT 2167.895 216.390 2168.065 216.870 ;
      LAYER li1 ;
        RECT 2168.235 216.560 2168.565 217.040 ;
        RECT 2168.735 216.390 2168.905 216.865 ;
        RECT 2169.075 216.560 2169.405 217.040 ;
        RECT 2169.575 216.390 2169.745 216.870 ;
      LAYER li1 ;
        RECT 2165.375 216.220 2168.065 216.390 ;
      LAYER li1 ;
        RECT 2168.325 216.220 2169.745 216.390 ;
        RECT 2170.005 216.315 2170.295 217.040 ;
        RECT 2170.855 216.240 2171.185 217.040 ;
      LAYER li1 ;
        RECT 2171.355 216.390 2171.525 216.870 ;
      LAYER li1 ;
        RECT 2171.695 216.560 2172.025 217.040 ;
      LAYER li1 ;
        RECT 2172.195 216.390 2172.365 216.870 ;
      LAYER li1 ;
        RECT 2172.535 216.560 2172.865 217.040 ;
      LAYER li1 ;
        RECT 2173.035 216.390 2173.205 216.870 ;
      LAYER li1 ;
        RECT 2173.375 216.560 2173.705 217.040 ;
      LAYER li1 ;
        RECT 2173.875 216.390 2174.045 216.870 ;
      LAYER li1 ;
        RECT 2174.215 216.560 2174.545 217.040 ;
        RECT 2174.715 216.390 2174.885 216.865 ;
        RECT 2175.055 216.560 2175.385 217.040 ;
        RECT 2175.555 216.390 2175.725 216.870 ;
      LAYER li1 ;
        RECT 2171.355 216.220 2174.045 216.390 ;
      LAYER li1 ;
        RECT 2174.305 216.220 2175.725 216.390 ;
        RECT 2175.985 216.315 2176.275 217.040 ;
        RECT 2176.835 216.240 2177.165 217.040 ;
      LAYER li1 ;
        RECT 2177.335 216.390 2177.505 216.870 ;
      LAYER li1 ;
        RECT 2177.675 216.560 2178.005 217.040 ;
      LAYER li1 ;
        RECT 2178.175 216.390 2178.345 216.870 ;
      LAYER li1 ;
        RECT 2178.515 216.560 2178.845 217.040 ;
      LAYER li1 ;
        RECT 2179.015 216.390 2179.185 216.870 ;
      LAYER li1 ;
        RECT 2179.355 216.560 2179.685 217.040 ;
      LAYER li1 ;
        RECT 2179.855 216.390 2180.025 216.870 ;
      LAYER li1 ;
        RECT 2180.195 216.560 2180.525 217.040 ;
        RECT 2180.695 216.390 2180.865 216.865 ;
        RECT 2181.035 216.560 2181.365 217.040 ;
        RECT 2181.535 216.390 2181.705 216.870 ;
      LAYER li1 ;
        RECT 2177.335 216.220 2180.025 216.390 ;
      LAYER li1 ;
        RECT 2180.285 216.220 2181.705 216.390 ;
        RECT 2181.965 216.315 2182.255 217.040 ;
        RECT 2182.815 216.240 2183.145 217.040 ;
      LAYER li1 ;
        RECT 2183.315 216.390 2183.485 216.870 ;
      LAYER li1 ;
        RECT 2183.655 216.560 2183.985 217.040 ;
      LAYER li1 ;
        RECT 2184.155 216.390 2184.325 216.870 ;
      LAYER li1 ;
        RECT 2184.495 216.560 2184.825 217.040 ;
      LAYER li1 ;
        RECT 2184.995 216.390 2185.165 216.870 ;
      LAYER li1 ;
        RECT 2185.335 216.560 2185.665 217.040 ;
      LAYER li1 ;
        RECT 2185.835 216.390 2186.005 216.870 ;
      LAYER li1 ;
        RECT 2186.175 216.560 2186.505 217.040 ;
        RECT 2186.675 216.390 2186.845 216.865 ;
        RECT 2187.015 216.560 2187.345 217.040 ;
        RECT 2187.515 216.390 2187.685 216.870 ;
      LAYER li1 ;
        RECT 2183.315 216.220 2186.005 216.390 ;
      LAYER li1 ;
        RECT 2186.265 216.220 2187.685 216.390 ;
        RECT 2187.945 216.315 2188.235 217.040 ;
        RECT 2188.795 216.240 2189.125 217.040 ;
      LAYER li1 ;
        RECT 2189.295 216.390 2189.465 216.870 ;
      LAYER li1 ;
        RECT 2189.635 216.560 2189.965 217.040 ;
      LAYER li1 ;
        RECT 2190.135 216.390 2190.305 216.870 ;
      LAYER li1 ;
        RECT 2190.475 216.560 2190.805 217.040 ;
      LAYER li1 ;
        RECT 2190.975 216.390 2191.145 216.870 ;
      LAYER li1 ;
        RECT 2191.315 216.560 2191.645 217.040 ;
      LAYER li1 ;
        RECT 2191.815 216.390 2191.985 216.870 ;
      LAYER li1 ;
        RECT 2192.155 216.560 2192.485 217.040 ;
        RECT 2192.655 216.390 2192.825 216.865 ;
        RECT 2192.995 216.560 2193.325 217.040 ;
        RECT 2193.495 216.390 2193.665 216.870 ;
      LAYER li1 ;
        RECT 2189.295 216.220 2191.985 216.390 ;
      LAYER li1 ;
        RECT 2192.245 216.220 2193.665 216.390 ;
        RECT 2193.925 216.315 2194.215 217.040 ;
        RECT 2194.775 216.240 2195.105 217.040 ;
      LAYER li1 ;
        RECT 2195.275 216.390 2195.445 216.870 ;
      LAYER li1 ;
        RECT 2195.615 216.560 2195.945 217.040 ;
      LAYER li1 ;
        RECT 2196.115 216.390 2196.285 216.870 ;
      LAYER li1 ;
        RECT 2196.455 216.560 2196.785 217.040 ;
      LAYER li1 ;
        RECT 2196.955 216.390 2197.125 216.870 ;
      LAYER li1 ;
        RECT 2197.295 216.560 2197.625 217.040 ;
      LAYER li1 ;
        RECT 2197.795 216.390 2197.965 216.870 ;
      LAYER li1 ;
        RECT 2198.135 216.560 2198.465 217.040 ;
        RECT 2198.635 216.390 2198.805 216.865 ;
        RECT 2198.975 216.560 2199.305 217.040 ;
        RECT 2199.475 216.390 2199.645 216.870 ;
      LAYER li1 ;
        RECT 2195.275 216.220 2197.965 216.390 ;
      LAYER li1 ;
        RECT 2198.225 216.220 2199.645 216.390 ;
        RECT 2199.905 216.315 2200.195 217.040 ;
        RECT 2205.885 216.315 2206.175 217.040 ;
        RECT 2235.785 216.315 2236.075 217.040 ;
        RECT 2236.635 216.240 2236.965 217.040 ;
      LAYER li1 ;
        RECT 2237.135 216.390 2237.305 216.870 ;
      LAYER li1 ;
        RECT 2237.475 216.560 2237.805 217.040 ;
      LAYER li1 ;
        RECT 2237.975 216.390 2238.145 216.870 ;
      LAYER li1 ;
        RECT 2238.315 216.560 2238.645 217.040 ;
      LAYER li1 ;
        RECT 2238.815 216.390 2238.985 216.870 ;
      LAYER li1 ;
        RECT 2239.155 216.560 2239.485 217.040 ;
      LAYER li1 ;
        RECT 2239.655 216.390 2239.825 216.870 ;
      LAYER li1 ;
        RECT 2239.995 216.560 2240.325 217.040 ;
        RECT 2240.495 216.390 2240.665 216.865 ;
        RECT 2240.835 216.560 2241.165 217.040 ;
        RECT 2241.335 216.390 2241.505 216.870 ;
      LAYER li1 ;
        RECT 2237.135 216.220 2239.825 216.390 ;
      LAYER li1 ;
        RECT 2240.085 216.220 2241.505 216.390 ;
        RECT 2241.765 216.315 2242.055 217.040 ;
        RECT 2242.615 216.240 2242.945 217.040 ;
      LAYER li1 ;
        RECT 2243.115 216.390 2243.285 216.870 ;
      LAYER li1 ;
        RECT 2243.455 216.560 2243.785 217.040 ;
      LAYER li1 ;
        RECT 2243.955 216.390 2244.125 216.870 ;
      LAYER li1 ;
        RECT 2244.295 216.560 2244.625 217.040 ;
      LAYER li1 ;
        RECT 2244.795 216.390 2244.965 216.870 ;
      LAYER li1 ;
        RECT 2245.135 216.560 2245.465 217.040 ;
      LAYER li1 ;
        RECT 2245.635 216.390 2245.805 216.870 ;
      LAYER li1 ;
        RECT 2245.975 216.560 2246.305 217.040 ;
        RECT 2246.475 216.390 2246.645 216.865 ;
        RECT 2246.815 216.560 2247.145 217.040 ;
        RECT 2247.315 216.390 2247.485 216.870 ;
      LAYER li1 ;
        RECT 2243.115 216.220 2245.805 216.390 ;
      LAYER li1 ;
        RECT 2246.065 216.220 2247.485 216.390 ;
        RECT 2247.745 216.315 2248.035 217.040 ;
        RECT 2248.595 216.240 2248.925 217.040 ;
      LAYER li1 ;
        RECT 2249.095 216.390 2249.265 216.870 ;
      LAYER li1 ;
        RECT 2249.435 216.560 2249.765 217.040 ;
      LAYER li1 ;
        RECT 2249.935 216.390 2250.105 216.870 ;
      LAYER li1 ;
        RECT 2250.275 216.560 2250.605 217.040 ;
      LAYER li1 ;
        RECT 2250.775 216.390 2250.945 216.870 ;
      LAYER li1 ;
        RECT 2251.115 216.560 2251.445 217.040 ;
      LAYER li1 ;
        RECT 2251.615 216.390 2251.785 216.870 ;
      LAYER li1 ;
        RECT 2251.955 216.560 2252.285 217.040 ;
        RECT 2252.455 216.390 2252.625 216.865 ;
        RECT 2252.795 216.560 2253.125 217.040 ;
        RECT 2253.295 216.390 2253.465 216.870 ;
      LAYER li1 ;
        RECT 2249.095 216.220 2251.785 216.390 ;
      LAYER li1 ;
        RECT 2252.045 216.220 2253.465 216.390 ;
        RECT 2253.725 216.315 2254.015 217.040 ;
        RECT 2254.575 216.240 2254.905 217.040 ;
      LAYER li1 ;
        RECT 2255.075 216.390 2255.245 216.870 ;
      LAYER li1 ;
        RECT 2255.415 216.560 2255.745 217.040 ;
      LAYER li1 ;
        RECT 2255.915 216.390 2256.085 216.870 ;
      LAYER li1 ;
        RECT 2256.255 216.560 2256.585 217.040 ;
      LAYER li1 ;
        RECT 2256.755 216.390 2256.925 216.870 ;
      LAYER li1 ;
        RECT 2257.095 216.560 2257.425 217.040 ;
      LAYER li1 ;
        RECT 2257.595 216.390 2257.765 216.870 ;
      LAYER li1 ;
        RECT 2257.935 216.560 2258.265 217.040 ;
        RECT 2258.435 216.390 2258.605 216.865 ;
        RECT 2258.775 216.560 2259.105 217.040 ;
        RECT 2259.275 216.390 2259.445 216.870 ;
      LAYER li1 ;
        RECT 2255.075 216.220 2257.765 216.390 ;
      LAYER li1 ;
        RECT 2258.025 216.220 2259.445 216.390 ;
        RECT 2259.705 216.315 2259.995 217.040 ;
        RECT 2260.555 216.240 2260.885 217.040 ;
      LAYER li1 ;
        RECT 2261.055 216.390 2261.225 216.870 ;
      LAYER li1 ;
        RECT 2261.395 216.560 2261.725 217.040 ;
      LAYER li1 ;
        RECT 2261.895 216.390 2262.065 216.870 ;
      LAYER li1 ;
        RECT 2262.235 216.560 2262.565 217.040 ;
      LAYER li1 ;
        RECT 2262.735 216.390 2262.905 216.870 ;
      LAYER li1 ;
        RECT 2263.075 216.560 2263.405 217.040 ;
      LAYER li1 ;
        RECT 2263.575 216.390 2263.745 216.870 ;
      LAYER li1 ;
        RECT 2263.915 216.560 2264.245 217.040 ;
        RECT 2264.415 216.390 2264.585 216.865 ;
        RECT 2264.755 216.560 2265.085 217.040 ;
        RECT 2265.255 216.390 2265.425 216.870 ;
      LAYER li1 ;
        RECT 2261.055 216.220 2263.745 216.390 ;
      LAYER li1 ;
        RECT 2264.005 216.220 2265.425 216.390 ;
        RECT 2265.685 216.315 2265.975 217.040 ;
        RECT 2266.535 216.240 2266.865 217.040 ;
      LAYER li1 ;
        RECT 2267.035 216.390 2267.205 216.870 ;
      LAYER li1 ;
        RECT 2267.375 216.560 2267.705 217.040 ;
      LAYER li1 ;
        RECT 2267.875 216.390 2268.045 216.870 ;
      LAYER li1 ;
        RECT 2268.215 216.560 2268.545 217.040 ;
      LAYER li1 ;
        RECT 2268.715 216.390 2268.885 216.870 ;
      LAYER li1 ;
        RECT 2269.055 216.560 2269.385 217.040 ;
      LAYER li1 ;
        RECT 2269.555 216.390 2269.725 216.870 ;
      LAYER li1 ;
        RECT 2269.895 216.560 2270.225 217.040 ;
        RECT 2270.395 216.390 2270.565 216.865 ;
        RECT 2270.735 216.560 2271.065 217.040 ;
        RECT 2271.235 216.390 2271.405 216.870 ;
      LAYER li1 ;
        RECT 2267.035 216.220 2269.725 216.390 ;
      LAYER li1 ;
        RECT 2269.985 216.220 2271.405 216.390 ;
        RECT 2271.665 216.315 2271.955 217.040 ;
      LAYER li1 ;
        RECT 670.435 215.680 670.690 216.220 ;
      LAYER li1 ;
        RECT 673.385 216.050 673.560 216.220 ;
        RECT 670.935 215.880 673.560 216.050 ;
        RECT 673.385 215.680 673.560 215.880 ;
      LAYER li1 ;
        RECT 673.740 215.850 675.330 216.050 ;
        RECT 676.415 215.680 676.670 216.220 ;
      LAYER li1 ;
        RECT 679.365 216.050 679.540 216.220 ;
        RECT 676.915 215.880 679.540 216.050 ;
        RECT 679.365 215.680 679.540 215.880 ;
      LAYER li1 ;
        RECT 679.720 215.850 681.310 216.050 ;
        RECT 682.395 215.680 682.650 216.220 ;
      LAYER li1 ;
        RECT 685.345 216.050 685.520 216.220 ;
        RECT 682.895 215.880 685.520 216.050 ;
        RECT 685.345 215.680 685.520 215.880 ;
      LAYER li1 ;
        RECT 685.700 215.850 687.290 216.050 ;
        RECT 688.375 215.680 688.630 216.220 ;
      LAYER li1 ;
        RECT 691.325 216.050 691.500 216.220 ;
        RECT 688.875 215.880 691.500 216.050 ;
        RECT 691.325 215.680 691.500 215.880 ;
      LAYER li1 ;
        RECT 691.680 215.850 693.270 216.050 ;
        RECT 694.355 215.680 694.610 216.220 ;
      LAYER li1 ;
        RECT 697.305 216.050 697.480 216.220 ;
        RECT 694.855 215.880 697.480 216.050 ;
        RECT 697.305 215.680 697.480 215.880 ;
      LAYER li1 ;
        RECT 697.660 215.850 699.250 216.050 ;
        RECT 700.335 215.680 700.590 216.220 ;
      LAYER li1 ;
        RECT 703.285 216.050 703.460 216.220 ;
        RECT 700.835 215.880 703.460 216.050 ;
        RECT 703.285 215.680 703.460 215.880 ;
      LAYER li1 ;
        RECT 703.640 215.850 705.230 216.050 ;
        RECT 706.315 215.680 706.570 216.220 ;
      LAYER li1 ;
        RECT 709.265 216.050 709.440 216.220 ;
        RECT 706.815 215.880 709.440 216.050 ;
        RECT 709.265 215.680 709.440 215.880 ;
      LAYER li1 ;
        RECT 709.620 215.850 711.210 216.050 ;
        RECT 712.295 215.680 712.550 216.220 ;
      LAYER li1 ;
        RECT 715.245 216.050 715.420 216.220 ;
        RECT 712.795 215.880 715.420 216.050 ;
        RECT 715.245 215.680 715.420 215.880 ;
      LAYER li1 ;
        RECT 715.600 215.850 717.190 216.050 ;
        RECT 718.275 215.680 718.530 216.220 ;
      LAYER li1 ;
        RECT 721.225 216.050 721.400 216.220 ;
        RECT 718.775 215.880 721.400 216.050 ;
        RECT 721.225 215.680 721.400 215.880 ;
      LAYER li1 ;
        RECT 721.580 215.850 723.170 216.050 ;
      LAYER li1 ;
        RECT 669.085 214.490 669.375 215.655 ;
        RECT 669.935 214.490 670.265 215.640 ;
      LAYER li1 ;
        RECT 670.435 215.510 673.125 215.680 ;
      LAYER li1 ;
        RECT 673.385 215.510 674.885 215.680 ;
      LAYER li1 ;
        RECT 670.435 214.660 670.605 215.510 ;
      LAYER li1 ;
        RECT 670.775 214.490 671.105 215.290 ;
      LAYER li1 ;
        RECT 671.275 214.660 671.445 215.510 ;
      LAYER li1 ;
        RECT 671.615 214.490 671.945 215.290 ;
      LAYER li1 ;
        RECT 672.115 214.660 672.285 215.510 ;
      LAYER li1 ;
        RECT 672.455 214.490 672.785 215.290 ;
      LAYER li1 ;
        RECT 672.955 214.660 673.125 215.510 ;
      LAYER li1 ;
        RECT 673.375 214.490 673.545 215.290 ;
        RECT 673.715 214.660 674.045 215.510 ;
        RECT 674.215 214.490 674.385 215.290 ;
        RECT 674.555 214.660 674.885 215.510 ;
        RECT 675.065 214.490 675.355 215.655 ;
        RECT 675.915 214.490 676.245 215.640 ;
      LAYER li1 ;
        RECT 676.415 215.510 679.105 215.680 ;
      LAYER li1 ;
        RECT 679.365 215.510 680.865 215.680 ;
      LAYER li1 ;
        RECT 676.415 214.660 676.585 215.510 ;
      LAYER li1 ;
        RECT 676.755 214.490 677.085 215.290 ;
      LAYER li1 ;
        RECT 677.255 214.660 677.425 215.510 ;
      LAYER li1 ;
        RECT 677.595 214.490 677.925 215.290 ;
      LAYER li1 ;
        RECT 678.095 214.660 678.265 215.510 ;
      LAYER li1 ;
        RECT 678.435 214.490 678.765 215.290 ;
      LAYER li1 ;
        RECT 678.935 214.660 679.105 215.510 ;
      LAYER li1 ;
        RECT 679.355 214.490 679.525 215.290 ;
        RECT 679.695 214.660 680.025 215.510 ;
        RECT 680.195 214.490 680.365 215.290 ;
        RECT 680.535 214.660 680.865 215.510 ;
        RECT 681.045 214.490 681.335 215.655 ;
        RECT 681.895 214.490 682.225 215.640 ;
      LAYER li1 ;
        RECT 682.395 215.510 685.085 215.680 ;
      LAYER li1 ;
        RECT 685.345 215.510 686.845 215.680 ;
      LAYER li1 ;
        RECT 682.395 214.660 682.565 215.510 ;
      LAYER li1 ;
        RECT 682.735 214.490 683.065 215.290 ;
      LAYER li1 ;
        RECT 683.235 214.660 683.405 215.510 ;
      LAYER li1 ;
        RECT 683.575 214.490 683.905 215.290 ;
      LAYER li1 ;
        RECT 684.075 214.660 684.245 215.510 ;
      LAYER li1 ;
        RECT 684.415 214.490 684.745 215.290 ;
      LAYER li1 ;
        RECT 684.915 214.660 685.085 215.510 ;
      LAYER li1 ;
        RECT 685.335 214.490 685.505 215.290 ;
        RECT 685.675 214.660 686.005 215.510 ;
        RECT 686.175 214.490 686.345 215.290 ;
        RECT 686.515 214.660 686.845 215.510 ;
        RECT 687.025 214.490 687.315 215.655 ;
        RECT 687.875 214.490 688.205 215.640 ;
      LAYER li1 ;
        RECT 688.375 215.510 691.065 215.680 ;
      LAYER li1 ;
        RECT 691.325 215.510 692.825 215.680 ;
      LAYER li1 ;
        RECT 688.375 214.660 688.545 215.510 ;
      LAYER li1 ;
        RECT 688.715 214.490 689.045 215.290 ;
      LAYER li1 ;
        RECT 689.215 214.660 689.385 215.510 ;
      LAYER li1 ;
        RECT 689.555 214.490 689.885 215.290 ;
      LAYER li1 ;
        RECT 690.055 214.660 690.225 215.510 ;
      LAYER li1 ;
        RECT 690.395 214.490 690.725 215.290 ;
      LAYER li1 ;
        RECT 690.895 214.660 691.065 215.510 ;
      LAYER li1 ;
        RECT 691.315 214.490 691.485 215.290 ;
        RECT 691.655 214.660 691.985 215.510 ;
        RECT 692.155 214.490 692.325 215.290 ;
        RECT 692.495 214.660 692.825 215.510 ;
        RECT 693.005 214.490 693.295 215.655 ;
        RECT 693.855 214.490 694.185 215.640 ;
      LAYER li1 ;
        RECT 694.355 215.510 697.045 215.680 ;
      LAYER li1 ;
        RECT 697.305 215.510 698.805 215.680 ;
      LAYER li1 ;
        RECT 694.355 214.660 694.525 215.510 ;
      LAYER li1 ;
        RECT 694.695 214.490 695.025 215.290 ;
      LAYER li1 ;
        RECT 695.195 214.660 695.365 215.510 ;
      LAYER li1 ;
        RECT 695.535 214.490 695.865 215.290 ;
      LAYER li1 ;
        RECT 696.035 214.660 696.205 215.510 ;
      LAYER li1 ;
        RECT 696.375 214.490 696.705 215.290 ;
      LAYER li1 ;
        RECT 696.875 214.660 697.045 215.510 ;
      LAYER li1 ;
        RECT 697.295 214.490 697.465 215.290 ;
        RECT 697.635 214.660 697.965 215.510 ;
        RECT 698.135 214.490 698.305 215.290 ;
        RECT 698.475 214.660 698.805 215.510 ;
        RECT 698.985 214.490 699.275 215.655 ;
        RECT 699.835 214.490 700.165 215.640 ;
      LAYER li1 ;
        RECT 700.335 215.510 703.025 215.680 ;
      LAYER li1 ;
        RECT 703.285 215.510 704.785 215.680 ;
      LAYER li1 ;
        RECT 700.335 214.660 700.505 215.510 ;
      LAYER li1 ;
        RECT 700.675 214.490 701.005 215.290 ;
      LAYER li1 ;
        RECT 701.175 214.660 701.345 215.510 ;
      LAYER li1 ;
        RECT 701.515 214.490 701.845 215.290 ;
      LAYER li1 ;
        RECT 702.015 214.660 702.185 215.510 ;
      LAYER li1 ;
        RECT 702.355 214.490 702.685 215.290 ;
      LAYER li1 ;
        RECT 702.855 214.660 703.025 215.510 ;
      LAYER li1 ;
        RECT 703.275 214.490 703.445 215.290 ;
        RECT 703.615 214.660 703.945 215.510 ;
        RECT 704.115 214.490 704.285 215.290 ;
        RECT 704.455 214.660 704.785 215.510 ;
        RECT 704.965 214.490 705.255 215.655 ;
        RECT 705.815 214.490 706.145 215.640 ;
      LAYER li1 ;
        RECT 706.315 215.510 709.005 215.680 ;
      LAYER li1 ;
        RECT 709.265 215.510 710.765 215.680 ;
      LAYER li1 ;
        RECT 706.315 214.660 706.485 215.510 ;
      LAYER li1 ;
        RECT 706.655 214.490 706.985 215.290 ;
      LAYER li1 ;
        RECT 707.155 214.660 707.325 215.510 ;
      LAYER li1 ;
        RECT 707.495 214.490 707.825 215.290 ;
      LAYER li1 ;
        RECT 707.995 214.660 708.165 215.510 ;
      LAYER li1 ;
        RECT 708.335 214.490 708.665 215.290 ;
      LAYER li1 ;
        RECT 708.835 214.660 709.005 215.510 ;
      LAYER li1 ;
        RECT 709.255 214.490 709.425 215.290 ;
        RECT 709.595 214.660 709.925 215.510 ;
        RECT 710.095 214.490 710.265 215.290 ;
        RECT 710.435 214.660 710.765 215.510 ;
        RECT 710.945 214.490 711.235 215.655 ;
        RECT 711.795 214.490 712.125 215.640 ;
      LAYER li1 ;
        RECT 712.295 215.510 714.985 215.680 ;
      LAYER li1 ;
        RECT 715.245 215.510 716.745 215.680 ;
      LAYER li1 ;
        RECT 712.295 214.660 712.465 215.510 ;
      LAYER li1 ;
        RECT 712.635 214.490 712.965 215.290 ;
      LAYER li1 ;
        RECT 713.135 214.660 713.305 215.510 ;
      LAYER li1 ;
        RECT 713.475 214.490 713.805 215.290 ;
      LAYER li1 ;
        RECT 713.975 214.660 714.145 215.510 ;
      LAYER li1 ;
        RECT 714.315 214.490 714.645 215.290 ;
      LAYER li1 ;
        RECT 714.815 214.660 714.985 215.510 ;
      LAYER li1 ;
        RECT 715.235 214.490 715.405 215.290 ;
        RECT 715.575 214.660 715.905 215.510 ;
        RECT 716.075 214.490 716.245 215.290 ;
        RECT 716.415 214.660 716.745 215.510 ;
        RECT 716.925 214.490 717.215 215.655 ;
        RECT 717.775 214.490 718.105 215.640 ;
      LAYER li1 ;
        RECT 718.275 215.510 720.965 215.680 ;
      LAYER li1 ;
        RECT 721.225 215.510 722.725 215.680 ;
      LAYER li1 ;
        RECT 718.275 214.660 718.445 215.510 ;
      LAYER li1 ;
        RECT 718.615 214.490 718.945 215.290 ;
      LAYER li1 ;
        RECT 719.115 214.660 719.285 215.510 ;
      LAYER li1 ;
        RECT 719.455 214.490 719.785 215.290 ;
      LAYER li1 ;
        RECT 719.955 214.660 720.125 215.510 ;
      LAYER li1 ;
        RECT 720.295 214.490 720.625 215.290 ;
      LAYER li1 ;
        RECT 720.795 214.660 720.965 215.510 ;
      LAYER li1 ;
        RECT 721.215 214.490 721.385 215.290 ;
        RECT 721.555 214.660 721.885 215.510 ;
        RECT 722.055 214.490 722.225 215.290 ;
        RECT 722.395 214.660 722.725 215.510 ;
        RECT 722.905 214.490 723.195 215.655 ;
      LAYER li1 ;
        RECT 726.770 214.925 727.120 216.175 ;
      LAYER li1 ;
        RECT 763.085 216.050 763.260 216.220 ;
        RECT 769.065 216.050 769.240 216.220 ;
        RECT 775.045 216.050 775.220 216.220 ;
        RECT 781.025 216.050 781.200 216.220 ;
        RECT 787.005 216.050 787.180 216.220 ;
        RECT 792.985 216.050 793.160 216.220 ;
        RECT 760.635 215.880 763.260 216.050 ;
        RECT 763.085 215.680 763.260 215.880 ;
      LAYER li1 ;
        RECT 763.440 215.850 765.030 216.050 ;
      LAYER li1 ;
        RECT 766.615 215.880 769.240 216.050 ;
        RECT 769.065 215.680 769.240 215.880 ;
      LAYER li1 ;
        RECT 769.420 215.850 771.010 216.050 ;
      LAYER li1 ;
        RECT 772.595 215.880 775.220 216.050 ;
        RECT 775.045 215.680 775.220 215.880 ;
      LAYER li1 ;
        RECT 775.400 215.850 776.990 216.050 ;
      LAYER li1 ;
        RECT 778.575 215.880 781.200 216.050 ;
        RECT 781.025 215.680 781.200 215.880 ;
      LAYER li1 ;
        RECT 781.380 215.850 782.970 216.050 ;
      LAYER li1 ;
        RECT 784.555 215.880 787.180 216.050 ;
        RECT 787.005 215.680 787.180 215.880 ;
      LAYER li1 ;
        RECT 787.360 215.850 788.950 216.050 ;
      LAYER li1 ;
        RECT 790.535 215.880 793.160 216.050 ;
        RECT 792.985 215.680 793.160 215.880 ;
      LAYER li1 ;
        RECT 793.340 215.850 794.930 216.050 ;
        RECT 2147.435 215.680 2147.690 216.220 ;
      LAYER li1 ;
        RECT 2150.385 216.050 2150.560 216.220 ;
        RECT 2147.935 215.880 2150.560 216.050 ;
        RECT 2150.385 215.680 2150.560 215.880 ;
      LAYER li1 ;
        RECT 2153.415 215.680 2153.670 216.220 ;
      LAYER li1 ;
        RECT 2156.365 216.050 2156.540 216.220 ;
        RECT 2153.915 215.880 2156.540 216.050 ;
        RECT 2156.365 215.680 2156.540 215.880 ;
      LAYER li1 ;
        RECT 2159.395 215.680 2159.650 216.220 ;
      LAYER li1 ;
        RECT 2162.345 216.050 2162.520 216.220 ;
        RECT 2159.895 215.880 2162.520 216.050 ;
        RECT 2162.345 215.680 2162.520 215.880 ;
      LAYER li1 ;
        RECT 2165.375 215.680 2165.630 216.220 ;
      LAYER li1 ;
        RECT 2168.325 216.050 2168.500 216.220 ;
        RECT 2165.875 215.880 2168.500 216.050 ;
        RECT 2168.325 215.680 2168.500 215.880 ;
      LAYER li1 ;
        RECT 2171.355 215.680 2171.610 216.220 ;
      LAYER li1 ;
        RECT 2174.305 216.050 2174.480 216.220 ;
        RECT 2171.855 215.880 2174.480 216.050 ;
        RECT 2174.305 215.680 2174.480 215.880 ;
      LAYER li1 ;
        RECT 2177.335 215.680 2177.590 216.220 ;
      LAYER li1 ;
        RECT 2180.285 216.050 2180.460 216.220 ;
        RECT 2177.835 215.880 2180.460 216.050 ;
        RECT 2180.285 215.680 2180.460 215.880 ;
      LAYER li1 ;
        RECT 2183.315 215.680 2183.570 216.220 ;
      LAYER li1 ;
        RECT 2186.265 216.050 2186.440 216.220 ;
        RECT 2183.815 215.880 2186.440 216.050 ;
        RECT 2186.265 215.680 2186.440 215.880 ;
      LAYER li1 ;
        RECT 2189.295 215.680 2189.550 216.220 ;
      LAYER li1 ;
        RECT 2192.245 216.050 2192.420 216.220 ;
        RECT 2189.795 215.880 2192.420 216.050 ;
        RECT 2192.245 215.680 2192.420 215.880 ;
      LAYER li1 ;
        RECT 2195.275 215.680 2195.530 216.220 ;
      LAYER li1 ;
        RECT 2198.225 216.050 2198.400 216.220 ;
        RECT 2195.775 215.880 2198.400 216.050 ;
        RECT 2198.225 215.680 2198.400 215.880 ;
      LAYER li1 ;
        RECT 723.365 214.490 728.710 214.925 ;
      LAYER li1 ;
        RECT 728.885 214.490 729.175 215.655 ;
        RECT 758.785 214.490 759.075 215.655 ;
        RECT 759.635 214.490 759.965 215.640 ;
        RECT 763.085 215.510 764.585 215.680 ;
        RECT 760.475 214.490 760.805 215.290 ;
        RECT 761.315 214.490 761.645 215.290 ;
        RECT 762.155 214.490 762.485 215.290 ;
        RECT 763.075 214.490 763.245 215.290 ;
        RECT 763.415 214.660 763.745 215.510 ;
        RECT 763.915 214.490 764.085 215.290 ;
        RECT 764.255 214.660 764.585 215.510 ;
        RECT 764.765 214.490 765.055 215.655 ;
        RECT 765.615 214.490 765.945 215.640 ;
        RECT 769.065 215.510 770.565 215.680 ;
        RECT 766.455 214.490 766.785 215.290 ;
        RECT 767.295 214.490 767.625 215.290 ;
        RECT 768.135 214.490 768.465 215.290 ;
        RECT 769.055 214.490 769.225 215.290 ;
        RECT 769.395 214.660 769.725 215.510 ;
        RECT 769.895 214.490 770.065 215.290 ;
        RECT 770.235 214.660 770.565 215.510 ;
        RECT 770.745 214.490 771.035 215.655 ;
        RECT 771.595 214.490 771.925 215.640 ;
        RECT 775.045 215.510 776.545 215.680 ;
        RECT 772.435 214.490 772.765 215.290 ;
        RECT 773.275 214.490 773.605 215.290 ;
        RECT 774.115 214.490 774.445 215.290 ;
        RECT 775.035 214.490 775.205 215.290 ;
        RECT 775.375 214.660 775.705 215.510 ;
        RECT 775.875 214.490 776.045 215.290 ;
        RECT 776.215 214.660 776.545 215.510 ;
        RECT 776.725 214.490 777.015 215.655 ;
        RECT 777.575 214.490 777.905 215.640 ;
        RECT 781.025 215.510 782.525 215.680 ;
        RECT 778.415 214.490 778.745 215.290 ;
        RECT 779.255 214.490 779.585 215.290 ;
        RECT 780.095 214.490 780.425 215.290 ;
        RECT 781.015 214.490 781.185 215.290 ;
        RECT 781.355 214.660 781.685 215.510 ;
        RECT 781.855 214.490 782.025 215.290 ;
        RECT 782.195 214.660 782.525 215.510 ;
        RECT 782.705 214.490 782.995 215.655 ;
        RECT 783.555 214.490 783.885 215.640 ;
        RECT 787.005 215.510 788.505 215.680 ;
        RECT 784.395 214.490 784.725 215.290 ;
        RECT 785.235 214.490 785.565 215.290 ;
        RECT 786.075 214.490 786.405 215.290 ;
        RECT 786.995 214.490 787.165 215.290 ;
        RECT 787.335 214.660 787.665 215.510 ;
        RECT 787.835 214.490 788.005 215.290 ;
        RECT 788.175 214.660 788.505 215.510 ;
        RECT 788.685 214.490 788.975 215.655 ;
        RECT 789.535 214.490 789.865 215.640 ;
        RECT 792.985 215.510 794.485 215.680 ;
        RECT 790.375 214.490 790.705 215.290 ;
        RECT 791.215 214.490 791.545 215.290 ;
        RECT 792.055 214.490 792.385 215.290 ;
        RECT 792.975 214.490 793.145 215.290 ;
        RECT 793.315 214.660 793.645 215.510 ;
        RECT 793.815 214.490 793.985 215.290 ;
        RECT 794.155 214.660 794.485 215.510 ;
        RECT 794.665 214.490 794.955 215.655 ;
        RECT 2146.085 214.490 2146.375 215.655 ;
        RECT 2146.935 214.490 2147.265 215.640 ;
      LAYER li1 ;
        RECT 2147.435 215.510 2150.125 215.680 ;
      LAYER li1 ;
        RECT 2150.385 215.510 2151.885 215.680 ;
      LAYER li1 ;
        RECT 2147.435 214.660 2147.605 215.510 ;
      LAYER li1 ;
        RECT 2147.775 214.490 2148.105 215.290 ;
      LAYER li1 ;
        RECT 2148.275 214.660 2148.445 215.510 ;
      LAYER li1 ;
        RECT 2148.615 214.490 2148.945 215.290 ;
      LAYER li1 ;
        RECT 2149.115 214.660 2149.285 215.510 ;
      LAYER li1 ;
        RECT 2149.455 214.490 2149.785 215.290 ;
      LAYER li1 ;
        RECT 2149.955 214.660 2150.125 215.510 ;
      LAYER li1 ;
        RECT 2150.375 214.490 2150.545 215.290 ;
        RECT 2150.715 214.660 2151.045 215.510 ;
        RECT 2151.215 214.490 2151.385 215.290 ;
        RECT 2151.555 214.660 2151.885 215.510 ;
        RECT 2152.065 214.490 2152.355 215.655 ;
        RECT 2152.915 214.490 2153.245 215.640 ;
      LAYER li1 ;
        RECT 2153.415 215.510 2156.105 215.680 ;
      LAYER li1 ;
        RECT 2156.365 215.510 2157.865 215.680 ;
      LAYER li1 ;
        RECT 2153.415 214.660 2153.585 215.510 ;
      LAYER li1 ;
        RECT 2153.755 214.490 2154.085 215.290 ;
      LAYER li1 ;
        RECT 2154.255 214.660 2154.425 215.510 ;
      LAYER li1 ;
        RECT 2154.595 214.490 2154.925 215.290 ;
      LAYER li1 ;
        RECT 2155.095 214.660 2155.265 215.510 ;
      LAYER li1 ;
        RECT 2155.435 214.490 2155.765 215.290 ;
      LAYER li1 ;
        RECT 2155.935 214.660 2156.105 215.510 ;
      LAYER li1 ;
        RECT 2156.355 214.490 2156.525 215.290 ;
        RECT 2156.695 214.660 2157.025 215.510 ;
        RECT 2157.195 214.490 2157.365 215.290 ;
        RECT 2157.535 214.660 2157.865 215.510 ;
        RECT 2158.045 214.490 2158.335 215.655 ;
        RECT 2158.895 214.490 2159.225 215.640 ;
      LAYER li1 ;
        RECT 2159.395 215.510 2162.085 215.680 ;
      LAYER li1 ;
        RECT 2162.345 215.510 2163.845 215.680 ;
      LAYER li1 ;
        RECT 2159.395 214.660 2159.565 215.510 ;
      LAYER li1 ;
        RECT 2159.735 214.490 2160.065 215.290 ;
      LAYER li1 ;
        RECT 2160.235 214.660 2160.405 215.510 ;
      LAYER li1 ;
        RECT 2160.575 214.490 2160.905 215.290 ;
      LAYER li1 ;
        RECT 2161.075 214.660 2161.245 215.510 ;
      LAYER li1 ;
        RECT 2161.415 214.490 2161.745 215.290 ;
      LAYER li1 ;
        RECT 2161.915 214.660 2162.085 215.510 ;
      LAYER li1 ;
        RECT 2162.335 214.490 2162.505 215.290 ;
        RECT 2162.675 214.660 2163.005 215.510 ;
        RECT 2163.175 214.490 2163.345 215.290 ;
        RECT 2163.515 214.660 2163.845 215.510 ;
        RECT 2164.025 214.490 2164.315 215.655 ;
        RECT 2164.875 214.490 2165.205 215.640 ;
      LAYER li1 ;
        RECT 2165.375 215.510 2168.065 215.680 ;
      LAYER li1 ;
        RECT 2168.325 215.510 2169.825 215.680 ;
      LAYER li1 ;
        RECT 2165.375 214.660 2165.545 215.510 ;
      LAYER li1 ;
        RECT 2165.715 214.490 2166.045 215.290 ;
      LAYER li1 ;
        RECT 2166.215 214.660 2166.385 215.510 ;
      LAYER li1 ;
        RECT 2166.555 214.490 2166.885 215.290 ;
      LAYER li1 ;
        RECT 2167.055 214.660 2167.225 215.510 ;
      LAYER li1 ;
        RECT 2167.395 214.490 2167.725 215.290 ;
      LAYER li1 ;
        RECT 2167.895 214.660 2168.065 215.510 ;
      LAYER li1 ;
        RECT 2168.315 214.490 2168.485 215.290 ;
        RECT 2168.655 214.660 2168.985 215.510 ;
        RECT 2169.155 214.490 2169.325 215.290 ;
        RECT 2169.495 214.660 2169.825 215.510 ;
        RECT 2170.005 214.490 2170.295 215.655 ;
        RECT 2170.855 214.490 2171.185 215.640 ;
      LAYER li1 ;
        RECT 2171.355 215.510 2174.045 215.680 ;
      LAYER li1 ;
        RECT 2174.305 215.510 2175.805 215.680 ;
      LAYER li1 ;
        RECT 2171.355 214.660 2171.525 215.510 ;
      LAYER li1 ;
        RECT 2171.695 214.490 2172.025 215.290 ;
      LAYER li1 ;
        RECT 2172.195 214.660 2172.365 215.510 ;
      LAYER li1 ;
        RECT 2172.535 214.490 2172.865 215.290 ;
      LAYER li1 ;
        RECT 2173.035 214.660 2173.205 215.510 ;
      LAYER li1 ;
        RECT 2173.375 214.490 2173.705 215.290 ;
      LAYER li1 ;
        RECT 2173.875 214.660 2174.045 215.510 ;
      LAYER li1 ;
        RECT 2174.295 214.490 2174.465 215.290 ;
        RECT 2174.635 214.660 2174.965 215.510 ;
        RECT 2175.135 214.490 2175.305 215.290 ;
        RECT 2175.475 214.660 2175.805 215.510 ;
        RECT 2175.985 214.490 2176.275 215.655 ;
        RECT 2176.835 214.490 2177.165 215.640 ;
      LAYER li1 ;
        RECT 2177.335 215.510 2180.025 215.680 ;
      LAYER li1 ;
        RECT 2180.285 215.510 2181.785 215.680 ;
      LAYER li1 ;
        RECT 2177.335 214.660 2177.505 215.510 ;
      LAYER li1 ;
        RECT 2177.675 214.490 2178.005 215.290 ;
      LAYER li1 ;
        RECT 2178.175 214.660 2178.345 215.510 ;
      LAYER li1 ;
        RECT 2178.515 214.490 2178.845 215.290 ;
      LAYER li1 ;
        RECT 2179.015 214.660 2179.185 215.510 ;
      LAYER li1 ;
        RECT 2179.355 214.490 2179.685 215.290 ;
      LAYER li1 ;
        RECT 2179.855 214.660 2180.025 215.510 ;
      LAYER li1 ;
        RECT 2180.275 214.490 2180.445 215.290 ;
        RECT 2180.615 214.660 2180.945 215.510 ;
        RECT 2181.115 214.490 2181.285 215.290 ;
        RECT 2181.455 214.660 2181.785 215.510 ;
        RECT 2181.965 214.490 2182.255 215.655 ;
        RECT 2182.815 214.490 2183.145 215.640 ;
      LAYER li1 ;
        RECT 2183.315 215.510 2186.005 215.680 ;
      LAYER li1 ;
        RECT 2186.265 215.510 2187.765 215.680 ;
      LAYER li1 ;
        RECT 2183.315 214.660 2183.485 215.510 ;
      LAYER li1 ;
        RECT 2183.655 214.490 2183.985 215.290 ;
      LAYER li1 ;
        RECT 2184.155 214.660 2184.325 215.510 ;
      LAYER li1 ;
        RECT 2184.495 214.490 2184.825 215.290 ;
      LAYER li1 ;
        RECT 2184.995 214.660 2185.165 215.510 ;
      LAYER li1 ;
        RECT 2185.335 214.490 2185.665 215.290 ;
      LAYER li1 ;
        RECT 2185.835 214.660 2186.005 215.510 ;
      LAYER li1 ;
        RECT 2186.255 214.490 2186.425 215.290 ;
        RECT 2186.595 214.660 2186.925 215.510 ;
        RECT 2187.095 214.490 2187.265 215.290 ;
        RECT 2187.435 214.660 2187.765 215.510 ;
        RECT 2187.945 214.490 2188.235 215.655 ;
        RECT 2188.795 214.490 2189.125 215.640 ;
      LAYER li1 ;
        RECT 2189.295 215.510 2191.985 215.680 ;
      LAYER li1 ;
        RECT 2192.245 215.510 2193.745 215.680 ;
      LAYER li1 ;
        RECT 2189.295 214.660 2189.465 215.510 ;
      LAYER li1 ;
        RECT 2189.635 214.490 2189.965 215.290 ;
      LAYER li1 ;
        RECT 2190.135 214.660 2190.305 215.510 ;
      LAYER li1 ;
        RECT 2190.475 214.490 2190.805 215.290 ;
      LAYER li1 ;
        RECT 2190.975 214.660 2191.145 215.510 ;
      LAYER li1 ;
        RECT 2191.315 214.490 2191.645 215.290 ;
      LAYER li1 ;
        RECT 2191.815 214.660 2191.985 215.510 ;
      LAYER li1 ;
        RECT 2192.235 214.490 2192.405 215.290 ;
        RECT 2192.575 214.660 2192.905 215.510 ;
        RECT 2193.075 214.490 2193.245 215.290 ;
        RECT 2193.415 214.660 2193.745 215.510 ;
        RECT 2193.925 214.490 2194.215 215.655 ;
        RECT 2194.775 214.490 2195.105 215.640 ;
      LAYER li1 ;
        RECT 2195.275 215.510 2197.965 215.680 ;
      LAYER li1 ;
        RECT 2198.225 215.510 2199.725 215.680 ;
      LAYER li1 ;
        RECT 2195.275 214.660 2195.445 215.510 ;
      LAYER li1 ;
        RECT 2195.615 214.490 2195.945 215.290 ;
      LAYER li1 ;
        RECT 2196.115 214.660 2196.285 215.510 ;
      LAYER li1 ;
        RECT 2196.455 214.490 2196.785 215.290 ;
      LAYER li1 ;
        RECT 2196.955 214.660 2197.125 215.510 ;
      LAYER li1 ;
        RECT 2197.295 214.490 2197.625 215.290 ;
      LAYER li1 ;
        RECT 2197.795 214.660 2197.965 215.510 ;
      LAYER li1 ;
        RECT 2198.215 214.490 2198.385 215.290 ;
        RECT 2198.555 214.660 2198.885 215.510 ;
        RECT 2199.055 214.490 2199.225 215.290 ;
        RECT 2199.395 214.660 2199.725 215.510 ;
        RECT 2199.905 214.490 2200.195 215.655 ;
      LAYER li1 ;
        RECT 2203.770 214.925 2204.120 216.175 ;
        RECT 2237.135 215.680 2237.390 216.220 ;
      LAYER li1 ;
        RECT 2240.085 216.050 2240.260 216.220 ;
        RECT 2237.635 215.880 2240.260 216.050 ;
        RECT 2240.085 215.680 2240.260 215.880 ;
      LAYER li1 ;
        RECT 2243.115 215.680 2243.370 216.220 ;
      LAYER li1 ;
        RECT 2246.065 216.050 2246.240 216.220 ;
        RECT 2243.615 215.880 2246.240 216.050 ;
        RECT 2246.065 215.680 2246.240 215.880 ;
      LAYER li1 ;
        RECT 2249.095 215.680 2249.350 216.220 ;
      LAYER li1 ;
        RECT 2252.045 216.050 2252.220 216.220 ;
        RECT 2249.595 215.880 2252.220 216.050 ;
        RECT 2252.045 215.680 2252.220 215.880 ;
      LAYER li1 ;
        RECT 2255.075 215.680 2255.330 216.220 ;
      LAYER li1 ;
        RECT 2258.025 216.050 2258.200 216.220 ;
        RECT 2255.575 215.880 2258.200 216.050 ;
        RECT 2258.025 215.680 2258.200 215.880 ;
      LAYER li1 ;
        RECT 2261.055 215.680 2261.310 216.220 ;
      LAYER li1 ;
        RECT 2264.005 216.050 2264.180 216.220 ;
        RECT 2261.555 215.880 2264.180 216.050 ;
        RECT 2264.005 215.680 2264.180 215.880 ;
      LAYER li1 ;
        RECT 2267.035 215.680 2267.290 216.220 ;
      LAYER li1 ;
        RECT 2269.985 216.050 2270.160 216.220 ;
        RECT 2267.535 215.880 2270.160 216.050 ;
        RECT 2269.985 215.680 2270.160 215.880 ;
      LAYER li1 ;
        RECT 2200.365 214.490 2205.710 214.925 ;
      LAYER li1 ;
        RECT 2205.885 214.490 2206.175 215.655 ;
        RECT 2235.785 214.490 2236.075 215.655 ;
        RECT 2236.635 214.490 2236.965 215.640 ;
      LAYER li1 ;
        RECT 2237.135 215.510 2239.825 215.680 ;
      LAYER li1 ;
        RECT 2240.085 215.510 2241.585 215.680 ;
      LAYER li1 ;
        RECT 2237.135 214.660 2237.305 215.510 ;
      LAYER li1 ;
        RECT 2237.475 214.490 2237.805 215.290 ;
      LAYER li1 ;
        RECT 2237.975 214.660 2238.145 215.510 ;
      LAYER li1 ;
        RECT 2238.315 214.490 2238.645 215.290 ;
      LAYER li1 ;
        RECT 2238.815 214.660 2238.985 215.510 ;
      LAYER li1 ;
        RECT 2239.155 214.490 2239.485 215.290 ;
      LAYER li1 ;
        RECT 2239.655 214.660 2239.825 215.510 ;
      LAYER li1 ;
        RECT 2240.075 214.490 2240.245 215.290 ;
        RECT 2240.415 214.660 2240.745 215.510 ;
        RECT 2240.915 214.490 2241.085 215.290 ;
        RECT 2241.255 214.660 2241.585 215.510 ;
        RECT 2241.765 214.490 2242.055 215.655 ;
        RECT 2242.615 214.490 2242.945 215.640 ;
      LAYER li1 ;
        RECT 2243.115 215.510 2245.805 215.680 ;
      LAYER li1 ;
        RECT 2246.065 215.510 2247.565 215.680 ;
      LAYER li1 ;
        RECT 2243.115 214.660 2243.285 215.510 ;
      LAYER li1 ;
        RECT 2243.455 214.490 2243.785 215.290 ;
      LAYER li1 ;
        RECT 2243.955 214.660 2244.125 215.510 ;
      LAYER li1 ;
        RECT 2244.295 214.490 2244.625 215.290 ;
      LAYER li1 ;
        RECT 2244.795 214.660 2244.965 215.510 ;
      LAYER li1 ;
        RECT 2245.135 214.490 2245.465 215.290 ;
      LAYER li1 ;
        RECT 2245.635 214.660 2245.805 215.510 ;
      LAYER li1 ;
        RECT 2246.055 214.490 2246.225 215.290 ;
        RECT 2246.395 214.660 2246.725 215.510 ;
        RECT 2246.895 214.490 2247.065 215.290 ;
        RECT 2247.235 214.660 2247.565 215.510 ;
        RECT 2247.745 214.490 2248.035 215.655 ;
        RECT 2248.595 214.490 2248.925 215.640 ;
      LAYER li1 ;
        RECT 2249.095 215.510 2251.785 215.680 ;
      LAYER li1 ;
        RECT 2252.045 215.510 2253.545 215.680 ;
      LAYER li1 ;
        RECT 2249.095 214.660 2249.265 215.510 ;
      LAYER li1 ;
        RECT 2249.435 214.490 2249.765 215.290 ;
      LAYER li1 ;
        RECT 2249.935 214.660 2250.105 215.510 ;
      LAYER li1 ;
        RECT 2250.275 214.490 2250.605 215.290 ;
      LAYER li1 ;
        RECT 2250.775 214.660 2250.945 215.510 ;
      LAYER li1 ;
        RECT 2251.115 214.490 2251.445 215.290 ;
      LAYER li1 ;
        RECT 2251.615 214.660 2251.785 215.510 ;
      LAYER li1 ;
        RECT 2252.035 214.490 2252.205 215.290 ;
        RECT 2252.375 214.660 2252.705 215.510 ;
        RECT 2252.875 214.490 2253.045 215.290 ;
        RECT 2253.215 214.660 2253.545 215.510 ;
        RECT 2253.725 214.490 2254.015 215.655 ;
        RECT 2254.575 214.490 2254.905 215.640 ;
      LAYER li1 ;
        RECT 2255.075 215.510 2257.765 215.680 ;
      LAYER li1 ;
        RECT 2258.025 215.510 2259.525 215.680 ;
      LAYER li1 ;
        RECT 2255.075 214.660 2255.245 215.510 ;
      LAYER li1 ;
        RECT 2255.415 214.490 2255.745 215.290 ;
      LAYER li1 ;
        RECT 2255.915 214.660 2256.085 215.510 ;
      LAYER li1 ;
        RECT 2256.255 214.490 2256.585 215.290 ;
      LAYER li1 ;
        RECT 2256.755 214.660 2256.925 215.510 ;
      LAYER li1 ;
        RECT 2257.095 214.490 2257.425 215.290 ;
      LAYER li1 ;
        RECT 2257.595 214.660 2257.765 215.510 ;
      LAYER li1 ;
        RECT 2258.015 214.490 2258.185 215.290 ;
        RECT 2258.355 214.660 2258.685 215.510 ;
        RECT 2258.855 214.490 2259.025 215.290 ;
        RECT 2259.195 214.660 2259.525 215.510 ;
        RECT 2259.705 214.490 2259.995 215.655 ;
        RECT 2260.555 214.490 2260.885 215.640 ;
      LAYER li1 ;
        RECT 2261.055 215.510 2263.745 215.680 ;
      LAYER li1 ;
        RECT 2264.005 215.510 2265.505 215.680 ;
      LAYER li1 ;
        RECT 2261.055 214.660 2261.225 215.510 ;
      LAYER li1 ;
        RECT 2261.395 214.490 2261.725 215.290 ;
      LAYER li1 ;
        RECT 2261.895 214.660 2262.065 215.510 ;
      LAYER li1 ;
        RECT 2262.235 214.490 2262.565 215.290 ;
      LAYER li1 ;
        RECT 2262.735 214.660 2262.905 215.510 ;
      LAYER li1 ;
        RECT 2263.075 214.490 2263.405 215.290 ;
      LAYER li1 ;
        RECT 2263.575 214.660 2263.745 215.510 ;
      LAYER li1 ;
        RECT 2263.995 214.490 2264.165 215.290 ;
        RECT 2264.335 214.660 2264.665 215.510 ;
        RECT 2264.835 214.490 2265.005 215.290 ;
        RECT 2265.175 214.660 2265.505 215.510 ;
        RECT 2265.685 214.490 2265.975 215.655 ;
        RECT 2266.535 214.490 2266.865 215.640 ;
      LAYER li1 ;
        RECT 2267.035 215.510 2269.725 215.680 ;
      LAYER li1 ;
        RECT 2269.985 215.510 2271.485 215.680 ;
      LAYER li1 ;
        RECT 2267.035 214.660 2267.205 215.510 ;
      LAYER li1 ;
        RECT 2267.375 214.490 2267.705 215.290 ;
      LAYER li1 ;
        RECT 2267.875 214.660 2268.045 215.510 ;
      LAYER li1 ;
        RECT 2268.215 214.490 2268.545 215.290 ;
      LAYER li1 ;
        RECT 2268.715 214.660 2268.885 215.510 ;
      LAYER li1 ;
        RECT 2269.055 214.490 2269.385 215.290 ;
      LAYER li1 ;
        RECT 2269.555 214.660 2269.725 215.510 ;
      LAYER li1 ;
        RECT 2269.975 214.490 2270.145 215.290 ;
        RECT 2270.315 214.660 2270.645 215.510 ;
        RECT 2270.815 214.490 2270.985 215.290 ;
        RECT 2271.155 214.660 2271.485 215.510 ;
        RECT 2271.665 214.490 2271.955 215.655 ;
        RECT 669.000 214.320 669.145 214.490 ;
        RECT 669.315 214.320 669.605 214.490 ;
        RECT 669.775 214.320 670.065 214.490 ;
        RECT 670.235 214.320 670.525 214.490 ;
        RECT 670.695 214.320 670.985 214.490 ;
        RECT 671.155 214.320 671.445 214.490 ;
        RECT 671.615 214.320 671.905 214.490 ;
        RECT 672.075 214.320 672.365 214.490 ;
        RECT 672.535 214.320 672.825 214.490 ;
        RECT 672.995 214.320 673.285 214.490 ;
        RECT 673.455 214.320 673.745 214.490 ;
        RECT 673.915 214.320 674.205 214.490 ;
        RECT 674.375 214.320 674.665 214.490 ;
        RECT 674.835 214.320 675.125 214.490 ;
        RECT 675.295 214.320 675.585 214.490 ;
        RECT 675.755 214.320 676.045 214.490 ;
        RECT 676.215 214.320 676.505 214.490 ;
        RECT 676.675 214.320 676.965 214.490 ;
        RECT 677.135 214.320 677.425 214.490 ;
        RECT 677.595 214.320 677.885 214.490 ;
        RECT 678.055 214.320 678.345 214.490 ;
        RECT 678.515 214.320 678.805 214.490 ;
        RECT 678.975 214.320 679.265 214.490 ;
        RECT 679.435 214.320 679.725 214.490 ;
        RECT 679.895 214.320 680.185 214.490 ;
        RECT 680.355 214.320 680.645 214.490 ;
        RECT 680.815 214.320 681.105 214.490 ;
        RECT 681.275 214.320 681.565 214.490 ;
        RECT 681.735 214.320 682.025 214.490 ;
        RECT 682.195 214.320 682.485 214.490 ;
        RECT 682.655 214.320 682.945 214.490 ;
        RECT 683.115 214.320 683.405 214.490 ;
        RECT 683.575 214.320 683.865 214.490 ;
        RECT 684.035 214.320 684.325 214.490 ;
        RECT 684.495 214.320 684.785 214.490 ;
        RECT 684.955 214.320 685.245 214.490 ;
        RECT 685.415 214.320 685.705 214.490 ;
        RECT 685.875 214.320 686.165 214.490 ;
        RECT 686.335 214.320 686.625 214.490 ;
        RECT 686.795 214.320 687.085 214.490 ;
        RECT 687.255 214.320 687.545 214.490 ;
        RECT 687.715 214.320 688.005 214.490 ;
        RECT 688.175 214.320 688.465 214.490 ;
        RECT 688.635 214.320 688.925 214.490 ;
        RECT 689.095 214.320 689.385 214.490 ;
        RECT 689.555 214.320 689.845 214.490 ;
        RECT 690.015 214.320 690.305 214.490 ;
        RECT 690.475 214.320 690.765 214.490 ;
        RECT 690.935 214.320 691.225 214.490 ;
        RECT 691.395 214.320 691.685 214.490 ;
        RECT 691.855 214.320 692.145 214.490 ;
        RECT 692.315 214.320 692.605 214.490 ;
        RECT 692.775 214.320 693.065 214.490 ;
        RECT 693.235 214.320 693.525 214.490 ;
        RECT 693.695 214.320 693.985 214.490 ;
        RECT 694.155 214.320 694.445 214.490 ;
        RECT 694.615 214.320 694.905 214.490 ;
        RECT 695.075 214.320 695.365 214.490 ;
        RECT 695.535 214.320 695.825 214.490 ;
        RECT 695.995 214.320 696.285 214.490 ;
        RECT 696.455 214.320 696.745 214.490 ;
        RECT 696.915 214.320 697.205 214.490 ;
        RECT 697.375 214.320 697.665 214.490 ;
        RECT 697.835 214.320 698.125 214.490 ;
        RECT 698.295 214.320 698.585 214.490 ;
        RECT 698.755 214.320 699.045 214.490 ;
        RECT 699.215 214.320 699.505 214.490 ;
        RECT 699.675 214.320 699.965 214.490 ;
        RECT 700.135 214.320 700.425 214.490 ;
        RECT 700.595 214.320 700.885 214.490 ;
        RECT 701.055 214.320 701.345 214.490 ;
        RECT 701.515 214.320 701.805 214.490 ;
        RECT 701.975 214.320 702.265 214.490 ;
        RECT 702.435 214.320 702.725 214.490 ;
        RECT 702.895 214.320 703.185 214.490 ;
        RECT 703.355 214.320 703.645 214.490 ;
        RECT 703.815 214.320 704.105 214.490 ;
        RECT 704.275 214.320 704.565 214.490 ;
        RECT 704.735 214.320 705.025 214.490 ;
        RECT 705.195 214.320 705.485 214.490 ;
        RECT 705.655 214.320 705.945 214.490 ;
        RECT 706.115 214.320 706.405 214.490 ;
        RECT 706.575 214.320 706.865 214.490 ;
        RECT 707.035 214.320 707.325 214.490 ;
        RECT 707.495 214.320 707.785 214.490 ;
        RECT 707.955 214.320 708.245 214.490 ;
        RECT 708.415 214.320 708.705 214.490 ;
        RECT 708.875 214.320 709.165 214.490 ;
        RECT 709.335 214.320 709.625 214.490 ;
        RECT 709.795 214.320 710.085 214.490 ;
        RECT 710.255 214.320 710.545 214.490 ;
        RECT 710.715 214.320 711.005 214.490 ;
        RECT 711.175 214.320 711.465 214.490 ;
        RECT 711.635 214.320 711.925 214.490 ;
        RECT 712.095 214.320 712.385 214.490 ;
        RECT 712.555 214.320 712.845 214.490 ;
        RECT 713.015 214.320 713.305 214.490 ;
        RECT 713.475 214.320 713.765 214.490 ;
        RECT 713.935 214.320 714.225 214.490 ;
        RECT 714.395 214.320 714.685 214.490 ;
        RECT 714.855 214.320 715.145 214.490 ;
        RECT 715.315 214.320 715.605 214.490 ;
        RECT 715.775 214.320 716.065 214.490 ;
        RECT 716.235 214.320 716.525 214.490 ;
        RECT 716.695 214.320 716.985 214.490 ;
        RECT 717.155 214.320 717.445 214.490 ;
        RECT 717.615 214.320 717.905 214.490 ;
        RECT 718.075 214.320 718.365 214.490 ;
        RECT 718.535 214.320 718.825 214.490 ;
        RECT 718.995 214.320 719.285 214.490 ;
        RECT 719.455 214.320 719.745 214.490 ;
        RECT 719.915 214.320 720.205 214.490 ;
        RECT 720.375 214.320 720.665 214.490 ;
        RECT 720.835 214.320 721.125 214.490 ;
        RECT 721.295 214.320 721.585 214.490 ;
        RECT 721.755 214.320 722.045 214.490 ;
        RECT 722.215 214.320 722.505 214.490 ;
        RECT 722.675 214.320 722.965 214.490 ;
        RECT 723.135 214.320 723.425 214.490 ;
        RECT 723.595 214.320 723.885 214.490 ;
        RECT 724.055 214.320 724.345 214.490 ;
        RECT 724.515 214.320 724.805 214.490 ;
        RECT 724.975 214.320 725.265 214.490 ;
        RECT 725.435 214.320 725.725 214.490 ;
        RECT 725.895 214.320 726.185 214.490 ;
        RECT 726.355 214.320 726.645 214.490 ;
        RECT 726.815 214.320 727.105 214.490 ;
        RECT 727.275 214.320 727.565 214.490 ;
        RECT 727.735 214.320 728.025 214.490 ;
        RECT 728.195 214.320 728.485 214.490 ;
        RECT 728.655 214.320 728.945 214.490 ;
        RECT 729.115 214.320 729.260 214.490 ;
        RECT 758.700 214.320 758.845 214.490 ;
        RECT 759.015 214.320 759.305 214.490 ;
        RECT 759.475 214.320 759.765 214.490 ;
        RECT 759.935 214.320 760.225 214.490 ;
        RECT 760.395 214.320 760.685 214.490 ;
        RECT 760.855 214.320 761.145 214.490 ;
        RECT 761.315 214.320 761.605 214.490 ;
        RECT 761.775 214.320 762.065 214.490 ;
        RECT 762.235 214.320 762.525 214.490 ;
        RECT 762.695 214.320 762.985 214.490 ;
        RECT 763.155 214.320 763.445 214.490 ;
        RECT 763.615 214.320 763.905 214.490 ;
        RECT 764.075 214.320 764.365 214.490 ;
        RECT 764.535 214.320 764.825 214.490 ;
        RECT 764.995 214.320 765.285 214.490 ;
        RECT 765.455 214.320 765.745 214.490 ;
        RECT 765.915 214.320 766.205 214.490 ;
        RECT 766.375 214.320 766.665 214.490 ;
        RECT 766.835 214.320 767.125 214.490 ;
        RECT 767.295 214.320 767.585 214.490 ;
        RECT 767.755 214.320 768.045 214.490 ;
        RECT 768.215 214.320 768.505 214.490 ;
        RECT 768.675 214.320 768.965 214.490 ;
        RECT 769.135 214.320 769.425 214.490 ;
        RECT 769.595 214.320 769.885 214.490 ;
        RECT 770.055 214.320 770.345 214.490 ;
        RECT 770.515 214.320 770.805 214.490 ;
        RECT 770.975 214.320 771.265 214.490 ;
        RECT 771.435 214.320 771.725 214.490 ;
        RECT 771.895 214.320 772.185 214.490 ;
        RECT 772.355 214.320 772.645 214.490 ;
        RECT 772.815 214.320 773.105 214.490 ;
        RECT 773.275 214.320 773.565 214.490 ;
        RECT 773.735 214.320 774.025 214.490 ;
        RECT 774.195 214.320 774.485 214.490 ;
        RECT 774.655 214.320 774.945 214.490 ;
        RECT 775.115 214.320 775.405 214.490 ;
        RECT 775.575 214.320 775.865 214.490 ;
        RECT 776.035 214.320 776.325 214.490 ;
        RECT 776.495 214.320 776.785 214.490 ;
        RECT 776.955 214.320 777.245 214.490 ;
        RECT 777.415 214.320 777.705 214.490 ;
        RECT 777.875 214.320 778.165 214.490 ;
        RECT 778.335 214.320 778.625 214.490 ;
        RECT 778.795 214.320 779.085 214.490 ;
        RECT 779.255 214.320 779.545 214.490 ;
        RECT 779.715 214.320 780.005 214.490 ;
        RECT 780.175 214.320 780.465 214.490 ;
        RECT 780.635 214.320 780.925 214.490 ;
        RECT 781.095 214.320 781.385 214.490 ;
        RECT 781.555 214.320 781.845 214.490 ;
        RECT 782.015 214.320 782.305 214.490 ;
        RECT 782.475 214.320 782.765 214.490 ;
        RECT 782.935 214.320 783.225 214.490 ;
        RECT 783.395 214.320 783.685 214.490 ;
        RECT 783.855 214.320 784.145 214.490 ;
        RECT 784.315 214.320 784.605 214.490 ;
        RECT 784.775 214.320 785.065 214.490 ;
        RECT 785.235 214.320 785.525 214.490 ;
        RECT 785.695 214.320 785.985 214.490 ;
        RECT 786.155 214.320 786.445 214.490 ;
        RECT 786.615 214.320 786.905 214.490 ;
        RECT 787.075 214.320 787.365 214.490 ;
        RECT 787.535 214.320 787.825 214.490 ;
        RECT 787.995 214.320 788.285 214.490 ;
        RECT 788.455 214.320 788.745 214.490 ;
        RECT 788.915 214.320 789.205 214.490 ;
        RECT 789.375 214.320 789.665 214.490 ;
        RECT 789.835 214.320 790.125 214.490 ;
        RECT 790.295 214.320 790.585 214.490 ;
        RECT 790.755 214.320 791.045 214.490 ;
        RECT 791.215 214.320 791.505 214.490 ;
        RECT 791.675 214.320 791.965 214.490 ;
        RECT 792.135 214.320 792.425 214.490 ;
        RECT 792.595 214.320 792.885 214.490 ;
        RECT 793.055 214.320 793.345 214.490 ;
        RECT 793.515 214.320 793.805 214.490 ;
        RECT 793.975 214.320 794.265 214.490 ;
        RECT 794.435 214.320 794.725 214.490 ;
        RECT 794.895 214.320 795.040 214.490 ;
        RECT 2146.000 214.320 2146.145 214.490 ;
        RECT 2146.315 214.320 2146.605 214.490 ;
        RECT 2146.775 214.320 2147.065 214.490 ;
        RECT 2147.235 214.320 2147.525 214.490 ;
        RECT 2147.695 214.320 2147.985 214.490 ;
        RECT 2148.155 214.320 2148.445 214.490 ;
        RECT 2148.615 214.320 2148.905 214.490 ;
        RECT 2149.075 214.320 2149.365 214.490 ;
        RECT 2149.535 214.320 2149.825 214.490 ;
        RECT 2149.995 214.320 2150.285 214.490 ;
        RECT 2150.455 214.320 2150.745 214.490 ;
        RECT 2150.915 214.320 2151.205 214.490 ;
        RECT 2151.375 214.320 2151.665 214.490 ;
        RECT 2151.835 214.320 2152.125 214.490 ;
        RECT 2152.295 214.320 2152.585 214.490 ;
        RECT 2152.755 214.320 2153.045 214.490 ;
        RECT 2153.215 214.320 2153.505 214.490 ;
        RECT 2153.675 214.320 2153.965 214.490 ;
        RECT 2154.135 214.320 2154.425 214.490 ;
        RECT 2154.595 214.320 2154.885 214.490 ;
        RECT 2155.055 214.320 2155.345 214.490 ;
        RECT 2155.515 214.320 2155.805 214.490 ;
        RECT 2155.975 214.320 2156.265 214.490 ;
        RECT 2156.435 214.320 2156.725 214.490 ;
        RECT 2156.895 214.320 2157.185 214.490 ;
        RECT 2157.355 214.320 2157.645 214.490 ;
        RECT 2157.815 214.320 2158.105 214.490 ;
        RECT 2158.275 214.320 2158.565 214.490 ;
        RECT 2158.735 214.320 2159.025 214.490 ;
        RECT 2159.195 214.320 2159.485 214.490 ;
        RECT 2159.655 214.320 2159.945 214.490 ;
        RECT 2160.115 214.320 2160.405 214.490 ;
        RECT 2160.575 214.320 2160.865 214.490 ;
        RECT 2161.035 214.320 2161.325 214.490 ;
        RECT 2161.495 214.320 2161.785 214.490 ;
        RECT 2161.955 214.320 2162.245 214.490 ;
        RECT 2162.415 214.320 2162.705 214.490 ;
        RECT 2162.875 214.320 2163.165 214.490 ;
        RECT 2163.335 214.320 2163.625 214.490 ;
        RECT 2163.795 214.320 2164.085 214.490 ;
        RECT 2164.255 214.320 2164.545 214.490 ;
        RECT 2164.715 214.320 2165.005 214.490 ;
        RECT 2165.175 214.320 2165.465 214.490 ;
        RECT 2165.635 214.320 2165.925 214.490 ;
        RECT 2166.095 214.320 2166.385 214.490 ;
        RECT 2166.555 214.320 2166.845 214.490 ;
        RECT 2167.015 214.320 2167.305 214.490 ;
        RECT 2167.475 214.320 2167.765 214.490 ;
        RECT 2167.935 214.320 2168.225 214.490 ;
        RECT 2168.395 214.320 2168.685 214.490 ;
        RECT 2168.855 214.320 2169.145 214.490 ;
        RECT 2169.315 214.320 2169.605 214.490 ;
        RECT 2169.775 214.320 2170.065 214.490 ;
        RECT 2170.235 214.320 2170.525 214.490 ;
        RECT 2170.695 214.320 2170.985 214.490 ;
        RECT 2171.155 214.320 2171.445 214.490 ;
        RECT 2171.615 214.320 2171.905 214.490 ;
        RECT 2172.075 214.320 2172.365 214.490 ;
        RECT 2172.535 214.320 2172.825 214.490 ;
        RECT 2172.995 214.320 2173.285 214.490 ;
        RECT 2173.455 214.320 2173.745 214.490 ;
        RECT 2173.915 214.320 2174.205 214.490 ;
        RECT 2174.375 214.320 2174.665 214.490 ;
        RECT 2174.835 214.320 2175.125 214.490 ;
        RECT 2175.295 214.320 2175.585 214.490 ;
        RECT 2175.755 214.320 2176.045 214.490 ;
        RECT 2176.215 214.320 2176.505 214.490 ;
        RECT 2176.675 214.320 2176.965 214.490 ;
        RECT 2177.135 214.320 2177.425 214.490 ;
        RECT 2177.595 214.320 2177.885 214.490 ;
        RECT 2178.055 214.320 2178.345 214.490 ;
        RECT 2178.515 214.320 2178.805 214.490 ;
        RECT 2178.975 214.320 2179.265 214.490 ;
        RECT 2179.435 214.320 2179.725 214.490 ;
        RECT 2179.895 214.320 2180.185 214.490 ;
        RECT 2180.355 214.320 2180.645 214.490 ;
        RECT 2180.815 214.320 2181.105 214.490 ;
        RECT 2181.275 214.320 2181.565 214.490 ;
        RECT 2181.735 214.320 2182.025 214.490 ;
        RECT 2182.195 214.320 2182.485 214.490 ;
        RECT 2182.655 214.320 2182.945 214.490 ;
        RECT 2183.115 214.320 2183.405 214.490 ;
        RECT 2183.575 214.320 2183.865 214.490 ;
        RECT 2184.035 214.320 2184.325 214.490 ;
        RECT 2184.495 214.320 2184.785 214.490 ;
        RECT 2184.955 214.320 2185.245 214.490 ;
        RECT 2185.415 214.320 2185.705 214.490 ;
        RECT 2185.875 214.320 2186.165 214.490 ;
        RECT 2186.335 214.320 2186.625 214.490 ;
        RECT 2186.795 214.320 2187.085 214.490 ;
        RECT 2187.255 214.320 2187.545 214.490 ;
        RECT 2187.715 214.320 2188.005 214.490 ;
        RECT 2188.175 214.320 2188.465 214.490 ;
        RECT 2188.635 214.320 2188.925 214.490 ;
        RECT 2189.095 214.320 2189.385 214.490 ;
        RECT 2189.555 214.320 2189.845 214.490 ;
        RECT 2190.015 214.320 2190.305 214.490 ;
        RECT 2190.475 214.320 2190.765 214.490 ;
        RECT 2190.935 214.320 2191.225 214.490 ;
        RECT 2191.395 214.320 2191.685 214.490 ;
        RECT 2191.855 214.320 2192.145 214.490 ;
        RECT 2192.315 214.320 2192.605 214.490 ;
        RECT 2192.775 214.320 2193.065 214.490 ;
        RECT 2193.235 214.320 2193.525 214.490 ;
        RECT 2193.695 214.320 2193.985 214.490 ;
        RECT 2194.155 214.320 2194.445 214.490 ;
        RECT 2194.615 214.320 2194.905 214.490 ;
        RECT 2195.075 214.320 2195.365 214.490 ;
        RECT 2195.535 214.320 2195.825 214.490 ;
        RECT 2195.995 214.320 2196.285 214.490 ;
        RECT 2196.455 214.320 2196.745 214.490 ;
        RECT 2196.915 214.320 2197.205 214.490 ;
        RECT 2197.375 214.320 2197.665 214.490 ;
        RECT 2197.835 214.320 2198.125 214.490 ;
        RECT 2198.295 214.320 2198.585 214.490 ;
        RECT 2198.755 214.320 2199.045 214.490 ;
        RECT 2199.215 214.320 2199.505 214.490 ;
        RECT 2199.675 214.320 2199.965 214.490 ;
        RECT 2200.135 214.320 2200.425 214.490 ;
        RECT 2200.595 214.320 2200.885 214.490 ;
        RECT 2201.055 214.320 2201.345 214.490 ;
        RECT 2201.515 214.320 2201.805 214.490 ;
        RECT 2201.975 214.320 2202.265 214.490 ;
        RECT 2202.435 214.320 2202.725 214.490 ;
        RECT 2202.895 214.320 2203.185 214.490 ;
        RECT 2203.355 214.320 2203.645 214.490 ;
        RECT 2203.815 214.320 2204.105 214.490 ;
        RECT 2204.275 214.320 2204.565 214.490 ;
        RECT 2204.735 214.320 2205.025 214.490 ;
        RECT 2205.195 214.320 2205.485 214.490 ;
        RECT 2205.655 214.320 2205.945 214.490 ;
        RECT 2206.115 214.320 2206.260 214.490 ;
        RECT 2235.700 214.320 2235.845 214.490 ;
        RECT 2236.015 214.320 2236.305 214.490 ;
        RECT 2236.475 214.320 2236.765 214.490 ;
        RECT 2236.935 214.320 2237.225 214.490 ;
        RECT 2237.395 214.320 2237.685 214.490 ;
        RECT 2237.855 214.320 2238.145 214.490 ;
        RECT 2238.315 214.320 2238.605 214.490 ;
        RECT 2238.775 214.320 2239.065 214.490 ;
        RECT 2239.235 214.320 2239.525 214.490 ;
        RECT 2239.695 214.320 2239.985 214.490 ;
        RECT 2240.155 214.320 2240.445 214.490 ;
        RECT 2240.615 214.320 2240.905 214.490 ;
        RECT 2241.075 214.320 2241.365 214.490 ;
        RECT 2241.535 214.320 2241.825 214.490 ;
        RECT 2241.995 214.320 2242.285 214.490 ;
        RECT 2242.455 214.320 2242.745 214.490 ;
        RECT 2242.915 214.320 2243.205 214.490 ;
        RECT 2243.375 214.320 2243.665 214.490 ;
        RECT 2243.835 214.320 2244.125 214.490 ;
        RECT 2244.295 214.320 2244.585 214.490 ;
        RECT 2244.755 214.320 2245.045 214.490 ;
        RECT 2245.215 214.320 2245.505 214.490 ;
        RECT 2245.675 214.320 2245.965 214.490 ;
        RECT 2246.135 214.320 2246.425 214.490 ;
        RECT 2246.595 214.320 2246.885 214.490 ;
        RECT 2247.055 214.320 2247.345 214.490 ;
        RECT 2247.515 214.320 2247.805 214.490 ;
        RECT 2247.975 214.320 2248.265 214.490 ;
        RECT 2248.435 214.320 2248.725 214.490 ;
        RECT 2248.895 214.320 2249.185 214.490 ;
        RECT 2249.355 214.320 2249.645 214.490 ;
        RECT 2249.815 214.320 2250.105 214.490 ;
        RECT 2250.275 214.320 2250.565 214.490 ;
        RECT 2250.735 214.320 2251.025 214.490 ;
        RECT 2251.195 214.320 2251.485 214.490 ;
        RECT 2251.655 214.320 2251.945 214.490 ;
        RECT 2252.115 214.320 2252.405 214.490 ;
        RECT 2252.575 214.320 2252.865 214.490 ;
        RECT 2253.035 214.320 2253.325 214.490 ;
        RECT 2253.495 214.320 2253.785 214.490 ;
        RECT 2253.955 214.320 2254.245 214.490 ;
        RECT 2254.415 214.320 2254.705 214.490 ;
        RECT 2254.875 214.320 2255.165 214.490 ;
        RECT 2255.335 214.320 2255.625 214.490 ;
        RECT 2255.795 214.320 2256.085 214.490 ;
        RECT 2256.255 214.320 2256.545 214.490 ;
        RECT 2256.715 214.320 2257.005 214.490 ;
        RECT 2257.175 214.320 2257.465 214.490 ;
        RECT 2257.635 214.320 2257.925 214.490 ;
        RECT 2258.095 214.320 2258.385 214.490 ;
        RECT 2258.555 214.320 2258.845 214.490 ;
        RECT 2259.015 214.320 2259.305 214.490 ;
        RECT 2259.475 214.320 2259.765 214.490 ;
        RECT 2259.935 214.320 2260.225 214.490 ;
        RECT 2260.395 214.320 2260.685 214.490 ;
        RECT 2260.855 214.320 2261.145 214.490 ;
        RECT 2261.315 214.320 2261.605 214.490 ;
        RECT 2261.775 214.320 2262.065 214.490 ;
        RECT 2262.235 214.320 2262.525 214.490 ;
        RECT 2262.695 214.320 2262.985 214.490 ;
        RECT 2263.155 214.320 2263.445 214.490 ;
        RECT 2263.615 214.320 2263.905 214.490 ;
        RECT 2264.075 214.320 2264.365 214.490 ;
        RECT 2264.535 214.320 2264.825 214.490 ;
        RECT 2264.995 214.320 2265.285 214.490 ;
        RECT 2265.455 214.320 2265.745 214.490 ;
        RECT 2265.915 214.320 2266.205 214.490 ;
        RECT 2266.375 214.320 2266.665 214.490 ;
        RECT 2266.835 214.320 2267.125 214.490 ;
        RECT 2267.295 214.320 2267.585 214.490 ;
        RECT 2267.755 214.320 2268.045 214.490 ;
        RECT 2268.215 214.320 2268.505 214.490 ;
        RECT 2268.675 214.320 2268.965 214.490 ;
        RECT 2269.135 214.320 2269.425 214.490 ;
        RECT 2269.595 214.320 2269.885 214.490 ;
        RECT 2270.055 214.320 2270.345 214.490 ;
        RECT 2270.515 214.320 2270.805 214.490 ;
        RECT 2270.975 214.320 2271.265 214.490 ;
        RECT 2271.435 214.320 2271.725 214.490 ;
        RECT 2271.895 214.320 2272.040 214.490 ;
        RECT 669.085 213.155 669.375 214.320 ;
      LAYER li1 ;
        RECT 669.545 213.885 674.890 214.320 ;
        RECT 672.950 212.635 673.300 213.885 ;
      LAYER li1 ;
        RECT 675.065 213.155 675.355 214.320 ;
        RECT 675.535 213.300 675.865 214.150 ;
        RECT 676.035 213.520 676.205 214.320 ;
        RECT 676.375 213.300 676.705 214.150 ;
        RECT 676.875 213.520 677.045 214.320 ;
      LAYER li1 ;
        RECT 677.295 213.300 677.465 214.150 ;
      LAYER li1 ;
        RECT 677.635 213.520 677.965 214.320 ;
      LAYER li1 ;
        RECT 678.135 213.300 678.305 214.150 ;
      LAYER li1 ;
        RECT 678.475 213.520 678.805 214.320 ;
      LAYER li1 ;
        RECT 678.975 213.300 679.145 214.150 ;
      LAYER li1 ;
        RECT 679.315 213.520 679.645 214.320 ;
      LAYER li1 ;
        RECT 679.815 213.300 679.985 214.150 ;
      LAYER li1 ;
        RECT 675.535 213.130 677.035 213.300 ;
      LAYER li1 ;
        RECT 677.295 213.130 679.985 213.300 ;
      LAYER li1 ;
        RECT 680.155 213.170 680.485 214.320 ;
        RECT 681.045 213.155 681.335 214.320 ;
        RECT 681.515 213.300 681.845 214.150 ;
        RECT 682.015 213.520 682.185 214.320 ;
        RECT 682.355 213.300 682.685 214.150 ;
        RECT 682.855 213.520 683.025 214.320 ;
      LAYER li1 ;
        RECT 683.275 213.300 683.445 214.150 ;
      LAYER li1 ;
        RECT 683.615 213.520 683.945 214.320 ;
      LAYER li1 ;
        RECT 684.115 213.300 684.285 214.150 ;
      LAYER li1 ;
        RECT 684.455 213.520 684.785 214.320 ;
      LAYER li1 ;
        RECT 684.955 213.300 685.125 214.150 ;
      LAYER li1 ;
        RECT 685.295 213.520 685.625 214.320 ;
      LAYER li1 ;
        RECT 685.795 213.300 685.965 214.150 ;
      LAYER li1 ;
        RECT 681.515 213.130 683.015 213.300 ;
      LAYER li1 ;
        RECT 683.275 213.130 685.965 213.300 ;
      LAYER li1 ;
        RECT 686.135 213.170 686.465 214.320 ;
        RECT 687.025 213.155 687.315 214.320 ;
        RECT 687.495 213.300 687.825 214.150 ;
        RECT 687.995 213.520 688.165 214.320 ;
        RECT 688.335 213.300 688.665 214.150 ;
        RECT 688.835 213.520 689.005 214.320 ;
      LAYER li1 ;
        RECT 689.255 213.300 689.425 214.150 ;
      LAYER li1 ;
        RECT 689.595 213.520 689.925 214.320 ;
      LAYER li1 ;
        RECT 690.095 213.300 690.265 214.150 ;
      LAYER li1 ;
        RECT 690.435 213.520 690.765 214.320 ;
      LAYER li1 ;
        RECT 690.935 213.300 691.105 214.150 ;
      LAYER li1 ;
        RECT 691.275 213.520 691.605 214.320 ;
      LAYER li1 ;
        RECT 691.775 213.300 691.945 214.150 ;
      LAYER li1 ;
        RECT 687.495 213.130 688.995 213.300 ;
      LAYER li1 ;
        RECT 689.255 213.130 691.945 213.300 ;
      LAYER li1 ;
        RECT 692.115 213.170 692.445 214.320 ;
        RECT 693.005 213.155 693.295 214.320 ;
        RECT 693.475 213.300 693.805 214.150 ;
        RECT 693.975 213.520 694.145 214.320 ;
        RECT 694.315 213.300 694.645 214.150 ;
        RECT 694.815 213.520 694.985 214.320 ;
      LAYER li1 ;
        RECT 695.235 213.300 695.405 214.150 ;
      LAYER li1 ;
        RECT 695.575 213.520 695.905 214.320 ;
      LAYER li1 ;
        RECT 696.075 213.300 696.245 214.150 ;
      LAYER li1 ;
        RECT 696.415 213.520 696.745 214.320 ;
      LAYER li1 ;
        RECT 696.915 213.300 697.085 214.150 ;
      LAYER li1 ;
        RECT 697.255 213.520 697.585 214.320 ;
      LAYER li1 ;
        RECT 697.755 213.300 697.925 214.150 ;
      LAYER li1 ;
        RECT 693.475 213.130 694.975 213.300 ;
      LAYER li1 ;
        RECT 695.235 213.130 697.925 213.300 ;
      LAYER li1 ;
        RECT 698.095 213.170 698.425 214.320 ;
        RECT 698.985 213.155 699.275 214.320 ;
        RECT 699.455 213.300 699.785 214.150 ;
        RECT 699.955 213.520 700.125 214.320 ;
        RECT 700.295 213.300 700.625 214.150 ;
        RECT 700.795 213.520 700.965 214.320 ;
      LAYER li1 ;
        RECT 701.215 213.300 701.385 214.150 ;
      LAYER li1 ;
        RECT 701.555 213.520 701.885 214.320 ;
      LAYER li1 ;
        RECT 702.055 213.300 702.225 214.150 ;
      LAYER li1 ;
        RECT 702.395 213.520 702.725 214.320 ;
      LAYER li1 ;
        RECT 702.895 213.300 703.065 214.150 ;
      LAYER li1 ;
        RECT 703.235 213.520 703.565 214.320 ;
      LAYER li1 ;
        RECT 703.735 213.300 703.905 214.150 ;
      LAYER li1 ;
        RECT 699.455 213.130 700.955 213.300 ;
      LAYER li1 ;
        RECT 701.215 213.130 703.905 213.300 ;
      LAYER li1 ;
        RECT 704.075 213.170 704.405 214.320 ;
        RECT 704.965 213.155 705.255 214.320 ;
        RECT 705.435 213.300 705.765 214.150 ;
        RECT 705.935 213.520 706.105 214.320 ;
        RECT 706.275 213.300 706.605 214.150 ;
        RECT 706.775 213.520 706.945 214.320 ;
      LAYER li1 ;
        RECT 707.195 213.300 707.365 214.150 ;
      LAYER li1 ;
        RECT 707.535 213.520 707.865 214.320 ;
      LAYER li1 ;
        RECT 708.035 213.300 708.205 214.150 ;
      LAYER li1 ;
        RECT 708.375 213.520 708.705 214.320 ;
      LAYER li1 ;
        RECT 708.875 213.300 709.045 214.150 ;
      LAYER li1 ;
        RECT 709.215 213.520 709.545 214.320 ;
      LAYER li1 ;
        RECT 709.715 213.300 709.885 214.150 ;
      LAYER li1 ;
        RECT 705.435 213.130 706.935 213.300 ;
      LAYER li1 ;
        RECT 707.195 213.130 709.885 213.300 ;
      LAYER li1 ;
        RECT 710.055 213.170 710.385 214.320 ;
        RECT 710.945 213.155 711.235 214.320 ;
        RECT 711.415 213.300 711.745 214.150 ;
        RECT 711.915 213.520 712.085 214.320 ;
        RECT 712.255 213.300 712.585 214.150 ;
        RECT 712.755 213.520 712.925 214.320 ;
      LAYER li1 ;
        RECT 713.175 213.300 713.345 214.150 ;
      LAYER li1 ;
        RECT 713.515 213.520 713.845 214.320 ;
      LAYER li1 ;
        RECT 714.015 213.300 714.185 214.150 ;
      LAYER li1 ;
        RECT 714.355 213.520 714.685 214.320 ;
      LAYER li1 ;
        RECT 714.855 213.300 715.025 214.150 ;
      LAYER li1 ;
        RECT 715.195 213.520 715.525 214.320 ;
      LAYER li1 ;
        RECT 715.695 213.300 715.865 214.150 ;
      LAYER li1 ;
        RECT 711.415 213.130 712.915 213.300 ;
      LAYER li1 ;
        RECT 713.175 213.130 715.865 213.300 ;
      LAYER li1 ;
        RECT 716.035 213.170 716.365 214.320 ;
        RECT 716.925 213.155 717.215 214.320 ;
        RECT 717.395 213.300 717.725 214.150 ;
        RECT 717.895 213.520 718.065 214.320 ;
        RECT 718.235 213.300 718.565 214.150 ;
        RECT 718.735 213.520 718.905 214.320 ;
      LAYER li1 ;
        RECT 719.155 213.300 719.325 214.150 ;
      LAYER li1 ;
        RECT 719.495 213.520 719.825 214.320 ;
      LAYER li1 ;
        RECT 719.995 213.300 720.165 214.150 ;
      LAYER li1 ;
        RECT 720.335 213.520 720.665 214.320 ;
      LAYER li1 ;
        RECT 720.835 213.300 721.005 214.150 ;
      LAYER li1 ;
        RECT 721.175 213.520 721.505 214.320 ;
      LAYER li1 ;
        RECT 721.675 213.300 721.845 214.150 ;
      LAYER li1 ;
        RECT 717.395 213.130 718.895 213.300 ;
      LAYER li1 ;
        RECT 719.155 213.130 721.845 213.300 ;
      LAYER li1 ;
        RECT 722.015 213.170 722.345 214.320 ;
        RECT 722.905 213.155 723.195 214.320 ;
        RECT 723.375 213.300 723.705 214.150 ;
        RECT 723.875 213.520 724.045 214.320 ;
        RECT 724.215 213.300 724.545 214.150 ;
        RECT 724.715 213.520 724.885 214.320 ;
      LAYER li1 ;
        RECT 725.135 213.300 725.305 214.150 ;
      LAYER li1 ;
        RECT 725.475 213.520 725.805 214.320 ;
      LAYER li1 ;
        RECT 725.975 213.300 726.145 214.150 ;
      LAYER li1 ;
        RECT 726.315 213.520 726.645 214.320 ;
      LAYER li1 ;
        RECT 726.815 213.300 726.985 214.150 ;
      LAYER li1 ;
        RECT 727.155 213.520 727.485 214.320 ;
      LAYER li1 ;
        RECT 727.655 213.300 727.825 214.150 ;
      LAYER li1 ;
        RECT 723.375 213.130 724.875 213.300 ;
      LAYER li1 ;
        RECT 725.135 213.130 727.825 213.300 ;
      LAYER li1 ;
        RECT 727.995 213.170 728.325 214.320 ;
        RECT 728.885 213.155 729.175 214.320 ;
        RECT 758.785 213.155 759.075 214.320 ;
      LAYER li1 ;
        RECT 759.245 213.885 764.590 214.320 ;
        RECT 675.580 212.760 676.680 212.960 ;
      LAYER li1 ;
        RECT 676.860 212.930 677.035 213.130 ;
        RECT 676.860 212.760 679.485 212.930 ;
        RECT 676.860 212.590 677.035 212.760 ;
      LAYER li1 ;
        RECT 679.730 212.590 679.985 213.130 ;
        RECT 681.560 212.760 682.660 212.960 ;
      LAYER li1 ;
        RECT 682.840 212.930 683.015 213.130 ;
        RECT 682.840 212.760 685.465 212.930 ;
        RECT 682.840 212.590 683.015 212.760 ;
      LAYER li1 ;
        RECT 685.710 212.590 685.965 213.130 ;
        RECT 687.540 212.760 688.640 212.960 ;
      LAYER li1 ;
        RECT 688.820 212.930 688.995 213.130 ;
        RECT 688.820 212.760 691.445 212.930 ;
        RECT 688.820 212.590 688.995 212.760 ;
      LAYER li1 ;
        RECT 691.690 212.590 691.945 213.130 ;
        RECT 693.520 212.760 694.620 212.960 ;
      LAYER li1 ;
        RECT 694.800 212.930 694.975 213.130 ;
        RECT 694.800 212.760 697.425 212.930 ;
        RECT 694.800 212.590 694.975 212.760 ;
      LAYER li1 ;
        RECT 697.670 212.590 697.925 213.130 ;
        RECT 699.500 212.760 700.600 212.960 ;
      LAYER li1 ;
        RECT 700.780 212.930 700.955 213.130 ;
        RECT 700.780 212.760 703.405 212.930 ;
        RECT 700.780 212.590 700.955 212.760 ;
      LAYER li1 ;
        RECT 703.650 212.590 703.905 213.130 ;
        RECT 705.480 212.760 706.580 212.960 ;
      LAYER li1 ;
        RECT 706.760 212.930 706.935 213.130 ;
        RECT 706.760 212.760 709.385 212.930 ;
        RECT 706.760 212.590 706.935 212.760 ;
      LAYER li1 ;
        RECT 709.630 212.590 709.885 213.130 ;
        RECT 711.460 212.760 712.560 212.960 ;
      LAYER li1 ;
        RECT 712.740 212.930 712.915 213.130 ;
        RECT 712.740 212.760 715.365 212.930 ;
        RECT 712.740 212.590 712.915 212.760 ;
      LAYER li1 ;
        RECT 715.610 212.590 715.865 213.130 ;
        RECT 717.440 212.760 718.540 212.960 ;
      LAYER li1 ;
        RECT 718.720 212.930 718.895 213.130 ;
        RECT 718.720 212.760 721.345 212.930 ;
        RECT 718.720 212.590 718.895 212.760 ;
      LAYER li1 ;
        RECT 721.590 212.590 721.845 213.130 ;
        RECT 723.420 212.760 724.520 212.960 ;
      LAYER li1 ;
        RECT 724.700 212.930 724.875 213.130 ;
        RECT 724.700 212.760 727.325 212.930 ;
        RECT 724.700 212.590 724.875 212.760 ;
      LAYER li1 ;
        RECT 727.570 212.590 727.825 213.130 ;
        RECT 762.650 212.635 763.000 213.885 ;
      LAYER li1 ;
        RECT 764.765 213.155 765.055 214.320 ;
        RECT 765.235 213.300 765.565 214.150 ;
        RECT 765.735 213.520 765.905 214.320 ;
        RECT 766.075 213.300 766.405 214.150 ;
        RECT 766.575 213.520 766.745 214.320 ;
      LAYER li1 ;
        RECT 766.995 213.300 767.165 214.150 ;
      LAYER li1 ;
        RECT 767.335 213.520 767.665 214.320 ;
      LAYER li1 ;
        RECT 767.835 213.300 768.005 214.150 ;
      LAYER li1 ;
        RECT 768.175 213.520 768.505 214.320 ;
      LAYER li1 ;
        RECT 768.675 213.300 768.845 214.150 ;
      LAYER li1 ;
        RECT 769.015 213.520 769.345 214.320 ;
      LAYER li1 ;
        RECT 769.515 213.300 769.685 214.150 ;
      LAYER li1 ;
        RECT 765.235 213.130 766.735 213.300 ;
      LAYER li1 ;
        RECT 766.995 213.130 769.685 213.300 ;
      LAYER li1 ;
        RECT 769.855 213.170 770.185 214.320 ;
        RECT 770.745 213.155 771.035 214.320 ;
        RECT 771.215 213.300 771.545 214.150 ;
        RECT 771.715 213.520 771.885 214.320 ;
        RECT 772.055 213.300 772.385 214.150 ;
        RECT 772.555 213.520 772.725 214.320 ;
      LAYER li1 ;
        RECT 772.975 213.300 773.145 214.150 ;
      LAYER li1 ;
        RECT 773.315 213.520 773.645 214.320 ;
      LAYER li1 ;
        RECT 773.815 213.300 773.985 214.150 ;
      LAYER li1 ;
        RECT 774.155 213.520 774.485 214.320 ;
      LAYER li1 ;
        RECT 774.655 213.300 774.825 214.150 ;
      LAYER li1 ;
        RECT 774.995 213.520 775.325 214.320 ;
      LAYER li1 ;
        RECT 775.495 213.300 775.665 214.150 ;
      LAYER li1 ;
        RECT 771.215 213.130 772.715 213.300 ;
      LAYER li1 ;
        RECT 772.975 213.130 775.665 213.300 ;
      LAYER li1 ;
        RECT 775.835 213.170 776.165 214.320 ;
        RECT 776.725 213.155 777.015 214.320 ;
        RECT 777.195 213.300 777.525 214.150 ;
        RECT 777.695 213.520 777.865 214.320 ;
        RECT 778.035 213.300 778.365 214.150 ;
        RECT 778.535 213.520 778.705 214.320 ;
      LAYER li1 ;
        RECT 778.955 213.300 779.125 214.150 ;
      LAYER li1 ;
        RECT 779.295 213.520 779.625 214.320 ;
      LAYER li1 ;
        RECT 779.795 213.300 779.965 214.150 ;
      LAYER li1 ;
        RECT 780.135 213.520 780.465 214.320 ;
      LAYER li1 ;
        RECT 780.635 213.300 780.805 214.150 ;
      LAYER li1 ;
        RECT 780.975 213.520 781.305 214.320 ;
      LAYER li1 ;
        RECT 781.475 213.300 781.645 214.150 ;
      LAYER li1 ;
        RECT 777.195 213.130 778.695 213.300 ;
      LAYER li1 ;
        RECT 778.955 213.130 781.645 213.300 ;
      LAYER li1 ;
        RECT 781.815 213.170 782.145 214.320 ;
        RECT 782.705 213.155 782.995 214.320 ;
        RECT 783.175 213.300 783.505 214.150 ;
        RECT 783.675 213.520 783.845 214.320 ;
        RECT 784.015 213.300 784.345 214.150 ;
        RECT 784.515 213.520 784.685 214.320 ;
      LAYER li1 ;
        RECT 784.935 213.300 785.105 214.150 ;
      LAYER li1 ;
        RECT 785.275 213.520 785.605 214.320 ;
      LAYER li1 ;
        RECT 785.775 213.300 785.945 214.150 ;
      LAYER li1 ;
        RECT 786.115 213.520 786.445 214.320 ;
      LAYER li1 ;
        RECT 786.615 213.300 786.785 214.150 ;
      LAYER li1 ;
        RECT 786.955 213.520 787.285 214.320 ;
      LAYER li1 ;
        RECT 787.455 213.300 787.625 214.150 ;
      LAYER li1 ;
        RECT 783.175 213.130 784.675 213.300 ;
      LAYER li1 ;
        RECT 784.935 213.130 787.625 213.300 ;
      LAYER li1 ;
        RECT 787.795 213.170 788.125 214.320 ;
        RECT 788.685 213.155 788.975 214.320 ;
        RECT 789.535 213.170 789.865 214.320 ;
        RECT 790.375 213.520 790.705 214.320 ;
        RECT 791.215 213.520 791.545 214.320 ;
        RECT 792.055 213.520 792.385 214.320 ;
        RECT 792.975 213.520 793.145 214.320 ;
        RECT 793.315 213.300 793.645 214.150 ;
        RECT 793.815 213.520 793.985 214.320 ;
        RECT 794.155 213.300 794.485 214.150 ;
        RECT 766.560 212.930 766.735 213.130 ;
        RECT 766.560 212.760 769.185 212.930 ;
        RECT 766.560 212.590 766.735 212.760 ;
      LAYER li1 ;
        RECT 769.430 212.590 769.685 213.130 ;
      LAYER li1 ;
        RECT 772.540 212.930 772.715 213.130 ;
        RECT 772.540 212.760 775.165 212.930 ;
        RECT 772.540 212.590 772.715 212.760 ;
      LAYER li1 ;
        RECT 775.410 212.590 775.665 213.130 ;
      LAYER li1 ;
        RECT 778.520 212.930 778.695 213.130 ;
        RECT 778.520 212.760 781.145 212.930 ;
        RECT 778.520 212.590 778.695 212.760 ;
      LAYER li1 ;
        RECT 781.390 212.590 781.645 213.130 ;
      LAYER li1 ;
        RECT 784.500 212.930 784.675 213.130 ;
        RECT 784.500 212.760 787.125 212.930 ;
        RECT 784.500 212.590 784.675 212.760 ;
      LAYER li1 ;
        RECT 787.370 212.590 787.625 213.130 ;
      LAYER li1 ;
        RECT 792.985 213.130 794.485 213.300 ;
        RECT 794.665 213.155 794.955 214.320 ;
        RECT 2146.085 213.155 2146.375 214.320 ;
      LAYER li1 ;
        RECT 2146.545 213.885 2151.890 214.320 ;
      LAYER li1 ;
        RECT 792.985 212.930 793.160 213.130 ;
        RECT 790.535 212.760 793.160 212.930 ;
      LAYER li1 ;
        RECT 793.340 212.760 794.440 212.960 ;
      LAYER li1 ;
        RECT 669.085 211.770 669.375 212.495 ;
        RECT 675.065 211.770 675.355 212.495 ;
        RECT 675.615 212.420 677.035 212.590 ;
      LAYER li1 ;
        RECT 677.295 212.420 679.985 212.590 ;
      LAYER li1 ;
        RECT 675.615 211.940 675.785 212.420 ;
        RECT 675.955 211.770 676.285 212.250 ;
        RECT 676.455 211.945 676.625 212.420 ;
        RECT 676.795 211.770 677.125 212.250 ;
      LAYER li1 ;
        RECT 677.295 211.940 677.465 212.420 ;
      LAYER li1 ;
        RECT 677.635 211.770 677.965 212.250 ;
      LAYER li1 ;
        RECT 678.135 211.940 678.305 212.420 ;
      LAYER li1 ;
        RECT 678.475 211.770 678.805 212.250 ;
      LAYER li1 ;
        RECT 678.975 211.940 679.145 212.420 ;
      LAYER li1 ;
        RECT 679.315 211.770 679.645 212.250 ;
      LAYER li1 ;
        RECT 679.815 211.940 679.985 212.420 ;
      LAYER li1 ;
        RECT 680.155 211.770 680.485 212.570 ;
        RECT 681.045 211.770 681.335 212.495 ;
        RECT 681.595 212.420 683.015 212.590 ;
      LAYER li1 ;
        RECT 683.275 212.420 685.965 212.590 ;
      LAYER li1 ;
        RECT 681.595 211.940 681.765 212.420 ;
        RECT 681.935 211.770 682.265 212.250 ;
        RECT 682.435 211.945 682.605 212.420 ;
        RECT 682.775 211.770 683.105 212.250 ;
      LAYER li1 ;
        RECT 683.275 211.940 683.445 212.420 ;
      LAYER li1 ;
        RECT 683.615 211.770 683.945 212.250 ;
      LAYER li1 ;
        RECT 684.115 211.940 684.285 212.420 ;
      LAYER li1 ;
        RECT 684.455 211.770 684.785 212.250 ;
      LAYER li1 ;
        RECT 684.955 211.940 685.125 212.420 ;
      LAYER li1 ;
        RECT 685.295 211.770 685.625 212.250 ;
      LAYER li1 ;
        RECT 685.795 211.940 685.965 212.420 ;
      LAYER li1 ;
        RECT 686.135 211.770 686.465 212.570 ;
        RECT 687.025 211.770 687.315 212.495 ;
        RECT 687.575 212.420 688.995 212.590 ;
      LAYER li1 ;
        RECT 689.255 212.420 691.945 212.590 ;
      LAYER li1 ;
        RECT 687.575 211.940 687.745 212.420 ;
        RECT 687.915 211.770 688.245 212.250 ;
        RECT 688.415 211.945 688.585 212.420 ;
        RECT 688.755 211.770 689.085 212.250 ;
      LAYER li1 ;
        RECT 689.255 211.940 689.425 212.420 ;
      LAYER li1 ;
        RECT 689.595 211.770 689.925 212.250 ;
      LAYER li1 ;
        RECT 690.095 211.940 690.265 212.420 ;
      LAYER li1 ;
        RECT 690.435 211.770 690.765 212.250 ;
      LAYER li1 ;
        RECT 690.935 211.940 691.105 212.420 ;
      LAYER li1 ;
        RECT 691.275 211.770 691.605 212.250 ;
      LAYER li1 ;
        RECT 691.775 211.940 691.945 212.420 ;
      LAYER li1 ;
        RECT 692.115 211.770 692.445 212.570 ;
        RECT 693.005 211.770 693.295 212.495 ;
        RECT 693.555 212.420 694.975 212.590 ;
      LAYER li1 ;
        RECT 695.235 212.420 697.925 212.590 ;
      LAYER li1 ;
        RECT 693.555 211.940 693.725 212.420 ;
        RECT 693.895 211.770 694.225 212.250 ;
        RECT 694.395 211.945 694.565 212.420 ;
        RECT 694.735 211.770 695.065 212.250 ;
      LAYER li1 ;
        RECT 695.235 211.940 695.405 212.420 ;
      LAYER li1 ;
        RECT 695.575 211.770 695.905 212.250 ;
      LAYER li1 ;
        RECT 696.075 211.940 696.245 212.420 ;
      LAYER li1 ;
        RECT 696.415 211.770 696.745 212.250 ;
      LAYER li1 ;
        RECT 696.915 211.940 697.085 212.420 ;
      LAYER li1 ;
        RECT 697.255 211.770 697.585 212.250 ;
      LAYER li1 ;
        RECT 697.755 211.940 697.925 212.420 ;
      LAYER li1 ;
        RECT 698.095 211.770 698.425 212.570 ;
        RECT 698.985 211.770 699.275 212.495 ;
        RECT 699.535 212.420 700.955 212.590 ;
      LAYER li1 ;
        RECT 701.215 212.420 703.905 212.590 ;
      LAYER li1 ;
        RECT 699.535 211.940 699.705 212.420 ;
        RECT 699.875 211.770 700.205 212.250 ;
        RECT 700.375 211.945 700.545 212.420 ;
        RECT 700.715 211.770 701.045 212.250 ;
      LAYER li1 ;
        RECT 701.215 211.940 701.385 212.420 ;
      LAYER li1 ;
        RECT 701.555 211.770 701.885 212.250 ;
      LAYER li1 ;
        RECT 702.055 211.940 702.225 212.420 ;
      LAYER li1 ;
        RECT 702.395 211.770 702.725 212.250 ;
      LAYER li1 ;
        RECT 702.895 211.940 703.065 212.420 ;
      LAYER li1 ;
        RECT 703.235 211.770 703.565 212.250 ;
      LAYER li1 ;
        RECT 703.735 211.940 703.905 212.420 ;
      LAYER li1 ;
        RECT 704.075 211.770 704.405 212.570 ;
        RECT 704.965 211.770 705.255 212.495 ;
        RECT 705.515 212.420 706.935 212.590 ;
      LAYER li1 ;
        RECT 707.195 212.420 709.885 212.590 ;
      LAYER li1 ;
        RECT 705.515 211.940 705.685 212.420 ;
        RECT 705.855 211.770 706.185 212.250 ;
        RECT 706.355 211.945 706.525 212.420 ;
        RECT 706.695 211.770 707.025 212.250 ;
      LAYER li1 ;
        RECT 707.195 211.940 707.365 212.420 ;
      LAYER li1 ;
        RECT 707.535 211.770 707.865 212.250 ;
      LAYER li1 ;
        RECT 708.035 211.940 708.205 212.420 ;
      LAYER li1 ;
        RECT 708.375 211.770 708.705 212.250 ;
      LAYER li1 ;
        RECT 708.875 211.940 709.045 212.420 ;
      LAYER li1 ;
        RECT 709.215 211.770 709.545 212.250 ;
      LAYER li1 ;
        RECT 709.715 211.940 709.885 212.420 ;
      LAYER li1 ;
        RECT 710.055 211.770 710.385 212.570 ;
        RECT 710.945 211.770 711.235 212.495 ;
        RECT 711.495 212.420 712.915 212.590 ;
      LAYER li1 ;
        RECT 713.175 212.420 715.865 212.590 ;
      LAYER li1 ;
        RECT 711.495 211.940 711.665 212.420 ;
        RECT 711.835 211.770 712.165 212.250 ;
        RECT 712.335 211.945 712.505 212.420 ;
        RECT 712.675 211.770 713.005 212.250 ;
      LAYER li1 ;
        RECT 713.175 211.940 713.345 212.420 ;
      LAYER li1 ;
        RECT 713.515 211.770 713.845 212.250 ;
      LAYER li1 ;
        RECT 714.015 211.940 714.185 212.420 ;
      LAYER li1 ;
        RECT 714.355 211.770 714.685 212.250 ;
      LAYER li1 ;
        RECT 714.855 211.940 715.025 212.420 ;
      LAYER li1 ;
        RECT 715.195 211.770 715.525 212.250 ;
      LAYER li1 ;
        RECT 715.695 211.940 715.865 212.420 ;
      LAYER li1 ;
        RECT 716.035 211.770 716.365 212.570 ;
        RECT 716.925 211.770 717.215 212.495 ;
        RECT 717.475 212.420 718.895 212.590 ;
      LAYER li1 ;
        RECT 719.155 212.420 721.845 212.590 ;
      LAYER li1 ;
        RECT 717.475 211.940 717.645 212.420 ;
        RECT 717.815 211.770 718.145 212.250 ;
        RECT 718.315 211.945 718.485 212.420 ;
        RECT 718.655 211.770 718.985 212.250 ;
      LAYER li1 ;
        RECT 719.155 211.940 719.325 212.420 ;
      LAYER li1 ;
        RECT 719.495 211.770 719.825 212.250 ;
      LAYER li1 ;
        RECT 719.995 211.940 720.165 212.420 ;
      LAYER li1 ;
        RECT 720.335 211.770 720.665 212.250 ;
      LAYER li1 ;
        RECT 720.835 211.940 721.005 212.420 ;
      LAYER li1 ;
        RECT 721.175 211.770 721.505 212.250 ;
      LAYER li1 ;
        RECT 721.675 211.940 721.845 212.420 ;
      LAYER li1 ;
        RECT 722.015 211.770 722.345 212.570 ;
        RECT 722.905 211.770 723.195 212.495 ;
        RECT 723.455 212.420 724.875 212.590 ;
      LAYER li1 ;
        RECT 725.135 212.420 727.825 212.590 ;
      LAYER li1 ;
        RECT 723.455 211.940 723.625 212.420 ;
        RECT 723.795 211.770 724.125 212.250 ;
        RECT 724.295 211.945 724.465 212.420 ;
        RECT 724.635 211.770 724.965 212.250 ;
      LAYER li1 ;
        RECT 725.135 211.940 725.305 212.420 ;
      LAYER li1 ;
        RECT 725.475 211.770 725.805 212.250 ;
      LAYER li1 ;
        RECT 725.975 211.940 726.145 212.420 ;
      LAYER li1 ;
        RECT 726.315 211.770 726.645 212.250 ;
      LAYER li1 ;
        RECT 726.815 211.940 726.985 212.420 ;
      LAYER li1 ;
        RECT 727.155 211.770 727.485 212.250 ;
      LAYER li1 ;
        RECT 727.655 211.940 727.825 212.420 ;
      LAYER li1 ;
        RECT 727.995 211.770 728.325 212.570 ;
        RECT 728.885 211.770 729.175 212.495 ;
        RECT 758.785 211.770 759.075 212.495 ;
        RECT 764.765 211.770 765.055 212.495 ;
        RECT 765.315 212.420 766.735 212.590 ;
      LAYER li1 ;
        RECT 766.995 212.420 769.685 212.590 ;
      LAYER li1 ;
        RECT 765.315 211.940 765.485 212.420 ;
        RECT 765.655 211.770 765.985 212.250 ;
        RECT 766.155 211.945 766.325 212.420 ;
        RECT 766.495 211.770 766.825 212.250 ;
      LAYER li1 ;
        RECT 766.995 211.940 767.165 212.420 ;
      LAYER li1 ;
        RECT 767.335 211.770 767.665 212.250 ;
      LAYER li1 ;
        RECT 767.835 211.940 768.005 212.420 ;
      LAYER li1 ;
        RECT 768.175 211.770 768.505 212.250 ;
      LAYER li1 ;
        RECT 768.675 211.940 768.845 212.420 ;
      LAYER li1 ;
        RECT 769.015 211.770 769.345 212.250 ;
      LAYER li1 ;
        RECT 769.515 211.940 769.685 212.420 ;
      LAYER li1 ;
        RECT 769.855 211.770 770.185 212.570 ;
        RECT 770.745 211.770 771.035 212.495 ;
        RECT 771.295 212.420 772.715 212.590 ;
      LAYER li1 ;
        RECT 772.975 212.420 775.665 212.590 ;
      LAYER li1 ;
        RECT 771.295 211.940 771.465 212.420 ;
        RECT 771.635 211.770 771.965 212.250 ;
        RECT 772.135 211.945 772.305 212.420 ;
        RECT 772.475 211.770 772.805 212.250 ;
      LAYER li1 ;
        RECT 772.975 211.940 773.145 212.420 ;
      LAYER li1 ;
        RECT 773.315 211.770 773.645 212.250 ;
      LAYER li1 ;
        RECT 773.815 211.940 773.985 212.420 ;
      LAYER li1 ;
        RECT 774.155 211.770 774.485 212.250 ;
      LAYER li1 ;
        RECT 774.655 211.940 774.825 212.420 ;
      LAYER li1 ;
        RECT 774.995 211.770 775.325 212.250 ;
      LAYER li1 ;
        RECT 775.495 211.940 775.665 212.420 ;
      LAYER li1 ;
        RECT 775.835 211.770 776.165 212.570 ;
        RECT 776.725 211.770 777.015 212.495 ;
        RECT 777.275 212.420 778.695 212.590 ;
      LAYER li1 ;
        RECT 778.955 212.420 781.645 212.590 ;
      LAYER li1 ;
        RECT 777.275 211.940 777.445 212.420 ;
        RECT 777.615 211.770 777.945 212.250 ;
        RECT 778.115 211.945 778.285 212.420 ;
        RECT 778.455 211.770 778.785 212.250 ;
      LAYER li1 ;
        RECT 778.955 211.940 779.125 212.420 ;
      LAYER li1 ;
        RECT 779.295 211.770 779.625 212.250 ;
      LAYER li1 ;
        RECT 779.795 211.940 779.965 212.420 ;
      LAYER li1 ;
        RECT 780.135 211.770 780.465 212.250 ;
      LAYER li1 ;
        RECT 780.635 211.940 780.805 212.420 ;
      LAYER li1 ;
        RECT 780.975 211.770 781.305 212.250 ;
      LAYER li1 ;
        RECT 781.475 211.940 781.645 212.420 ;
      LAYER li1 ;
        RECT 781.815 211.770 782.145 212.570 ;
        RECT 782.705 211.770 782.995 212.495 ;
        RECT 783.255 212.420 784.675 212.590 ;
      LAYER li1 ;
        RECT 784.935 212.420 787.625 212.590 ;
      LAYER li1 ;
        RECT 792.985 212.590 793.160 212.760 ;
      LAYER li1 ;
        RECT 2149.950 212.635 2150.300 213.885 ;
      LAYER li1 ;
        RECT 2152.065 213.155 2152.355 214.320 ;
        RECT 2152.535 213.300 2152.865 214.150 ;
        RECT 2153.035 213.520 2153.205 214.320 ;
        RECT 2153.375 213.300 2153.705 214.150 ;
        RECT 2153.875 213.520 2154.045 214.320 ;
        RECT 2154.635 213.520 2154.965 214.320 ;
        RECT 2155.475 213.520 2155.805 214.320 ;
        RECT 2156.315 213.520 2156.645 214.320 ;
        RECT 2152.535 213.130 2154.035 213.300 ;
        RECT 2157.155 213.170 2157.485 214.320 ;
        RECT 2158.045 213.155 2158.335 214.320 ;
        RECT 2158.515 213.300 2158.845 214.150 ;
        RECT 2159.015 213.520 2159.185 214.320 ;
        RECT 2159.355 213.300 2159.685 214.150 ;
        RECT 2159.855 213.520 2160.025 214.320 ;
        RECT 2160.615 213.520 2160.945 214.320 ;
        RECT 2161.455 213.520 2161.785 214.320 ;
        RECT 2162.295 213.520 2162.625 214.320 ;
        RECT 2158.515 213.130 2160.015 213.300 ;
        RECT 2163.135 213.170 2163.465 214.320 ;
        RECT 2164.025 213.155 2164.315 214.320 ;
        RECT 2164.495 213.300 2164.825 214.150 ;
        RECT 2164.995 213.520 2165.165 214.320 ;
        RECT 2165.335 213.300 2165.665 214.150 ;
        RECT 2165.835 213.520 2166.005 214.320 ;
        RECT 2166.595 213.520 2166.925 214.320 ;
        RECT 2167.435 213.520 2167.765 214.320 ;
        RECT 2168.275 213.520 2168.605 214.320 ;
        RECT 2164.495 213.130 2165.995 213.300 ;
        RECT 2169.115 213.170 2169.445 214.320 ;
        RECT 2170.005 213.155 2170.295 214.320 ;
        RECT 2170.475 213.300 2170.805 214.150 ;
        RECT 2170.975 213.520 2171.145 214.320 ;
        RECT 2171.315 213.300 2171.645 214.150 ;
        RECT 2171.815 213.520 2171.985 214.320 ;
        RECT 2172.575 213.520 2172.905 214.320 ;
        RECT 2173.415 213.520 2173.745 214.320 ;
        RECT 2174.255 213.520 2174.585 214.320 ;
        RECT 2170.475 213.130 2171.975 213.300 ;
        RECT 2175.095 213.170 2175.425 214.320 ;
        RECT 2175.985 213.155 2176.275 214.320 ;
        RECT 2176.455 213.300 2176.785 214.150 ;
        RECT 2176.955 213.520 2177.125 214.320 ;
        RECT 2177.295 213.300 2177.625 214.150 ;
        RECT 2177.795 213.520 2177.965 214.320 ;
        RECT 2178.555 213.520 2178.885 214.320 ;
        RECT 2179.395 213.520 2179.725 214.320 ;
        RECT 2180.235 213.520 2180.565 214.320 ;
        RECT 2176.455 213.130 2177.955 213.300 ;
        RECT 2181.075 213.170 2181.405 214.320 ;
        RECT 2181.965 213.155 2182.255 214.320 ;
        RECT 2182.435 213.300 2182.765 214.150 ;
        RECT 2182.935 213.520 2183.105 214.320 ;
        RECT 2183.275 213.300 2183.605 214.150 ;
        RECT 2183.775 213.520 2183.945 214.320 ;
        RECT 2184.535 213.520 2184.865 214.320 ;
        RECT 2185.375 213.520 2185.705 214.320 ;
        RECT 2186.215 213.520 2186.545 214.320 ;
        RECT 2182.435 213.130 2183.935 213.300 ;
        RECT 2187.055 213.170 2187.385 214.320 ;
        RECT 2187.945 213.155 2188.235 214.320 ;
        RECT 2188.415 213.300 2188.745 214.150 ;
        RECT 2188.915 213.520 2189.085 214.320 ;
        RECT 2189.255 213.300 2189.585 214.150 ;
        RECT 2189.755 213.520 2189.925 214.320 ;
        RECT 2190.515 213.520 2190.845 214.320 ;
        RECT 2191.355 213.520 2191.685 214.320 ;
        RECT 2192.195 213.520 2192.525 214.320 ;
        RECT 2188.415 213.130 2189.915 213.300 ;
        RECT 2193.035 213.170 2193.365 214.320 ;
        RECT 2193.925 213.155 2194.215 214.320 ;
        RECT 2194.395 213.300 2194.725 214.150 ;
        RECT 2194.895 213.520 2195.065 214.320 ;
        RECT 2195.235 213.300 2195.565 214.150 ;
        RECT 2195.735 213.520 2195.905 214.320 ;
        RECT 2196.495 213.520 2196.825 214.320 ;
        RECT 2197.335 213.520 2197.665 214.320 ;
        RECT 2198.175 213.520 2198.505 214.320 ;
        RECT 2194.395 213.130 2195.895 213.300 ;
        RECT 2199.015 213.170 2199.345 214.320 ;
        RECT 2199.905 213.155 2200.195 214.320 ;
        RECT 2200.375 213.300 2200.705 214.150 ;
        RECT 2200.875 213.520 2201.045 214.320 ;
        RECT 2201.215 213.300 2201.545 214.150 ;
        RECT 2201.715 213.520 2201.885 214.320 ;
        RECT 2202.475 213.520 2202.805 214.320 ;
        RECT 2203.315 213.520 2203.645 214.320 ;
        RECT 2204.155 213.520 2204.485 214.320 ;
        RECT 2200.375 213.130 2201.875 213.300 ;
        RECT 2204.995 213.170 2205.325 214.320 ;
        RECT 2205.885 213.155 2206.175 214.320 ;
        RECT 2235.785 213.155 2236.075 214.320 ;
      LAYER li1 ;
        RECT 2236.245 213.885 2241.590 214.320 ;
        RECT 2152.580 212.760 2153.680 212.960 ;
      LAYER li1 ;
        RECT 2153.860 212.930 2154.035 213.130 ;
        RECT 2153.860 212.760 2156.485 212.930 ;
      LAYER li1 ;
        RECT 2158.560 212.760 2159.660 212.960 ;
      LAYER li1 ;
        RECT 2159.840 212.930 2160.015 213.130 ;
        RECT 2159.840 212.760 2162.465 212.930 ;
      LAYER li1 ;
        RECT 2164.540 212.760 2165.640 212.960 ;
      LAYER li1 ;
        RECT 2165.820 212.930 2165.995 213.130 ;
        RECT 2165.820 212.760 2168.445 212.930 ;
      LAYER li1 ;
        RECT 2170.520 212.760 2171.620 212.960 ;
      LAYER li1 ;
        RECT 2171.800 212.930 2171.975 213.130 ;
        RECT 2171.800 212.760 2174.425 212.930 ;
      LAYER li1 ;
        RECT 2176.500 212.760 2177.600 212.960 ;
      LAYER li1 ;
        RECT 2177.780 212.930 2177.955 213.130 ;
        RECT 2177.780 212.760 2180.405 212.930 ;
      LAYER li1 ;
        RECT 2182.480 212.760 2183.580 212.960 ;
      LAYER li1 ;
        RECT 2183.760 212.930 2183.935 213.130 ;
        RECT 2183.760 212.760 2186.385 212.930 ;
      LAYER li1 ;
        RECT 2188.460 212.760 2189.560 212.960 ;
      LAYER li1 ;
        RECT 2189.740 212.930 2189.915 213.130 ;
        RECT 2189.740 212.760 2192.365 212.930 ;
      LAYER li1 ;
        RECT 2194.440 212.760 2195.540 212.960 ;
      LAYER li1 ;
        RECT 2195.720 212.930 2195.895 213.130 ;
        RECT 2195.720 212.760 2198.345 212.930 ;
      LAYER li1 ;
        RECT 2200.420 212.760 2201.520 212.960 ;
      LAYER li1 ;
        RECT 2201.700 212.930 2201.875 213.130 ;
        RECT 2201.700 212.760 2204.325 212.930 ;
        RECT 2153.860 212.590 2154.035 212.760 ;
        RECT 2159.840 212.590 2160.015 212.760 ;
        RECT 2165.820 212.590 2165.995 212.760 ;
        RECT 2171.800 212.590 2171.975 212.760 ;
        RECT 2177.780 212.590 2177.955 212.760 ;
        RECT 2183.760 212.590 2183.935 212.760 ;
        RECT 2189.740 212.590 2189.915 212.760 ;
        RECT 2195.720 212.590 2195.895 212.760 ;
        RECT 2201.700 212.590 2201.875 212.760 ;
      LAYER li1 ;
        RECT 2239.650 212.635 2240.000 213.885 ;
      LAYER li1 ;
        RECT 2241.765 213.155 2242.055 214.320 ;
        RECT 2242.235 213.300 2242.565 214.150 ;
        RECT 2242.735 213.520 2242.905 214.320 ;
        RECT 2243.075 213.300 2243.405 214.150 ;
        RECT 2243.575 213.520 2243.745 214.320 ;
        RECT 2244.335 213.520 2244.665 214.320 ;
        RECT 2245.175 213.520 2245.505 214.320 ;
        RECT 2246.015 213.520 2246.345 214.320 ;
        RECT 2242.235 213.130 2243.735 213.300 ;
        RECT 2246.855 213.170 2247.185 214.320 ;
        RECT 2247.745 213.155 2248.035 214.320 ;
        RECT 2248.215 213.300 2248.545 214.150 ;
        RECT 2248.715 213.520 2248.885 214.320 ;
        RECT 2249.055 213.300 2249.385 214.150 ;
        RECT 2249.555 213.520 2249.725 214.320 ;
        RECT 2250.315 213.520 2250.645 214.320 ;
        RECT 2251.155 213.520 2251.485 214.320 ;
        RECT 2251.995 213.520 2252.325 214.320 ;
        RECT 2248.215 213.130 2249.715 213.300 ;
        RECT 2252.835 213.170 2253.165 214.320 ;
        RECT 2253.725 213.155 2254.015 214.320 ;
        RECT 2254.195 213.300 2254.525 214.150 ;
        RECT 2254.695 213.520 2254.865 214.320 ;
        RECT 2255.035 213.300 2255.365 214.150 ;
        RECT 2255.535 213.520 2255.705 214.320 ;
        RECT 2256.295 213.520 2256.625 214.320 ;
        RECT 2257.135 213.520 2257.465 214.320 ;
        RECT 2257.975 213.520 2258.305 214.320 ;
        RECT 2254.195 213.130 2255.695 213.300 ;
        RECT 2258.815 213.170 2259.145 214.320 ;
        RECT 2259.705 213.155 2259.995 214.320 ;
        RECT 2260.175 213.300 2260.505 214.150 ;
        RECT 2260.675 213.520 2260.845 214.320 ;
        RECT 2261.015 213.300 2261.345 214.150 ;
        RECT 2261.515 213.520 2261.685 214.320 ;
        RECT 2262.275 213.520 2262.605 214.320 ;
        RECT 2263.115 213.520 2263.445 214.320 ;
        RECT 2263.955 213.520 2264.285 214.320 ;
        RECT 2260.175 213.130 2261.675 213.300 ;
        RECT 2264.795 213.170 2265.125 214.320 ;
        RECT 2265.685 213.155 2265.975 214.320 ;
        RECT 2266.535 213.170 2266.865 214.320 ;
      LAYER li1 ;
        RECT 2267.035 213.300 2267.205 214.150 ;
      LAYER li1 ;
        RECT 2267.375 213.520 2267.705 214.320 ;
      LAYER li1 ;
        RECT 2267.875 213.300 2268.045 214.150 ;
      LAYER li1 ;
        RECT 2268.215 213.520 2268.545 214.320 ;
      LAYER li1 ;
        RECT 2268.715 213.300 2268.885 214.150 ;
      LAYER li1 ;
        RECT 2269.055 213.520 2269.385 214.320 ;
      LAYER li1 ;
        RECT 2269.555 213.300 2269.725 214.150 ;
      LAYER li1 ;
        RECT 2269.975 213.520 2270.145 214.320 ;
        RECT 2270.315 213.300 2270.645 214.150 ;
        RECT 2270.815 213.520 2270.985 214.320 ;
        RECT 2271.155 213.300 2271.485 214.150 ;
      LAYER li1 ;
        RECT 2242.280 212.760 2243.380 212.960 ;
      LAYER li1 ;
        RECT 2243.560 212.930 2243.735 213.130 ;
        RECT 2243.560 212.760 2246.185 212.930 ;
      LAYER li1 ;
        RECT 2248.260 212.760 2249.360 212.960 ;
      LAYER li1 ;
        RECT 2249.540 212.930 2249.715 213.130 ;
        RECT 2249.540 212.760 2252.165 212.930 ;
      LAYER li1 ;
        RECT 2254.240 212.760 2255.340 212.960 ;
      LAYER li1 ;
        RECT 2255.520 212.930 2255.695 213.130 ;
        RECT 2255.520 212.760 2258.145 212.930 ;
      LAYER li1 ;
        RECT 2260.220 212.760 2261.320 212.960 ;
      LAYER li1 ;
        RECT 2261.500 212.930 2261.675 213.130 ;
      LAYER li1 ;
        RECT 2267.035 213.130 2269.725 213.300 ;
      LAYER li1 ;
        RECT 2269.985 213.130 2271.485 213.300 ;
        RECT 2271.665 213.155 2271.955 214.320 ;
        RECT 2261.500 212.760 2264.125 212.930 ;
        RECT 2243.560 212.590 2243.735 212.760 ;
        RECT 2249.540 212.590 2249.715 212.760 ;
        RECT 2255.520 212.590 2255.695 212.760 ;
        RECT 2261.500 212.590 2261.675 212.760 ;
        RECT 783.255 211.940 783.425 212.420 ;
        RECT 783.595 211.770 783.925 212.250 ;
        RECT 784.095 211.945 784.265 212.420 ;
        RECT 784.435 211.770 784.765 212.250 ;
      LAYER li1 ;
        RECT 784.935 211.940 785.105 212.420 ;
      LAYER li1 ;
        RECT 785.275 211.770 785.605 212.250 ;
      LAYER li1 ;
        RECT 785.775 211.940 785.945 212.420 ;
      LAYER li1 ;
        RECT 786.115 211.770 786.445 212.250 ;
      LAYER li1 ;
        RECT 786.615 211.940 786.785 212.420 ;
      LAYER li1 ;
        RECT 786.955 211.770 787.285 212.250 ;
      LAYER li1 ;
        RECT 787.455 211.940 787.625 212.420 ;
      LAYER li1 ;
        RECT 787.795 211.770 788.125 212.570 ;
        RECT 788.685 211.770 788.975 212.495 ;
        RECT 789.535 211.770 789.865 212.570 ;
        RECT 792.985 212.420 794.405 212.590 ;
        RECT 790.375 211.770 790.705 212.250 ;
        RECT 791.215 211.770 791.545 212.250 ;
        RECT 792.055 211.770 792.385 212.250 ;
        RECT 792.895 211.770 793.225 212.250 ;
        RECT 793.395 211.945 793.565 212.420 ;
        RECT 793.735 211.770 794.065 212.250 ;
        RECT 794.235 211.940 794.405 212.420 ;
        RECT 794.665 211.770 794.955 212.495 ;
        RECT 2146.085 211.770 2146.375 212.495 ;
        RECT 2152.065 211.770 2152.355 212.495 ;
        RECT 2152.615 212.420 2154.035 212.590 ;
        RECT 2152.615 211.940 2152.785 212.420 ;
        RECT 2152.955 211.770 2153.285 212.250 ;
        RECT 2153.455 211.945 2153.625 212.420 ;
        RECT 2153.795 211.770 2154.125 212.250 ;
        RECT 2154.635 211.770 2154.965 212.250 ;
        RECT 2155.475 211.770 2155.805 212.250 ;
        RECT 2156.315 211.770 2156.645 212.250 ;
        RECT 2157.155 211.770 2157.485 212.570 ;
        RECT 2158.045 211.770 2158.335 212.495 ;
        RECT 2158.595 212.420 2160.015 212.590 ;
        RECT 2158.595 211.940 2158.765 212.420 ;
        RECT 2158.935 211.770 2159.265 212.250 ;
        RECT 2159.435 211.945 2159.605 212.420 ;
        RECT 2159.775 211.770 2160.105 212.250 ;
        RECT 2160.615 211.770 2160.945 212.250 ;
        RECT 2161.455 211.770 2161.785 212.250 ;
        RECT 2162.295 211.770 2162.625 212.250 ;
        RECT 2163.135 211.770 2163.465 212.570 ;
        RECT 2164.025 211.770 2164.315 212.495 ;
        RECT 2164.575 212.420 2165.995 212.590 ;
        RECT 2164.575 211.940 2164.745 212.420 ;
        RECT 2164.915 211.770 2165.245 212.250 ;
        RECT 2165.415 211.945 2165.585 212.420 ;
        RECT 2165.755 211.770 2166.085 212.250 ;
        RECT 2166.595 211.770 2166.925 212.250 ;
        RECT 2167.435 211.770 2167.765 212.250 ;
        RECT 2168.275 211.770 2168.605 212.250 ;
        RECT 2169.115 211.770 2169.445 212.570 ;
        RECT 2170.005 211.770 2170.295 212.495 ;
        RECT 2170.555 212.420 2171.975 212.590 ;
        RECT 2170.555 211.940 2170.725 212.420 ;
        RECT 2170.895 211.770 2171.225 212.250 ;
        RECT 2171.395 211.945 2171.565 212.420 ;
        RECT 2171.735 211.770 2172.065 212.250 ;
        RECT 2172.575 211.770 2172.905 212.250 ;
        RECT 2173.415 211.770 2173.745 212.250 ;
        RECT 2174.255 211.770 2174.585 212.250 ;
        RECT 2175.095 211.770 2175.425 212.570 ;
        RECT 2175.985 211.770 2176.275 212.495 ;
        RECT 2176.535 212.420 2177.955 212.590 ;
        RECT 2176.535 211.940 2176.705 212.420 ;
        RECT 2176.875 211.770 2177.205 212.250 ;
        RECT 2177.375 211.945 2177.545 212.420 ;
        RECT 2177.715 211.770 2178.045 212.250 ;
        RECT 2178.555 211.770 2178.885 212.250 ;
        RECT 2179.395 211.770 2179.725 212.250 ;
        RECT 2180.235 211.770 2180.565 212.250 ;
        RECT 2181.075 211.770 2181.405 212.570 ;
        RECT 2181.965 211.770 2182.255 212.495 ;
        RECT 2182.515 212.420 2183.935 212.590 ;
        RECT 2182.515 211.940 2182.685 212.420 ;
        RECT 2182.855 211.770 2183.185 212.250 ;
        RECT 2183.355 211.945 2183.525 212.420 ;
        RECT 2183.695 211.770 2184.025 212.250 ;
        RECT 2184.535 211.770 2184.865 212.250 ;
        RECT 2185.375 211.770 2185.705 212.250 ;
        RECT 2186.215 211.770 2186.545 212.250 ;
        RECT 2187.055 211.770 2187.385 212.570 ;
        RECT 2187.945 211.770 2188.235 212.495 ;
        RECT 2188.495 212.420 2189.915 212.590 ;
        RECT 2188.495 211.940 2188.665 212.420 ;
        RECT 2188.835 211.770 2189.165 212.250 ;
        RECT 2189.335 211.945 2189.505 212.420 ;
        RECT 2189.675 211.770 2190.005 212.250 ;
        RECT 2190.515 211.770 2190.845 212.250 ;
        RECT 2191.355 211.770 2191.685 212.250 ;
        RECT 2192.195 211.770 2192.525 212.250 ;
        RECT 2193.035 211.770 2193.365 212.570 ;
        RECT 2193.925 211.770 2194.215 212.495 ;
        RECT 2194.475 212.420 2195.895 212.590 ;
        RECT 2194.475 211.940 2194.645 212.420 ;
        RECT 2194.815 211.770 2195.145 212.250 ;
        RECT 2195.315 211.945 2195.485 212.420 ;
        RECT 2195.655 211.770 2195.985 212.250 ;
        RECT 2196.495 211.770 2196.825 212.250 ;
        RECT 2197.335 211.770 2197.665 212.250 ;
        RECT 2198.175 211.770 2198.505 212.250 ;
        RECT 2199.015 211.770 2199.345 212.570 ;
        RECT 2199.905 211.770 2200.195 212.495 ;
        RECT 2200.455 212.420 2201.875 212.590 ;
        RECT 2200.455 211.940 2200.625 212.420 ;
        RECT 2200.795 211.770 2201.125 212.250 ;
        RECT 2201.295 211.945 2201.465 212.420 ;
        RECT 2201.635 211.770 2201.965 212.250 ;
        RECT 2202.475 211.770 2202.805 212.250 ;
        RECT 2203.315 211.770 2203.645 212.250 ;
        RECT 2204.155 211.770 2204.485 212.250 ;
        RECT 2204.995 211.770 2205.325 212.570 ;
        RECT 2205.885 211.770 2206.175 212.495 ;
        RECT 2235.785 211.770 2236.075 212.495 ;
        RECT 2241.765 211.770 2242.055 212.495 ;
        RECT 2242.315 212.420 2243.735 212.590 ;
        RECT 2242.315 211.940 2242.485 212.420 ;
        RECT 2242.655 211.770 2242.985 212.250 ;
        RECT 2243.155 211.945 2243.325 212.420 ;
        RECT 2243.495 211.770 2243.825 212.250 ;
        RECT 2244.335 211.770 2244.665 212.250 ;
        RECT 2245.175 211.770 2245.505 212.250 ;
        RECT 2246.015 211.770 2246.345 212.250 ;
        RECT 2246.855 211.770 2247.185 212.570 ;
        RECT 2247.745 211.770 2248.035 212.495 ;
        RECT 2248.295 212.420 2249.715 212.590 ;
        RECT 2248.295 211.940 2248.465 212.420 ;
        RECT 2248.635 211.770 2248.965 212.250 ;
        RECT 2249.135 211.945 2249.305 212.420 ;
        RECT 2249.475 211.770 2249.805 212.250 ;
        RECT 2250.315 211.770 2250.645 212.250 ;
        RECT 2251.155 211.770 2251.485 212.250 ;
        RECT 2251.995 211.770 2252.325 212.250 ;
        RECT 2252.835 211.770 2253.165 212.570 ;
        RECT 2253.725 211.770 2254.015 212.495 ;
        RECT 2254.275 212.420 2255.695 212.590 ;
        RECT 2254.275 211.940 2254.445 212.420 ;
        RECT 2254.615 211.770 2254.945 212.250 ;
        RECT 2255.115 211.945 2255.285 212.420 ;
        RECT 2255.455 211.770 2255.785 212.250 ;
        RECT 2256.295 211.770 2256.625 212.250 ;
        RECT 2257.135 211.770 2257.465 212.250 ;
        RECT 2257.975 211.770 2258.305 212.250 ;
        RECT 2258.815 211.770 2259.145 212.570 ;
        RECT 2259.705 211.770 2259.995 212.495 ;
        RECT 2260.255 212.420 2261.675 212.590 ;
      LAYER li1 ;
        RECT 2267.035 212.590 2267.290 213.130 ;
      LAYER li1 ;
        RECT 2269.985 212.930 2270.160 213.130 ;
        RECT 2267.535 212.760 2270.160 212.930 ;
        RECT 2269.985 212.590 2270.160 212.760 ;
        RECT 2260.255 211.940 2260.425 212.420 ;
        RECT 2260.595 211.770 2260.925 212.250 ;
        RECT 2261.095 211.945 2261.265 212.420 ;
        RECT 2261.435 211.770 2261.765 212.250 ;
        RECT 2262.275 211.770 2262.605 212.250 ;
        RECT 2263.115 211.770 2263.445 212.250 ;
        RECT 2263.955 211.770 2264.285 212.250 ;
        RECT 2264.795 211.770 2265.125 212.570 ;
        RECT 2265.685 211.770 2265.975 212.495 ;
        RECT 2266.535 211.770 2266.865 212.570 ;
      LAYER li1 ;
        RECT 2267.035 212.420 2269.725 212.590 ;
      LAYER li1 ;
        RECT 2269.985 212.420 2271.405 212.590 ;
      LAYER li1 ;
        RECT 2267.035 211.940 2267.205 212.420 ;
      LAYER li1 ;
        RECT 2267.375 211.770 2267.705 212.250 ;
      LAYER li1 ;
        RECT 2267.875 211.940 2268.045 212.420 ;
      LAYER li1 ;
        RECT 2268.215 211.770 2268.545 212.250 ;
      LAYER li1 ;
        RECT 2268.715 211.940 2268.885 212.420 ;
      LAYER li1 ;
        RECT 2269.055 211.770 2269.385 212.250 ;
      LAYER li1 ;
        RECT 2269.555 211.940 2269.725 212.420 ;
      LAYER li1 ;
        RECT 2269.895 211.770 2270.225 212.250 ;
        RECT 2270.395 211.945 2270.565 212.420 ;
        RECT 2270.735 211.770 2271.065 212.250 ;
        RECT 2271.235 211.940 2271.405 212.420 ;
        RECT 2271.665 211.770 2271.955 212.495 ;
        RECT 669.000 211.600 669.145 211.770 ;
        RECT 669.315 211.600 669.460 211.770 ;
        RECT 674.980 211.600 675.125 211.770 ;
        RECT 675.295 211.600 675.585 211.770 ;
        RECT 675.755 211.600 676.045 211.770 ;
        RECT 676.215 211.600 676.505 211.770 ;
        RECT 676.675 211.600 676.965 211.770 ;
        RECT 677.135 211.600 677.425 211.770 ;
        RECT 677.595 211.600 677.885 211.770 ;
        RECT 678.055 211.600 678.345 211.770 ;
        RECT 678.515 211.600 678.805 211.770 ;
        RECT 678.975 211.600 679.265 211.770 ;
        RECT 679.435 211.600 679.725 211.770 ;
        RECT 679.895 211.600 680.185 211.770 ;
        RECT 680.355 211.600 680.645 211.770 ;
        RECT 680.815 211.600 681.105 211.770 ;
        RECT 681.275 211.600 681.565 211.770 ;
        RECT 681.735 211.600 682.025 211.770 ;
        RECT 682.195 211.600 682.485 211.770 ;
        RECT 682.655 211.600 682.945 211.770 ;
        RECT 683.115 211.600 683.405 211.770 ;
        RECT 683.575 211.600 683.865 211.770 ;
        RECT 684.035 211.600 684.325 211.770 ;
        RECT 684.495 211.600 684.785 211.770 ;
        RECT 684.955 211.600 685.245 211.770 ;
        RECT 685.415 211.600 685.705 211.770 ;
        RECT 685.875 211.600 686.165 211.770 ;
        RECT 686.335 211.600 686.625 211.770 ;
        RECT 686.795 211.600 687.085 211.770 ;
        RECT 687.255 211.600 687.545 211.770 ;
        RECT 687.715 211.600 688.005 211.770 ;
        RECT 688.175 211.600 688.465 211.770 ;
        RECT 688.635 211.600 688.925 211.770 ;
        RECT 689.095 211.600 689.385 211.770 ;
        RECT 689.555 211.600 689.845 211.770 ;
        RECT 690.015 211.600 690.305 211.770 ;
        RECT 690.475 211.600 690.765 211.770 ;
        RECT 690.935 211.600 691.225 211.770 ;
        RECT 691.395 211.600 691.685 211.770 ;
        RECT 691.855 211.600 692.145 211.770 ;
        RECT 692.315 211.600 692.605 211.770 ;
        RECT 692.775 211.600 693.065 211.770 ;
        RECT 693.235 211.600 693.525 211.770 ;
        RECT 693.695 211.600 693.985 211.770 ;
        RECT 694.155 211.600 694.445 211.770 ;
        RECT 694.615 211.600 694.905 211.770 ;
        RECT 695.075 211.600 695.365 211.770 ;
        RECT 695.535 211.600 695.825 211.770 ;
        RECT 695.995 211.600 696.285 211.770 ;
        RECT 696.455 211.600 696.745 211.770 ;
        RECT 696.915 211.600 697.205 211.770 ;
        RECT 697.375 211.600 697.665 211.770 ;
        RECT 697.835 211.600 698.125 211.770 ;
        RECT 698.295 211.600 698.585 211.770 ;
        RECT 698.755 211.600 699.045 211.770 ;
        RECT 699.215 211.600 699.505 211.770 ;
        RECT 699.675 211.600 699.965 211.770 ;
        RECT 700.135 211.600 700.425 211.770 ;
        RECT 700.595 211.600 700.885 211.770 ;
        RECT 701.055 211.600 701.345 211.770 ;
        RECT 701.515 211.600 701.805 211.770 ;
        RECT 701.975 211.600 702.265 211.770 ;
        RECT 702.435 211.600 702.725 211.770 ;
        RECT 702.895 211.600 703.185 211.770 ;
        RECT 703.355 211.600 703.645 211.770 ;
        RECT 703.815 211.600 704.105 211.770 ;
        RECT 704.275 211.600 704.565 211.770 ;
        RECT 704.735 211.600 705.025 211.770 ;
        RECT 705.195 211.600 705.485 211.770 ;
        RECT 705.655 211.600 705.945 211.770 ;
        RECT 706.115 211.600 706.405 211.770 ;
        RECT 706.575 211.600 706.865 211.770 ;
        RECT 707.035 211.600 707.325 211.770 ;
        RECT 707.495 211.600 707.785 211.770 ;
        RECT 707.955 211.600 708.245 211.770 ;
        RECT 708.415 211.600 708.705 211.770 ;
        RECT 708.875 211.600 709.165 211.770 ;
        RECT 709.335 211.600 709.625 211.770 ;
        RECT 709.795 211.600 710.085 211.770 ;
        RECT 710.255 211.600 710.545 211.770 ;
        RECT 710.715 211.600 711.005 211.770 ;
        RECT 711.175 211.600 711.465 211.770 ;
        RECT 711.635 211.600 711.925 211.770 ;
        RECT 712.095 211.600 712.385 211.770 ;
        RECT 712.555 211.600 712.845 211.770 ;
        RECT 713.015 211.600 713.305 211.770 ;
        RECT 713.475 211.600 713.765 211.770 ;
        RECT 713.935 211.600 714.225 211.770 ;
        RECT 714.395 211.600 714.685 211.770 ;
        RECT 714.855 211.600 715.145 211.770 ;
        RECT 715.315 211.600 715.605 211.770 ;
        RECT 715.775 211.600 716.065 211.770 ;
        RECT 716.235 211.600 716.525 211.770 ;
        RECT 716.695 211.600 716.985 211.770 ;
        RECT 717.155 211.600 717.445 211.770 ;
        RECT 717.615 211.600 717.905 211.770 ;
        RECT 718.075 211.600 718.365 211.770 ;
        RECT 718.535 211.600 718.825 211.770 ;
        RECT 718.995 211.600 719.285 211.770 ;
        RECT 719.455 211.600 719.745 211.770 ;
        RECT 719.915 211.600 720.205 211.770 ;
        RECT 720.375 211.600 720.665 211.770 ;
        RECT 720.835 211.600 721.125 211.770 ;
        RECT 721.295 211.600 721.585 211.770 ;
        RECT 721.755 211.600 722.045 211.770 ;
        RECT 722.215 211.600 722.505 211.770 ;
        RECT 722.675 211.600 722.965 211.770 ;
        RECT 723.135 211.600 723.425 211.770 ;
        RECT 723.595 211.600 723.885 211.770 ;
        RECT 724.055 211.600 724.345 211.770 ;
        RECT 724.515 211.600 724.805 211.770 ;
        RECT 724.975 211.600 725.265 211.770 ;
        RECT 725.435 211.600 725.725 211.770 ;
        RECT 725.895 211.600 726.185 211.770 ;
        RECT 726.355 211.600 726.645 211.770 ;
        RECT 726.815 211.600 727.105 211.770 ;
        RECT 727.275 211.600 727.565 211.770 ;
        RECT 727.735 211.600 728.025 211.770 ;
        RECT 728.195 211.600 728.485 211.770 ;
        RECT 728.655 211.600 728.945 211.770 ;
        RECT 729.115 211.600 729.260 211.770 ;
        RECT 758.700 211.600 758.845 211.770 ;
        RECT 759.015 211.600 759.160 211.770 ;
        RECT 764.680 211.600 764.825 211.770 ;
        RECT 764.995 211.600 765.285 211.770 ;
        RECT 765.455 211.600 765.745 211.770 ;
        RECT 765.915 211.600 766.205 211.770 ;
        RECT 766.375 211.600 766.665 211.770 ;
        RECT 766.835 211.600 767.125 211.770 ;
        RECT 767.295 211.600 767.585 211.770 ;
        RECT 767.755 211.600 768.045 211.770 ;
        RECT 768.215 211.600 768.505 211.770 ;
        RECT 768.675 211.600 768.965 211.770 ;
        RECT 769.135 211.600 769.425 211.770 ;
        RECT 769.595 211.600 769.885 211.770 ;
        RECT 770.055 211.600 770.345 211.770 ;
        RECT 770.515 211.600 770.805 211.770 ;
        RECT 770.975 211.600 771.265 211.770 ;
        RECT 771.435 211.600 771.725 211.770 ;
        RECT 771.895 211.600 772.185 211.770 ;
        RECT 772.355 211.600 772.645 211.770 ;
        RECT 772.815 211.600 773.105 211.770 ;
        RECT 773.275 211.600 773.565 211.770 ;
        RECT 773.735 211.600 774.025 211.770 ;
        RECT 774.195 211.600 774.485 211.770 ;
        RECT 774.655 211.600 774.945 211.770 ;
        RECT 775.115 211.600 775.405 211.770 ;
        RECT 775.575 211.600 775.865 211.770 ;
        RECT 776.035 211.600 776.325 211.770 ;
        RECT 776.495 211.600 776.785 211.770 ;
        RECT 776.955 211.600 777.245 211.770 ;
        RECT 777.415 211.600 777.705 211.770 ;
        RECT 777.875 211.600 778.165 211.770 ;
        RECT 778.335 211.600 778.625 211.770 ;
        RECT 778.795 211.600 779.085 211.770 ;
        RECT 779.255 211.600 779.545 211.770 ;
        RECT 779.715 211.600 780.005 211.770 ;
        RECT 780.175 211.600 780.465 211.770 ;
        RECT 780.635 211.600 780.925 211.770 ;
        RECT 781.095 211.600 781.385 211.770 ;
        RECT 781.555 211.600 781.845 211.770 ;
        RECT 782.015 211.600 782.305 211.770 ;
        RECT 782.475 211.600 782.765 211.770 ;
        RECT 782.935 211.600 783.225 211.770 ;
        RECT 783.395 211.600 783.685 211.770 ;
        RECT 783.855 211.600 784.145 211.770 ;
        RECT 784.315 211.600 784.605 211.770 ;
        RECT 784.775 211.600 785.065 211.770 ;
        RECT 785.235 211.600 785.525 211.770 ;
        RECT 785.695 211.600 785.985 211.770 ;
        RECT 786.155 211.600 786.445 211.770 ;
        RECT 786.615 211.600 786.905 211.770 ;
        RECT 787.075 211.600 787.365 211.770 ;
        RECT 787.535 211.600 787.825 211.770 ;
        RECT 787.995 211.600 788.285 211.770 ;
        RECT 788.455 211.600 788.745 211.770 ;
        RECT 788.915 211.600 789.205 211.770 ;
        RECT 789.375 211.600 789.665 211.770 ;
        RECT 789.835 211.600 790.125 211.770 ;
        RECT 790.295 211.600 790.585 211.770 ;
        RECT 790.755 211.600 791.045 211.770 ;
        RECT 791.215 211.600 791.505 211.770 ;
        RECT 791.675 211.600 791.965 211.770 ;
        RECT 792.135 211.600 792.425 211.770 ;
        RECT 792.595 211.600 792.885 211.770 ;
        RECT 793.055 211.600 793.345 211.770 ;
        RECT 793.515 211.600 793.805 211.770 ;
        RECT 793.975 211.600 794.265 211.770 ;
        RECT 794.435 211.600 794.725 211.770 ;
        RECT 794.895 211.600 795.040 211.770 ;
        RECT 2146.000 211.600 2146.145 211.770 ;
        RECT 2146.315 211.600 2146.460 211.770 ;
        RECT 2151.980 211.600 2152.125 211.770 ;
        RECT 2152.295 211.600 2152.585 211.770 ;
        RECT 2152.755 211.600 2153.045 211.770 ;
        RECT 2153.215 211.600 2153.505 211.770 ;
        RECT 2153.675 211.600 2153.965 211.770 ;
        RECT 2154.135 211.600 2154.425 211.770 ;
        RECT 2154.595 211.600 2154.885 211.770 ;
        RECT 2155.055 211.600 2155.345 211.770 ;
        RECT 2155.515 211.600 2155.805 211.770 ;
        RECT 2155.975 211.600 2156.265 211.770 ;
        RECT 2156.435 211.600 2156.725 211.770 ;
        RECT 2156.895 211.600 2157.185 211.770 ;
        RECT 2157.355 211.600 2157.645 211.770 ;
        RECT 2157.815 211.600 2158.105 211.770 ;
        RECT 2158.275 211.600 2158.565 211.770 ;
        RECT 2158.735 211.600 2159.025 211.770 ;
        RECT 2159.195 211.600 2159.485 211.770 ;
        RECT 2159.655 211.600 2159.945 211.770 ;
        RECT 2160.115 211.600 2160.405 211.770 ;
        RECT 2160.575 211.600 2160.865 211.770 ;
        RECT 2161.035 211.600 2161.325 211.770 ;
        RECT 2161.495 211.600 2161.785 211.770 ;
        RECT 2161.955 211.600 2162.245 211.770 ;
        RECT 2162.415 211.600 2162.705 211.770 ;
        RECT 2162.875 211.600 2163.165 211.770 ;
        RECT 2163.335 211.600 2163.625 211.770 ;
        RECT 2163.795 211.600 2164.085 211.770 ;
        RECT 2164.255 211.600 2164.545 211.770 ;
        RECT 2164.715 211.600 2165.005 211.770 ;
        RECT 2165.175 211.600 2165.465 211.770 ;
        RECT 2165.635 211.600 2165.925 211.770 ;
        RECT 2166.095 211.600 2166.385 211.770 ;
        RECT 2166.555 211.600 2166.845 211.770 ;
        RECT 2167.015 211.600 2167.305 211.770 ;
        RECT 2167.475 211.600 2167.765 211.770 ;
        RECT 2167.935 211.600 2168.225 211.770 ;
        RECT 2168.395 211.600 2168.685 211.770 ;
        RECT 2168.855 211.600 2169.145 211.770 ;
        RECT 2169.315 211.600 2169.605 211.770 ;
        RECT 2169.775 211.600 2170.065 211.770 ;
        RECT 2170.235 211.600 2170.525 211.770 ;
        RECT 2170.695 211.600 2170.985 211.770 ;
        RECT 2171.155 211.600 2171.445 211.770 ;
        RECT 2171.615 211.600 2171.905 211.770 ;
        RECT 2172.075 211.600 2172.365 211.770 ;
        RECT 2172.535 211.600 2172.825 211.770 ;
        RECT 2172.995 211.600 2173.285 211.770 ;
        RECT 2173.455 211.600 2173.745 211.770 ;
        RECT 2173.915 211.600 2174.205 211.770 ;
        RECT 2174.375 211.600 2174.665 211.770 ;
        RECT 2174.835 211.600 2175.125 211.770 ;
        RECT 2175.295 211.600 2175.585 211.770 ;
        RECT 2175.755 211.600 2176.045 211.770 ;
        RECT 2176.215 211.600 2176.505 211.770 ;
        RECT 2176.675 211.600 2176.965 211.770 ;
        RECT 2177.135 211.600 2177.425 211.770 ;
        RECT 2177.595 211.600 2177.885 211.770 ;
        RECT 2178.055 211.600 2178.345 211.770 ;
        RECT 2178.515 211.600 2178.805 211.770 ;
        RECT 2178.975 211.600 2179.265 211.770 ;
        RECT 2179.435 211.600 2179.725 211.770 ;
        RECT 2179.895 211.600 2180.185 211.770 ;
        RECT 2180.355 211.600 2180.645 211.770 ;
        RECT 2180.815 211.600 2181.105 211.770 ;
        RECT 2181.275 211.600 2181.565 211.770 ;
        RECT 2181.735 211.600 2182.025 211.770 ;
        RECT 2182.195 211.600 2182.485 211.770 ;
        RECT 2182.655 211.600 2182.945 211.770 ;
        RECT 2183.115 211.600 2183.405 211.770 ;
        RECT 2183.575 211.600 2183.865 211.770 ;
        RECT 2184.035 211.600 2184.325 211.770 ;
        RECT 2184.495 211.600 2184.785 211.770 ;
        RECT 2184.955 211.600 2185.245 211.770 ;
        RECT 2185.415 211.600 2185.705 211.770 ;
        RECT 2185.875 211.600 2186.165 211.770 ;
        RECT 2186.335 211.600 2186.625 211.770 ;
        RECT 2186.795 211.600 2187.085 211.770 ;
        RECT 2187.255 211.600 2187.545 211.770 ;
        RECT 2187.715 211.600 2188.005 211.770 ;
        RECT 2188.175 211.600 2188.465 211.770 ;
        RECT 2188.635 211.600 2188.925 211.770 ;
        RECT 2189.095 211.600 2189.385 211.770 ;
        RECT 2189.555 211.600 2189.845 211.770 ;
        RECT 2190.015 211.600 2190.305 211.770 ;
        RECT 2190.475 211.600 2190.765 211.770 ;
        RECT 2190.935 211.600 2191.225 211.770 ;
        RECT 2191.395 211.600 2191.685 211.770 ;
        RECT 2191.855 211.600 2192.145 211.770 ;
        RECT 2192.315 211.600 2192.605 211.770 ;
        RECT 2192.775 211.600 2193.065 211.770 ;
        RECT 2193.235 211.600 2193.525 211.770 ;
        RECT 2193.695 211.600 2193.985 211.770 ;
        RECT 2194.155 211.600 2194.445 211.770 ;
        RECT 2194.615 211.600 2194.905 211.770 ;
        RECT 2195.075 211.600 2195.365 211.770 ;
        RECT 2195.535 211.600 2195.825 211.770 ;
        RECT 2195.995 211.600 2196.285 211.770 ;
        RECT 2196.455 211.600 2196.745 211.770 ;
        RECT 2196.915 211.600 2197.205 211.770 ;
        RECT 2197.375 211.600 2197.665 211.770 ;
        RECT 2197.835 211.600 2198.125 211.770 ;
        RECT 2198.295 211.600 2198.585 211.770 ;
        RECT 2198.755 211.600 2199.045 211.770 ;
        RECT 2199.215 211.600 2199.505 211.770 ;
        RECT 2199.675 211.600 2199.965 211.770 ;
        RECT 2200.135 211.600 2200.425 211.770 ;
        RECT 2200.595 211.600 2200.885 211.770 ;
        RECT 2201.055 211.600 2201.345 211.770 ;
        RECT 2201.515 211.600 2201.805 211.770 ;
        RECT 2201.975 211.600 2202.265 211.770 ;
        RECT 2202.435 211.600 2202.725 211.770 ;
        RECT 2202.895 211.600 2203.185 211.770 ;
        RECT 2203.355 211.600 2203.645 211.770 ;
        RECT 2203.815 211.600 2204.105 211.770 ;
        RECT 2204.275 211.600 2204.565 211.770 ;
        RECT 2204.735 211.600 2205.025 211.770 ;
        RECT 2205.195 211.600 2205.485 211.770 ;
        RECT 2205.655 211.600 2205.945 211.770 ;
        RECT 2206.115 211.600 2206.260 211.770 ;
        RECT 2235.700 211.600 2235.845 211.770 ;
        RECT 2236.015 211.600 2236.160 211.770 ;
        RECT 2241.680 211.600 2241.825 211.770 ;
        RECT 2241.995 211.600 2242.285 211.770 ;
        RECT 2242.455 211.600 2242.745 211.770 ;
        RECT 2242.915 211.600 2243.205 211.770 ;
        RECT 2243.375 211.600 2243.665 211.770 ;
        RECT 2243.835 211.600 2244.125 211.770 ;
        RECT 2244.295 211.600 2244.585 211.770 ;
        RECT 2244.755 211.600 2245.045 211.770 ;
        RECT 2245.215 211.600 2245.505 211.770 ;
        RECT 2245.675 211.600 2245.965 211.770 ;
        RECT 2246.135 211.600 2246.425 211.770 ;
        RECT 2246.595 211.600 2246.885 211.770 ;
        RECT 2247.055 211.600 2247.345 211.770 ;
        RECT 2247.515 211.600 2247.805 211.770 ;
        RECT 2247.975 211.600 2248.265 211.770 ;
        RECT 2248.435 211.600 2248.725 211.770 ;
        RECT 2248.895 211.600 2249.185 211.770 ;
        RECT 2249.355 211.600 2249.645 211.770 ;
        RECT 2249.815 211.600 2250.105 211.770 ;
        RECT 2250.275 211.600 2250.565 211.770 ;
        RECT 2250.735 211.600 2251.025 211.770 ;
        RECT 2251.195 211.600 2251.485 211.770 ;
        RECT 2251.655 211.600 2251.945 211.770 ;
        RECT 2252.115 211.600 2252.405 211.770 ;
        RECT 2252.575 211.600 2252.865 211.770 ;
        RECT 2253.035 211.600 2253.325 211.770 ;
        RECT 2253.495 211.600 2253.785 211.770 ;
        RECT 2253.955 211.600 2254.245 211.770 ;
        RECT 2254.415 211.600 2254.705 211.770 ;
        RECT 2254.875 211.600 2255.165 211.770 ;
        RECT 2255.335 211.600 2255.625 211.770 ;
        RECT 2255.795 211.600 2256.085 211.770 ;
        RECT 2256.255 211.600 2256.545 211.770 ;
        RECT 2256.715 211.600 2257.005 211.770 ;
        RECT 2257.175 211.600 2257.465 211.770 ;
        RECT 2257.635 211.600 2257.925 211.770 ;
        RECT 2258.095 211.600 2258.385 211.770 ;
        RECT 2258.555 211.600 2258.845 211.770 ;
        RECT 2259.015 211.600 2259.305 211.770 ;
        RECT 2259.475 211.600 2259.765 211.770 ;
        RECT 2259.935 211.600 2260.225 211.770 ;
        RECT 2260.395 211.600 2260.685 211.770 ;
        RECT 2260.855 211.600 2261.145 211.770 ;
        RECT 2261.315 211.600 2261.605 211.770 ;
        RECT 2261.775 211.600 2262.065 211.770 ;
        RECT 2262.235 211.600 2262.525 211.770 ;
        RECT 2262.695 211.600 2262.985 211.770 ;
        RECT 2263.155 211.600 2263.445 211.770 ;
        RECT 2263.615 211.600 2263.905 211.770 ;
        RECT 2264.075 211.600 2264.365 211.770 ;
        RECT 2264.535 211.600 2264.825 211.770 ;
        RECT 2264.995 211.600 2265.285 211.770 ;
        RECT 2265.455 211.600 2265.745 211.770 ;
        RECT 2265.915 211.600 2266.205 211.770 ;
        RECT 2266.375 211.600 2266.665 211.770 ;
        RECT 2266.835 211.600 2267.125 211.770 ;
        RECT 2267.295 211.600 2267.585 211.770 ;
        RECT 2267.755 211.600 2268.045 211.770 ;
        RECT 2268.215 211.600 2268.505 211.770 ;
        RECT 2268.675 211.600 2268.965 211.770 ;
        RECT 2269.135 211.600 2269.425 211.770 ;
        RECT 2269.595 211.600 2269.885 211.770 ;
        RECT 2270.055 211.600 2270.345 211.770 ;
        RECT 2270.515 211.600 2270.805 211.770 ;
        RECT 2270.975 211.600 2271.265 211.770 ;
        RECT 2271.435 211.600 2271.725 211.770 ;
        RECT 2271.895 211.600 2272.040 211.770 ;
      LAYER mcon ;
        RECT 3381.350 3603.580 3382.200 3603.750 ;
        RECT 3384.750 3602.670 3384.920 3603.760 ;
        RECT 203.075 3009.260 203.245 3010.350 ;
        RECT 205.795 3010.170 206.645 3010.340 ;
        RECT 203.075 3003.280 203.245 3004.370 ;
        RECT 205.795 3004.190 206.645 3004.360 ;
        RECT 203.075 2997.300 203.245 2998.390 ;
        RECT 205.795 2998.210 206.645 2998.380 ;
        RECT 203.075 2991.320 203.245 2992.410 ;
        RECT 205.795 2992.230 206.645 2992.400 ;
        RECT 203.075 2985.340 203.245 2986.430 ;
        RECT 205.795 2986.250 206.645 2986.420 ;
        RECT 3381.690 2237.180 3381.860 2238.270 ;
        RECT 202.845 1725.495 203.695 1725.665 ;
        RECT 206.245 1725.985 206.415 1727.075 ;
        RECT 203.185 1721.355 203.355 1722.445 ;
        RECT 205.905 1722.265 206.755 1722.435 ;
        RECT 202.845 1719.515 203.695 1719.685 ;
        RECT 206.245 1720.005 206.415 1721.095 ;
        RECT 203.185 1715.375 203.355 1716.465 ;
        RECT 205.905 1716.285 206.755 1716.455 ;
        RECT 202.845 1713.535 203.695 1713.705 ;
        RECT 206.245 1714.025 206.415 1715.115 ;
        RECT 203.185 1709.395 203.355 1710.485 ;
        RECT 205.905 1710.305 206.755 1710.475 ;
        RECT 202.845 1707.555 203.695 1707.725 ;
        RECT 206.245 1708.045 206.415 1709.135 ;
        RECT 203.185 1703.415 203.355 1704.505 ;
        RECT 205.905 1704.325 206.755 1704.495 ;
        RECT 202.845 1701.575 203.695 1701.745 ;
        RECT 206.245 1702.065 206.415 1703.155 ;
        RECT 203.185 1697.435 203.355 1698.525 ;
        RECT 205.905 1698.345 206.755 1698.515 ;
        RECT 203.185 1691.455 203.355 1692.545 ;
        RECT 205.905 1692.365 206.755 1692.535 ;
        RECT 203.185 1685.475 203.355 1686.565 ;
        RECT 205.905 1686.385 206.755 1686.555 ;
        RECT 203.185 1679.495 203.355 1680.585 ;
        RECT 205.905 1680.405 206.755 1680.575 ;
        RECT 203.185 1673.515 203.355 1674.605 ;
        RECT 205.905 1674.425 206.755 1674.595 ;
        RECT 670.520 215.510 670.690 216.360 ;
        RECT 674.240 215.850 675.330 216.020 ;
        RECT 676.500 215.510 676.670 216.360 ;
        RECT 680.220 215.850 681.310 216.020 ;
        RECT 682.480 215.510 682.650 216.360 ;
        RECT 686.200 215.850 687.290 216.020 ;
        RECT 688.460 215.510 688.630 216.360 ;
        RECT 692.180 215.850 693.270 216.020 ;
        RECT 694.440 215.510 694.610 216.360 ;
        RECT 698.160 215.850 699.250 216.020 ;
        RECT 700.420 215.510 700.590 216.360 ;
        RECT 704.140 215.850 705.230 216.020 ;
        RECT 706.400 215.510 706.570 216.360 ;
        RECT 710.120 215.850 711.210 216.020 ;
        RECT 712.380 215.510 712.550 216.360 ;
        RECT 716.100 215.850 717.190 216.020 ;
        RECT 718.360 215.510 718.530 216.360 ;
        RECT 722.080 215.850 723.170 216.020 ;
        RECT 763.940 215.850 765.030 216.020 ;
        RECT 769.920 215.850 771.010 216.020 ;
        RECT 775.900 215.850 776.990 216.020 ;
        RECT 781.880 215.850 782.970 216.020 ;
        RECT 787.860 215.850 788.950 216.020 ;
        RECT 793.840 215.850 794.930 216.020 ;
        RECT 2147.520 215.510 2147.690 216.360 ;
        RECT 2153.500 215.510 2153.670 216.360 ;
        RECT 2159.480 215.510 2159.650 216.360 ;
        RECT 2165.460 215.510 2165.630 216.360 ;
        RECT 2171.440 215.510 2171.610 216.360 ;
        RECT 2177.420 215.510 2177.590 216.360 ;
        RECT 2183.400 215.510 2183.570 216.360 ;
        RECT 2189.380 215.510 2189.550 216.360 ;
        RECT 2195.360 215.510 2195.530 216.360 ;
        RECT 2237.220 215.510 2237.390 216.360 ;
        RECT 2243.200 215.510 2243.370 216.360 ;
        RECT 2249.180 215.510 2249.350 216.360 ;
        RECT 2255.160 215.510 2255.330 216.360 ;
        RECT 2261.140 215.510 2261.310 216.360 ;
        RECT 2267.120 215.510 2267.290 216.360 ;
        RECT 675.590 212.790 676.680 212.960 ;
        RECT 679.730 212.450 679.900 213.300 ;
        RECT 681.570 212.790 682.660 212.960 ;
        RECT 685.710 212.450 685.880 213.300 ;
        RECT 687.550 212.790 688.640 212.960 ;
        RECT 691.690 212.450 691.860 213.300 ;
        RECT 693.530 212.790 694.620 212.960 ;
        RECT 697.670 212.450 697.840 213.300 ;
        RECT 699.510 212.790 700.600 212.960 ;
        RECT 703.650 212.450 703.820 213.300 ;
        RECT 705.490 212.790 706.580 212.960 ;
        RECT 709.630 212.450 709.800 213.300 ;
        RECT 711.470 212.790 712.560 212.960 ;
        RECT 715.610 212.450 715.780 213.300 ;
        RECT 717.450 212.790 718.540 212.960 ;
        RECT 721.590 212.450 721.760 213.300 ;
        RECT 723.430 212.790 724.520 212.960 ;
        RECT 727.570 212.450 727.740 213.300 ;
        RECT 769.430 212.450 769.600 213.300 ;
        RECT 775.410 212.450 775.580 213.300 ;
        RECT 781.390 212.450 781.560 213.300 ;
        RECT 787.370 212.450 787.540 213.300 ;
        RECT 793.340 212.790 794.430 212.960 ;
        RECT 2152.590 212.790 2153.680 212.960 ;
        RECT 2158.570 212.790 2159.660 212.960 ;
        RECT 2164.550 212.790 2165.640 212.960 ;
        RECT 2170.530 212.790 2171.620 212.960 ;
        RECT 2176.510 212.790 2177.600 212.960 ;
        RECT 2182.490 212.790 2183.580 212.960 ;
        RECT 2188.470 212.790 2189.560 212.960 ;
        RECT 2194.450 212.790 2195.540 212.960 ;
        RECT 2200.430 212.790 2201.520 212.960 ;
        RECT 2242.290 212.790 2243.380 212.960 ;
        RECT 2248.270 212.790 2249.360 212.960 ;
        RECT 2254.250 212.790 2255.340 212.960 ;
        RECT 2260.230 212.790 2261.320 212.960 ;
        RECT 2267.120 212.450 2267.290 213.300 ;
      LAYER met1 ;
        RECT 3370.800 3603.550 3371.060 3603.870 ;
        RECT 3370.640 3603.250 3370.780 3603.275 ;
        RECT 3370.520 3602.930 3370.780 3603.250 ;
        RECT 203.035 3009.200 203.295 3010.410 ;
        RECT 205.735 3010.120 206.705 3010.380 ;
        RECT 217.615 3010.140 217.875 3010.460 ;
        RECT 203.035 3003.220 203.295 3004.430 ;
        RECT 205.735 3004.140 206.705 3004.400 ;
        RECT 203.035 2997.240 203.295 2998.450 ;
        RECT 205.735 2998.160 206.705 2998.420 ;
        RECT 203.035 2991.260 203.295 2992.470 ;
        RECT 205.735 2992.180 206.705 2992.440 ;
        RECT 203.035 2985.280 203.295 2986.490 ;
        RECT 205.735 2986.200 206.705 2986.460 ;
        RECT 206.205 1725.925 206.465 1727.135 ;
        RECT 217.615 1726.770 217.755 3010.140 ;
        RECT 217.495 1726.450 217.755 1726.770 ;
        RECT 217.895 3009.520 218.155 3009.840 ;
        RECT 217.895 1725.800 218.035 3009.520 ;
        RECT 202.785 1725.445 203.755 1725.705 ;
        RECT 217.775 1725.480 218.035 1725.800 ;
        RECT 218.735 3004.160 218.995 3004.480 ;
        RECT 203.145 1721.295 203.405 1722.505 ;
        RECT 205.845 1722.215 206.815 1722.475 ;
        RECT 217.475 1722.235 217.735 1722.555 ;
        RECT 206.205 1719.945 206.465 1721.155 ;
        RECT 202.785 1719.465 203.755 1719.725 ;
        RECT 203.145 1715.315 203.405 1716.525 ;
        RECT 205.845 1716.235 206.815 1716.495 ;
        RECT 206.205 1713.965 206.465 1715.175 ;
        RECT 202.785 1713.485 203.755 1713.745 ;
        RECT 203.145 1709.335 203.405 1710.545 ;
        RECT 205.845 1710.255 206.815 1710.515 ;
        RECT 206.205 1707.985 206.465 1709.195 ;
        RECT 202.785 1707.505 203.755 1707.765 ;
        RECT 203.145 1703.355 203.405 1704.565 ;
        RECT 205.845 1704.275 206.815 1704.535 ;
        RECT 206.205 1702.005 206.465 1703.215 ;
        RECT 202.785 1701.525 203.755 1701.785 ;
        RECT 203.145 1697.375 203.405 1698.585 ;
        RECT 205.845 1698.295 206.815 1698.555 ;
        RECT 203.145 1691.395 203.405 1692.605 ;
        RECT 205.845 1692.315 206.815 1692.575 ;
        RECT 203.145 1685.415 203.405 1686.625 ;
        RECT 205.845 1686.335 206.815 1686.595 ;
        RECT 203.145 1679.435 203.405 1680.645 ;
        RECT 205.845 1680.355 206.815 1680.615 ;
        RECT 203.145 1673.455 203.405 1674.665 ;
        RECT 205.845 1674.375 206.815 1674.635 ;
        RECT 217.475 230.980 217.615 1722.235 ;
        RECT 217.755 1721.615 218.015 1721.935 ;
        RECT 217.755 231.260 217.895 1721.615 ;
        RECT 218.735 1720.790 218.875 3004.160 ;
        RECT 218.615 1720.470 218.875 1720.790 ;
        RECT 219.015 3003.540 219.275 3003.860 ;
        RECT 219.015 1719.820 219.155 3003.540 ;
        RECT 218.895 1719.500 219.155 1719.820 ;
        RECT 219.855 2998.180 220.115 2998.500 ;
        RECT 218.595 1716.255 218.855 1716.575 ;
        RECT 218.595 231.820 218.735 1716.255 ;
        RECT 218.875 1715.635 219.135 1715.955 ;
        RECT 218.875 232.100 219.015 1715.635 ;
        RECT 219.855 1714.810 219.995 2998.180 ;
        RECT 219.735 1714.490 219.995 1714.810 ;
        RECT 220.135 2997.560 220.395 2997.880 ;
        RECT 220.135 1713.840 220.275 2997.560 ;
        RECT 220.015 1713.520 220.275 1713.840 ;
        RECT 220.975 2992.200 221.235 2992.520 ;
        RECT 219.715 1710.275 219.975 1710.595 ;
        RECT 219.715 232.660 219.855 1710.275 ;
        RECT 219.995 1709.655 220.255 1709.975 ;
        RECT 219.995 232.940 220.135 1709.655 ;
        RECT 220.975 1708.830 221.115 2992.200 ;
        RECT 220.855 1708.510 221.115 1708.830 ;
        RECT 221.255 2991.580 221.515 2991.900 ;
        RECT 221.255 1707.860 221.395 2991.580 ;
        RECT 221.135 1707.540 221.395 1707.860 ;
        RECT 222.095 2986.220 222.355 2986.540 ;
        RECT 220.835 1704.295 221.095 1704.615 ;
        RECT 220.835 233.500 220.975 1704.295 ;
        RECT 221.115 1703.675 221.375 1703.995 ;
        RECT 221.115 233.780 221.255 1703.675 ;
        RECT 222.095 1702.850 222.235 2986.220 ;
        RECT 221.975 1702.530 222.235 1702.850 ;
        RECT 222.375 2985.600 222.635 2985.920 ;
        RECT 222.375 1701.880 222.515 2985.600 ;
        RECT 3370.640 2236.995 3370.780 3602.930 ;
        RECT 3370.920 2237.965 3371.060 3603.550 ;
        RECT 3381.290 3603.530 3382.260 3603.790 ;
        RECT 3384.700 3602.610 3384.960 3603.820 ;
        RECT 3370.920 2237.645 3371.180 2237.965 ;
        RECT 3381.640 2237.120 3381.900 2238.330 ;
        RECT 3370.640 2236.675 3370.900 2236.995 ;
        RECT 3384.350 2236.640 3385.320 2236.900 ;
        RECT 222.255 1701.560 222.515 1701.880 ;
        RECT 221.955 1698.315 222.215 1698.635 ;
        RECT 221.955 234.340 222.095 1698.315 ;
        RECT 222.235 1697.695 222.495 1698.015 ;
        RECT 222.235 234.620 222.375 1697.695 ;
        RECT 223.075 1692.335 223.335 1692.655 ;
        RECT 223.075 235.180 223.215 1692.335 ;
        RECT 223.355 1691.715 223.615 1692.035 ;
        RECT 223.355 235.460 223.495 1691.715 ;
        RECT 224.195 1686.355 224.455 1686.675 ;
        RECT 224.195 236.020 224.335 1686.355 ;
        RECT 224.475 1685.735 224.735 1686.055 ;
        RECT 224.475 236.300 224.615 1685.735 ;
        RECT 225.315 1680.375 225.575 1680.695 ;
        RECT 225.315 236.860 225.455 1680.375 ;
        RECT 225.595 1679.755 225.855 1680.075 ;
        RECT 225.595 237.140 225.735 1679.755 ;
        RECT 226.435 1674.395 226.695 1674.715 ;
        RECT 226.435 237.700 226.575 1674.395 ;
        RECT 226.715 1673.775 226.975 1674.095 ;
        RECT 226.715 237.980 226.855 1673.775 ;
        RECT 2147.490 238.120 2147.810 238.240 ;
        RECT 670.490 237.980 670.810 238.100 ;
        RECT 226.715 237.840 670.810 237.980 ;
        RECT 674.705 237.980 706.345 238.120 ;
        RECT 674.705 237.860 675.025 237.980 ;
        RECT 675.850 237.700 676.170 237.820 ;
        RECT 226.435 237.560 676.170 237.700 ;
        RECT 679.715 237.700 706.065 237.840 ;
        RECT 679.715 237.580 680.035 237.700 ;
        RECT 676.470 237.140 676.790 237.260 ;
        RECT 225.595 237.000 676.790 237.140 ;
        RECT 680.685 237.140 705.505 237.280 ;
        RECT 680.685 237.020 681.005 237.140 ;
        RECT 681.830 236.860 682.150 236.980 ;
        RECT 225.315 236.720 682.150 236.860 ;
        RECT 685.695 236.860 705.225 237.000 ;
        RECT 685.695 236.740 686.015 236.860 ;
        RECT 682.450 236.300 682.770 236.420 ;
        RECT 224.475 236.160 682.770 236.300 ;
        RECT 686.665 236.300 704.665 236.440 ;
        RECT 686.665 236.180 686.985 236.300 ;
        RECT 687.810 236.020 688.130 236.140 ;
        RECT 224.195 235.880 688.130 236.020 ;
        RECT 691.675 236.020 704.385 236.160 ;
        RECT 691.675 235.900 691.995 236.020 ;
        RECT 688.430 235.460 688.750 235.580 ;
        RECT 223.355 235.320 688.750 235.460 ;
        RECT 692.645 235.460 703.825 235.600 ;
        RECT 692.645 235.340 692.965 235.460 ;
        RECT 693.790 235.180 694.110 235.300 ;
        RECT 223.075 235.040 694.110 235.180 ;
        RECT 697.655 235.180 703.545 235.320 ;
        RECT 697.655 235.060 697.975 235.180 ;
        RECT 694.410 234.620 694.730 234.740 ;
        RECT 222.235 234.480 694.730 234.620 ;
        RECT 698.625 234.620 703.255 234.760 ;
        RECT 698.625 234.500 698.945 234.620 ;
        RECT 699.770 234.340 700.090 234.460 ;
        RECT 221.955 234.200 700.090 234.340 ;
        RECT 700.390 233.780 700.710 233.900 ;
        RECT 221.115 233.640 700.710 233.780 ;
        RECT 220.835 233.360 702.925 233.500 ;
        RECT 219.995 232.800 702.630 232.940 ;
        RECT 219.715 232.520 702.310 232.660 ;
        RECT 218.875 231.960 702.015 232.100 ;
        RECT 218.595 231.680 701.735 231.820 ;
        RECT 217.755 231.120 701.435 231.260 ;
        RECT 217.475 230.840 701.155 230.980 ;
        RECT 701.015 230.420 701.155 230.840 ;
        RECT 701.295 230.700 701.435 231.120 ;
        RECT 701.595 230.980 701.735 231.680 ;
        RECT 701.875 231.260 702.015 231.960 ;
        RECT 702.170 231.540 702.310 232.520 ;
        RECT 702.490 231.820 702.630 232.800 ;
        RECT 702.785 232.100 702.925 233.360 ;
        RECT 703.115 233.080 703.255 234.620 ;
        RECT 703.405 233.360 703.545 235.180 ;
        RECT 703.685 233.640 703.825 235.460 ;
        RECT 704.245 233.920 704.385 236.020 ;
        RECT 704.525 234.200 704.665 236.300 ;
        RECT 705.085 234.480 705.225 236.860 ;
        RECT 705.365 234.760 705.505 237.140 ;
        RECT 705.925 235.040 706.065 237.700 ;
        RECT 706.205 235.320 706.345 237.980 ;
        RECT 778.015 237.980 2147.810 238.120 ;
        RECT 778.015 235.320 778.155 237.980 ;
        RECT 2152.850 237.840 2153.170 237.960 ;
        RECT 706.205 235.180 778.155 235.320 ;
        RECT 778.295 237.700 2153.170 237.840 ;
        RECT 778.295 235.040 778.435 237.700 ;
        RECT 2153.470 237.280 2153.790 237.400 ;
        RECT 705.925 234.900 778.435 235.040 ;
        RECT 778.855 237.140 2153.790 237.280 ;
        RECT 778.855 234.760 778.995 237.140 ;
        RECT 2158.830 237.000 2159.150 237.120 ;
        RECT 705.365 234.620 778.995 234.760 ;
        RECT 779.135 236.860 2159.150 237.000 ;
        RECT 779.135 234.480 779.275 236.860 ;
        RECT 2159.450 236.440 2159.770 236.560 ;
        RECT 705.085 234.340 779.275 234.480 ;
        RECT 779.695 236.300 2159.770 236.440 ;
        RECT 779.695 234.200 779.835 236.300 ;
        RECT 2164.810 236.160 2165.130 236.280 ;
        RECT 704.525 234.060 779.835 234.200 ;
        RECT 779.975 236.020 2165.130 236.160 ;
        RECT 779.975 233.920 780.115 236.020 ;
        RECT 2165.430 235.600 2165.750 235.720 ;
        RECT 704.245 233.780 780.115 233.920 ;
        RECT 780.535 235.460 2165.750 235.600 ;
        RECT 780.535 233.640 780.675 235.460 ;
        RECT 2170.790 235.320 2171.110 235.440 ;
        RECT 703.685 233.500 780.675 233.640 ;
        RECT 780.815 235.180 2171.110 235.320 ;
        RECT 780.815 233.360 780.955 235.180 ;
        RECT 2171.410 234.760 2171.730 234.880 ;
        RECT 703.405 233.220 780.955 233.360 ;
        RECT 781.375 234.620 2171.730 234.760 ;
        RECT 781.375 233.080 781.515 234.620 ;
        RECT 2176.770 234.480 2177.090 234.600 ;
        RECT 703.115 232.940 781.515 233.080 ;
        RECT 781.655 234.340 2177.090 234.480 ;
        RECT 781.655 232.800 781.795 234.340 ;
        RECT 2177.390 233.920 2177.710 234.040 ;
        RECT 703.635 232.660 781.795 232.800 ;
        RECT 782.215 233.780 2177.710 233.920 ;
        RECT 703.635 232.540 703.955 232.660 ;
        RECT 782.215 232.520 782.355 233.780 ;
        RECT 2182.750 233.640 2183.070 233.760 ;
        RECT 704.485 232.380 782.355 232.520 ;
        RECT 782.495 233.500 2183.070 233.640 ;
        RECT 704.485 232.260 704.805 232.380 ;
        RECT 782.495 232.240 782.635 233.500 ;
        RECT 2183.370 233.080 2183.690 233.200 ;
        RECT 705.750 232.100 706.070 232.220 ;
        RECT 702.785 231.960 706.070 232.100 ;
        RECT 709.615 232.100 782.635 232.240 ;
        RECT 783.055 232.940 2183.690 233.080 ;
        RECT 709.615 231.980 709.935 232.100 ;
        RECT 783.055 231.960 783.195 232.940 ;
        RECT 2188.730 232.800 2189.050 232.920 ;
        RECT 706.370 231.820 706.690 231.940 ;
        RECT 702.490 231.680 706.690 231.820 ;
        RECT 710.585 231.820 783.195 231.960 ;
        RECT 783.335 232.660 2189.050 232.800 ;
        RECT 710.585 231.700 710.905 231.820 ;
        RECT 783.335 231.680 783.475 232.660 ;
        RECT 2189.350 232.240 2189.670 232.360 ;
        RECT 711.730 231.540 712.050 231.660 ;
        RECT 702.170 231.400 712.050 231.540 ;
        RECT 715.595 231.540 783.475 231.680 ;
        RECT 783.895 232.100 2189.670 232.240 ;
        RECT 715.595 231.420 715.915 231.540 ;
        RECT 783.895 231.400 784.035 232.100 ;
        RECT 2194.710 231.960 2195.030 232.080 ;
        RECT 712.350 231.260 712.670 231.380 ;
        RECT 701.875 231.120 712.670 231.260 ;
        RECT 716.445 231.260 784.035 231.400 ;
        RECT 784.175 231.820 2195.030 231.960 ;
        RECT 716.445 231.140 716.765 231.260 ;
        RECT 784.175 231.120 784.315 231.820 ;
        RECT 2195.330 231.400 2195.650 231.520 ;
        RECT 717.710 230.980 718.030 231.100 ;
        RECT 701.595 230.840 718.030 230.980 ;
        RECT 721.575 230.980 784.315 231.120 ;
        RECT 784.735 231.260 2195.650 231.400 ;
        RECT 721.575 230.860 721.895 230.980 ;
        RECT 784.735 230.840 784.875 231.260 ;
        RECT 2200.690 231.120 2201.010 231.240 ;
        RECT 718.330 230.700 718.650 230.820 ;
        RECT 701.295 230.560 718.650 230.700 ;
        RECT 722.545 230.700 784.875 230.840 ;
        RECT 785.015 230.980 2201.010 231.120 ;
        RECT 722.545 230.580 722.865 230.700 ;
        RECT 785.015 230.560 785.155 230.980 ;
        RECT 723.690 230.420 724.010 230.540 ;
        RECT 701.015 230.280 724.010 230.420 ;
        RECT 727.555 230.420 785.155 230.560 ;
        RECT 727.555 230.300 727.875 230.420 ;
        RECT 2237.190 225.520 2237.510 225.640 ;
        RECT 764.405 225.380 2237.510 225.520 ;
        RECT 764.405 225.260 764.725 225.380 ;
        RECT 2242.550 225.240 2242.870 225.360 ;
        RECT 769.415 225.100 2242.870 225.240 ;
        RECT 769.415 224.980 769.735 225.100 ;
        RECT 2243.170 224.680 2243.490 224.800 ;
        RECT 770.385 224.540 2243.490 224.680 ;
        RECT 770.385 224.420 770.705 224.540 ;
        RECT 2248.530 224.400 2248.850 224.520 ;
        RECT 775.395 224.260 2248.850 224.400 ;
        RECT 775.395 224.140 775.715 224.260 ;
        RECT 2249.150 223.840 2249.470 223.960 ;
        RECT 776.245 223.700 2249.470 223.840 ;
        RECT 776.245 223.580 776.565 223.700 ;
        RECT 2254.510 223.560 2254.830 223.680 ;
        RECT 781.375 223.420 2254.830 223.560 ;
        RECT 781.375 223.300 781.695 223.420 ;
        RECT 2255.130 223.000 2255.450 223.120 ;
        RECT 782.345 222.860 2255.450 223.000 ;
        RECT 782.345 222.740 782.665 222.860 ;
        RECT 2260.490 222.720 2260.810 222.840 ;
        RECT 787.355 222.580 2260.810 222.720 ;
        RECT 787.355 222.460 787.675 222.580 ;
        RECT 2261.110 222.160 2261.430 222.280 ;
        RECT 788.205 222.020 2261.430 222.160 ;
        RECT 788.205 221.900 788.525 222.020 ;
        RECT 2266.470 221.600 2266.790 221.720 ;
        RECT 793.335 221.460 2266.790 221.600 ;
        RECT 793.335 221.340 793.655 221.460 ;
        RECT 2267.090 221.040 2267.410 221.160 ;
        RECT 794.305 220.900 2267.410 221.040 ;
        RECT 794.305 220.780 794.625 220.900 ;
        RECT 670.470 215.450 670.730 216.420 ;
        RECT 674.180 215.810 675.390 216.070 ;
        RECT 676.450 215.450 676.710 216.420 ;
        RECT 680.160 215.810 681.370 216.070 ;
        RECT 682.430 215.450 682.690 216.420 ;
        RECT 686.140 215.810 687.350 216.070 ;
        RECT 688.410 215.450 688.670 216.420 ;
        RECT 692.120 215.810 693.330 216.070 ;
        RECT 694.390 215.450 694.650 216.420 ;
        RECT 698.100 215.810 699.310 216.070 ;
        RECT 700.370 215.450 700.630 216.420 ;
        RECT 704.080 215.810 705.290 216.070 ;
        RECT 706.350 215.450 706.610 216.420 ;
        RECT 710.060 215.810 711.270 216.070 ;
        RECT 712.330 215.450 712.590 216.420 ;
        RECT 716.040 215.810 717.250 216.070 ;
        RECT 718.310 215.450 718.570 216.420 ;
        RECT 722.020 215.810 723.230 216.070 ;
        RECT 763.880 215.810 765.090 216.070 ;
        RECT 769.860 215.810 771.070 216.070 ;
        RECT 775.840 215.810 777.050 216.070 ;
        RECT 781.820 215.810 783.030 216.070 ;
        RECT 787.800 215.810 789.010 216.070 ;
        RECT 793.780 215.810 794.990 216.070 ;
        RECT 2147.470 215.450 2147.730 216.420 ;
        RECT 2153.450 215.450 2153.710 216.420 ;
        RECT 2159.430 215.450 2159.690 216.420 ;
        RECT 2165.410 215.450 2165.670 216.420 ;
        RECT 2171.390 215.450 2171.650 216.420 ;
        RECT 2177.370 215.450 2177.630 216.420 ;
        RECT 2183.350 215.450 2183.610 216.420 ;
        RECT 2189.330 215.450 2189.590 216.420 ;
        RECT 2195.310 215.450 2195.570 216.420 ;
        RECT 2237.170 215.450 2237.430 216.420 ;
        RECT 2243.150 215.450 2243.410 216.420 ;
        RECT 2249.130 215.450 2249.390 216.420 ;
        RECT 2255.110 215.450 2255.370 216.420 ;
        RECT 2261.090 215.450 2261.350 216.420 ;
        RECT 2267.070 215.450 2267.330 216.420 ;
        RECT 675.530 212.750 676.740 213.010 ;
        RECT 679.680 212.390 679.940 213.360 ;
        RECT 681.510 212.750 682.720 213.010 ;
        RECT 685.660 212.390 685.920 213.360 ;
        RECT 687.490 212.750 688.700 213.010 ;
        RECT 691.640 212.390 691.900 213.360 ;
        RECT 693.470 212.750 694.680 213.010 ;
        RECT 697.620 212.390 697.880 213.360 ;
        RECT 699.450 212.750 700.660 213.010 ;
        RECT 703.600 212.390 703.860 213.360 ;
        RECT 705.430 212.750 706.640 213.010 ;
        RECT 709.580 212.390 709.840 213.360 ;
        RECT 711.410 212.750 712.620 213.010 ;
        RECT 715.560 212.390 715.820 213.360 ;
        RECT 717.390 212.750 718.600 213.010 ;
        RECT 721.540 212.390 721.800 213.360 ;
        RECT 723.370 212.750 724.580 213.010 ;
        RECT 727.520 212.390 727.780 213.360 ;
        RECT 769.380 212.390 769.640 213.360 ;
        RECT 775.360 212.390 775.620 213.360 ;
        RECT 781.340 212.390 781.600 213.360 ;
        RECT 787.320 212.390 787.580 213.360 ;
        RECT 793.280 212.750 794.490 213.010 ;
        RECT 2152.530 212.750 2153.740 213.010 ;
        RECT 2158.510 212.750 2159.720 213.010 ;
        RECT 2164.490 212.750 2165.700 213.010 ;
        RECT 2170.470 212.750 2171.680 213.010 ;
        RECT 2176.450 212.750 2177.660 213.010 ;
        RECT 2182.430 212.750 2183.640 213.010 ;
        RECT 2188.410 212.750 2189.620 213.010 ;
        RECT 2194.390 212.750 2195.600 213.010 ;
        RECT 2200.370 212.750 2201.580 213.010 ;
        RECT 2242.230 212.750 2243.440 213.010 ;
        RECT 2248.210 212.750 2249.420 213.010 ;
        RECT 2254.190 212.750 2255.400 213.010 ;
        RECT 2260.170 212.750 2261.380 213.010 ;
        RECT 2267.080 212.390 2267.340 213.360 ;
      LAYER via ;
        RECT 3370.800 3603.580 3371.060 3603.840 ;
        RECT 3370.520 3602.960 3370.780 3603.220 ;
        RECT 203.035 3009.260 203.295 3010.350 ;
        RECT 205.795 3010.120 206.645 3010.380 ;
        RECT 217.615 3010.170 217.875 3010.430 ;
        RECT 203.035 3003.280 203.295 3004.370 ;
        RECT 205.795 3004.140 206.645 3004.400 ;
        RECT 203.035 2997.300 203.295 2998.390 ;
        RECT 205.795 2998.160 206.645 2998.420 ;
        RECT 203.035 2991.320 203.295 2992.410 ;
        RECT 205.795 2992.180 206.645 2992.440 ;
        RECT 203.035 2985.340 203.295 2986.430 ;
        RECT 205.795 2986.200 206.645 2986.460 ;
        RECT 206.205 1725.985 206.465 1727.075 ;
        RECT 217.495 1726.480 217.755 1726.740 ;
        RECT 217.895 3009.550 218.155 3009.810 ;
        RECT 202.845 1725.445 203.695 1725.705 ;
        RECT 217.775 1725.510 218.035 1725.770 ;
        RECT 218.735 3004.190 218.995 3004.450 ;
        RECT 203.145 1721.355 203.405 1722.445 ;
        RECT 205.905 1722.215 206.755 1722.475 ;
        RECT 217.475 1722.265 217.735 1722.525 ;
        RECT 206.205 1720.005 206.465 1721.095 ;
        RECT 202.845 1719.465 203.695 1719.725 ;
        RECT 203.145 1715.805 203.405 1716.465 ;
        RECT 205.905 1716.235 206.755 1716.495 ;
        RECT 203.145 1715.375 203.405 1715.665 ;
        RECT 206.205 1714.025 206.465 1715.115 ;
        RECT 202.845 1713.485 203.695 1713.745 ;
        RECT 203.145 1709.395 203.405 1710.485 ;
        RECT 205.905 1710.255 206.755 1710.515 ;
        RECT 206.205 1708.045 206.465 1709.135 ;
        RECT 202.845 1707.505 203.695 1707.765 ;
        RECT 203.145 1703.415 203.405 1704.505 ;
        RECT 205.905 1704.275 206.755 1704.535 ;
        RECT 206.205 1702.065 206.465 1703.155 ;
        RECT 202.845 1701.525 203.695 1701.785 ;
        RECT 203.145 1697.435 203.405 1698.525 ;
        RECT 205.905 1698.295 206.755 1698.555 ;
        RECT 203.145 1691.455 203.405 1692.545 ;
        RECT 205.905 1692.315 206.755 1692.575 ;
        RECT 203.145 1685.475 203.405 1686.565 ;
        RECT 205.905 1686.335 206.755 1686.595 ;
        RECT 203.145 1679.495 203.405 1680.585 ;
        RECT 205.905 1680.355 206.755 1680.615 ;
        RECT 203.145 1673.515 203.405 1674.605 ;
        RECT 205.905 1674.375 206.755 1674.635 ;
        RECT 217.755 1721.645 218.015 1721.905 ;
        RECT 218.615 1720.500 218.875 1720.760 ;
        RECT 219.015 3003.570 219.275 3003.830 ;
        RECT 218.895 1719.530 219.155 1719.790 ;
        RECT 219.855 2998.210 220.115 2998.470 ;
        RECT 218.595 1716.285 218.855 1716.545 ;
        RECT 218.875 1715.665 219.135 1715.925 ;
        RECT 219.735 1714.520 219.995 1714.780 ;
        RECT 220.135 2997.590 220.395 2997.850 ;
        RECT 220.015 1713.550 220.275 1713.810 ;
        RECT 220.975 2992.230 221.235 2992.490 ;
        RECT 219.715 1710.305 219.975 1710.565 ;
        RECT 219.995 1709.685 220.255 1709.945 ;
        RECT 220.855 1708.540 221.115 1708.800 ;
        RECT 221.255 2991.610 221.515 2991.870 ;
        RECT 221.135 1707.570 221.395 1707.830 ;
        RECT 222.095 2986.250 222.355 2986.510 ;
        RECT 220.835 1704.325 221.095 1704.585 ;
        RECT 221.115 1703.705 221.375 1703.965 ;
        RECT 221.975 1702.560 222.235 1702.820 ;
        RECT 222.375 2985.630 222.635 2985.890 ;
        RECT 3381.350 3603.530 3382.200 3603.790 ;
        RECT 3384.700 3602.670 3384.960 3603.760 ;
        RECT 3370.920 2237.675 3371.180 2237.935 ;
        RECT 3381.640 2237.180 3381.900 2238.270 ;
        RECT 3370.640 2236.705 3370.900 2236.965 ;
        RECT 3384.410 2236.640 3385.260 2236.900 ;
        RECT 222.255 1701.590 222.515 1701.850 ;
        RECT 221.955 1698.345 222.215 1698.605 ;
        RECT 222.235 1697.725 222.495 1697.985 ;
        RECT 223.075 1692.365 223.335 1692.625 ;
        RECT 223.355 1691.745 223.615 1692.005 ;
        RECT 224.195 1686.385 224.455 1686.645 ;
        RECT 224.475 1685.765 224.735 1686.025 ;
        RECT 225.315 1680.405 225.575 1680.665 ;
        RECT 225.595 1679.785 225.855 1680.045 ;
        RECT 226.435 1674.425 226.695 1674.685 ;
        RECT 226.715 1673.805 226.975 1674.065 ;
        RECT 670.520 237.840 670.780 238.100 ;
        RECT 674.735 237.860 674.995 238.120 ;
        RECT 675.880 237.560 676.140 237.820 ;
        RECT 679.745 237.580 680.005 237.840 ;
        RECT 676.500 237.000 676.760 237.260 ;
        RECT 680.715 237.020 680.975 237.280 ;
        RECT 681.860 236.720 682.120 236.980 ;
        RECT 685.725 236.740 685.985 237.000 ;
        RECT 682.480 236.160 682.740 236.420 ;
        RECT 686.695 236.180 686.955 236.440 ;
        RECT 687.840 235.880 688.100 236.140 ;
        RECT 691.705 235.900 691.965 236.160 ;
        RECT 688.460 235.320 688.720 235.580 ;
        RECT 692.675 235.340 692.935 235.600 ;
        RECT 693.820 235.040 694.080 235.300 ;
        RECT 697.685 235.060 697.945 235.320 ;
        RECT 694.440 234.480 694.700 234.740 ;
        RECT 698.655 234.500 698.915 234.760 ;
        RECT 699.800 234.200 700.060 234.460 ;
        RECT 700.420 233.640 700.680 233.900 ;
        RECT 2147.520 237.980 2147.780 238.240 ;
        RECT 2152.880 237.700 2153.140 237.960 ;
        RECT 2153.500 237.140 2153.760 237.400 ;
        RECT 2158.860 236.860 2159.120 237.120 ;
        RECT 2159.480 236.300 2159.740 236.560 ;
        RECT 2164.840 236.020 2165.100 236.280 ;
        RECT 2165.460 235.460 2165.720 235.720 ;
        RECT 2170.820 235.180 2171.080 235.440 ;
        RECT 2171.440 234.620 2171.700 234.880 ;
        RECT 2176.800 234.340 2177.060 234.600 ;
        RECT 703.665 232.540 703.925 232.800 ;
        RECT 2177.420 233.780 2177.680 234.040 ;
        RECT 704.515 232.260 704.775 232.520 ;
        RECT 2182.780 233.500 2183.040 233.760 ;
        RECT 705.780 231.960 706.040 232.220 ;
        RECT 709.645 231.980 709.905 232.240 ;
        RECT 2183.400 232.940 2183.660 233.200 ;
        RECT 706.400 231.680 706.660 231.940 ;
        RECT 710.615 231.700 710.875 231.960 ;
        RECT 2188.760 232.660 2189.020 232.920 ;
        RECT 711.760 231.400 712.020 231.660 ;
        RECT 715.625 231.420 715.885 231.680 ;
        RECT 2189.380 232.100 2189.640 232.360 ;
        RECT 712.380 231.120 712.640 231.380 ;
        RECT 716.475 231.140 716.735 231.400 ;
        RECT 2194.740 231.820 2195.000 232.080 ;
        RECT 717.740 230.840 718.000 231.100 ;
        RECT 721.605 230.860 721.865 231.120 ;
        RECT 2195.360 231.260 2195.620 231.520 ;
        RECT 718.360 230.560 718.620 230.820 ;
        RECT 722.575 230.580 722.835 230.840 ;
        RECT 2200.720 230.980 2200.980 231.240 ;
        RECT 723.720 230.280 723.980 230.540 ;
        RECT 727.585 230.300 727.845 230.560 ;
        RECT 764.435 225.260 764.695 225.520 ;
        RECT 2237.220 225.380 2237.480 225.640 ;
        RECT 769.445 224.980 769.705 225.240 ;
        RECT 2242.580 225.100 2242.840 225.360 ;
        RECT 770.415 224.420 770.675 224.680 ;
        RECT 2243.200 224.540 2243.460 224.800 ;
        RECT 775.425 224.140 775.685 224.400 ;
        RECT 2248.560 224.260 2248.820 224.520 ;
        RECT 776.275 223.580 776.535 223.840 ;
        RECT 2249.180 223.700 2249.440 223.960 ;
        RECT 781.405 223.300 781.665 223.560 ;
        RECT 2254.540 223.420 2254.800 223.680 ;
        RECT 782.375 222.740 782.635 223.000 ;
        RECT 2255.160 222.860 2255.420 223.120 ;
        RECT 787.385 222.460 787.645 222.720 ;
        RECT 2260.520 222.580 2260.780 222.840 ;
        RECT 788.235 221.900 788.495 222.160 ;
        RECT 2261.140 222.020 2261.400 222.280 ;
        RECT 793.365 221.340 793.625 221.600 ;
        RECT 2266.500 221.460 2266.760 221.720 ;
        RECT 794.335 220.780 794.595 221.040 ;
        RECT 2267.120 220.900 2267.380 221.160 ;
        RECT 670.470 215.510 670.730 216.360 ;
        RECT 674.240 215.810 675.330 216.070 ;
        RECT 676.450 215.510 676.710 216.360 ;
        RECT 680.220 215.810 681.310 216.070 ;
        RECT 682.430 215.510 682.690 216.360 ;
        RECT 686.200 215.810 687.290 216.070 ;
        RECT 688.410 215.510 688.670 216.360 ;
        RECT 692.180 215.810 693.270 216.070 ;
        RECT 694.390 215.510 694.650 216.360 ;
        RECT 698.160 215.810 699.250 216.070 ;
        RECT 700.370 215.510 700.630 216.360 ;
        RECT 704.140 215.810 705.230 216.070 ;
        RECT 706.350 215.510 706.610 216.360 ;
        RECT 710.120 215.810 711.210 216.070 ;
        RECT 712.330 215.510 712.590 216.360 ;
        RECT 716.100 215.810 717.190 216.070 ;
        RECT 718.310 215.510 718.570 216.360 ;
        RECT 722.080 215.810 723.170 216.070 ;
        RECT 763.940 215.810 765.030 216.070 ;
        RECT 769.920 215.810 771.010 216.070 ;
        RECT 775.900 215.810 776.990 216.070 ;
        RECT 781.880 215.810 782.970 216.070 ;
        RECT 787.860 215.810 788.950 216.070 ;
        RECT 793.840 215.810 794.930 216.070 ;
        RECT 2147.470 215.510 2147.730 216.360 ;
        RECT 2153.450 215.510 2153.710 216.360 ;
        RECT 2159.430 215.510 2159.690 216.360 ;
        RECT 2165.410 215.510 2165.670 216.360 ;
        RECT 2171.390 215.510 2171.650 216.360 ;
        RECT 2177.370 215.510 2177.630 216.360 ;
        RECT 2183.350 215.510 2183.610 216.360 ;
        RECT 2189.330 215.510 2189.590 216.360 ;
        RECT 2195.310 215.510 2195.570 216.360 ;
        RECT 2237.170 215.510 2237.430 216.360 ;
        RECT 2243.150 215.510 2243.410 216.360 ;
        RECT 2249.130 215.510 2249.390 216.360 ;
        RECT 2255.110 215.510 2255.370 216.360 ;
        RECT 2261.090 215.510 2261.350 216.360 ;
        RECT 2267.070 215.510 2267.330 216.360 ;
        RECT 675.590 212.750 676.680 213.010 ;
        RECT 679.680 212.450 679.940 213.300 ;
        RECT 681.570 212.750 682.660 213.010 ;
        RECT 685.660 212.450 685.920 213.300 ;
        RECT 687.550 212.750 688.640 213.010 ;
        RECT 691.640 212.450 691.900 213.300 ;
        RECT 693.530 212.750 694.620 213.010 ;
        RECT 697.620 212.450 697.880 213.300 ;
        RECT 699.510 212.750 700.600 213.010 ;
        RECT 703.600 212.450 703.860 213.300 ;
        RECT 705.490 212.750 706.580 213.010 ;
        RECT 709.580 212.450 709.840 213.300 ;
        RECT 711.470 212.750 712.560 213.010 ;
        RECT 715.560 212.450 715.820 213.300 ;
        RECT 717.450 212.750 718.540 213.010 ;
        RECT 721.540 212.450 721.800 213.300 ;
        RECT 723.430 212.750 724.520 213.010 ;
        RECT 727.520 212.450 727.780 213.300 ;
        RECT 769.380 212.450 769.640 213.300 ;
        RECT 775.360 212.450 775.620 213.300 ;
        RECT 781.340 212.450 781.600 213.300 ;
        RECT 787.320 212.450 787.580 213.300 ;
        RECT 793.340 212.750 794.430 213.010 ;
        RECT 2152.590 212.750 2153.680 213.010 ;
        RECT 2158.570 212.750 2159.660 213.010 ;
        RECT 2164.550 212.750 2165.640 213.010 ;
        RECT 2170.530 212.750 2171.620 213.010 ;
        RECT 2176.510 212.750 2177.600 213.010 ;
        RECT 2182.490 212.750 2183.580 213.010 ;
        RECT 2188.470 212.750 2189.560 213.010 ;
        RECT 2194.450 212.750 2195.540 213.010 ;
        RECT 2200.430 212.750 2201.520 213.010 ;
        RECT 2242.290 212.750 2243.380 213.010 ;
        RECT 2248.270 212.750 2249.360 213.010 ;
        RECT 2254.250 212.750 2255.340 213.010 ;
        RECT 2260.230 212.750 2261.320 213.010 ;
        RECT 2267.080 212.450 2267.340 213.300 ;
      LAYER met2 ;
        RECT 3370.770 3603.720 3371.090 3603.840 ;
        RECT 3381.350 3603.720 3382.200 3603.820 ;
        RECT 3370.330 3603.580 3382.200 3603.720 ;
        RECT 3381.350 3603.500 3382.200 3603.580 ;
        RECT 3370.490 3603.100 3370.810 3603.220 ;
        RECT 3384.670 3603.100 3384.990 3603.760 ;
        RECT 3370.330 3602.960 3384.990 3603.100 ;
        RECT 3384.670 3602.670 3384.990 3602.960 ;
        RECT 203.005 3009.690 203.325 3010.350 ;
        RECT 205.795 3010.310 206.645 3010.410 ;
        RECT 217.585 3010.310 217.905 3010.430 ;
        RECT 205.795 3010.170 221.600 3010.310 ;
        RECT 205.795 3010.090 206.645 3010.170 ;
        RECT 217.865 3009.690 218.185 3009.810 ;
        RECT 203.005 3009.550 221.600 3009.690 ;
        RECT 203.005 3009.260 203.325 3009.550 ;
        RECT 203.005 3003.710 203.325 3004.370 ;
        RECT 205.795 3004.330 206.645 3004.430 ;
        RECT 218.705 3004.330 219.025 3004.450 ;
        RECT 205.795 3004.190 221.600 3004.330 ;
        RECT 205.795 3004.110 206.645 3004.190 ;
        RECT 218.985 3003.710 219.305 3003.830 ;
        RECT 203.005 3003.570 221.600 3003.710 ;
        RECT 203.005 3003.280 203.325 3003.570 ;
        RECT 203.005 2997.730 203.325 2998.390 ;
        RECT 205.795 2998.350 206.645 2998.450 ;
        RECT 219.825 2998.350 220.145 2998.470 ;
        RECT 205.795 2998.210 221.600 2998.350 ;
        RECT 205.795 2998.130 206.645 2998.210 ;
        RECT 220.105 2997.730 220.425 2997.850 ;
        RECT 203.005 2997.590 221.600 2997.730 ;
        RECT 203.005 2997.300 203.325 2997.590 ;
        RECT 203.005 2991.750 203.325 2992.410 ;
        RECT 205.795 2992.370 206.645 2992.470 ;
        RECT 220.945 2992.370 221.265 2992.490 ;
        RECT 205.795 2992.230 221.675 2992.370 ;
        RECT 205.795 2992.150 206.645 2992.230 ;
        RECT 221.225 2991.750 221.545 2991.870 ;
        RECT 203.005 2991.610 221.675 2991.750 ;
        RECT 203.005 2991.320 203.325 2991.610 ;
        RECT 203.005 2985.770 203.325 2986.430 ;
        RECT 205.795 2986.390 206.645 2986.490 ;
        RECT 222.065 2986.390 222.385 2986.510 ;
        RECT 205.795 2986.250 222.720 2986.390 ;
        RECT 205.795 2986.170 206.645 2986.250 ;
        RECT 222.345 2985.770 222.665 2985.890 ;
        RECT 203.005 2985.630 222.720 2985.770 ;
        RECT 203.005 2985.340 203.325 2985.630 ;
        RECT 3370.890 2237.815 3371.210 2237.935 ;
        RECT 3381.610 2237.815 3381.930 2238.270 ;
        RECT 3365.990 2237.675 3381.930 2237.815 ;
        RECT 3381.610 2237.180 3381.930 2237.675 ;
        RECT 3370.610 2236.845 3370.930 2236.965 ;
        RECT 3384.410 2236.845 3385.260 2236.930 ;
        RECT 3365.990 2236.705 3385.260 2236.845 ;
        RECT 3384.410 2236.610 3385.260 2236.705 ;
        RECT 206.175 1726.620 206.495 1727.075 ;
        RECT 217.465 1726.620 217.785 1726.740 ;
        RECT 206.175 1726.480 223.740 1726.620 ;
        RECT 206.175 1725.985 206.495 1726.480 ;
        RECT 202.845 1725.650 203.695 1725.735 ;
        RECT 217.745 1725.650 218.065 1725.770 ;
        RECT 202.845 1725.510 223.740 1725.650 ;
        RECT 202.845 1725.415 203.695 1725.510 ;
        RECT 203.115 1721.785 203.435 1722.445 ;
        RECT 205.905 1722.405 206.755 1722.505 ;
        RECT 217.445 1722.405 217.765 1722.525 ;
        RECT 205.905 1722.265 223.740 1722.405 ;
        RECT 205.905 1722.185 206.755 1722.265 ;
        RECT 217.725 1721.785 218.045 1721.905 ;
        RECT 203.115 1721.645 223.740 1721.785 ;
        RECT 203.115 1721.355 203.435 1721.645 ;
        RECT 206.175 1720.640 206.495 1721.095 ;
        RECT 218.585 1720.640 218.905 1720.760 ;
        RECT 206.175 1720.500 223.740 1720.640 ;
        RECT 206.175 1720.005 206.495 1720.500 ;
        RECT 202.845 1719.670 203.695 1719.755 ;
        RECT 218.865 1719.670 219.185 1719.790 ;
        RECT 202.845 1719.530 223.740 1719.670 ;
        RECT 202.845 1719.435 203.695 1719.530 ;
        RECT 203.115 1715.805 203.435 1716.465 ;
        RECT 205.905 1716.425 206.755 1716.525 ;
        RECT 218.565 1716.425 218.885 1716.545 ;
        RECT 205.905 1716.285 223.740 1716.425 ;
        RECT 205.905 1716.205 206.755 1716.285 ;
        RECT 218.845 1715.805 219.165 1715.925 ;
        RECT 202.845 1715.665 223.740 1715.805 ;
        RECT 203.115 1715.375 203.435 1715.665 ;
        RECT 206.175 1714.660 206.495 1715.115 ;
        RECT 219.705 1714.660 220.025 1714.780 ;
        RECT 206.175 1714.520 223.740 1714.660 ;
        RECT 206.175 1714.025 206.495 1714.520 ;
        RECT 202.845 1713.690 203.695 1713.775 ;
        RECT 219.985 1713.690 220.305 1713.810 ;
        RECT 202.845 1713.550 223.740 1713.690 ;
        RECT 202.845 1713.455 203.695 1713.550 ;
        RECT 203.115 1709.825 203.435 1710.485 ;
        RECT 205.905 1710.445 206.755 1710.545 ;
        RECT 219.685 1710.445 220.005 1710.565 ;
        RECT 205.905 1710.305 223.740 1710.445 ;
        RECT 205.905 1710.225 206.755 1710.305 ;
        RECT 219.965 1709.825 220.285 1709.945 ;
        RECT 203.115 1709.685 223.740 1709.825 ;
        RECT 203.115 1709.395 203.435 1709.685 ;
        RECT 206.175 1708.680 206.495 1709.135 ;
        RECT 220.825 1708.680 221.145 1708.800 ;
        RECT 206.175 1708.540 223.740 1708.680 ;
        RECT 206.175 1708.045 206.495 1708.540 ;
        RECT 202.845 1707.710 203.695 1707.795 ;
        RECT 221.105 1707.710 221.425 1707.830 ;
        RECT 202.845 1707.570 223.740 1707.710 ;
        RECT 202.845 1707.475 203.695 1707.570 ;
        RECT 203.115 1703.845 203.435 1704.505 ;
        RECT 205.905 1704.465 206.755 1704.565 ;
        RECT 220.805 1704.465 221.125 1704.585 ;
        RECT 205.905 1704.325 223.740 1704.465 ;
        RECT 205.905 1704.245 206.755 1704.325 ;
        RECT 221.085 1703.845 221.405 1703.965 ;
        RECT 203.115 1703.705 223.740 1703.845 ;
        RECT 203.115 1703.415 203.435 1703.705 ;
        RECT 206.175 1702.700 206.495 1703.155 ;
        RECT 221.945 1702.700 222.265 1702.820 ;
        RECT 206.175 1702.560 223.740 1702.700 ;
        RECT 206.175 1702.065 206.495 1702.560 ;
        RECT 202.845 1701.730 203.695 1701.815 ;
        RECT 222.225 1701.730 222.545 1701.850 ;
        RECT 202.845 1701.590 223.740 1701.730 ;
        RECT 202.845 1701.495 203.695 1701.590 ;
        RECT 203.115 1697.865 203.435 1698.525 ;
        RECT 205.905 1698.485 206.755 1698.585 ;
        RECT 221.925 1698.485 222.245 1698.605 ;
        RECT 205.905 1698.345 223.740 1698.485 ;
        RECT 205.905 1698.265 206.755 1698.345 ;
        RECT 222.205 1697.865 222.525 1697.985 ;
        RECT 203.115 1697.725 223.740 1697.865 ;
        RECT 203.115 1697.435 203.435 1697.725 ;
        RECT 203.115 1691.885 203.435 1692.545 ;
        RECT 205.905 1692.505 206.755 1692.605 ;
        RECT 223.045 1692.505 223.365 1692.625 ;
        RECT 205.905 1692.365 223.745 1692.505 ;
        RECT 205.905 1692.285 206.755 1692.365 ;
        RECT 223.325 1691.885 223.645 1692.005 ;
        RECT 203.115 1691.745 223.745 1691.885 ;
        RECT 203.115 1691.455 203.435 1691.745 ;
        RECT 203.115 1685.905 203.435 1686.565 ;
        RECT 205.905 1686.525 206.755 1686.625 ;
        RECT 224.165 1686.525 224.485 1686.645 ;
        RECT 205.905 1686.385 224.805 1686.525 ;
        RECT 205.905 1686.305 206.755 1686.385 ;
        RECT 224.445 1685.905 224.765 1686.025 ;
        RECT 203.115 1685.765 224.805 1685.905 ;
        RECT 203.115 1685.475 203.435 1685.765 ;
        RECT 203.115 1679.925 203.435 1680.585 ;
        RECT 205.905 1680.545 206.755 1680.645 ;
        RECT 225.285 1680.545 225.605 1680.665 ;
        RECT 205.905 1680.405 226.030 1680.545 ;
        RECT 205.905 1680.325 206.755 1680.405 ;
        RECT 225.565 1679.925 225.885 1680.045 ;
        RECT 203.115 1679.785 226.030 1679.925 ;
        RECT 203.115 1679.495 203.435 1679.785 ;
        RECT 203.115 1673.945 203.435 1674.605 ;
        RECT 205.905 1674.565 206.755 1674.665 ;
        RECT 226.405 1674.565 226.725 1674.685 ;
        RECT 205.905 1674.425 227.100 1674.565 ;
        RECT 205.905 1674.345 206.755 1674.425 ;
        RECT 226.685 1673.945 227.005 1674.065 ;
        RECT 203.115 1673.805 227.100 1673.945 ;
        RECT 203.115 1673.515 203.435 1673.805 ;
        RECT 2147.520 238.270 2147.660 238.365 ;
        RECT 670.520 238.130 670.660 238.225 ;
        RECT 674.735 238.150 674.875 238.225 ;
        RECT 670.520 237.810 670.780 238.130 ;
        RECT 674.735 237.830 674.995 238.150 ;
        RECT 2147.520 237.950 2147.780 238.270 ;
        RECT 2152.880 237.990 2153.020 238.050 ;
        RECT 675.880 237.850 676.020 237.900 ;
        RECT 679.745 237.870 679.885 237.925 ;
        RECT 670.520 216.360 670.660 237.810 ;
        RECT 670.440 215.510 670.760 216.360 ;
        RECT 674.735 216.100 674.875 237.830 ;
        RECT 675.880 237.530 676.140 237.850 ;
        RECT 679.745 237.550 680.005 237.870 ;
        RECT 674.240 215.780 675.330 216.100 ;
        RECT 675.880 213.040 676.020 237.530 ;
        RECT 676.500 237.290 676.640 237.400 ;
        RECT 676.500 236.970 676.760 237.290 ;
        RECT 676.500 216.360 676.640 236.970 ;
        RECT 676.420 215.510 676.740 216.360 ;
        RECT 679.745 213.300 679.885 237.550 ;
        RECT 680.715 237.310 680.855 237.400 ;
        RECT 680.715 236.990 680.975 237.310 ;
        RECT 681.860 237.010 682.000 237.050 ;
        RECT 685.725 237.030 685.865 237.085 ;
        RECT 680.715 216.100 680.855 236.990 ;
        RECT 681.860 236.690 682.120 237.010 ;
        RECT 685.725 236.710 685.985 237.030 ;
        RECT 680.220 215.780 681.310 216.100 ;
        RECT 675.590 212.720 676.680 213.040 ;
        RECT 679.650 212.450 679.970 213.300 ;
        RECT 681.860 213.040 682.000 236.690 ;
        RECT 682.480 236.450 682.620 236.545 ;
        RECT 682.480 236.130 682.740 236.450 ;
        RECT 682.480 216.360 682.620 236.130 ;
        RECT 682.400 215.510 682.720 216.360 ;
        RECT 685.725 213.300 685.865 236.710 ;
        RECT 686.695 236.470 686.835 236.520 ;
        RECT 686.695 236.150 686.955 236.470 ;
        RECT 687.840 236.170 687.980 236.235 ;
        RECT 691.705 236.190 691.845 236.260 ;
        RECT 686.695 216.100 686.835 236.150 ;
        RECT 687.840 235.850 688.100 236.170 ;
        RECT 691.705 235.870 691.965 236.190 ;
        RECT 686.200 215.780 687.290 216.100 ;
        RECT 681.570 212.720 682.660 213.040 ;
        RECT 685.630 212.450 685.950 213.300 ;
        RECT 687.840 213.040 687.980 235.850 ;
        RECT 688.460 235.610 688.600 235.815 ;
        RECT 688.460 235.290 688.720 235.610 ;
        RECT 688.460 216.360 688.600 235.290 ;
        RECT 688.380 215.510 688.700 216.360 ;
        RECT 691.705 213.300 691.845 235.870 ;
        RECT 692.675 235.630 692.815 235.695 ;
        RECT 692.675 235.310 692.935 235.630 ;
        RECT 693.820 235.330 693.960 235.450 ;
        RECT 697.685 235.350 697.825 235.470 ;
        RECT 692.675 216.100 692.815 235.310 ;
        RECT 693.820 235.010 694.080 235.330 ;
        RECT 697.685 235.030 697.945 235.350 ;
        RECT 692.180 215.780 693.270 216.100 ;
        RECT 687.550 212.720 688.640 213.040 ;
        RECT 691.610 212.450 691.930 213.300 ;
        RECT 693.820 213.040 693.960 235.010 ;
        RECT 694.440 234.770 694.580 234.870 ;
        RECT 694.440 234.450 694.700 234.770 ;
        RECT 694.440 216.360 694.580 234.450 ;
        RECT 694.360 215.510 694.680 216.360 ;
        RECT 697.685 213.300 697.825 235.030 ;
        RECT 698.655 234.790 698.795 234.905 ;
        RECT 698.655 234.470 698.915 234.790 ;
        RECT 699.800 234.490 699.940 234.515 ;
        RECT 698.655 216.100 698.795 234.470 ;
        RECT 699.800 234.170 700.060 234.490 ;
        RECT 698.160 215.780 699.250 216.100 ;
        RECT 693.530 212.720 694.620 213.040 ;
        RECT 697.590 212.450 697.910 213.300 ;
        RECT 699.800 213.040 699.940 234.170 ;
        RECT 700.420 233.930 700.560 234.060 ;
        RECT 700.420 233.610 700.680 233.930 ;
        RECT 700.420 216.360 700.560 233.610 ;
        RECT 703.665 232.830 703.805 232.890 ;
        RECT 703.665 232.510 703.925 232.830 ;
        RECT 704.635 232.550 704.775 232.680 ;
        RECT 700.340 215.510 700.660 216.360 ;
        RECT 703.665 213.300 703.805 232.510 ;
        RECT 704.515 232.230 704.775 232.550 ;
        RECT 704.635 216.100 704.775 232.230 ;
        RECT 705.780 232.250 705.920 232.315 ;
        RECT 709.645 232.270 709.785 232.310 ;
        RECT 705.780 231.930 706.040 232.250 ;
        RECT 706.400 231.970 706.540 232.150 ;
        RECT 704.140 215.780 705.230 216.100 ;
        RECT 699.510 212.720 700.600 213.040 ;
        RECT 703.570 212.450 703.890 213.300 ;
        RECT 705.780 213.040 705.920 231.930 ;
        RECT 706.400 231.650 706.660 231.970 ;
        RECT 709.645 231.950 709.905 232.270 ;
        RECT 710.615 231.990 710.755 232.190 ;
        RECT 706.400 216.360 706.540 231.650 ;
        RECT 706.320 215.510 706.640 216.360 ;
        RECT 709.645 213.300 709.785 231.950 ;
        RECT 710.615 231.670 710.875 231.990 ;
        RECT 711.760 231.690 711.900 231.750 ;
        RECT 715.625 231.710 715.765 231.780 ;
        RECT 710.615 216.100 710.755 231.670 ;
        RECT 711.760 231.370 712.020 231.690 ;
        RECT 712.380 231.410 712.520 231.505 ;
        RECT 710.120 215.780 711.210 216.100 ;
        RECT 705.490 212.720 706.580 213.040 ;
        RECT 709.550 212.450 709.870 213.300 ;
        RECT 711.760 213.040 711.900 231.370 ;
        RECT 712.380 231.090 712.640 231.410 ;
        RECT 715.625 231.390 715.885 231.710 ;
        RECT 716.595 231.430 716.735 231.525 ;
        RECT 712.380 216.360 712.520 231.090 ;
        RECT 712.300 215.510 712.620 216.360 ;
        RECT 715.625 213.300 715.765 231.390 ;
        RECT 716.475 231.110 716.735 231.430 ;
        RECT 716.595 216.100 716.735 231.110 ;
        RECT 717.740 231.130 717.880 232.345 ;
        RECT 717.740 230.810 718.000 231.130 ;
        RECT 718.360 230.850 718.500 232.345 ;
        RECT 721.605 231.150 721.745 232.345 ;
        RECT 716.100 215.780 717.190 216.100 ;
        RECT 711.470 212.720 712.560 213.040 ;
        RECT 715.530 212.450 715.850 213.300 ;
        RECT 717.740 213.040 717.880 230.810 ;
        RECT 718.360 230.530 718.620 230.850 ;
        RECT 721.605 230.830 721.865 231.150 ;
        RECT 722.575 230.870 722.715 232.345 ;
        RECT 718.360 216.360 718.500 230.530 ;
        RECT 718.280 215.510 718.600 216.360 ;
        RECT 721.605 213.300 721.745 230.830 ;
        RECT 722.575 230.550 722.835 230.870 ;
        RECT 723.720 230.570 723.860 232.345 ;
        RECT 727.585 230.590 727.725 232.345 ;
        RECT 722.575 216.100 722.715 230.550 ;
        RECT 723.720 230.250 723.980 230.570 ;
        RECT 727.585 230.270 727.845 230.590 ;
        RECT 722.080 215.780 723.170 216.100 ;
        RECT 717.450 212.720 718.540 213.040 ;
        RECT 721.510 212.450 721.830 213.300 ;
        RECT 723.720 213.040 723.860 230.250 ;
        RECT 727.585 213.300 727.725 230.270 ;
        RECT 764.435 225.550 764.575 232.345 ;
        RECT 764.435 225.230 764.695 225.550 ;
        RECT 769.445 225.270 769.585 232.345 ;
        RECT 764.435 216.100 764.575 225.230 ;
        RECT 769.445 224.950 769.705 225.270 ;
        RECT 763.940 215.780 765.030 216.100 ;
        RECT 769.445 213.300 769.585 224.950 ;
        RECT 770.415 224.710 770.555 232.345 ;
        RECT 770.415 224.390 770.675 224.710 ;
        RECT 775.425 224.430 775.565 232.345 ;
        RECT 770.415 216.100 770.555 224.390 ;
        RECT 775.425 224.110 775.685 224.430 ;
        RECT 769.920 215.780 771.010 216.100 ;
        RECT 775.425 213.300 775.565 224.110 ;
        RECT 776.395 223.870 776.535 232.345 ;
        RECT 776.275 223.550 776.535 223.870 ;
        RECT 776.395 216.100 776.535 223.550 ;
        RECT 781.405 223.590 781.545 232.345 ;
        RECT 781.405 223.270 781.665 223.590 ;
        RECT 775.900 215.780 776.990 216.100 ;
        RECT 781.405 213.300 781.545 223.270 ;
        RECT 782.375 223.030 782.515 232.345 ;
        RECT 782.375 222.710 782.635 223.030 ;
        RECT 787.385 222.750 787.525 232.345 ;
        RECT 782.375 216.100 782.515 222.710 ;
        RECT 787.385 222.430 787.645 222.750 ;
        RECT 781.880 215.780 782.970 216.100 ;
        RECT 787.385 213.300 787.525 222.430 ;
        RECT 788.355 222.190 788.495 232.345 ;
        RECT 788.235 221.870 788.495 222.190 ;
        RECT 788.355 216.100 788.495 221.870 ;
        RECT 793.365 221.630 793.505 232.345 ;
        RECT 793.365 221.310 793.625 221.630 ;
        RECT 787.860 215.780 788.950 216.100 ;
        RECT 793.365 214.240 793.505 221.310 ;
        RECT 794.335 221.070 794.475 232.345 ;
        RECT 794.335 220.750 794.595 221.070 ;
        RECT 794.335 216.100 794.475 220.750 ;
        RECT 2147.520 216.360 2147.660 237.950 ;
        RECT 2152.880 237.670 2153.140 237.990 ;
        RECT 793.840 215.780 794.930 216.100 ;
        RECT 2147.440 215.510 2147.760 216.360 ;
        RECT 793.365 214.100 794.140 214.240 ;
        RECT 723.430 212.720 724.520 213.040 ;
        RECT 727.490 212.450 727.810 213.300 ;
        RECT 769.350 212.450 769.670 213.300 ;
        RECT 775.330 212.450 775.650 213.300 ;
        RECT 781.310 212.450 781.630 213.300 ;
        RECT 787.290 212.450 787.610 213.300 ;
        RECT 794.000 213.040 794.140 214.100 ;
        RECT 2152.880 213.040 2153.020 237.670 ;
        RECT 2153.500 237.430 2153.640 237.525 ;
        RECT 2153.500 237.110 2153.760 237.430 ;
        RECT 2158.860 237.150 2159.000 237.235 ;
        RECT 2153.500 216.360 2153.640 237.110 ;
        RECT 2158.860 236.830 2159.120 237.150 ;
        RECT 2153.420 215.510 2153.740 216.360 ;
        RECT 2158.860 213.040 2159.000 236.830 ;
        RECT 2159.480 236.590 2159.620 236.705 ;
        RECT 2159.480 236.270 2159.740 236.590 ;
        RECT 2164.840 236.310 2164.980 236.395 ;
        RECT 2159.480 216.360 2159.620 236.270 ;
        RECT 2164.840 235.990 2165.100 236.310 ;
        RECT 2159.400 215.510 2159.720 216.360 ;
        RECT 2164.840 213.040 2164.980 235.990 ;
        RECT 2165.460 235.750 2165.600 235.815 ;
        RECT 2165.460 235.430 2165.720 235.750 ;
        RECT 2170.820 235.470 2170.960 235.540 ;
        RECT 2165.460 216.360 2165.600 235.430 ;
        RECT 2170.820 235.150 2171.080 235.470 ;
        RECT 2165.380 215.510 2165.700 216.360 ;
        RECT 2170.820 213.040 2170.960 235.150 ;
        RECT 2171.440 234.910 2171.580 234.990 ;
        RECT 2171.440 234.590 2171.700 234.910 ;
        RECT 2176.800 234.630 2176.940 234.675 ;
        RECT 2171.440 216.360 2171.580 234.590 ;
        RECT 2176.800 234.310 2177.060 234.630 ;
        RECT 2171.360 215.510 2171.680 216.360 ;
        RECT 2176.800 213.040 2176.940 234.310 ;
        RECT 2177.420 234.070 2177.560 234.180 ;
        RECT 2177.420 233.750 2177.680 234.070 ;
        RECT 2182.780 233.790 2182.920 233.845 ;
        RECT 2177.420 216.360 2177.560 233.750 ;
        RECT 2182.780 233.470 2183.040 233.790 ;
        RECT 2177.340 215.510 2177.660 216.360 ;
        RECT 2182.780 213.040 2182.920 233.470 ;
        RECT 2183.400 233.230 2183.540 233.310 ;
        RECT 2183.400 232.910 2183.660 233.230 ;
        RECT 2188.760 232.950 2188.900 233.000 ;
        RECT 2183.400 216.360 2183.540 232.910 ;
        RECT 2188.760 232.630 2189.020 232.950 ;
        RECT 2183.320 215.510 2183.640 216.360 ;
        RECT 2188.760 213.040 2188.900 232.630 ;
        RECT 2189.380 232.390 2189.520 232.485 ;
        RECT 2189.380 232.070 2189.640 232.390 ;
        RECT 2194.740 232.110 2194.880 232.485 ;
        RECT 2189.380 216.360 2189.520 232.070 ;
        RECT 2194.740 231.790 2195.000 232.110 ;
        RECT 2189.300 215.510 2189.620 216.360 ;
        RECT 2194.740 213.040 2194.880 231.790 ;
        RECT 2195.360 231.550 2195.500 232.485 ;
        RECT 2195.360 231.230 2195.620 231.550 ;
        RECT 2200.720 231.270 2200.860 232.485 ;
        RECT 2195.360 216.360 2195.500 231.230 ;
        RECT 2200.720 230.950 2200.980 231.270 ;
        RECT 2195.280 215.510 2195.600 216.360 ;
        RECT 2200.720 213.040 2200.860 230.950 ;
        RECT 2237.220 225.670 2237.360 232.485 ;
        RECT 2237.220 225.350 2237.480 225.670 ;
        RECT 2242.580 225.390 2242.720 232.485 ;
        RECT 2237.220 216.360 2237.360 225.350 ;
        RECT 2242.580 225.070 2242.840 225.390 ;
        RECT 2237.140 215.510 2237.460 216.360 ;
        RECT 2242.580 213.040 2242.720 225.070 ;
        RECT 2243.200 224.830 2243.340 232.485 ;
        RECT 2243.200 224.510 2243.460 224.830 ;
        RECT 2248.560 224.550 2248.700 232.485 ;
        RECT 2243.200 216.360 2243.340 224.510 ;
        RECT 2248.560 224.230 2248.820 224.550 ;
        RECT 2243.120 215.510 2243.440 216.360 ;
        RECT 2248.560 213.040 2248.700 224.230 ;
        RECT 2249.180 223.990 2249.320 232.485 ;
        RECT 2249.180 223.670 2249.440 223.990 ;
        RECT 2254.540 223.710 2254.680 232.485 ;
        RECT 2249.180 216.360 2249.320 223.670 ;
        RECT 2254.540 223.390 2254.800 223.710 ;
        RECT 2249.100 215.510 2249.420 216.360 ;
        RECT 2254.540 213.040 2254.680 223.390 ;
        RECT 2255.160 223.150 2255.300 232.485 ;
        RECT 2255.160 222.830 2255.420 223.150 ;
        RECT 2260.520 222.870 2260.660 232.485 ;
        RECT 2255.160 216.360 2255.300 222.830 ;
        RECT 2260.520 222.550 2260.780 222.870 ;
        RECT 2255.080 215.510 2255.400 216.360 ;
        RECT 2260.520 213.040 2260.660 222.550 ;
        RECT 2261.140 222.310 2261.280 232.485 ;
        RECT 2261.140 221.990 2261.400 222.310 ;
        RECT 2261.140 216.360 2261.280 221.990 ;
        RECT 2266.500 221.750 2266.640 232.485 ;
        RECT 2266.500 221.430 2266.760 221.750 ;
        RECT 2261.060 215.510 2261.380 216.360 ;
        RECT 2266.500 214.170 2266.640 221.430 ;
        RECT 2267.120 221.190 2267.260 232.485 ;
        RECT 2267.120 220.870 2267.380 221.190 ;
        RECT 2267.120 216.360 2267.260 220.870 ;
        RECT 2267.040 215.510 2267.360 216.360 ;
        RECT 2266.500 214.030 2267.275 214.170 ;
        RECT 2267.135 213.300 2267.275 214.030 ;
        RECT 793.340 212.720 794.430 213.040 ;
        RECT 2152.590 212.720 2153.680 213.040 ;
        RECT 2158.570 212.720 2159.660 213.040 ;
        RECT 2164.550 212.720 2165.640 213.040 ;
        RECT 2170.530 212.720 2171.620 213.040 ;
        RECT 2176.510 212.720 2177.600 213.040 ;
        RECT 2182.490 212.720 2183.580 213.040 ;
        RECT 2188.470 212.720 2189.560 213.040 ;
        RECT 2194.450 212.720 2195.540 213.040 ;
        RECT 2200.430 212.720 2201.520 213.040 ;
        RECT 2242.290 212.720 2243.380 213.040 ;
        RECT 2248.270 212.720 2249.360 213.040 ;
        RECT 2254.250 212.720 2255.340 213.040 ;
        RECT 2260.230 212.720 2261.320 213.040 ;
        RECT 2267.050 212.450 2267.370 213.300 ;
  END
END gpio_signal_buffering_alt
END LIBRARY

