magic
tech sky130A
magscale 1 2
timestamp 1686151263
<< checkpaint >>
rect 675396 121665 678085 122078
rect 675258 117277 678085 121665
rect 674508 115475 678085 117277
rect 674508 114693 678023 115475
rect 674516 114683 678023 114693
rect 674516 114672 678018 114683
rect 674516 103443 677084 114672
rect 674514 103440 677086 103443
rect 674514 103439 677088 103440
rect 674509 103379 677091 103439
rect 674509 100863 677215 103379
rect 674512 100696 677215 100863
rect 674516 99196 677084 100696
<< metal1 >>
rect 675768 115959 675774 116011
rect 675826 115959 675832 116011
rect 675682 113371 675734 115709
rect 675586 112665 675638 112671
rect 675586 112487 675638 112493
rect 675490 109630 675542 109636
rect 675490 109452 675542 109458
rect 675492 101631 675540 109452
rect 675588 108347 675636 112487
rect 675682 109050 675734 113199
rect 675586 108341 675638 108347
rect 675586 108163 675638 108169
rect 675490 101625 675542 101631
rect 675490 101567 675542 101573
rect 675492 100265 675540 101567
rect 675588 100462 675636 108163
rect 675586 100456 675638 100462
rect 675586 100278 675638 100284
rect 675588 100265 675636 100278
rect 675682 99896 675734 108866
rect 675776 102183 675824 115959
rect 675774 102177 675826 102183
rect 675774 102119 675826 102125
<< via1 >>
rect 675774 115959 675826 116011
rect 675682 113199 675734 113371
rect 675586 112493 675638 112665
rect 675490 109458 675542 109630
rect 675682 108866 675734 109050
rect 675586 108169 675638 108341
rect 675490 101573 675542 101625
rect 675586 100284 675638 100456
rect 675774 102125 675826 102177
<< metal2 >>
rect 675774 116011 675826 116017
rect 676698 116015 676758 116024
rect 675826 115961 676698 116009
rect 675774 115953 675826 115959
rect 676698 115946 676758 115955
rect 675676 113311 675682 113371
rect 675407 113255 675682 113311
rect 675676 113199 675682 113255
rect 675734 113311 675740 113371
rect 675734 113255 675887 113311
rect 675734 113199 675740 113255
rect 675407 112665 675887 112667
rect 675407 112611 675586 112665
rect 675580 112493 675586 112611
rect 675638 112611 675887 112665
rect 675638 112493 675644 112611
rect 675407 109630 675887 109631
rect 675407 109575 675490 109630
rect 675484 109458 675490 109575
rect 675542 109575 675887 109630
rect 675542 109458 675548 109575
rect 675676 108866 675682 109050
rect 675734 108866 675740 109050
rect 675407 108341 675887 108343
rect 675407 108287 675586 108341
rect 675580 108169 675586 108287
rect 675638 108287 675887 108341
rect 675638 108169 675644 108287
rect 675407 102177 675887 102179
rect 675407 102125 675774 102177
rect 675826 102125 675887 102177
rect 675407 102123 675887 102125
rect 675407 101625 675887 101627
rect 675407 101573 675490 101625
rect 675542 101573 675887 101625
rect 675407 101571 675887 101573
rect 675580 100339 675586 100456
rect 675407 100284 675586 100339
rect 675638 100339 675644 100456
rect 675638 100284 675887 100339
rect 675407 100283 675887 100284
<< via2 >>
rect 676698 115955 676758 116015
<< metal3 >>
rect 676696 116020 676756 117658
rect 676693 116015 676763 116020
rect 676693 115955 676698 116015
rect 676758 115955 676763 116015
rect 676693 115950 676763 115955
rect 676696 115943 676756 115950
<< properties >>
string flatten true
<< end >>
