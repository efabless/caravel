magic
tech sky130A
magscale 1 2
timestamp 1666277172
<< checkpaint >>
rect 39764 415548 677806 997846
<< metal3 >>
tri 81502 983518 82144 984160 se
rect 82144 984060 87144 997762
rect 82144 983518 86502 984060
rect 81502 982718 86502 983518
tri 86502 983418 87144 984060 nw
rect 133544 983518 138544 997772
rect 133502 983382 138544 983518
rect 184944 983518 189944 997736
rect 221000 995620 235279 997736
rect 221000 993820 221400 995620
rect 234879 993820 235279 995620
rect 221000 993420 235279 993820
tri 221000 983518 230902 993420 ne
rect 230902 983518 235279 993420
rect 235579 984141 237779 997736
tri 235579 983518 236202 984141 ne
rect 236202 983518 237779 984141
rect 237978 984242 240178 997736
tri 237978 983868 238352 984242 ne
rect 238352 983868 240178 984242
rect 240478 995620 254800 997736
rect 240478 993820 240878 995620
rect 254357 993820 254800 995620
rect 240478 992116 254800 993820
rect 240478 984242 246202 992116
tri 240478 983868 240852 984242 ne
rect 240852 983868 246202 984242
tri 237779 983518 238129 983868 sw
tri 238352 983518 238702 983868 ne
rect 238702 983518 240178 983868
tri 240178 983518 240528 983868 sw
tri 240852 983518 241202 983868 ne
rect 184944 983452 190502 983518
rect 133502 982718 138502 983382
rect 185502 982718 190502 983452
rect 230902 982718 235902 983518
rect 236202 982718 238402 983518
rect 238702 982718 240902 983518
rect 241202 982718 246202 983868
tri 246202 983518 254800 992116 nw
rect 273600 995620 287879 997754
rect 273600 993820 274000 995620
rect 287479 993820 287879 995620
rect 273600 992520 287879 993820
tri 273600 983518 282602 992520 ne
rect 282602 983795 287879 992520
rect 282602 982718 287602 983795
tri 287602 983518 287879 983795 nw
rect 288179 983795 290379 997754
tri 287979 983518 288179 983718 se
rect 288179 983518 290102 983795
tri 290102 983518 290379 983795 nw
rect 290578 983694 292778 997754
tri 290402 983518 290578 983694 se
rect 290578 983518 292602 983694
tri 292602 983518 292778 983694 nw
rect 293078 995620 307400 997754
rect 293078 993820 293478 995620
rect 306957 993820 307400 995620
rect 293078 993016 307400 993820
rect 293078 983518 297902 993016
tri 297902 983518 307400 993016 nw
rect 375400 995620 389679 997722
rect 375400 993820 375800 995620
rect 389279 993820 389679 995620
rect 375400 992420 389679 993820
tri 375400 983518 384302 992420 ne
rect 384302 983895 389679 992420
rect 287902 982718 290102 983518
rect 290402 982718 292602 983518
rect 292902 982718 297902 983518
rect 384302 982718 389302 983895
tri 389302 983518 389679 983895 nw
rect 389979 983895 392179 997722
tri 389699 983518 389979 983798 se
rect 389979 983794 392078 983895
tri 392078 983794 392179 983895 nw
rect 392378 983794 394578 997722
rect 389979 983518 391802 983794
tri 391802 983518 392078 983794 nw
tri 392102 983518 392378 983794 se
rect 392378 983518 394302 983794
tri 394302 983518 394578 983794 nw
rect 394878 995620 409200 997722
rect 394878 993820 395278 995620
rect 408757 993820 409200 995620
rect 394878 993116 409200 993820
rect 394878 983518 399602 993116
tri 399602 983518 409200 993116 nw
rect 478744 983518 483744 997704
rect 389602 982718 391802 983518
rect 392102 982718 394302 983518
rect 394602 982718 399602 983518
rect 478702 983384 483744 983518
rect 530144 984064 535144 997792
tri 530144 983506 530702 984064 ne
rect 530702 983518 535144 984064
tri 535144 983518 535702 984076 sw
rect 478702 982718 483702 983384
rect 530702 982718 535702 983518
rect 575700 983678 580479 995092
tri 575700 983476 575902 983678 ne
rect 575902 983518 580479 983678
tri 580479 983518 580702 983741 sw
rect 575902 982718 580702 983518
rect 585678 983700 590458 995092
tri 585678 983476 585902 983700 ne
rect 585902 983518 590458 983700
tri 590458 983518 590702 983762 sw
rect 631944 983518 636944 997846
rect 585902 982718 590702 983518
rect 631902 983374 636944 983518
rect 631902 982718 636902 983374
rect 39764 963960 63464 965144
tri 63464 963960 64648 965144 sw
rect 39764 960144 65308 963960
tri 63325 958961 64508 960144 ne
rect 64508 958960 65308 960144
rect 649308 961656 650108 961702
rect 649308 956702 677806 961656
rect 650016 956656 677806 956702
rect 64508 926940 65308 927360
rect 46756 922560 65308 926940
rect 46756 922151 64552 922560
rect 649308 922502 650108 923302
tri 650108 922502 650908 923302 sw
rect 649308 918502 670780 922502
tri 649926 917700 650728 918502 ne
rect 650728 917700 670780 918502
rect 64508 916900 65308 917361
rect 46756 912560 65308 916900
rect 46756 912100 64560 912560
rect 649308 912449 650108 913302
tri 650108 912449 650961 913302 sw
rect 649308 908502 670788 912449
tri 649934 907660 650776 908502 ne
rect 650776 907660 670788 908502
tri 64006 842458 64508 842960 se
rect 64508 842458 65308 842960
rect 49892 838160 65308 842458
rect 49892 837678 64152 838160
tri 64152 837678 64634 838160 nw
rect 649308 833301 650108 834080
tri 64027 832479 64508 832960 se
rect 64508 832479 65308 832960
rect 49892 828160 65308 832479
rect 649308 829280 667192 833301
rect 649858 828521 667192 829280
rect 49892 828159 64634 828160
rect 49892 827699 64174 828159
tri 64174 827699 64634 828159 nw
rect 649308 823322 650108 824080
rect 649308 819280 667192 823322
rect 649858 818542 667192 819280
rect 649308 518701 650108 518748
rect 649308 513948 667116 518701
rect 650058 513921 667116 513948
rect 649308 508722 650108 508748
rect 649308 503948 667124 508722
rect 650066 503942 667124 503948
tri 63960 497858 64508 498406 se
rect 64508 497858 65308 498406
rect 52228 493606 65308 497858
rect 52228 493078 64012 493606
tri 64012 493078 64540 493606 nw
tri 63982 487879 64508 488405 se
rect 64508 487879 65308 488406
rect 52236 483606 65308 487879
rect 52236 483099 64041 483606
tri 64041 483099 64548 483606 nw
rect 649308 474700 650108 474948
rect 649308 470148 670778 474700
rect 650042 469900 670778 470148
rect 649308 464649 650108 464948
rect 649308 460148 670778 464649
rect 650042 459860 670778 460148
tri 63842 455740 64508 456406 se
rect 64508 455740 65308 456406
rect 46742 451606 65308 455740
rect 46742 450951 63927 451606
tri 63927 450951 64582 451606 nw
tri 63802 445700 64508 446406 se
rect 64508 445700 65308 446406
rect 46768 441606 65308 445700
rect 46768 440900 63858 441606
tri 63858 440900 64564 441606 nw
rect 650068 430348 663976 430501
rect 649308 425562 663976 430348
rect 649308 425548 650108 425562
rect 650058 420348 663966 420522
rect 649308 415742 663966 420348
rect 649308 415548 650108 415742
<< via3 >>
rect 221400 993820 234879 995620
rect 240878 993820 254357 995620
rect 274000 993820 287479 995620
rect 293478 993820 306957 995620
rect 375800 993820 389279 995620
rect 395278 993820 408757 995620
<< metal4 >>
rect 221000 995620 235279 996020
rect 221000 993820 221400 995620
rect 234879 993820 235279 995620
rect 221000 993420 235279 993820
tri 221000 983518 230902 993420 ne
rect 230902 983518 235279 993420
rect 240478 995620 254757 996020
rect 240478 993820 240878 995620
rect 254357 993820 254757 995620
rect 273600 995620 287879 996020
rect 273600 993820 274000 995620
rect 287479 993820 287879 995620
rect 240478 992116 254800 993820
rect 240478 984242 246202 992116
tri 240478 983518 241202 984242 ne
rect 230902 982718 235902 983518
rect 241202 982718 246202 984242
tri 246202 983518 254800 992116 nw
rect 273600 992520 287879 993820
tri 273600 983518 282602 992520 ne
rect 282602 983795 287879 992520
rect 282602 982718 287602 983795
tri 287602 983518 287879 983795 nw
rect 293078 995620 307357 996020
rect 293078 993820 293478 995620
rect 306957 993820 307357 995620
rect 375400 995620 389679 996020
rect 375400 993820 375800 995620
rect 389279 993820 389679 995620
rect 293078 993016 307400 993820
rect 293078 983518 297902 993016
tri 297902 983518 307400 993016 nw
rect 375400 992420 389679 993820
tri 375400 983518 384302 992420 ne
rect 384302 983895 389679 992420
rect 292902 982718 297902 983518
rect 384302 982718 389302 983895
tri 389302 983518 389679 983895 nw
rect 394878 995620 409157 996020
rect 394878 993820 395278 995620
rect 408757 993820 409157 995620
rect 394878 993116 409200 993820
rect 394878 983518 399602 993116
tri 399602 983518 409200 993116 nw
rect 394602 982718 399602 983518
<< via4 >>
rect 221400 993820 234879 995620
rect 240878 993820 254357 995620
rect 274000 993820 287479 995620
rect 293478 993820 306957 995620
rect 375800 993820 389279 995620
rect 395278 993820 408757 995620
<< metal5 >>
rect 221000 995620 235279 996020
rect 221000 993820 221400 995620
rect 234879 993820 235279 995620
rect 221000 993420 235279 993820
tri 221000 983518 230902 993420 ne
rect 230902 983518 235279 993420
rect 240478 995620 254757 996020
rect 240478 993820 240878 995620
rect 254357 993820 254757 995620
rect 273600 995620 287879 996020
rect 273600 993820 274000 995620
rect 287479 993820 287879 995620
rect 240478 992116 254800 993820
rect 240478 984242 246202 992116
tri 240478 983518 241202 984242 ne
rect 230902 982718 235902 983518
rect 241202 982718 246202 984242
tri 246202 983518 254800 992116 nw
rect 273600 992520 287879 993820
tri 273600 983518 282602 992520 ne
rect 282602 983795 287879 992520
rect 282602 982718 287602 983795
tri 287602 983518 287879 983795 nw
rect 293078 995620 307357 996020
rect 293078 993820 293478 995620
rect 306957 993820 307357 995620
rect 375400 995620 389679 996020
rect 375400 993820 375800 995620
rect 389279 993820 389679 995620
rect 293078 993016 307400 993820
rect 293078 983518 297902 993016
tri 297902 983518 307400 993016 nw
rect 375400 992420 389679 993820
tri 375400 983518 384302 992420 ne
rect 384302 983895 389679 992420
rect 292902 982718 297902 983518
rect 384302 982718 389302 983895
tri 389302 983518 389679 983895 nw
rect 394878 995620 409157 996020
rect 394878 993820 395278 995620
rect 408757 993820 409157 995620
rect 394878 993116 409200 993820
rect 394878 983518 399602 993116
tri 399602 983518 409200 993116 nw
rect 394602 982718 399602 983518
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
