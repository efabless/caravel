magic
tech sky130A
magscale 1 2
timestamp 1667138844
<< isosubstrate >>
rect 1096 1592 2678 4514
<< viali >>
rect 3433 11849 3467 11883
rect 9137 11781 9171 11815
rect 1409 11713 1443 11747
rect 1593 11713 1627 11747
rect 7941 11713 7975 11747
rect 8769 11713 8803 11747
rect 1685 11645 1719 11679
rect 3617 11645 3651 11679
rect 3801 11645 3835 11679
rect 5917 11645 5951 11679
rect 6193 11645 6227 11679
rect 6347 11645 6381 11679
rect 8493 11645 8527 11679
rect 8953 11645 8987 11679
rect 9443 11645 9477 11679
rect 9597 11645 9631 11679
rect 9873 11645 9907 11679
rect 10057 11645 10091 11679
rect 1225 11577 1259 11611
rect 1961 11577 1995 11611
rect 3985 11577 4019 11611
rect 9689 11577 9723 11611
rect 5089 11509 5123 11543
rect 6561 11509 6595 11543
rect 9229 11509 9263 11543
rect 1593 11305 1627 11339
rect 2145 11305 2179 11339
rect 5929 11237 5963 11271
rect 7389 11237 7423 11271
rect 1225 11169 1259 11203
rect 1318 11169 1352 11203
rect 3433 11169 3467 11203
rect 3525 11169 3559 11203
rect 5365 11169 5399 11203
rect 7573 11169 7607 11203
rect 9413 11169 9447 11203
rect 3893 11101 3927 11135
rect 6193 11101 6227 11135
rect 6929 11101 6963 11135
rect 7113 11101 7147 11135
rect 7941 11101 7975 11135
rect 7297 11033 7331 11067
rect 9977 11033 10011 11067
rect 6837 10965 6871 10999
rect 1409 10761 1443 10795
rect 6009 10761 6043 10795
rect 8769 10761 8803 10795
rect 9965 10761 9999 10795
rect 3433 10693 3467 10727
rect 4261 10625 4295 10659
rect 9321 10625 9355 10659
rect 9505 10625 9539 10659
rect 1225 10557 1259 10591
rect 1379 10557 1413 10591
rect 1685 10557 1719 10591
rect 3801 10557 3835 10591
rect 3894 10557 3928 10591
rect 6101 10557 6135 10591
rect 6469 10557 6503 10591
rect 7941 10557 7975 10591
rect 8505 10557 8539 10591
rect 9689 10557 9723 10591
rect 1961 10489 1995 10523
rect 4537 10489 4571 10523
rect 9873 10489 9907 10523
rect 3709 10421 3743 10455
rect 4169 10421 4203 10455
rect 1409 10217 1443 10251
rect 3433 10217 3467 10251
rect 5929 10217 5963 10251
rect 9597 10149 9631 10183
rect 1593 10081 1627 10115
rect 5365 10081 5399 10115
rect 6285 10081 6319 10115
rect 8861 10081 8895 10115
rect 9872 10081 9906 10115
rect 9965 10081 9999 10115
rect 1685 10013 1719 10047
rect 1961 10013 1995 10047
rect 3525 10013 3559 10047
rect 3893 10013 3927 10047
rect 7021 10013 7055 10047
rect 7389 10013 7423 10047
rect 6929 9877 6963 9911
rect 9425 9877 9459 9911
rect 1409 9605 1443 9639
rect 9689 9605 9723 9639
rect 3433 9537 3467 9571
rect 4261 9537 4295 9571
rect 6837 9537 6871 9571
rect 8585 9537 8619 9571
rect 9229 9537 9263 9571
rect 1593 9469 1627 9503
rect 3617 9469 3651 9503
rect 3893 9469 3927 9503
rect 5733 9469 5767 9503
rect 6561 9469 6595 9503
rect 8983 9469 9017 9503
rect 9137 9469 9171 9503
rect 9413 9469 9447 9503
rect 9873 9469 9907 9503
rect 3157 9401 3191 9435
rect 9597 9401 9631 9435
rect 1685 9333 1719 9367
rect 3709 9333 3743 9367
rect 6297 9333 6331 9367
rect 8769 9333 8803 9367
rect 10057 9333 10091 9367
rect 1317 9129 1351 9163
rect 2145 9061 2179 9095
rect 1409 8993 1443 9027
rect 3985 8993 4019 9027
rect 4077 8993 4111 9027
rect 6009 8993 6043 9027
rect 6745 8993 6779 9027
rect 6929 8993 6963 9027
rect 7022 8993 7056 9027
rect 8217 8993 8251 9027
rect 9689 8993 9723 9027
rect 1593 8925 1627 8959
rect 7297 8925 7331 8959
rect 10057 8925 10091 8959
rect 7481 8857 7515 8891
rect 2697 8789 2731 8823
rect 6193 8789 6227 8823
rect 7652 8789 7686 8823
rect 1501 8585 1535 8619
rect 4261 8585 4295 8619
rect 3433 8449 3467 8483
rect 1685 8381 1719 8415
rect 3617 8381 3651 8415
rect 4353 8381 4387 8415
rect 4537 8381 4571 8415
rect 4813 8381 4847 8415
rect 6561 8381 6595 8415
rect 8585 8381 8619 8415
rect 8769 8381 8803 8415
rect 8953 8381 8987 8415
rect 9229 8381 9263 8415
rect 9322 8381 9356 8415
rect 9689 8381 9723 8415
rect 9873 8381 9907 8415
rect 1409 8313 1443 8347
rect 4721 8313 4755 8347
rect 9137 8313 9171 8347
rect 9597 8313 9631 8347
rect 10057 8313 10091 8347
rect 7665 8245 7699 8279
rect 1501 8041 1535 8075
rect 6837 8041 6871 8075
rect 1409 7973 1443 8007
rect 3341 7973 3375 8007
rect 1685 7905 1719 7939
rect 3893 7905 3927 7939
rect 5365 7905 5399 7939
rect 6929 7905 6963 7939
rect 7297 7905 7331 7939
rect 8769 7905 8803 7939
rect 3525 7837 3559 7871
rect 6285 7837 6319 7871
rect 9505 7837 9539 7871
rect 9781 7769 9815 7803
rect 5925 7701 5959 7735
rect 9329 7701 9363 7735
rect 9965 7701 9999 7735
rect 1409 7497 1443 7531
rect 8953 7497 8987 7531
rect 9229 7429 9263 7463
rect 3617 7361 3651 7395
rect 7941 7361 7975 7395
rect 1500 7293 1534 7327
rect 1593 7293 1627 7327
rect 3433 7293 3467 7327
rect 4353 7293 4387 7327
rect 6561 7293 6595 7327
rect 8585 7293 8619 7327
rect 8861 7293 8895 7327
rect 9505 7293 9539 7327
rect 9781 7293 9815 7327
rect 4445 7225 4479 7259
rect 9689 7225 9723 7259
rect 2145 7157 2179 7191
rect 4261 7157 4295 7191
rect 5641 7157 5675 7191
rect 9965 7157 9999 7191
rect 6929 6953 6963 6987
rect 9137 6953 9171 6987
rect 1409 6885 1443 6919
rect 1685 6817 1719 6851
rect 3433 6817 3467 6851
rect 3525 6817 3559 6851
rect 5365 6817 5399 6851
rect 7113 6817 7147 6851
rect 7481 6817 7515 6851
rect 8953 6817 8987 6851
rect 3893 6749 3927 6783
rect 6193 6749 6227 6783
rect 6837 6749 6871 6783
rect 9689 6749 9723 6783
rect 9873 6749 9907 6783
rect 1501 6613 1535 6647
rect 5929 6613 5963 6647
rect 9513 6613 9547 6647
rect 10057 6613 10091 6647
rect 5365 6409 5399 6443
rect 8769 6341 8803 6375
rect 9137 6341 9171 6375
rect 1685 6273 1719 6307
rect 3893 6273 3927 6307
rect 5825 6273 5859 6307
rect 9965 6273 9999 6307
rect 1409 6205 1443 6239
rect 3617 6205 3651 6239
rect 5457 6205 5491 6239
rect 7297 6205 7331 6239
rect 8033 6205 8067 6239
rect 8217 6205 8251 6239
rect 9137 6205 9171 6239
rect 9505 6205 9539 6239
rect 1961 6137 1995 6171
rect 8493 6137 8527 6171
rect 8585 6137 8619 6171
rect 1501 6069 1535 6103
rect 3433 6069 3467 6103
rect 7857 6069 7891 6103
rect 1409 5865 1443 5899
rect 7665 5865 7699 5899
rect 1961 5797 1995 5831
rect 4261 5797 4295 5831
rect 6561 5797 6595 5831
rect 9689 5797 9723 5831
rect 1501 5729 1535 5763
rect 3617 5729 3651 5763
rect 4169 5729 4203 5763
rect 6193 5729 6227 5763
rect 8585 5729 8619 5763
rect 10057 5729 10091 5763
rect 1685 5661 1719 5695
rect 3801 5661 3835 5695
rect 3985 5661 4019 5695
rect 6009 5661 6043 5695
rect 6377 5661 6411 5695
rect 9413 5661 9447 5695
rect 3433 5593 3467 5627
rect 8769 5593 8803 5627
rect 9505 5593 9539 5627
rect 9689 5525 9723 5559
rect 3525 5321 3559 5355
rect 5917 5321 5951 5355
rect 10057 5321 10091 5355
rect 3801 5185 3835 5219
rect 8033 5185 8067 5219
rect 3341 5117 3375 5151
rect 3495 5117 3529 5151
rect 6101 5117 6135 5151
rect 8309 5117 8343 5151
rect 4077 5049 4111 5083
rect 5825 5049 5859 5083
rect 5549 4981 5583 5015
rect 3985 4777 4019 4811
rect 4169 4777 4203 4811
rect 6929 4777 6963 4811
rect 7573 4777 7607 4811
rect 8125 4777 8159 4811
rect 10057 4777 10091 4811
rect 3433 4641 3467 4675
rect 4261 4641 4295 4675
rect 6193 4641 6227 4675
rect 7143 4641 7177 4675
rect 7297 4641 7331 4675
rect 7483 4641 7517 4675
rect 7757 4641 7791 4675
rect 7911 4641 7945 4675
rect 8309 4641 8343 4675
rect 4353 4573 4387 4607
rect 4721 4573 4755 4607
rect 8585 4573 8619 4607
rect 6753 4437 6787 4471
rect 5365 4233 5399 4267
rect 5733 4233 5767 4267
rect 3341 4097 3375 4131
rect 5089 4097 5123 4131
rect 6929 4097 6963 4131
rect 7389 4097 7423 4131
rect 5181 4029 5215 4063
rect 5335 4029 5369 4063
rect 6285 4029 6319 4063
rect 6837 4029 6871 4063
rect 3617 3961 3651 3995
rect 6653 3961 6687 3995
rect 7205 3961 7239 3995
rect 6561 3893 6595 3927
rect 3341 3689 3375 3723
rect 6009 3689 6043 3723
rect 7205 3689 7239 3723
rect 8493 3689 8527 3723
rect 9965 3689 9999 3723
rect 4813 3621 4847 3655
rect 5089 3553 5123 3587
rect 5917 3553 5951 3587
rect 8125 3553 8159 3587
rect 8401 3553 8435 3587
rect 8861 3553 8895 3587
rect 9045 3553 9079 3587
rect 9229 3553 9263 3587
rect 9505 3553 9539 3587
rect 9873 3553 9907 3587
rect 5733 3485 5767 3519
rect 9321 3485 9355 3519
rect 5181 3349 5215 3383
rect 9689 3349 9723 3383
rect 3341 3145 3375 3179
rect 5273 3145 5307 3179
rect 10057 3145 10091 3179
rect 5733 3077 5767 3111
rect 5089 3009 5123 3043
rect 7389 3009 7423 3043
rect 5917 2941 5951 2975
rect 8033 2941 8067 2975
rect 8493 2941 8527 2975
rect 4813 2873 4847 2907
rect 5365 2873 5399 2907
rect 4261 2601 4295 2635
rect 5273 2601 5307 2635
rect 5549 2601 5583 2635
rect 6009 2601 6043 2635
rect 8401 2601 8435 2635
rect 8677 2601 8711 2635
rect 9413 2601 9447 2635
rect 9781 2601 9815 2635
rect 3801 2533 3835 2567
rect 4169 2533 4203 2567
rect 5825 2533 5859 2567
rect 9137 2533 9171 2567
rect 3433 2465 3467 2499
rect 4629 2465 4663 2499
rect 4905 2465 4939 2499
rect 5365 2465 5399 2499
rect 5641 2465 5675 2499
rect 5917 2465 5951 2499
rect 6561 2465 6595 2499
rect 8493 2465 8527 2499
rect 8769 2465 8803 2499
rect 9505 2465 9539 2499
rect 9873 2465 9907 2499
rect 4445 2397 4479 2431
rect 8125 2329 8159 2363
rect 3525 2261 3559 2295
rect 3893 2261 3927 2295
rect 4997 2261 5031 2295
rect 9045 2261 9079 2295
rect 3893 2057 3927 2091
rect 4261 2057 4295 2091
rect 4813 2057 4847 2091
rect 5365 2057 5399 2091
rect 5457 2057 5491 2091
rect 5825 2057 5859 2091
rect 6009 2057 6043 2091
rect 4537 1989 4571 2023
rect 5089 1989 5123 2023
rect 6929 1989 6963 2023
rect 9413 1921 9447 1955
rect 3801 1853 3835 1887
rect 4077 1853 4111 1887
rect 4629 1853 4663 1887
rect 4905 1853 4939 1887
rect 5181 1853 5215 1887
rect 7941 1853 7975 1887
rect 9781 1853 9815 1887
rect 3433 1785 3467 1819
rect 3525 1717 3559 1751
rect 4077 1513 4111 1547
rect 5181 1513 5215 1547
rect 8125 1513 8159 1547
rect 9229 1445 9263 1479
rect 9413 1445 9447 1479
rect 9689 1445 9723 1479
rect 3893 1377 3927 1411
rect 6101 1377 6135 1411
rect 6285 1377 6319 1411
rect 8585 1377 8619 1411
rect 9873 1377 9907 1411
rect 3341 1309 3375 1343
rect 8769 1309 8803 1343
rect 9597 1241 9631 1275
rect 3525 1173 3559 1207
rect 8309 1173 8343 1207
rect 8861 1173 8895 1207
rect 9045 1173 9079 1207
rect 1501 969 1535 1003
rect 2513 969 2547 1003
rect 2881 969 2915 1003
rect 3065 969 3099 1003
rect 3249 969 3283 1003
rect 3709 969 3743 1003
rect 3985 969 4019 1003
rect 5089 969 5123 1003
rect 9229 969 9263 1003
rect 9689 969 9723 1003
rect 1685 901 1719 935
rect 2329 901 2363 935
rect 3433 901 3467 935
rect 6193 901 6227 935
rect 7665 901 7699 935
rect 1409 765 1443 799
rect 1869 765 1903 799
rect 2605 765 2639 799
rect 6009 765 6043 799
rect 8585 765 8619 799
rect 8769 765 8803 799
rect 9597 765 9631 799
rect 2145 697 2179 731
rect 9873 697 9907 731
rect 6377 629 6411 663
rect 9045 629 9079 663
<< metal1 >>
rect 1026 12384 1032 12436
rect 1084 12424 1090 12436
rect 8754 12424 8760 12436
rect 1084 12396 8760 12424
rect 1084 12384 1090 12396
rect 8754 12384 8760 12396
rect 8812 12384 8818 12436
rect 2406 12180 2412 12232
rect 2464 12220 2470 12232
rect 6178 12220 6184 12232
rect 2464 12192 6184 12220
rect 2464 12180 2470 12192
rect 6178 12180 6184 12192
rect 6236 12180 6242 12232
rect 3694 12112 3700 12164
rect 3752 12152 3758 12164
rect 7098 12152 7104 12164
rect 3752 12124 7104 12152
rect 3752 12112 3758 12124
rect 7098 12112 7104 12124
rect 7156 12112 7162 12164
rect 5902 12044 5908 12096
rect 5960 12084 5966 12096
rect 10502 12084 10508 12096
rect 5960 12056 10508 12084
rect 5960 12044 5966 12056
rect 10502 12044 10508 12056
rect 10560 12044 10566 12096
rect 920 11994 10396 12016
rect 920 11942 2566 11994
rect 2618 11942 2630 11994
rect 2682 11942 2694 11994
rect 2746 11942 2758 11994
rect 2810 11942 2822 11994
rect 2874 11942 7566 11994
rect 7618 11942 7630 11994
rect 7682 11942 7694 11994
rect 7746 11942 7758 11994
rect 7810 11942 7822 11994
rect 7874 11942 10396 11994
rect 920 11920 10396 11942
rect 3421 11883 3479 11889
rect 1320 11852 3372 11880
rect 1320 11744 1348 11852
rect 3344 11812 3372 11852
rect 3421 11849 3433 11883
rect 3467 11880 3479 11883
rect 9306 11880 9312 11892
rect 3467 11852 9312 11880
rect 3467 11849 3479 11852
rect 3421 11843 3479 11849
rect 9306 11840 9312 11852
rect 9364 11840 9370 11892
rect 5442 11812 5448 11824
rect 1596 11784 1808 11812
rect 3344 11784 5448 11812
rect 1596 11753 1624 11784
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 1320 11716 1409 11744
rect 1397 11713 1409 11716
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 1581 11747 1639 11753
rect 1581 11713 1593 11747
rect 1627 11713 1639 11747
rect 1780 11744 1808 11784
rect 5442 11772 5448 11784
rect 5500 11772 5506 11824
rect 5534 11772 5540 11824
rect 5592 11812 5598 11824
rect 9125 11815 9183 11821
rect 9125 11812 9137 11815
rect 5592 11784 9137 11812
rect 5592 11772 5598 11784
rect 9125 11781 9137 11784
rect 9171 11781 9183 11815
rect 9125 11775 9183 11781
rect 7926 11744 7932 11756
rect 1780 11716 6132 11744
rect 1581 11707 1639 11713
rect 1670 11676 1676 11688
rect 1631 11648 1676 11676
rect 1670 11636 1676 11648
rect 1728 11636 1734 11688
rect 3510 11636 3516 11688
rect 3568 11676 3574 11688
rect 3605 11679 3663 11685
rect 3605 11676 3617 11679
rect 3568 11648 3617 11676
rect 3568 11636 3574 11648
rect 3605 11645 3617 11648
rect 3651 11645 3663 11679
rect 3605 11639 3663 11645
rect 1210 11608 1216 11620
rect 1171 11580 1216 11608
rect 1210 11568 1216 11580
rect 1268 11568 1274 11620
rect 1946 11608 1952 11620
rect 1907 11580 1952 11608
rect 1946 11568 1952 11580
rect 2004 11568 2010 11620
rect 2406 11568 2412 11620
rect 2464 11568 2470 11620
rect 3620 11608 3648 11639
rect 3694 11636 3700 11688
rect 3752 11676 3758 11688
rect 3789 11679 3847 11685
rect 3789 11676 3801 11679
rect 3752 11648 3801 11676
rect 3752 11636 3758 11648
rect 3789 11645 3801 11648
rect 3835 11645 3847 11679
rect 3789 11639 3847 11645
rect 4062 11636 4068 11688
rect 4120 11676 4126 11688
rect 5902 11676 5908 11688
rect 4120 11648 5580 11676
rect 5863 11648 5908 11676
rect 4120 11636 4126 11648
rect 3878 11608 3884 11620
rect 3344 11580 3556 11608
rect 3620 11580 3884 11608
rect 1578 11500 1584 11552
rect 1636 11540 1642 11552
rect 3344 11540 3372 11580
rect 1636 11512 3372 11540
rect 3528 11540 3556 11580
rect 3878 11568 3884 11580
rect 3936 11568 3942 11620
rect 3973 11611 4031 11617
rect 3973 11577 3985 11611
rect 4019 11608 4031 11611
rect 4890 11608 4896 11620
rect 4019 11580 4896 11608
rect 4019 11577 4031 11580
rect 3973 11571 4031 11577
rect 4890 11568 4896 11580
rect 4948 11568 4954 11620
rect 4154 11540 4160 11552
rect 3528 11512 4160 11540
rect 1636 11500 1642 11512
rect 4154 11500 4160 11512
rect 4212 11500 4218 11552
rect 5077 11543 5135 11549
rect 5077 11509 5089 11543
rect 5123 11540 5135 11543
rect 5442 11540 5448 11552
rect 5123 11512 5448 11540
rect 5123 11509 5135 11512
rect 5077 11503 5135 11509
rect 5442 11500 5448 11512
rect 5500 11500 5506 11552
rect 5552 11540 5580 11648
rect 5902 11636 5908 11648
rect 5960 11636 5966 11688
rect 6104 11608 6132 11716
rect 6196 11716 6960 11744
rect 7887 11716 7932 11744
rect 6196 11688 6224 11716
rect 6178 11636 6184 11688
rect 6236 11676 6242 11688
rect 6362 11685 6368 11688
rect 6335 11679 6368 11685
rect 6236 11648 6281 11676
rect 6236 11636 6242 11648
rect 6335 11645 6347 11679
rect 6335 11639 6368 11645
rect 6362 11636 6368 11639
rect 6420 11636 6426 11688
rect 6932 11676 6960 11716
rect 7926 11704 7932 11716
rect 7984 11704 7990 11756
rect 8754 11744 8760 11756
rect 8036 11716 8616 11744
rect 8715 11716 8760 11744
rect 8036 11676 8064 11716
rect 8478 11676 8484 11688
rect 6932 11648 8064 11676
rect 8439 11648 8484 11676
rect 8478 11636 8484 11648
rect 8536 11636 8542 11688
rect 8588 11676 8616 11716
rect 8754 11704 8760 11716
rect 8812 11704 8818 11756
rect 9950 11744 9956 11756
rect 8956 11716 9956 11744
rect 8956 11685 8984 11716
rect 9950 11704 9956 11716
rect 10008 11704 10014 11756
rect 8941 11679 8999 11685
rect 8941 11676 8953 11679
rect 8588 11648 8953 11676
rect 8941 11645 8953 11648
rect 8987 11645 8999 11679
rect 8941 11639 8999 11645
rect 9431 11679 9489 11685
rect 9431 11645 9443 11679
rect 9477 11645 9489 11679
rect 9431 11639 9489 11645
rect 9585 11679 9643 11685
rect 9585 11645 9597 11679
rect 9631 11676 9643 11679
rect 9858 11676 9864 11688
rect 9631 11648 9864 11676
rect 9631 11645 9643 11648
rect 9585 11639 9643 11645
rect 8110 11608 8116 11620
rect 6104 11580 8116 11608
rect 8110 11568 8116 11580
rect 8168 11608 8174 11620
rect 9446 11608 9474 11639
rect 9858 11636 9864 11648
rect 9916 11636 9922 11688
rect 10045 11679 10103 11685
rect 10045 11645 10057 11679
rect 10091 11676 10103 11679
rect 10226 11676 10232 11688
rect 10091 11648 10232 11676
rect 10091 11645 10103 11648
rect 10045 11639 10103 11645
rect 10226 11636 10232 11648
rect 10284 11636 10290 11688
rect 8168 11580 9474 11608
rect 9677 11611 9735 11617
rect 8168 11568 8174 11580
rect 9677 11577 9689 11611
rect 9723 11608 9735 11611
rect 9766 11608 9772 11620
rect 9723 11580 9772 11608
rect 9723 11577 9735 11580
rect 9677 11571 9735 11577
rect 9766 11568 9772 11580
rect 9824 11568 9830 11620
rect 6454 11540 6460 11552
rect 5552 11512 6460 11540
rect 6454 11500 6460 11512
rect 6512 11500 6518 11552
rect 6549 11543 6607 11549
rect 6549 11509 6561 11543
rect 6595 11540 6607 11543
rect 6914 11540 6920 11552
rect 6595 11512 6920 11540
rect 6595 11509 6607 11512
rect 6549 11503 6607 11509
rect 6914 11500 6920 11512
rect 6972 11500 6978 11552
rect 7006 11500 7012 11552
rect 7064 11540 7070 11552
rect 9030 11540 9036 11552
rect 7064 11512 9036 11540
rect 7064 11500 7070 11512
rect 9030 11500 9036 11512
rect 9088 11500 9094 11552
rect 9214 11540 9220 11552
rect 9175 11512 9220 11540
rect 9214 11500 9220 11512
rect 9272 11500 9278 11552
rect 920 11450 10396 11472
rect 920 11398 5066 11450
rect 5118 11398 5130 11450
rect 5182 11398 5194 11450
rect 5246 11398 5258 11450
rect 5310 11398 5322 11450
rect 5374 11398 10396 11450
rect 920 11376 10396 11398
rect 1578 11336 1584 11348
rect 1539 11308 1584 11336
rect 1578 11296 1584 11308
rect 1636 11296 1642 11348
rect 2133 11339 2191 11345
rect 2133 11305 2145 11339
rect 2179 11336 2191 11339
rect 2179 11308 16574 11336
rect 2179 11305 2191 11308
rect 2133 11299 2191 11305
rect 4246 11228 4252 11280
rect 4304 11228 4310 11280
rect 5917 11271 5975 11277
rect 5917 11237 5929 11271
rect 5963 11268 5975 11271
rect 7006 11268 7012 11280
rect 5963 11240 7012 11268
rect 5963 11237 5975 11240
rect 5917 11231 5975 11237
rect 7006 11228 7012 11240
rect 7064 11228 7070 11280
rect 7098 11228 7104 11280
rect 7156 11268 7162 11280
rect 7377 11271 7435 11277
rect 7377 11268 7389 11271
rect 7156 11240 7389 11268
rect 7156 11228 7162 11240
rect 7377 11237 7389 11240
rect 7423 11237 7435 11271
rect 9214 11268 9220 11280
rect 9062 11240 9220 11268
rect 7377 11231 7435 11237
rect 9214 11228 9220 11240
rect 9272 11228 9278 11280
rect 1210 11200 1216 11212
rect 1171 11172 1216 11200
rect 1210 11160 1216 11172
rect 1268 11160 1274 11212
rect 1306 11203 1364 11209
rect 1306 11169 1318 11203
rect 1352 11169 1364 11203
rect 1306 11163 1364 11169
rect 1026 11092 1032 11144
rect 1084 11132 1090 11144
rect 1320 11132 1348 11163
rect 1762 11160 1768 11212
rect 1820 11200 1826 11212
rect 2406 11200 2412 11212
rect 1820 11172 2412 11200
rect 1820 11160 1826 11172
rect 2406 11160 2412 11172
rect 2464 11160 2470 11212
rect 3421 11203 3479 11209
rect 3421 11169 3433 11203
rect 3467 11169 3479 11203
rect 3421 11163 3479 11169
rect 3513 11203 3571 11209
rect 3513 11169 3525 11203
rect 3559 11200 3571 11203
rect 3559 11172 4016 11200
rect 3559 11169 3571 11172
rect 3513 11163 3571 11169
rect 1084 11104 1348 11132
rect 1084 11092 1090 11104
rect 3436 11064 3464 11163
rect 3786 11092 3792 11144
rect 3844 11132 3850 11144
rect 3881 11135 3939 11141
rect 3881 11132 3893 11135
rect 3844 11104 3893 11132
rect 3844 11092 3850 11104
rect 3881 11101 3893 11104
rect 3927 11101 3939 11135
rect 3988 11132 4016 11172
rect 4890 11160 4896 11212
rect 4948 11200 4954 11212
rect 5353 11203 5411 11209
rect 5353 11200 5365 11203
rect 4948 11172 5365 11200
rect 4948 11160 4954 11172
rect 5353 11169 5365 11172
rect 5399 11169 5411 11203
rect 5353 11163 5411 11169
rect 6822 11160 6828 11212
rect 6880 11200 6886 11212
rect 7561 11203 7619 11209
rect 6880 11172 7236 11200
rect 6880 11160 6886 11172
rect 4522 11132 4528 11144
rect 3988 11104 4528 11132
rect 3881 11095 3939 11101
rect 4522 11092 4528 11104
rect 4580 11092 4586 11144
rect 6178 11132 6184 11144
rect 6139 11104 6184 11132
rect 6178 11092 6184 11104
rect 6236 11092 6242 11144
rect 6454 11092 6460 11144
rect 6512 11132 6518 11144
rect 6917 11135 6975 11141
rect 6917 11132 6929 11135
rect 6512 11104 6929 11132
rect 6512 11092 6518 11104
rect 6917 11101 6929 11104
rect 6963 11101 6975 11135
rect 7098 11132 7104 11144
rect 7059 11104 7104 11132
rect 6917 11095 6975 11101
rect 7098 11092 7104 11104
rect 7156 11092 7162 11144
rect 7208 11132 7236 11172
rect 7561 11169 7573 11203
rect 7607 11200 7619 11203
rect 7607 11172 8064 11200
rect 7607 11169 7619 11172
rect 7561 11163 7619 11169
rect 7929 11135 7987 11141
rect 7929 11132 7941 11135
rect 7208 11104 7941 11132
rect 7929 11101 7941 11104
rect 7975 11101 7987 11135
rect 8036 11132 8064 11172
rect 9122 11160 9128 11212
rect 9180 11200 9186 11212
rect 9401 11203 9459 11209
rect 9401 11200 9413 11203
rect 9180 11172 9413 11200
rect 9180 11160 9186 11172
rect 9401 11169 9413 11172
rect 9447 11169 9459 11203
rect 9401 11163 9459 11169
rect 8386 11132 8392 11144
rect 8036 11104 8392 11132
rect 7929 11095 7987 11101
rect 8386 11092 8392 11104
rect 8444 11092 8450 11144
rect 16546 11076 16574 11308
rect 3436 11036 3648 11064
rect 1486 10956 1492 11008
rect 1544 10996 1550 11008
rect 3510 10996 3516 11008
rect 1544 10968 3516 10996
rect 1544 10956 1550 10968
rect 3510 10956 3516 10968
rect 3568 10956 3574 11008
rect 3620 10996 3648 11036
rect 5718 11024 5724 11076
rect 5776 11064 5782 11076
rect 7285 11067 7343 11073
rect 7285 11064 7297 11067
rect 5776 11036 7297 11064
rect 5776 11024 5782 11036
rect 7285 11033 7297 11036
rect 7331 11033 7343 11067
rect 7285 11027 7343 11033
rect 9965 11067 10023 11073
rect 9965 11033 9977 11067
rect 10011 11064 10023 11067
rect 10410 11064 10416 11076
rect 10011 11036 10416 11064
rect 10011 11033 10023 11036
rect 9965 11027 10023 11033
rect 10410 11024 10416 11036
rect 10468 11024 10474 11076
rect 16546 11036 16580 11076
rect 16574 11024 16580 11036
rect 16632 11024 16638 11076
rect 4430 10996 4436 11008
rect 3620 10968 4436 10996
rect 4430 10956 4436 10968
rect 4488 10956 4494 11008
rect 4522 10956 4528 11008
rect 4580 10996 4586 11008
rect 4798 10996 4804 11008
rect 4580 10968 4804 10996
rect 4580 10956 4586 10968
rect 4798 10956 4804 10968
rect 4856 10956 4862 11008
rect 6825 10999 6883 11005
rect 6825 10965 6837 10999
rect 6871 10996 6883 10999
rect 7190 10996 7196 11008
rect 6871 10968 7196 10996
rect 6871 10965 6883 10968
rect 6825 10959 6883 10965
rect 7190 10956 7196 10968
rect 7248 10956 7254 11008
rect 920 10906 10396 10928
rect 920 10854 2566 10906
rect 2618 10854 2630 10906
rect 2682 10854 2694 10906
rect 2746 10854 2758 10906
rect 2810 10854 2822 10906
rect 2874 10854 7566 10906
rect 7618 10854 7630 10906
rect 7682 10854 7694 10906
rect 7746 10854 7758 10906
rect 7810 10854 7822 10906
rect 7874 10854 10396 10906
rect 920 10832 10396 10854
rect 1397 10795 1455 10801
rect 1397 10761 1409 10795
rect 1443 10792 1455 10795
rect 4246 10792 4252 10804
rect 1443 10764 4252 10792
rect 1443 10761 1455 10764
rect 1397 10755 1455 10761
rect 4246 10752 4252 10764
rect 4304 10752 4310 10804
rect 4706 10752 4712 10804
rect 4764 10792 4770 10804
rect 5902 10792 5908 10804
rect 4764 10764 5908 10792
rect 4764 10752 4770 10764
rect 5902 10752 5908 10764
rect 5960 10752 5966 10804
rect 5997 10795 6055 10801
rect 5997 10761 6009 10795
rect 6043 10792 6055 10795
rect 6178 10792 6184 10804
rect 6043 10764 6184 10792
rect 6043 10761 6055 10764
rect 5997 10755 6055 10761
rect 6178 10752 6184 10764
rect 6236 10752 6242 10804
rect 6454 10752 6460 10804
rect 6512 10792 6518 10804
rect 8757 10795 8815 10801
rect 8757 10792 8769 10795
rect 6512 10764 8769 10792
rect 6512 10752 6518 10764
rect 8757 10761 8769 10764
rect 8803 10761 8815 10795
rect 9950 10792 9956 10804
rect 9911 10764 9956 10792
rect 8757 10755 8815 10761
rect 9950 10752 9956 10764
rect 10008 10752 10014 10804
rect 3421 10727 3479 10733
rect 3421 10693 3433 10727
rect 3467 10724 3479 10727
rect 3467 10696 4384 10724
rect 3467 10693 3479 10696
rect 3421 10687 3479 10693
rect 4249 10659 4307 10665
rect 4249 10656 4261 10659
rect 1688 10628 4261 10656
rect 1688 10600 1716 10628
rect 4249 10625 4261 10628
rect 4295 10625 4307 10659
rect 4356 10656 4384 10696
rect 7374 10684 7380 10736
rect 7432 10724 7438 10736
rect 7432 10696 9536 10724
rect 7432 10684 7438 10696
rect 6730 10656 6736 10668
rect 4356 10628 6736 10656
rect 4249 10619 4307 10625
rect 6730 10616 6736 10628
rect 6788 10616 6794 10668
rect 9306 10656 9312 10668
rect 9267 10628 9312 10656
rect 9306 10616 9312 10628
rect 9364 10616 9370 10668
rect 9508 10665 9536 10696
rect 9493 10659 9551 10665
rect 9493 10625 9505 10659
rect 9539 10625 9551 10659
rect 9493 10619 9551 10625
rect 1210 10588 1216 10600
rect 1171 10560 1216 10588
rect 1210 10548 1216 10560
rect 1268 10548 1274 10600
rect 1367 10591 1425 10597
rect 1367 10557 1379 10591
rect 1413 10588 1425 10591
rect 1486 10588 1492 10600
rect 1413 10560 1492 10588
rect 1413 10557 1425 10560
rect 1367 10551 1425 10557
rect 1486 10548 1492 10560
rect 1544 10548 1550 10600
rect 1670 10588 1676 10600
rect 1631 10560 1676 10588
rect 1670 10548 1676 10560
rect 1728 10548 1734 10600
rect 3694 10588 3700 10600
rect 3344 10560 3700 10588
rect 1949 10523 2007 10529
rect 1949 10489 1961 10523
rect 1995 10520 2007 10523
rect 2038 10520 2044 10532
rect 1995 10492 2044 10520
rect 1995 10489 2007 10492
rect 1949 10483 2007 10489
rect 2038 10480 2044 10492
rect 2096 10480 2102 10532
rect 2148 10492 2438 10520
rect 1486 10412 1492 10464
rect 1544 10452 1550 10464
rect 2148 10452 2176 10492
rect 1544 10424 2176 10452
rect 1544 10412 1550 10424
rect 2958 10412 2964 10464
rect 3016 10452 3022 10464
rect 3344 10452 3372 10560
rect 3694 10548 3700 10560
rect 3752 10588 3758 10600
rect 3789 10591 3847 10597
rect 3789 10588 3801 10591
rect 3752 10560 3801 10588
rect 3752 10548 3758 10560
rect 3789 10557 3801 10560
rect 3835 10557 3847 10591
rect 3789 10551 3847 10557
rect 3882 10591 3940 10597
rect 3882 10557 3894 10591
rect 3928 10588 3940 10591
rect 4062 10588 4068 10600
rect 3928 10560 4068 10588
rect 3928 10557 3940 10560
rect 3882 10551 3940 10557
rect 3418 10480 3424 10532
rect 3476 10520 3482 10532
rect 3896 10520 3924 10551
rect 4062 10548 4068 10560
rect 4120 10548 4126 10600
rect 5626 10548 5632 10600
rect 5684 10548 5690 10600
rect 6086 10588 6092 10600
rect 6047 10560 6092 10588
rect 6086 10548 6092 10560
rect 6144 10548 6150 10600
rect 6454 10588 6460 10600
rect 6415 10560 6460 10588
rect 6454 10548 6460 10560
rect 6512 10548 6518 10600
rect 7929 10591 7987 10597
rect 7929 10557 7941 10591
rect 7975 10557 7987 10591
rect 7929 10551 7987 10557
rect 8493 10591 8551 10597
rect 8493 10557 8505 10591
rect 8539 10588 8551 10591
rect 9214 10588 9220 10600
rect 8539 10560 9220 10588
rect 8539 10557 8551 10560
rect 8493 10551 8551 10557
rect 3476 10492 3924 10520
rect 4525 10523 4583 10529
rect 3476 10480 3482 10492
rect 4525 10489 4537 10523
rect 4571 10520 4583 10523
rect 4571 10492 4936 10520
rect 4571 10489 4583 10492
rect 4525 10483 4583 10489
rect 3016 10424 3372 10452
rect 3697 10455 3755 10461
rect 3016 10412 3022 10424
rect 3697 10421 3709 10455
rect 3743 10452 3755 10455
rect 4062 10452 4068 10464
rect 3743 10424 4068 10452
rect 3743 10421 3755 10424
rect 3697 10415 3755 10421
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 4157 10455 4215 10461
rect 4157 10421 4169 10455
rect 4203 10452 4215 10455
rect 4706 10452 4712 10464
rect 4203 10424 4712 10452
rect 4203 10421 4215 10424
rect 4157 10415 4215 10421
rect 4706 10412 4712 10424
rect 4764 10412 4770 10464
rect 4908 10452 4936 10492
rect 6914 10480 6920 10532
rect 6972 10480 6978 10532
rect 7944 10520 7972 10551
rect 9214 10548 9220 10560
rect 9272 10548 9278 10600
rect 9677 10591 9735 10597
rect 9677 10557 9689 10591
rect 9723 10588 9735 10591
rect 9950 10588 9956 10600
rect 9723 10560 9956 10588
rect 9723 10557 9735 10560
rect 9677 10551 9735 10557
rect 9950 10548 9956 10560
rect 10008 10548 10014 10600
rect 9861 10523 9919 10529
rect 9861 10520 9873 10523
rect 7944 10492 9873 10520
rect 9861 10489 9873 10492
rect 9907 10489 9919 10523
rect 9861 10483 9919 10489
rect 7374 10452 7380 10464
rect 4908 10424 7380 10452
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 7466 10412 7472 10464
rect 7524 10452 7530 10464
rect 9950 10452 9956 10464
rect 7524 10424 9956 10452
rect 7524 10412 7530 10424
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 920 10362 10396 10384
rect 920 10310 5066 10362
rect 5118 10310 5130 10362
rect 5182 10310 5194 10362
rect 5246 10310 5258 10362
rect 5310 10310 5322 10362
rect 5374 10310 10396 10362
rect 920 10288 10396 10310
rect 1397 10251 1455 10257
rect 1397 10217 1409 10251
rect 1443 10248 1455 10251
rect 2222 10248 2228 10260
rect 1443 10220 2228 10248
rect 1443 10217 1455 10220
rect 1397 10211 1455 10217
rect 2222 10208 2228 10220
rect 2280 10208 2286 10260
rect 2958 10248 2964 10260
rect 2332 10220 2964 10248
rect 1210 10140 1216 10192
rect 1268 10180 1274 10192
rect 2332 10180 2360 10220
rect 2958 10208 2964 10220
rect 3016 10208 3022 10260
rect 3421 10251 3479 10257
rect 3421 10217 3433 10251
rect 3467 10248 3479 10251
rect 5917 10251 5975 10257
rect 3467 10220 5488 10248
rect 3467 10217 3479 10220
rect 3421 10211 3479 10217
rect 1268 10152 2360 10180
rect 1268 10140 1274 10152
rect 4154 10140 4160 10192
rect 4212 10180 4218 10192
rect 4212 10152 4278 10180
rect 4212 10140 4218 10152
rect 1486 10072 1492 10124
rect 1544 10112 1550 10124
rect 1581 10115 1639 10121
rect 1581 10112 1593 10115
rect 1544 10084 1593 10112
rect 1544 10072 1550 10084
rect 1581 10081 1593 10084
rect 1627 10081 1639 10115
rect 5353 10115 5411 10121
rect 3082 10084 4016 10112
rect 1581 10075 1639 10081
rect 1670 10044 1676 10056
rect 1583 10016 1676 10044
rect 1670 10004 1676 10016
rect 1728 10004 1734 10056
rect 1946 10044 1952 10056
rect 1907 10016 1952 10044
rect 1946 10004 1952 10016
rect 2004 10004 2010 10056
rect 3513 10047 3571 10053
rect 3513 10013 3525 10047
rect 3559 10013 3571 10047
rect 3878 10044 3884 10056
rect 3839 10016 3884 10044
rect 3513 10007 3571 10013
rect 1688 9908 1716 10004
rect 2130 9908 2136 9920
rect 1688 9880 2136 9908
rect 2130 9868 2136 9880
rect 2188 9868 2194 9920
rect 2314 9868 2320 9920
rect 2372 9908 2378 9920
rect 3234 9908 3240 9920
rect 2372 9880 3240 9908
rect 2372 9868 2378 9880
rect 3234 9868 3240 9880
rect 3292 9868 3298 9920
rect 3528 9908 3556 10007
rect 3878 10004 3884 10016
rect 3936 10004 3942 10056
rect 3988 10044 4016 10084
rect 5353 10081 5365 10115
rect 5399 10081 5411 10115
rect 5460 10112 5488 10220
rect 5917 10217 5929 10251
rect 5963 10248 5975 10251
rect 9674 10248 9680 10260
rect 5963 10220 9680 10248
rect 5963 10217 5975 10220
rect 5917 10211 5975 10217
rect 9674 10208 9680 10220
rect 9732 10208 9738 10260
rect 9766 10208 9772 10260
rect 9824 10208 9830 10260
rect 9585 10183 9643 10189
rect 9585 10180 9597 10183
rect 8510 10152 9597 10180
rect 9585 10149 9597 10152
rect 9631 10149 9643 10183
rect 9784 10180 9812 10208
rect 9585 10143 9643 10149
rect 9692 10152 9812 10180
rect 6273 10115 6331 10121
rect 6273 10112 6285 10115
rect 5460 10084 6285 10112
rect 5353 10075 5411 10081
rect 6273 10081 6285 10084
rect 6319 10081 6331 10115
rect 6273 10075 6331 10081
rect 4522 10044 4528 10056
rect 3988 10016 4528 10044
rect 4522 10004 4528 10016
rect 4580 10004 4586 10056
rect 5368 10044 5396 10075
rect 6362 10072 6368 10124
rect 6420 10112 6426 10124
rect 6420 10084 7144 10112
rect 6420 10072 6426 10084
rect 5534 10044 5540 10056
rect 5368 10016 5540 10044
rect 5534 10004 5540 10016
rect 5592 10004 5598 10056
rect 6914 10004 6920 10056
rect 6972 10044 6978 10056
rect 7009 10047 7067 10053
rect 7009 10044 7021 10047
rect 6972 10016 7021 10044
rect 6972 10004 6978 10016
rect 7009 10013 7021 10016
rect 7055 10013 7067 10047
rect 7116 10044 7144 10084
rect 7190 10072 7196 10124
rect 7248 10112 7254 10124
rect 8849 10115 8907 10121
rect 7248 10084 7420 10112
rect 7248 10072 7254 10084
rect 7282 10044 7288 10056
rect 7116 10016 7288 10044
rect 7009 10007 7067 10013
rect 7282 10004 7288 10016
rect 7340 10004 7346 10056
rect 7392 10053 7420 10084
rect 8849 10081 8861 10115
rect 8895 10112 8907 10115
rect 9692 10112 9720 10152
rect 8895 10084 9720 10112
rect 9860 10115 9918 10121
rect 8895 10081 8907 10084
rect 8849 10075 8907 10081
rect 9860 10081 9872 10115
rect 9906 10081 9918 10115
rect 9860 10075 9918 10081
rect 7377 10047 7435 10053
rect 7377 10013 7389 10047
rect 7423 10044 7435 10047
rect 8018 10044 8024 10056
rect 7423 10016 8024 10044
rect 7423 10013 7435 10016
rect 7377 10007 7435 10013
rect 8018 10004 8024 10016
rect 8076 10004 8082 10056
rect 9876 10044 9904 10075
rect 9950 10072 9956 10124
rect 10008 10112 10014 10124
rect 10778 10112 10784 10124
rect 10008 10084 10784 10112
rect 10008 10072 10014 10084
rect 10778 10072 10784 10084
rect 10836 10072 10842 10124
rect 10226 10044 10232 10056
rect 9876 10016 10232 10044
rect 10226 10004 10232 10016
rect 10284 10004 10290 10056
rect 6546 9936 6552 9988
rect 6604 9976 6610 9988
rect 7098 9976 7104 9988
rect 6604 9948 7104 9976
rect 6604 9936 6610 9948
rect 7098 9936 7104 9948
rect 7156 9936 7162 9988
rect 9766 9976 9772 9988
rect 9324 9948 9772 9976
rect 4246 9908 4252 9920
rect 3528 9880 4252 9908
rect 4246 9868 4252 9880
rect 4304 9868 4310 9920
rect 4522 9868 4528 9920
rect 4580 9908 4586 9920
rect 6178 9908 6184 9920
rect 4580 9880 6184 9908
rect 4580 9868 4586 9880
rect 6178 9868 6184 9880
rect 6236 9868 6242 9920
rect 6917 9911 6975 9917
rect 6917 9877 6929 9911
rect 6963 9908 6975 9911
rect 9324 9908 9352 9948
rect 9766 9936 9772 9948
rect 9824 9936 9830 9988
rect 6963 9880 9352 9908
rect 9413 9911 9471 9917
rect 6963 9877 6975 9880
rect 6917 9871 6975 9877
rect 9413 9877 9425 9911
rect 9459 9908 9471 9911
rect 10134 9908 10140 9920
rect 9459 9880 10140 9908
rect 9459 9877 9471 9880
rect 9413 9871 9471 9877
rect 10134 9868 10140 9880
rect 10192 9868 10198 9920
rect 920 9818 10396 9840
rect 920 9766 2566 9818
rect 2618 9766 2630 9818
rect 2682 9766 2694 9818
rect 2746 9766 2758 9818
rect 2810 9766 2822 9818
rect 2874 9766 7566 9818
rect 7618 9766 7630 9818
rect 7682 9766 7694 9818
rect 7746 9766 7758 9818
rect 7810 9766 7822 9818
rect 7874 9766 10396 9818
rect 920 9744 10396 9766
rect 1946 9664 1952 9716
rect 2004 9704 2010 9716
rect 6546 9704 6552 9716
rect 2004 9676 6552 9704
rect 2004 9664 2010 9676
rect 6546 9664 6552 9676
rect 6604 9664 6610 9716
rect 6656 9676 7880 9704
rect 1397 9639 1455 9645
rect 1397 9605 1409 9639
rect 1443 9636 1455 9639
rect 1443 9608 1992 9636
rect 1443 9605 1455 9608
rect 1397 9599 1455 9605
rect 1854 9568 1860 9580
rect 1780 9540 1860 9568
rect 1581 9503 1639 9509
rect 1581 9469 1593 9503
rect 1627 9500 1639 9503
rect 1670 9500 1676 9512
rect 1627 9472 1676 9500
rect 1627 9469 1639 9472
rect 1581 9463 1639 9469
rect 1670 9460 1676 9472
rect 1728 9460 1734 9512
rect 1780 9376 1808 9540
rect 1854 9528 1860 9540
rect 1912 9528 1918 9580
rect 1964 9500 1992 9608
rect 5442 9596 5448 9648
rect 5500 9636 5506 9648
rect 6656 9636 6684 9676
rect 5500 9608 6684 9636
rect 7852 9636 7880 9676
rect 9674 9636 9680 9648
rect 7852 9608 9536 9636
rect 9635 9608 9680 9636
rect 5500 9596 5506 9608
rect 2130 9528 2136 9580
rect 2188 9568 2194 9580
rect 3421 9571 3479 9577
rect 3421 9568 3433 9571
rect 2188 9540 3433 9568
rect 2188 9528 2194 9540
rect 3421 9537 3433 9540
rect 3467 9537 3479 9571
rect 3421 9531 3479 9537
rect 3694 9528 3700 9580
rect 3752 9568 3758 9580
rect 4249 9571 4307 9577
rect 4249 9568 4261 9571
rect 3752 9540 4261 9568
rect 3752 9528 3758 9540
rect 4249 9537 4261 9540
rect 4295 9537 4307 9571
rect 4249 9531 4307 9537
rect 6362 9528 6368 9580
rect 6420 9568 6426 9580
rect 6825 9571 6883 9577
rect 6825 9568 6837 9571
rect 6420 9540 6837 9568
rect 6420 9528 6426 9540
rect 6825 9537 6837 9540
rect 6871 9537 6883 9571
rect 6825 9531 6883 9537
rect 8478 9528 8484 9580
rect 8536 9568 8542 9580
rect 8573 9571 8631 9577
rect 8573 9568 8585 9571
rect 8536 9540 8585 9568
rect 8536 9528 8542 9540
rect 8573 9537 8585 9540
rect 8619 9537 8631 9571
rect 8573 9531 8631 9537
rect 9217 9571 9275 9577
rect 9217 9537 9229 9571
rect 9263 9568 9275 9571
rect 9306 9568 9312 9580
rect 9263 9540 9312 9568
rect 9263 9537 9275 9540
rect 9217 9531 9275 9537
rect 9306 9528 9312 9540
rect 9364 9528 9370 9580
rect 9508 9568 9536 9608
rect 9674 9596 9680 9608
rect 9732 9596 9738 9648
rect 16850 9636 16856 9648
rect 12406 9608 16856 9636
rect 12406 9568 12434 9608
rect 16850 9596 16856 9608
rect 16908 9596 16914 9648
rect 9508 9540 12434 9568
rect 1872 9472 1992 9500
rect 1578 9324 1584 9376
rect 1636 9364 1642 9376
rect 1673 9367 1731 9373
rect 1673 9364 1685 9367
rect 1636 9336 1685 9364
rect 1636 9324 1642 9336
rect 1673 9333 1685 9336
rect 1719 9333 1731 9367
rect 1673 9327 1731 9333
rect 1762 9324 1768 9376
rect 1820 9324 1826 9376
rect 1872 9364 1900 9472
rect 3510 9460 3516 9512
rect 3568 9500 3574 9512
rect 3605 9503 3663 9509
rect 3605 9500 3617 9503
rect 3568 9472 3617 9500
rect 3568 9460 3574 9472
rect 3605 9469 3617 9472
rect 3651 9469 3663 9503
rect 3878 9500 3884 9512
rect 3839 9472 3884 9500
rect 3605 9463 3663 9469
rect 3878 9460 3884 9472
rect 3936 9460 3942 9512
rect 5718 9500 5724 9512
rect 5679 9472 5724 9500
rect 5718 9460 5724 9472
rect 5776 9460 5782 9512
rect 6546 9500 6552 9512
rect 6507 9472 6552 9500
rect 6546 9460 6552 9472
rect 6604 9460 6610 9512
rect 8846 9460 8852 9512
rect 8904 9500 8910 9512
rect 8971 9503 9029 9509
rect 8971 9500 8983 9503
rect 8904 9472 8983 9500
rect 8904 9460 8910 9472
rect 8971 9469 8983 9472
rect 9017 9469 9029 9503
rect 8971 9463 9029 9469
rect 9122 9460 9128 9512
rect 9180 9500 9186 9512
rect 9401 9503 9459 9509
rect 9401 9500 9413 9503
rect 9180 9472 9413 9500
rect 9180 9460 9186 9472
rect 9401 9469 9413 9472
rect 9447 9469 9459 9503
rect 9858 9500 9864 9512
rect 9819 9472 9864 9500
rect 9401 9463 9459 9469
rect 9858 9460 9864 9472
rect 9916 9460 9922 9512
rect 2866 9432 2872 9444
rect 2714 9404 2872 9432
rect 2866 9392 2872 9404
rect 2924 9392 2930 9444
rect 3142 9432 3148 9444
rect 3103 9404 3148 9432
rect 3142 9392 3148 9404
rect 3200 9432 3206 9444
rect 3786 9432 3792 9444
rect 3200 9404 3792 9432
rect 3200 9392 3206 9404
rect 3786 9392 3792 9404
rect 3844 9392 3850 9444
rect 4706 9392 4712 9444
rect 4764 9392 4770 9444
rect 5736 9404 7314 9432
rect 5736 9376 5764 9404
rect 8202 9392 8208 9444
rect 8260 9432 8266 9444
rect 9585 9435 9643 9441
rect 9585 9432 9597 9435
rect 8260 9404 9597 9432
rect 8260 9392 8266 9404
rect 9585 9401 9597 9404
rect 9631 9401 9643 9435
rect 19794 9432 19800 9444
rect 9585 9395 9643 9401
rect 16546 9404 19800 9432
rect 2314 9364 2320 9376
rect 1872 9336 2320 9364
rect 2314 9324 2320 9336
rect 2372 9324 2378 9376
rect 3697 9367 3755 9373
rect 3697 9333 3709 9367
rect 3743 9364 3755 9367
rect 5442 9364 5448 9376
rect 3743 9336 5448 9364
rect 3743 9333 3755 9336
rect 3697 9327 3755 9333
rect 5442 9324 5448 9336
rect 5500 9324 5506 9376
rect 5718 9324 5724 9376
rect 5776 9324 5782 9376
rect 6285 9367 6343 9373
rect 6285 9333 6297 9367
rect 6331 9364 6343 9367
rect 8294 9364 8300 9376
rect 6331 9336 8300 9364
rect 6331 9333 6343 9336
rect 6285 9327 6343 9333
rect 8294 9324 8300 9336
rect 8352 9324 8358 9376
rect 8754 9364 8760 9376
rect 8715 9336 8760 9364
rect 8754 9324 8760 9336
rect 8812 9324 8818 9376
rect 8846 9324 8852 9376
rect 8904 9364 8910 9376
rect 9306 9364 9312 9376
rect 8904 9336 9312 9364
rect 8904 9324 8910 9336
rect 9306 9324 9312 9336
rect 9364 9324 9370 9376
rect 10045 9367 10103 9373
rect 10045 9333 10057 9367
rect 10091 9364 10103 9367
rect 10594 9364 10600 9376
rect 10091 9336 10600 9364
rect 10091 9333 10103 9336
rect 10045 9327 10103 9333
rect 10594 9324 10600 9336
rect 10652 9324 10658 9376
rect 920 9274 10396 9296
rect 920 9222 5066 9274
rect 5118 9222 5130 9274
rect 5182 9222 5194 9274
rect 5246 9222 5258 9274
rect 5310 9222 5322 9274
rect 5374 9222 10396 9274
rect 920 9200 10396 9222
rect 1305 9163 1363 9169
rect 1305 9129 1317 9163
rect 1351 9160 1363 9163
rect 6546 9160 6552 9172
rect 1351 9132 6552 9160
rect 1351 9129 1363 9132
rect 1305 9123 1363 9129
rect 6546 9120 6552 9132
rect 6604 9120 6610 9172
rect 8938 9120 8944 9172
rect 8996 9160 9002 9172
rect 16546 9160 16574 9404
rect 19794 9392 19800 9404
rect 19852 9392 19858 9444
rect 8996 9132 16574 9160
rect 8996 9120 9002 9132
rect 2038 9052 2044 9104
rect 2096 9092 2102 9104
rect 2133 9095 2191 9101
rect 2133 9092 2145 9095
rect 2096 9064 2145 9092
rect 2096 9052 2102 9064
rect 2133 9061 2145 9064
rect 2179 9092 2191 9095
rect 3694 9092 3700 9104
rect 2179 9064 3700 9092
rect 2179 9061 2191 9064
rect 2133 9055 2191 9061
rect 3694 9052 3700 9064
rect 3752 9052 3758 9104
rect 3878 9052 3884 9104
rect 3936 9092 3942 9104
rect 5534 9092 5540 9104
rect 3936 9064 5540 9092
rect 3936 9052 3942 9064
rect 5534 9052 5540 9064
rect 5592 9052 5598 9104
rect 6178 9052 6184 9104
rect 6236 9092 6242 9104
rect 8478 9092 8484 9104
rect 6236 9064 8484 9092
rect 6236 9052 6242 9064
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 2958 9024 2964 9036
rect 1443 8996 2964 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 2958 8984 2964 8996
rect 3016 8984 3022 9036
rect 3326 8984 3332 9036
rect 3384 9024 3390 9036
rect 3786 9024 3792 9036
rect 3384 8996 3792 9024
rect 3384 8984 3390 8996
rect 3786 8984 3792 8996
rect 3844 8984 3850 9036
rect 3970 9024 3976 9036
rect 3931 8996 3976 9024
rect 3970 8984 3976 8996
rect 4028 8984 4034 9036
rect 4065 9027 4123 9033
rect 4065 8993 4077 9027
rect 4111 8993 4123 9027
rect 4065 8987 4123 8993
rect 5997 9027 6055 9033
rect 5997 8993 6009 9027
rect 6043 9024 6055 9027
rect 6546 9024 6552 9036
rect 6043 8996 6552 9024
rect 6043 8993 6055 8996
rect 5997 8987 6055 8993
rect 1578 8956 1584 8968
rect 1539 8928 1584 8956
rect 1578 8916 1584 8928
rect 1636 8916 1642 8968
rect 1762 8916 1768 8968
rect 1820 8956 1826 8968
rect 4080 8956 4108 8987
rect 6546 8984 6552 8996
rect 6604 8984 6610 9036
rect 6730 9024 6736 9036
rect 6691 8996 6736 9024
rect 6730 8984 6736 8996
rect 6788 8984 6794 9036
rect 6932 9033 6960 9064
rect 8478 9052 8484 9064
rect 8536 9052 8542 9104
rect 8754 9052 8760 9104
rect 8812 9052 8818 9104
rect 6917 9027 6975 9033
rect 6917 8993 6929 9027
rect 6963 8993 6975 9027
rect 6917 8987 6975 8993
rect 7010 9027 7068 9033
rect 7010 8993 7022 9027
rect 7056 8993 7068 9027
rect 8202 9024 8208 9036
rect 8163 8996 8208 9024
rect 7010 8987 7068 8993
rect 1820 8928 4108 8956
rect 1820 8916 1826 8928
rect 4246 8916 4252 8968
rect 4304 8956 4310 8968
rect 4706 8956 4712 8968
rect 4304 8928 4712 8956
rect 4304 8916 4310 8928
rect 4706 8916 4712 8928
rect 4764 8916 4770 8968
rect 6178 8916 6184 8968
rect 6236 8956 6242 8968
rect 6236 8928 6592 8956
rect 6236 8916 6242 8928
rect 3786 8848 3792 8900
rect 3844 8888 3850 8900
rect 6564 8888 6592 8928
rect 6638 8916 6644 8968
rect 6696 8956 6702 8968
rect 7024 8956 7052 8987
rect 8202 8984 8208 8996
rect 8260 8984 8266 9036
rect 9677 9027 9735 9033
rect 9677 8993 9689 9027
rect 9723 9024 9735 9027
rect 9766 9024 9772 9036
rect 9723 8996 9772 9024
rect 9723 8993 9735 8996
rect 9677 8987 9735 8993
rect 9766 8984 9772 8996
rect 9824 9024 9830 9036
rect 10318 9024 10324 9036
rect 9824 8996 10324 9024
rect 9824 8984 9830 8996
rect 10318 8984 10324 8996
rect 10376 8984 10382 9036
rect 7282 8956 7288 8968
rect 6696 8928 7052 8956
rect 7243 8928 7288 8956
rect 6696 8916 6702 8928
rect 7282 8916 7288 8928
rect 7340 8916 7346 8968
rect 10042 8956 10048 8968
rect 10003 8928 10048 8956
rect 10042 8916 10048 8928
rect 10100 8916 10106 8968
rect 7469 8891 7527 8897
rect 7469 8888 7481 8891
rect 3844 8860 6500 8888
rect 6564 8860 7481 8888
rect 3844 8848 3850 8860
rect 2685 8823 2743 8829
rect 2685 8789 2697 8823
rect 2731 8820 2743 8823
rect 3326 8820 3332 8832
rect 2731 8792 3332 8820
rect 2731 8789 2743 8792
rect 2685 8783 2743 8789
rect 3326 8780 3332 8792
rect 3384 8780 3390 8832
rect 3878 8780 3884 8832
rect 3936 8820 3942 8832
rect 6181 8823 6239 8829
rect 6181 8820 6193 8823
rect 3936 8792 6193 8820
rect 3936 8780 3942 8792
rect 6181 8789 6193 8792
rect 6227 8789 6239 8823
rect 6472 8820 6500 8860
rect 7469 8857 7481 8860
rect 7515 8888 7527 8891
rect 7515 8860 8800 8888
rect 7515 8857 7527 8860
rect 7469 8851 7527 8857
rect 6730 8820 6736 8832
rect 6472 8792 6736 8820
rect 6181 8783 6239 8789
rect 6730 8780 6736 8792
rect 6788 8780 6794 8832
rect 7006 8780 7012 8832
rect 7064 8820 7070 8832
rect 7640 8823 7698 8829
rect 7640 8820 7652 8823
rect 7064 8792 7652 8820
rect 7064 8780 7070 8792
rect 7640 8789 7652 8792
rect 7686 8789 7698 8823
rect 8772 8820 8800 8860
rect 16666 8820 16672 8832
rect 8772 8792 16672 8820
rect 7640 8783 7698 8789
rect 16666 8780 16672 8792
rect 16724 8780 16730 8832
rect 920 8730 10396 8752
rect 920 8678 2566 8730
rect 2618 8678 2630 8730
rect 2682 8678 2694 8730
rect 2746 8678 2758 8730
rect 2810 8678 2822 8730
rect 2874 8678 7566 8730
rect 7618 8678 7630 8730
rect 7682 8678 7694 8730
rect 7746 8678 7758 8730
rect 7810 8678 7822 8730
rect 7874 8678 10396 8730
rect 920 8656 10396 8678
rect 1489 8619 1547 8625
rect 1489 8585 1501 8619
rect 1535 8616 1547 8619
rect 1762 8616 1768 8628
rect 1535 8588 1768 8616
rect 1535 8585 1547 8588
rect 1489 8579 1547 8585
rect 1762 8576 1768 8588
rect 1820 8576 1826 8628
rect 3142 8576 3148 8628
rect 3200 8616 3206 8628
rect 4249 8619 4307 8625
rect 4249 8616 4261 8619
rect 3200 8588 4261 8616
rect 3200 8576 3206 8588
rect 4249 8585 4261 8588
rect 4295 8585 4307 8619
rect 4249 8579 4307 8585
rect 5350 8576 5356 8628
rect 5408 8616 5414 8628
rect 5408 8588 9260 8616
rect 5408 8576 5414 8588
rect 3234 8508 3240 8560
rect 3292 8548 3298 8560
rect 3292 8520 4108 8548
rect 3292 8508 3298 8520
rect 3421 8483 3479 8489
rect 3421 8449 3433 8483
rect 3467 8480 3479 8483
rect 3970 8480 3976 8492
rect 3467 8452 3976 8480
rect 3467 8449 3479 8452
rect 3421 8443 3479 8449
rect 3970 8440 3976 8452
rect 4028 8440 4034 8492
rect 4080 8480 4108 8520
rect 8478 8508 8484 8560
rect 8536 8548 8542 8560
rect 9122 8548 9128 8560
rect 8536 8520 9128 8548
rect 8536 8508 8542 8520
rect 4080 8452 4568 8480
rect 1118 8372 1124 8424
rect 1176 8412 1182 8424
rect 1673 8415 1731 8421
rect 1673 8412 1685 8415
rect 1176 8384 1685 8412
rect 1176 8372 1182 8384
rect 1673 8381 1685 8384
rect 1719 8381 1731 8415
rect 1673 8375 1731 8381
rect 3142 8372 3148 8424
rect 3200 8412 3206 8424
rect 4540 8421 4568 8452
rect 5994 8440 6000 8492
rect 6052 8480 6058 8492
rect 8662 8480 8668 8492
rect 6052 8452 8668 8480
rect 6052 8440 6058 8452
rect 8662 8440 8668 8452
rect 8720 8440 8726 8492
rect 3605 8415 3663 8421
rect 3605 8412 3617 8415
rect 3200 8384 3617 8412
rect 3200 8372 3206 8384
rect 3605 8381 3617 8384
rect 3651 8381 3663 8415
rect 4341 8415 4399 8421
rect 4341 8412 4353 8415
rect 3605 8375 3663 8381
rect 3712 8384 4353 8412
rect 1397 8347 1455 8353
rect 1397 8313 1409 8347
rect 1443 8313 1455 8347
rect 1397 8307 1455 8313
rect 1412 8276 1440 8307
rect 3234 8304 3240 8356
rect 3292 8344 3298 8356
rect 3712 8344 3740 8384
rect 4341 8381 4353 8384
rect 4387 8381 4399 8415
rect 4341 8375 4399 8381
rect 4525 8415 4583 8421
rect 4525 8381 4537 8415
rect 4571 8381 4583 8415
rect 4801 8415 4859 8421
rect 4801 8412 4813 8415
rect 4525 8375 4583 8381
rect 4632 8384 4813 8412
rect 3292 8316 3740 8344
rect 3292 8304 3298 8316
rect 4246 8304 4252 8356
rect 4304 8344 4310 8356
rect 4632 8344 4660 8384
rect 4801 8381 4813 8384
rect 4847 8381 4859 8415
rect 4801 8375 4859 8381
rect 6178 8372 6184 8424
rect 6236 8412 6242 8424
rect 6549 8415 6607 8421
rect 6549 8412 6561 8415
rect 6236 8384 6561 8412
rect 6236 8372 6242 8384
rect 6549 8381 6561 8384
rect 6595 8381 6607 8415
rect 8570 8412 8576 8424
rect 8531 8384 8576 8412
rect 6549 8375 6607 8381
rect 8570 8372 8576 8384
rect 8628 8372 8634 8424
rect 8956 8421 8984 8520
rect 9122 8508 9128 8520
rect 9180 8508 9186 8560
rect 9232 8480 9260 8588
rect 9490 8508 9496 8560
rect 9548 8548 9554 8560
rect 9674 8548 9680 8560
rect 9548 8520 9680 8548
rect 9548 8508 9554 8520
rect 9674 8508 9680 8520
rect 9732 8508 9738 8560
rect 9232 8452 10180 8480
rect 8757 8415 8815 8421
rect 8757 8381 8769 8415
rect 8803 8381 8815 8415
rect 8757 8375 8815 8381
rect 8941 8415 8999 8421
rect 8941 8381 8953 8415
rect 8987 8381 8999 8415
rect 9214 8412 9220 8424
rect 9175 8384 9220 8412
rect 8941 8375 8999 8381
rect 4304 8316 4660 8344
rect 4709 8347 4767 8353
rect 4304 8304 4310 8316
rect 4709 8313 4721 8347
rect 4755 8344 4767 8347
rect 4890 8344 4896 8356
rect 4755 8316 4896 8344
rect 4755 8313 4767 8316
rect 4709 8307 4767 8313
rect 4890 8304 4896 8316
rect 4948 8304 4954 8356
rect 6638 8304 6644 8356
rect 6696 8344 6702 8356
rect 8772 8344 8800 8375
rect 9214 8372 9220 8384
rect 9272 8372 9278 8424
rect 9306 8372 9312 8424
rect 9364 8412 9370 8424
rect 9364 8384 9409 8412
rect 9364 8372 9370 8384
rect 9674 8372 9680 8424
rect 9732 8412 9738 8424
rect 9861 8415 9919 8421
rect 9732 8384 9777 8412
rect 9732 8372 9738 8384
rect 9861 8381 9873 8415
rect 9907 8412 9919 8415
rect 9950 8412 9956 8424
rect 9907 8384 9956 8412
rect 9907 8381 9919 8384
rect 9861 8375 9919 8381
rect 9950 8372 9956 8384
rect 10008 8372 10014 8424
rect 9122 8344 9128 8356
rect 6696 8316 8800 8344
rect 9083 8316 9128 8344
rect 6696 8304 6702 8316
rect 9122 8304 9128 8316
rect 9180 8304 9186 8356
rect 9582 8344 9588 8356
rect 9543 8316 9588 8344
rect 9582 8304 9588 8316
rect 9640 8304 9646 8356
rect 9766 8304 9772 8356
rect 9824 8344 9830 8356
rect 10045 8347 10103 8353
rect 10045 8344 10057 8347
rect 9824 8316 10057 8344
rect 9824 8304 9830 8316
rect 10045 8313 10057 8316
rect 10091 8313 10103 8347
rect 10152 8344 10180 8452
rect 11238 8372 11244 8424
rect 11296 8412 11302 8424
rect 19610 8412 19616 8424
rect 11296 8384 19616 8412
rect 11296 8372 11302 8384
rect 19610 8372 19616 8384
rect 19668 8372 19674 8424
rect 16758 8344 16764 8356
rect 10152 8316 16764 8344
rect 10045 8307 10103 8313
rect 16758 8304 16764 8316
rect 16816 8304 16822 8356
rect 5718 8276 5724 8288
rect 1412 8248 5724 8276
rect 5718 8236 5724 8248
rect 5776 8236 5782 8288
rect 5902 8236 5908 8288
rect 5960 8276 5966 8288
rect 6546 8276 6552 8288
rect 5960 8248 6552 8276
rect 5960 8236 5966 8248
rect 6546 8236 6552 8248
rect 6604 8236 6610 8288
rect 7653 8279 7711 8285
rect 7653 8245 7665 8279
rect 7699 8276 7711 8279
rect 12342 8276 12348 8288
rect 7699 8248 12348 8276
rect 7699 8245 7711 8248
rect 7653 8239 7711 8245
rect 12342 8236 12348 8248
rect 12400 8236 12406 8288
rect 920 8186 10396 8208
rect 920 8134 5066 8186
rect 5118 8134 5130 8186
rect 5182 8134 5194 8186
rect 5246 8134 5258 8186
rect 5310 8134 5322 8186
rect 5374 8134 10396 8186
rect 920 8112 10396 8134
rect 1489 8075 1547 8081
rect 1489 8041 1501 8075
rect 1535 8072 1547 8075
rect 3418 8072 3424 8084
rect 1535 8044 3424 8072
rect 1535 8041 1547 8044
rect 1489 8035 1547 8041
rect 3418 8032 3424 8044
rect 3476 8032 3482 8084
rect 6822 8072 6828 8084
rect 6783 8044 6828 8072
rect 6822 8032 6828 8044
rect 6880 8032 6886 8084
rect 7282 8032 7288 8084
rect 7340 8072 7346 8084
rect 7340 8044 7604 8072
rect 7340 8032 7346 8044
rect 1397 8007 1455 8013
rect 1397 7973 1409 8007
rect 1443 8004 1455 8007
rect 1762 8004 1768 8016
rect 1443 7976 1768 8004
rect 1443 7973 1455 7976
rect 1397 7967 1455 7973
rect 1762 7964 1768 7976
rect 1820 8004 1826 8016
rect 2406 8004 2412 8016
rect 1820 7976 2412 8004
rect 1820 7964 1826 7976
rect 2406 7964 2412 7976
rect 2464 7964 2470 8016
rect 3329 8007 3387 8013
rect 3329 7973 3341 8007
rect 3375 8004 3387 8007
rect 3510 8004 3516 8016
rect 3375 7976 3516 8004
rect 3375 7973 3387 7976
rect 3329 7967 3387 7973
rect 3510 7964 3516 7976
rect 3568 7964 3574 8016
rect 4246 7964 4252 8016
rect 4304 7964 4310 8016
rect 7576 8004 7604 8044
rect 7926 8032 7932 8084
rect 7984 8072 7990 8084
rect 16942 8072 16948 8084
rect 7984 8044 16948 8072
rect 7984 8032 7990 8044
rect 16942 8032 16948 8044
rect 17000 8032 17006 8084
rect 7576 7976 7682 8004
rect 9232 7976 16574 8004
rect 1673 7939 1731 7945
rect 1673 7905 1685 7939
rect 1719 7936 1731 7939
rect 3418 7936 3424 7948
rect 1719 7908 3424 7936
rect 1719 7905 1731 7908
rect 1673 7899 1731 7905
rect 3418 7896 3424 7908
rect 3476 7936 3482 7948
rect 3694 7936 3700 7948
rect 3476 7908 3700 7936
rect 3476 7896 3482 7908
rect 3694 7896 3700 7908
rect 3752 7896 3758 7948
rect 3878 7936 3884 7948
rect 3839 7908 3884 7936
rect 3878 7896 3884 7908
rect 3936 7896 3942 7948
rect 4890 7896 4896 7948
rect 4948 7936 4954 7948
rect 5353 7939 5411 7945
rect 5353 7936 5365 7939
rect 4948 7908 5365 7936
rect 4948 7896 4954 7908
rect 5353 7905 5365 7908
rect 5399 7905 5411 7939
rect 5353 7899 5411 7905
rect 5442 7896 5448 7948
rect 5500 7936 5506 7948
rect 6917 7939 6975 7945
rect 6917 7936 6929 7939
rect 5500 7908 6929 7936
rect 5500 7896 5506 7908
rect 6917 7905 6929 7908
rect 6963 7905 6975 7939
rect 6917 7899 6975 7905
rect 7098 7896 7104 7948
rect 7156 7936 7162 7948
rect 7285 7939 7343 7945
rect 7285 7936 7297 7939
rect 7156 7908 7297 7936
rect 7156 7896 7162 7908
rect 7285 7905 7297 7908
rect 7331 7905 7343 7939
rect 7285 7899 7343 7905
rect 8757 7939 8815 7945
rect 8757 7905 8769 7939
rect 8803 7936 8815 7939
rect 9122 7936 9128 7948
rect 8803 7908 9128 7936
rect 8803 7905 8815 7908
rect 8757 7899 8815 7905
rect 9122 7896 9128 7908
rect 9180 7896 9186 7948
rect 3510 7868 3516 7880
rect 3471 7840 3516 7868
rect 3510 7828 3516 7840
rect 3568 7828 3574 7880
rect 6273 7871 6331 7877
rect 6273 7837 6285 7871
rect 6319 7868 6331 7871
rect 6362 7868 6368 7880
rect 6319 7840 6368 7868
rect 6319 7837 6331 7840
rect 6273 7831 6331 7837
rect 6362 7828 6368 7840
rect 6420 7828 6426 7880
rect 9232 7800 9260 7976
rect 12342 7896 12348 7948
rect 12400 7936 12406 7948
rect 14090 7936 14096 7948
rect 12400 7908 14096 7936
rect 12400 7904 12434 7908
rect 12400 7896 12406 7904
rect 14090 7896 14096 7908
rect 14148 7896 14154 7948
rect 9490 7868 9496 7880
rect 9451 7840 9496 7868
rect 9490 7828 9496 7840
rect 9548 7828 9554 7880
rect 8220 7772 9260 7800
rect 1486 7692 1492 7744
rect 1544 7732 1550 7744
rect 3234 7732 3240 7744
rect 1544 7704 3240 7732
rect 1544 7692 1550 7704
rect 3234 7692 3240 7704
rect 3292 7692 3298 7744
rect 5902 7692 5908 7744
rect 5960 7741 5966 7744
rect 5960 7732 5971 7741
rect 5960 7704 6005 7732
rect 5960 7695 5971 7704
rect 5960 7692 5966 7695
rect 6270 7692 6276 7744
rect 6328 7732 6334 7744
rect 6822 7732 6828 7744
rect 6328 7704 6828 7732
rect 6328 7692 6334 7704
rect 6822 7692 6828 7704
rect 6880 7692 6886 7744
rect 7282 7692 7288 7744
rect 7340 7732 7346 7744
rect 8220 7732 8248 7772
rect 9582 7760 9588 7812
rect 9640 7800 9646 7812
rect 9769 7803 9827 7809
rect 9769 7800 9781 7803
rect 9640 7772 9781 7800
rect 9640 7760 9646 7772
rect 9769 7769 9781 7772
rect 9815 7769 9827 7803
rect 9769 7763 9827 7769
rect 7340 7704 8248 7732
rect 7340 7692 7346 7704
rect 8754 7692 8760 7744
rect 8812 7732 8818 7744
rect 9317 7735 9375 7741
rect 9317 7732 9329 7735
rect 8812 7704 9329 7732
rect 8812 7692 8818 7704
rect 9317 7701 9329 7704
rect 9363 7701 9375 7735
rect 9950 7732 9956 7744
rect 9911 7704 9956 7732
rect 9317 7695 9375 7701
rect 9950 7692 9956 7704
rect 10008 7692 10014 7744
rect 920 7642 10396 7664
rect 920 7590 2566 7642
rect 2618 7590 2630 7642
rect 2682 7590 2694 7642
rect 2746 7590 2758 7642
rect 2810 7590 2822 7642
rect 2874 7590 7566 7642
rect 7618 7590 7630 7642
rect 7682 7590 7694 7642
rect 7746 7590 7758 7642
rect 7810 7590 7822 7642
rect 7874 7590 10396 7642
rect 920 7568 10396 7590
rect 1397 7531 1455 7537
rect 1397 7497 1409 7531
rect 1443 7528 1455 7531
rect 4246 7528 4252 7540
rect 1443 7500 4252 7528
rect 1443 7497 1455 7500
rect 1397 7491 1455 7497
rect 4246 7488 4252 7500
rect 4304 7488 4310 7540
rect 8941 7531 8999 7537
rect 8941 7497 8953 7531
rect 8987 7528 8999 7531
rect 9122 7528 9128 7540
rect 8987 7500 9128 7528
rect 8987 7497 8999 7500
rect 8941 7491 8999 7497
rect 9122 7488 9128 7500
rect 9180 7488 9186 7540
rect 4062 7420 4068 7472
rect 4120 7460 4126 7472
rect 5994 7460 6000 7472
rect 4120 7432 6000 7460
rect 4120 7420 4126 7432
rect 5994 7420 6000 7432
rect 6052 7420 6058 7472
rect 8570 7420 8576 7472
rect 8628 7460 8634 7472
rect 9217 7463 9275 7469
rect 9217 7460 9229 7463
rect 8628 7432 9229 7460
rect 8628 7420 8634 7432
rect 9217 7429 9229 7432
rect 9263 7429 9275 7463
rect 9217 7423 9275 7429
rect 9582 7420 9588 7472
rect 9640 7460 9646 7472
rect 10226 7460 10232 7472
rect 9640 7432 10232 7460
rect 9640 7420 9646 7432
rect 10226 7420 10232 7432
rect 10284 7420 10290 7472
rect 13538 7460 13544 7472
rect 12406 7432 13544 7460
rect 3234 7352 3240 7404
rect 3292 7392 3298 7404
rect 3605 7395 3663 7401
rect 3605 7392 3617 7395
rect 3292 7364 3617 7392
rect 3292 7352 3298 7364
rect 3605 7361 3617 7364
rect 3651 7361 3663 7395
rect 3605 7355 3663 7361
rect 4246 7352 4252 7404
rect 4304 7392 4310 7404
rect 4522 7392 4528 7404
rect 4304 7364 4528 7392
rect 4304 7352 4310 7364
rect 4522 7352 4528 7364
rect 4580 7352 4586 7404
rect 7929 7395 7987 7401
rect 7929 7361 7941 7395
rect 7975 7392 7987 7395
rect 12406 7392 12434 7432
rect 13538 7420 13544 7432
rect 13596 7420 13602 7472
rect 7975 7364 12434 7392
rect 16546 7392 16574 7976
rect 20162 7392 20168 7404
rect 16546 7364 20168 7392
rect 7975 7361 7987 7364
rect 7929 7355 7987 7361
rect 20162 7352 20168 7364
rect 20220 7352 20226 7404
rect 1486 7324 1492 7336
rect 1447 7296 1492 7324
rect 1486 7284 1492 7296
rect 1544 7284 1550 7336
rect 1578 7284 1584 7336
rect 1636 7324 1642 7336
rect 1636 7296 1681 7324
rect 1636 7284 1642 7296
rect 3326 7284 3332 7336
rect 3384 7324 3390 7336
rect 3421 7327 3479 7333
rect 3421 7324 3433 7327
rect 3384 7296 3433 7324
rect 3384 7284 3390 7296
rect 3421 7293 3433 7296
rect 3467 7293 3479 7327
rect 3421 7287 3479 7293
rect 3694 7284 3700 7336
rect 3752 7324 3758 7336
rect 4341 7327 4399 7333
rect 4341 7324 4353 7327
rect 3752 7296 4353 7324
rect 3752 7284 3758 7296
rect 4341 7293 4353 7296
rect 4387 7324 4399 7327
rect 5442 7324 5448 7336
rect 4387 7296 5448 7324
rect 4387 7293 4399 7296
rect 4341 7287 4399 7293
rect 5442 7284 5448 7296
rect 5500 7284 5506 7336
rect 5626 7284 5632 7336
rect 5684 7324 5690 7336
rect 6270 7324 6276 7336
rect 5684 7296 6276 7324
rect 5684 7284 5690 7296
rect 6270 7284 6276 7296
rect 6328 7284 6334 7336
rect 6549 7327 6607 7333
rect 6549 7293 6561 7327
rect 6595 7324 6607 7327
rect 7006 7324 7012 7336
rect 6595 7296 7012 7324
rect 6595 7293 6607 7296
rect 6549 7287 6607 7293
rect 7006 7284 7012 7296
rect 7064 7284 7070 7336
rect 8570 7324 8576 7336
rect 8531 7296 8576 7324
rect 8570 7284 8576 7296
rect 8628 7284 8634 7336
rect 8662 7284 8668 7336
rect 8720 7326 8726 7336
rect 8849 7327 8907 7333
rect 8720 7318 8800 7326
rect 8849 7318 8861 7327
rect 8720 7298 8861 7318
rect 8720 7284 8726 7298
rect 8772 7293 8861 7298
rect 8895 7324 8907 7327
rect 8956 7324 9076 7334
rect 8895 7318 9168 7324
rect 8895 7306 9260 7318
rect 8895 7296 8984 7306
rect 9048 7296 9260 7306
rect 8895 7293 8907 7296
rect 8772 7290 8907 7293
rect 9140 7290 9260 7296
rect 8849 7287 8907 7290
rect 4433 7259 4491 7265
rect 4433 7225 4445 7259
rect 4479 7256 4491 7259
rect 7098 7256 7104 7268
rect 4479 7228 7104 7256
rect 4479 7225 4491 7228
rect 4433 7219 4491 7225
rect 7098 7216 7104 7228
rect 7156 7216 7162 7268
rect 9232 7256 9260 7290
rect 9490 7284 9496 7336
rect 9548 7324 9554 7336
rect 9769 7327 9827 7333
rect 9548 7296 9593 7324
rect 9548 7284 9554 7296
rect 9769 7293 9781 7327
rect 9815 7324 9827 7327
rect 10226 7324 10232 7336
rect 9815 7296 10232 7324
rect 9815 7293 9827 7296
rect 9769 7287 9827 7293
rect 10226 7284 10232 7296
rect 10284 7284 10290 7336
rect 9677 7259 9735 7265
rect 9232 7228 9536 7256
rect 2130 7188 2136 7200
rect 2091 7160 2136 7188
rect 2130 7148 2136 7160
rect 2188 7148 2194 7200
rect 4154 7148 4160 7200
rect 4212 7188 4218 7200
rect 4249 7191 4307 7197
rect 4249 7188 4261 7191
rect 4212 7160 4261 7188
rect 4212 7148 4218 7160
rect 4249 7157 4261 7160
rect 4295 7188 4307 7191
rect 4614 7188 4620 7200
rect 4295 7160 4620 7188
rect 4295 7157 4307 7160
rect 4249 7151 4307 7157
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 5626 7188 5632 7200
rect 5587 7160 5632 7188
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 9508 7188 9536 7228
rect 9677 7225 9689 7259
rect 9723 7256 9735 7259
rect 10594 7256 10600 7268
rect 9723 7228 10600 7256
rect 9723 7225 9735 7228
rect 9677 7219 9735 7225
rect 10594 7216 10600 7228
rect 10652 7216 10658 7268
rect 9953 7191 10011 7197
rect 9953 7188 9965 7191
rect 9508 7160 9965 7188
rect 9953 7157 9965 7160
rect 9999 7157 10011 7191
rect 9953 7151 10011 7157
rect 920 7098 10396 7120
rect 920 7046 5066 7098
rect 5118 7046 5130 7098
rect 5182 7046 5194 7098
rect 5246 7046 5258 7098
rect 5310 7046 5322 7098
rect 5374 7046 10396 7098
rect 11054 7080 11060 7132
rect 11112 7120 11118 7132
rect 19886 7120 19892 7132
rect 11112 7092 19892 7120
rect 11112 7080 11118 7092
rect 19886 7080 19892 7092
rect 19944 7080 19950 7132
rect 920 7024 10396 7046
rect 13630 7012 13636 7064
rect 13688 7052 13694 7064
rect 20254 7052 20260 7064
rect 13688 7024 20260 7052
rect 13688 7012 13694 7024
rect 20254 7012 20260 7024
rect 20312 7012 20318 7064
rect 1578 6944 1584 6996
rect 1636 6984 1642 6996
rect 3694 6984 3700 6996
rect 1636 6956 3700 6984
rect 1636 6944 1642 6956
rect 3694 6944 3700 6956
rect 3752 6944 3758 6996
rect 6270 6944 6276 6996
rect 6328 6984 6334 6996
rect 6917 6987 6975 6993
rect 6917 6984 6929 6987
rect 6328 6956 6929 6984
rect 6328 6944 6334 6956
rect 6917 6953 6929 6956
rect 6963 6953 6975 6987
rect 6917 6947 6975 6953
rect 9125 6987 9183 6993
rect 9125 6953 9137 6987
rect 9171 6984 9183 6987
rect 9306 6984 9312 6996
rect 9171 6956 9312 6984
rect 9171 6953 9183 6956
rect 9125 6947 9183 6953
rect 9306 6944 9312 6956
rect 9364 6944 9370 6996
rect 1397 6919 1455 6925
rect 1397 6885 1409 6919
rect 1443 6916 1455 6919
rect 2406 6916 2412 6928
rect 1443 6888 2412 6916
rect 1443 6885 1455 6888
rect 1397 6879 1455 6885
rect 2406 6876 2412 6888
rect 2464 6876 2470 6928
rect 4522 6876 4528 6928
rect 4580 6876 4586 6928
rect 5994 6876 6000 6928
rect 6052 6916 6058 6928
rect 6052 6888 6500 6916
rect 6052 6876 6058 6888
rect 1670 6848 1676 6860
rect 1631 6820 1676 6848
rect 1670 6808 1676 6820
rect 1728 6808 1734 6860
rect 3418 6848 3424 6860
rect 3379 6820 3424 6848
rect 3418 6808 3424 6820
rect 3476 6808 3482 6860
rect 3513 6851 3571 6857
rect 3513 6817 3525 6851
rect 3559 6848 3571 6851
rect 3559 6820 4016 6848
rect 3559 6817 3571 6820
rect 3513 6811 3571 6817
rect 3878 6780 3884 6792
rect 3839 6752 3884 6780
rect 3878 6740 3884 6752
rect 3936 6740 3942 6792
rect 3988 6780 4016 6820
rect 4890 6808 4896 6860
rect 4948 6848 4954 6860
rect 5353 6851 5411 6857
rect 5353 6848 5365 6851
rect 4948 6820 5365 6848
rect 4948 6808 4954 6820
rect 5353 6817 5365 6820
rect 5399 6817 5411 6851
rect 5353 6811 5411 6817
rect 4154 6780 4160 6792
rect 3988 6752 4160 6780
rect 4154 6740 4160 6752
rect 4212 6740 4218 6792
rect 6178 6780 6184 6792
rect 6139 6752 6184 6780
rect 6178 6740 6184 6752
rect 6236 6740 6242 6792
rect 6472 6712 6500 6888
rect 8110 6876 8116 6928
rect 8168 6876 8174 6928
rect 9214 6876 9220 6928
rect 9272 6916 9278 6928
rect 10226 6916 10232 6928
rect 9272 6888 10232 6916
rect 9272 6876 9278 6888
rect 10226 6876 10232 6888
rect 10284 6876 10290 6928
rect 7098 6808 7104 6860
rect 7156 6848 7162 6860
rect 7156 6820 7201 6848
rect 7156 6808 7162 6820
rect 7374 6808 7380 6860
rect 7432 6848 7438 6860
rect 7469 6851 7527 6857
rect 7469 6848 7481 6851
rect 7432 6820 7481 6848
rect 7432 6808 7438 6820
rect 7469 6817 7481 6820
rect 7515 6817 7527 6851
rect 7469 6811 7527 6817
rect 8941 6851 8999 6857
rect 8941 6817 8953 6851
rect 8987 6848 8999 6851
rect 9766 6848 9772 6860
rect 8987 6820 9772 6848
rect 8987 6817 8999 6820
rect 8941 6811 8999 6817
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 19334 6848 19340 6860
rect 16546 6820 19340 6848
rect 6825 6783 6883 6789
rect 6825 6749 6837 6783
rect 6871 6780 6883 6783
rect 7190 6780 7196 6792
rect 6871 6752 7196 6780
rect 6871 6749 6883 6752
rect 6825 6743 6883 6749
rect 7190 6740 7196 6752
rect 7248 6740 7254 6792
rect 9490 6740 9496 6792
rect 9548 6780 9554 6792
rect 9677 6783 9735 6789
rect 9677 6780 9689 6783
rect 9548 6752 9689 6780
rect 9548 6740 9554 6752
rect 9677 6749 9689 6752
rect 9723 6749 9735 6783
rect 9677 6743 9735 6749
rect 9861 6783 9919 6789
rect 9861 6749 9873 6783
rect 9907 6780 9919 6783
rect 10226 6780 10232 6792
rect 9907 6752 10232 6780
rect 9907 6749 9919 6752
rect 9861 6743 9919 6749
rect 10226 6740 10232 6752
rect 10284 6740 10290 6792
rect 16546 6712 16574 6820
rect 19334 6808 19340 6820
rect 19392 6808 19398 6860
rect 6472 6684 7052 6712
rect 1489 6647 1547 6653
rect 1489 6613 1501 6647
rect 1535 6644 1547 6647
rect 2038 6644 2044 6656
rect 1535 6616 2044 6644
rect 1535 6613 1547 6616
rect 1489 6607 1547 6613
rect 2038 6604 2044 6616
rect 2096 6604 2102 6656
rect 5917 6647 5975 6653
rect 5917 6613 5929 6647
rect 5963 6644 5975 6647
rect 6270 6644 6276 6656
rect 5963 6616 6276 6644
rect 5963 6613 5975 6616
rect 5917 6607 5975 6613
rect 6270 6604 6276 6616
rect 6328 6604 6334 6656
rect 7024 6644 7052 6684
rect 8404 6684 16574 6712
rect 8404 6644 8432 6684
rect 7024 6616 8432 6644
rect 8570 6604 8576 6656
rect 8628 6644 8634 6656
rect 9501 6647 9559 6653
rect 9501 6644 9513 6647
rect 8628 6616 9513 6644
rect 8628 6604 8634 6616
rect 9501 6613 9513 6616
rect 9547 6613 9559 6647
rect 9501 6607 9559 6613
rect 10045 6647 10103 6653
rect 10045 6613 10057 6647
rect 10091 6644 10103 6647
rect 10091 6616 10456 6644
rect 10091 6613 10103 6616
rect 10045 6607 10103 6613
rect 920 6554 10396 6576
rect 920 6502 2566 6554
rect 2618 6502 2630 6554
rect 2682 6502 2694 6554
rect 2746 6502 2758 6554
rect 2810 6502 2822 6554
rect 2874 6502 7566 6554
rect 7618 6502 7630 6554
rect 7682 6502 7694 6554
rect 7746 6502 7758 6554
rect 7810 6502 7822 6554
rect 7874 6502 10396 6554
rect 920 6480 10396 6502
rect 1670 6400 1676 6452
rect 1728 6440 1734 6452
rect 4246 6440 4252 6452
rect 1728 6412 4252 6440
rect 1728 6400 1734 6412
rect 4246 6400 4252 6412
rect 4304 6400 4310 6452
rect 5353 6443 5411 6449
rect 5353 6409 5365 6443
rect 5399 6440 5411 6443
rect 6178 6440 6184 6452
rect 5399 6412 6184 6440
rect 5399 6409 5411 6412
rect 5353 6403 5411 6409
rect 6178 6400 6184 6412
rect 6236 6400 6242 6452
rect 10428 6440 10456 6616
rect 8956 6412 10456 6440
rect 7834 6332 7840 6384
rect 7892 6372 7898 6384
rect 8757 6375 8815 6381
rect 8757 6372 8769 6375
rect 7892 6344 8769 6372
rect 7892 6332 7898 6344
rect 8757 6341 8769 6344
rect 8803 6341 8815 6375
rect 8757 6335 8815 6341
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6304 1731 6307
rect 2958 6304 2964 6316
rect 1719 6276 2964 6304
rect 1719 6273 1731 6276
rect 1673 6267 1731 6273
rect 2958 6264 2964 6276
rect 3016 6304 3022 6316
rect 3881 6307 3939 6313
rect 3016 6276 3648 6304
rect 3016 6264 3022 6276
rect 3620 6248 3648 6276
rect 3881 6273 3893 6307
rect 3927 6304 3939 6307
rect 5810 6304 5816 6316
rect 3927 6276 5816 6304
rect 3927 6273 3939 6276
rect 3881 6267 3939 6273
rect 5810 6264 5816 6276
rect 5868 6264 5874 6316
rect 8662 6264 8668 6316
rect 8720 6304 8726 6316
rect 8956 6304 8984 6412
rect 9030 6332 9036 6384
rect 9088 6372 9094 6384
rect 9125 6375 9183 6381
rect 9125 6372 9137 6375
rect 9088 6344 9137 6372
rect 9088 6332 9094 6344
rect 9125 6341 9137 6344
rect 9171 6341 9183 6375
rect 9125 6335 9183 6341
rect 9950 6304 9956 6316
rect 8720 6276 8984 6304
rect 9048 6276 9536 6304
rect 9911 6276 9956 6304
rect 8720 6264 8726 6276
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 1578 6236 1584 6248
rect 1443 6208 1584 6236
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 1578 6196 1584 6208
rect 1636 6196 1642 6248
rect 3602 6236 3608 6248
rect 3563 6208 3608 6236
rect 3602 6196 3608 6208
rect 3660 6196 3666 6248
rect 5445 6239 5503 6245
rect 5445 6205 5457 6239
rect 5491 6236 5503 6239
rect 5718 6236 5724 6248
rect 5491 6208 5724 6236
rect 5491 6205 5503 6208
rect 5445 6199 5503 6205
rect 5718 6196 5724 6208
rect 5776 6196 5782 6248
rect 7282 6236 7288 6248
rect 7243 6208 7288 6236
rect 7282 6196 7288 6208
rect 7340 6196 7346 6248
rect 7742 6196 7748 6248
rect 7800 6236 7806 6248
rect 8021 6239 8079 6245
rect 8021 6236 8033 6239
rect 7800 6208 8033 6236
rect 7800 6196 7806 6208
rect 8021 6205 8033 6208
rect 8067 6205 8079 6239
rect 8021 6199 8079 6205
rect 8205 6239 8263 6245
rect 8205 6205 8217 6239
rect 8251 6205 8263 6239
rect 9048 6236 9076 6276
rect 8864 6234 9076 6236
rect 8205 6199 8263 6205
rect 8496 6208 9076 6234
rect 9125 6239 9183 6245
rect 8496 6206 8892 6208
rect 1949 6171 2007 6177
rect 1949 6137 1961 6171
rect 1995 6137 2007 6171
rect 1949 6131 2007 6137
rect 1486 6100 1492 6112
rect 1447 6072 1492 6100
rect 1486 6060 1492 6072
rect 1544 6060 1550 6112
rect 1964 6100 1992 6131
rect 2958 6128 2964 6180
rect 3016 6128 3022 6180
rect 3970 6168 3976 6180
rect 3252 6140 3976 6168
rect 3252 6100 3280 6140
rect 3970 6128 3976 6140
rect 4028 6128 4034 6180
rect 7006 6168 7012 6180
rect 4264 6140 4370 6168
rect 6946 6140 7012 6168
rect 3418 6100 3424 6112
rect 1964 6072 3280 6100
rect 3379 6072 3424 6100
rect 3418 6060 3424 6072
rect 3476 6060 3482 6112
rect 3694 6060 3700 6112
rect 3752 6100 3758 6112
rect 4264 6100 4292 6140
rect 7006 6128 7012 6140
rect 7064 6128 7070 6180
rect 7834 6100 7840 6112
rect 7892 6109 7898 6112
rect 3752 6072 4292 6100
rect 7803 6072 7840 6100
rect 3752 6060 3758 6072
rect 7834 6060 7840 6072
rect 7892 6063 7903 6109
rect 8220 6100 8248 6199
rect 8496 6177 8524 6206
rect 9125 6205 9137 6239
rect 9171 6236 9183 6239
rect 9398 6236 9404 6248
rect 9171 6208 9404 6236
rect 9171 6205 9183 6208
rect 9125 6199 9183 6205
rect 9398 6196 9404 6208
rect 9456 6196 9462 6248
rect 9508 6245 9536 6276
rect 9950 6264 9956 6276
rect 10008 6264 10014 6316
rect 19702 6304 19708 6316
rect 16546 6276 19708 6304
rect 9493 6239 9551 6245
rect 9493 6205 9505 6239
rect 9539 6205 9551 6239
rect 16546 6236 16574 6276
rect 19702 6264 19708 6276
rect 19760 6264 19766 6316
rect 9493 6199 9551 6205
rect 12406 6208 16574 6236
rect 8481 6171 8539 6177
rect 8481 6137 8493 6171
rect 8527 6137 8539 6171
rect 8481 6131 8539 6137
rect 8573 6171 8631 6177
rect 8573 6137 8585 6171
rect 8619 6168 8631 6171
rect 9214 6168 9220 6180
rect 8619 6140 9220 6168
rect 8619 6137 8631 6140
rect 8573 6131 8631 6137
rect 9214 6128 9220 6140
rect 9272 6128 9278 6180
rect 9582 6168 9588 6180
rect 9324 6140 9588 6168
rect 9324 6100 9352 6140
rect 9582 6128 9588 6140
rect 9640 6128 9646 6180
rect 8220 6072 9352 6100
rect 7892 6060 7898 6063
rect 9398 6060 9404 6112
rect 9456 6100 9462 6112
rect 12406 6100 12434 6208
rect 19426 6100 19432 6112
rect 9456 6072 12434 6100
rect 16546 6072 19432 6100
rect 9456 6060 9462 6072
rect 920 6010 10396 6032
rect 920 5958 5066 6010
rect 5118 5958 5130 6010
rect 5182 5958 5194 6010
rect 5246 5958 5258 6010
rect 5310 5958 5322 6010
rect 5374 5958 10396 6010
rect 920 5936 10396 5958
rect 1394 5896 1400 5908
rect 1355 5868 1400 5896
rect 1394 5856 1400 5868
rect 1452 5856 1458 5908
rect 3878 5896 3884 5908
rect 1964 5868 3884 5896
rect 1964 5837 1992 5868
rect 3878 5856 3884 5868
rect 3936 5856 3942 5908
rect 7653 5899 7711 5905
rect 7653 5865 7665 5899
rect 7699 5896 7711 5899
rect 16546 5896 16574 6072
rect 19426 6060 19432 6072
rect 19484 6060 19490 6112
rect 7699 5868 16574 5896
rect 7699 5865 7711 5868
rect 7653 5859 7711 5865
rect 1949 5831 2007 5837
rect 1949 5797 1961 5831
rect 1995 5797 2007 5831
rect 1949 5791 2007 5797
rect 2958 5788 2964 5840
rect 3016 5788 3022 5840
rect 3326 5788 3332 5840
rect 3384 5828 3390 5840
rect 4249 5831 4307 5837
rect 4249 5828 4261 5831
rect 3384 5800 4261 5828
rect 3384 5788 3390 5800
rect 4249 5797 4261 5800
rect 4295 5797 4307 5831
rect 4249 5791 4307 5797
rect 6549 5831 6607 5837
rect 6549 5797 6561 5831
rect 6595 5828 6607 5831
rect 7282 5828 7288 5840
rect 6595 5800 7288 5828
rect 6595 5797 6607 5800
rect 6549 5791 6607 5797
rect 7282 5788 7288 5800
rect 7340 5788 7346 5840
rect 9677 5831 9735 5837
rect 9677 5797 9689 5831
rect 9723 5828 9735 5831
rect 9858 5828 9864 5840
rect 9723 5800 9864 5828
rect 9723 5797 9735 5800
rect 9677 5791 9735 5797
rect 9858 5788 9864 5800
rect 9916 5788 9922 5840
rect 1489 5763 1547 5769
rect 1489 5729 1501 5763
rect 1535 5729 1547 5763
rect 1489 5723 1547 5729
rect 3605 5763 3663 5769
rect 3605 5729 3617 5763
rect 3651 5760 3663 5763
rect 4062 5760 4068 5772
rect 3651 5732 4068 5760
rect 3651 5729 3663 5732
rect 3605 5723 3663 5729
rect 1504 5624 1532 5723
rect 4062 5720 4068 5732
rect 4120 5720 4126 5772
rect 4157 5763 4215 5769
rect 4157 5729 4169 5763
rect 4203 5760 4215 5763
rect 4890 5760 4896 5772
rect 4203 5732 4896 5760
rect 4203 5729 4215 5732
rect 4157 5723 4215 5729
rect 4890 5720 4896 5732
rect 4948 5720 4954 5772
rect 5350 5720 5356 5772
rect 5408 5760 5414 5772
rect 6181 5763 6239 5769
rect 5408 5732 6132 5760
rect 5408 5720 5414 5732
rect 1670 5692 1676 5704
rect 1631 5664 1676 5692
rect 1670 5652 1676 5664
rect 1728 5652 1734 5704
rect 1780 5664 3096 5692
rect 1780 5624 1808 5664
rect 3068 5636 3096 5664
rect 3694 5652 3700 5704
rect 3752 5692 3758 5704
rect 3789 5695 3847 5701
rect 3789 5692 3801 5695
rect 3752 5664 3801 5692
rect 3752 5652 3758 5664
rect 3789 5661 3801 5664
rect 3835 5661 3847 5695
rect 3970 5692 3976 5704
rect 3931 5664 3976 5692
rect 3789 5655 3847 5661
rect 3970 5652 3976 5664
rect 4028 5652 4034 5704
rect 4080 5692 4108 5720
rect 5074 5692 5080 5704
rect 4080 5664 5080 5692
rect 5074 5652 5080 5664
rect 5132 5652 5138 5704
rect 5994 5692 6000 5704
rect 5955 5664 6000 5692
rect 5994 5652 6000 5664
rect 6052 5652 6058 5704
rect 6104 5692 6132 5732
rect 6181 5729 6193 5763
rect 6227 5760 6239 5763
rect 7098 5760 7104 5772
rect 6227 5732 7104 5760
rect 6227 5729 6239 5732
rect 6181 5723 6239 5729
rect 7098 5720 7104 5732
rect 7156 5720 7162 5772
rect 8573 5763 8631 5769
rect 8573 5729 8585 5763
rect 8619 5760 8631 5763
rect 8754 5760 8760 5772
rect 8619 5732 8760 5760
rect 8619 5729 8631 5732
rect 8573 5723 8631 5729
rect 8754 5720 8760 5732
rect 8812 5720 8818 5772
rect 9030 5720 9036 5772
rect 9088 5760 9094 5772
rect 9490 5760 9496 5772
rect 9088 5732 9496 5760
rect 9088 5720 9094 5732
rect 9490 5720 9496 5732
rect 9548 5720 9554 5772
rect 10045 5763 10103 5769
rect 10045 5729 10057 5763
rect 10091 5760 10103 5763
rect 10410 5760 10416 5772
rect 10091 5732 10416 5760
rect 10091 5729 10103 5732
rect 10045 5723 10103 5729
rect 10410 5720 10416 5732
rect 10468 5720 10474 5772
rect 6365 5695 6423 5701
rect 6365 5692 6377 5695
rect 6104 5664 6377 5692
rect 6365 5661 6377 5664
rect 6411 5692 6423 5695
rect 7282 5692 7288 5704
rect 6411 5664 7288 5692
rect 6411 5661 6423 5664
rect 6365 5655 6423 5661
rect 7282 5652 7288 5664
rect 7340 5652 7346 5704
rect 7374 5652 7380 5704
rect 7432 5692 7438 5704
rect 9398 5692 9404 5704
rect 7432 5664 8800 5692
rect 9359 5664 9404 5692
rect 7432 5652 7438 5664
rect 1504 5596 1808 5624
rect 3050 5584 3056 5636
rect 3108 5584 3114 5636
rect 3421 5627 3479 5633
rect 3421 5593 3433 5627
rect 3467 5624 3479 5627
rect 5350 5624 5356 5636
rect 3467 5596 5356 5624
rect 3467 5593 3479 5596
rect 3421 5587 3479 5593
rect 5350 5584 5356 5596
rect 5408 5584 5414 5636
rect 7742 5584 7748 5636
rect 7800 5624 7806 5636
rect 8662 5624 8668 5636
rect 7800 5596 8668 5624
rect 7800 5584 7806 5596
rect 8662 5584 8668 5596
rect 8720 5584 8726 5636
rect 8772 5633 8800 5664
rect 9398 5652 9404 5664
rect 9456 5652 9462 5704
rect 9582 5692 9588 5704
rect 9508 5664 9588 5692
rect 9508 5633 9536 5664
rect 9582 5652 9588 5664
rect 9640 5652 9646 5704
rect 9766 5652 9772 5704
rect 9824 5692 9830 5704
rect 10134 5692 10140 5704
rect 9824 5664 10140 5692
rect 9824 5652 9830 5664
rect 10134 5652 10140 5664
rect 10192 5652 10198 5704
rect 13814 5652 13820 5704
rect 13872 5692 13878 5704
rect 17034 5692 17040 5704
rect 13872 5664 17040 5692
rect 13872 5652 13878 5664
rect 17034 5652 17040 5664
rect 17092 5652 17098 5704
rect 8757 5627 8815 5633
rect 8757 5593 8769 5627
rect 8803 5593 8815 5627
rect 8757 5587 8815 5593
rect 9493 5627 9551 5633
rect 9493 5593 9505 5627
rect 9539 5593 9551 5627
rect 10226 5624 10232 5636
rect 9493 5587 9551 5593
rect 9600 5596 10232 5624
rect 1670 5516 1676 5568
rect 1728 5556 1734 5568
rect 2130 5556 2136 5568
rect 1728 5528 2136 5556
rect 1728 5516 1734 5528
rect 2130 5516 2136 5528
rect 2188 5556 2194 5568
rect 3326 5556 3332 5568
rect 2188 5528 3332 5556
rect 2188 5516 2194 5528
rect 3326 5516 3332 5528
rect 3384 5516 3390 5568
rect 7282 5516 7288 5568
rect 7340 5556 7346 5568
rect 9600 5556 9628 5596
rect 10226 5584 10232 5596
rect 10284 5584 10290 5636
rect 11146 5584 11152 5636
rect 11204 5624 11210 5636
rect 16666 5624 16672 5636
rect 11204 5596 16672 5624
rect 11204 5584 11210 5596
rect 16666 5584 16672 5596
rect 16724 5584 16730 5636
rect 7340 5528 9628 5556
rect 9677 5559 9735 5565
rect 7340 5516 7346 5528
rect 9677 5525 9689 5559
rect 9723 5556 9735 5559
rect 10134 5556 10140 5568
rect 9723 5528 10140 5556
rect 9723 5525 9735 5528
rect 9677 5519 9735 5525
rect 10134 5516 10140 5528
rect 10192 5516 10198 5568
rect 13446 5516 13452 5568
rect 13504 5556 13510 5568
rect 16942 5556 16948 5568
rect 13504 5528 16948 5556
rect 13504 5516 13510 5528
rect 16942 5516 16948 5528
rect 17000 5516 17006 5568
rect 920 5466 10396 5488
rect 920 5414 2566 5466
rect 2618 5414 2630 5466
rect 2682 5414 2694 5466
rect 2746 5414 2758 5466
rect 2810 5414 2822 5466
rect 2874 5414 7566 5466
rect 7618 5414 7630 5466
rect 7682 5414 7694 5466
rect 7746 5414 7758 5466
rect 7810 5414 7822 5466
rect 7874 5414 10396 5466
rect 920 5392 10396 5414
rect 14090 5380 14096 5432
rect 14148 5420 14154 5432
rect 19518 5420 19524 5432
rect 14148 5392 19524 5420
rect 14148 5380 14154 5392
rect 19518 5380 19524 5392
rect 19576 5380 19582 5432
rect 2038 5312 2044 5364
rect 2096 5352 2102 5364
rect 2774 5352 2780 5364
rect 2096 5324 2780 5352
rect 2096 5312 2102 5324
rect 2774 5312 2780 5324
rect 2832 5312 2838 5364
rect 3513 5355 3571 5361
rect 3513 5321 3525 5355
rect 3559 5352 3571 5355
rect 4522 5352 4528 5364
rect 3559 5324 4528 5352
rect 3559 5321 3571 5324
rect 3513 5315 3571 5321
rect 4522 5312 4528 5324
rect 4580 5312 4586 5364
rect 5905 5355 5963 5361
rect 5905 5321 5917 5355
rect 5951 5352 5963 5355
rect 6638 5352 6644 5364
rect 5951 5324 6644 5352
rect 5951 5321 5963 5324
rect 5905 5315 5963 5321
rect 6638 5312 6644 5324
rect 6696 5312 6702 5364
rect 10045 5355 10103 5361
rect 10045 5321 10057 5355
rect 10091 5352 10103 5355
rect 11238 5352 11244 5364
rect 10091 5324 11244 5352
rect 10091 5321 10103 5324
rect 10045 5315 10103 5321
rect 11238 5312 11244 5324
rect 11296 5312 11302 5364
rect 20070 5352 20076 5364
rect 12406 5324 20076 5352
rect 5626 5244 5632 5296
rect 5684 5284 5690 5296
rect 12406 5284 12434 5324
rect 20070 5312 20076 5324
rect 20128 5312 20134 5364
rect 5684 5256 12434 5284
rect 5684 5244 5690 5256
rect 1762 5176 1768 5228
rect 1820 5216 1826 5228
rect 2498 5216 2504 5228
rect 1820 5188 2504 5216
rect 1820 5176 1826 5188
rect 2498 5176 2504 5188
rect 2556 5176 2562 5228
rect 3602 5176 3608 5228
rect 3660 5216 3666 5228
rect 3789 5219 3847 5225
rect 3789 5216 3801 5219
rect 3660 5188 3801 5216
rect 3660 5176 3666 5188
rect 3789 5185 3801 5188
rect 3835 5216 3847 5219
rect 5994 5216 6000 5228
rect 3835 5188 6000 5216
rect 3835 5185 3847 5188
rect 3789 5179 3847 5185
rect 5994 5176 6000 5188
rect 6052 5176 6058 5228
rect 8021 5219 8079 5225
rect 8021 5185 8033 5219
rect 8067 5216 8079 5219
rect 16574 5216 16580 5228
rect 8067 5188 16580 5216
rect 8067 5185 8079 5188
rect 8021 5179 8079 5185
rect 16574 5176 16580 5188
rect 16632 5176 16638 5228
rect 2958 5108 2964 5160
rect 3016 5148 3022 5160
rect 3329 5151 3387 5157
rect 3329 5148 3341 5151
rect 3016 5120 3341 5148
rect 3016 5108 3022 5120
rect 3329 5117 3341 5120
rect 3375 5117 3387 5151
rect 3329 5111 3387 5117
rect 3483 5151 3541 5157
rect 3483 5117 3495 5151
rect 3529 5148 3541 5151
rect 3694 5148 3700 5160
rect 3529 5120 3700 5148
rect 3529 5117 3541 5120
rect 3483 5111 3541 5117
rect 3694 5108 3700 5120
rect 3752 5108 3758 5160
rect 5902 5108 5908 5160
rect 5960 5148 5966 5160
rect 6089 5151 6147 5157
rect 6089 5148 6101 5151
rect 5960 5120 6101 5148
rect 5960 5108 5966 5120
rect 6089 5117 6101 5120
rect 6135 5117 6147 5151
rect 8294 5148 8300 5160
rect 8255 5120 8300 5148
rect 6089 5111 6147 5117
rect 8294 5108 8300 5120
rect 8352 5108 8358 5160
rect 4065 5083 4123 5089
rect 4065 5049 4077 5083
rect 4111 5080 4123 5083
rect 4111 5052 4292 5080
rect 4111 5049 4123 5052
rect 4065 5043 4123 5049
rect 4264 5012 4292 5052
rect 4522 5040 4528 5092
rect 4580 5040 4586 5092
rect 5813 5083 5871 5089
rect 5813 5080 5825 5083
rect 5368 5052 5825 5080
rect 4890 5012 4896 5024
rect 4264 4984 4896 5012
rect 4890 4972 4896 4984
rect 4948 4972 4954 5024
rect 5074 4972 5080 5024
rect 5132 5012 5138 5024
rect 5368 5012 5396 5052
rect 5813 5049 5825 5052
rect 5859 5049 5871 5083
rect 5813 5043 5871 5049
rect 6546 5040 6552 5092
rect 6604 5080 6610 5092
rect 8570 5080 8576 5092
rect 6604 5052 8576 5080
rect 6604 5040 6610 5052
rect 8570 5040 8576 5052
rect 8628 5040 8634 5092
rect 8754 5040 8760 5092
rect 8812 5080 8818 5092
rect 17310 5080 17316 5092
rect 8812 5052 12434 5080
rect 8812 5040 8818 5052
rect 5132 4984 5396 5012
rect 5537 5015 5595 5021
rect 5132 4972 5138 4984
rect 5537 4981 5549 5015
rect 5583 5012 5595 5015
rect 5626 5012 5632 5024
rect 5583 4984 5632 5012
rect 5583 4981 5595 4984
rect 5537 4975 5595 4981
rect 5626 4972 5632 4984
rect 5684 4972 5690 5024
rect 8294 4972 8300 5024
rect 8352 5012 8358 5024
rect 8846 5012 8852 5024
rect 8352 4984 8852 5012
rect 8352 4972 8358 4984
rect 8846 4972 8852 4984
rect 8904 4972 8910 5024
rect 12406 5012 12434 5052
rect 16546 5052 17316 5080
rect 16546 5012 16574 5052
rect 17310 5040 17316 5052
rect 17368 5040 17374 5092
rect 12406 4984 16574 5012
rect 3036 4922 10396 4944
rect 3036 4870 5066 4922
rect 5118 4870 5130 4922
rect 5182 4870 5194 4922
rect 5246 4870 5258 4922
rect 5310 4870 5322 4922
rect 5374 4870 10396 4922
rect 3036 4848 10396 4870
rect 3878 4768 3884 4820
rect 3936 4808 3942 4820
rect 3973 4811 4031 4817
rect 3973 4808 3985 4811
rect 3936 4780 3985 4808
rect 3936 4768 3942 4780
rect 3973 4777 3985 4780
rect 4019 4777 4031 4811
rect 4154 4808 4160 4820
rect 4115 4780 4160 4808
rect 3973 4771 4031 4777
rect 4154 4768 4160 4780
rect 4212 4768 4218 4820
rect 4246 4768 4252 4820
rect 4304 4768 4310 4820
rect 4522 4768 4528 4820
rect 4580 4808 4586 4820
rect 4982 4808 4988 4820
rect 4580 4780 4988 4808
rect 4580 4768 4586 4780
rect 4982 4768 4988 4780
rect 5040 4768 5046 4820
rect 6917 4811 6975 4817
rect 6917 4777 6929 4811
rect 6963 4808 6975 4811
rect 7006 4808 7012 4820
rect 6963 4780 7012 4808
rect 6963 4777 6975 4780
rect 6917 4771 6975 4777
rect 7006 4768 7012 4780
rect 7064 4768 7070 4820
rect 7374 4768 7380 4820
rect 7432 4808 7438 4820
rect 7561 4811 7619 4817
rect 7561 4808 7573 4811
rect 7432 4780 7573 4808
rect 7432 4768 7438 4780
rect 7561 4777 7573 4780
rect 7607 4777 7619 4811
rect 8110 4808 8116 4820
rect 8071 4780 8116 4808
rect 7561 4771 7619 4777
rect 8110 4768 8116 4780
rect 8168 4768 8174 4820
rect 9398 4768 9404 4820
rect 9456 4808 9462 4820
rect 10045 4811 10103 4817
rect 10045 4808 10057 4811
rect 9456 4780 10057 4808
rect 9456 4768 9462 4780
rect 10045 4777 10057 4780
rect 10091 4777 10103 4811
rect 10045 4771 10103 4777
rect 1302 4700 1308 4752
rect 1360 4740 1366 4752
rect 3602 4740 3608 4752
rect 1360 4712 3608 4740
rect 1360 4700 1366 4712
rect 3602 4700 3608 4712
rect 3660 4700 3666 4752
rect 2222 4632 2228 4684
rect 2280 4672 2286 4684
rect 2866 4672 2872 4684
rect 2280 4644 2872 4672
rect 2280 4632 2286 4644
rect 2866 4632 2872 4644
rect 2924 4632 2930 4684
rect 3418 4672 3424 4684
rect 3379 4644 3424 4672
rect 3418 4632 3424 4644
rect 3476 4632 3482 4684
rect 4264 4681 4292 4768
rect 5350 4700 5356 4752
rect 5408 4700 5414 4752
rect 5994 4700 6000 4752
rect 6052 4740 6058 4752
rect 6052 4712 8340 4740
rect 6052 4700 6058 4712
rect 4249 4675 4307 4681
rect 4249 4641 4261 4675
rect 4295 4672 4307 4675
rect 4614 4672 4620 4684
rect 4295 4644 4620 4672
rect 4295 4641 4307 4644
rect 4249 4635 4307 4641
rect 4614 4632 4620 4644
rect 4672 4632 4678 4684
rect 6181 4675 6239 4681
rect 6181 4641 6193 4675
rect 6227 4672 6239 4675
rect 6546 4672 6552 4684
rect 6227 4644 6552 4672
rect 6227 4641 6239 4644
rect 6181 4635 6239 4641
rect 6546 4632 6552 4644
rect 6604 4632 6610 4684
rect 7098 4632 7104 4684
rect 7156 4681 7162 4684
rect 7156 4675 7189 4681
rect 7177 4641 7189 4675
rect 7156 4635 7189 4641
rect 7156 4632 7162 4635
rect 7282 4632 7288 4684
rect 7340 4672 7346 4684
rect 7471 4675 7529 4681
rect 7340 4644 7385 4672
rect 7340 4632 7346 4644
rect 7471 4641 7483 4675
rect 7517 4672 7529 4675
rect 7745 4675 7803 4681
rect 7517 4644 7604 4672
rect 7517 4641 7529 4644
rect 7471 4635 7529 4641
rect 4338 4604 4344 4616
rect 4299 4576 4344 4604
rect 4338 4564 4344 4576
rect 4396 4564 4402 4616
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4604 4767 4607
rect 4890 4604 4896 4616
rect 4755 4576 4896 4604
rect 4755 4573 4767 4576
rect 4709 4567 4767 4573
rect 4890 4564 4896 4576
rect 4948 4564 4954 4616
rect 7576 4536 7604 4644
rect 7745 4641 7757 4675
rect 7791 4641 7803 4675
rect 7745 4635 7803 4641
rect 7899 4675 7957 4681
rect 7899 4641 7911 4675
rect 7945 4672 7957 4675
rect 8110 4672 8116 4684
rect 7945 4644 8116 4672
rect 7945 4641 7957 4644
rect 7899 4635 7957 4641
rect 7760 4604 7788 4635
rect 8110 4632 8116 4644
rect 8168 4632 8174 4684
rect 8312 4681 8340 4712
rect 9582 4700 9588 4752
rect 9640 4700 9646 4752
rect 8297 4675 8355 4681
rect 8297 4641 8309 4675
rect 8343 4641 8355 4675
rect 8297 4635 8355 4641
rect 8573 4607 8631 4613
rect 7760 4576 8248 4604
rect 8110 4536 8116 4548
rect 6472 4508 8116 4536
rect 2682 4428 2688 4480
rect 2740 4468 2746 4480
rect 6472 4468 6500 4508
rect 8110 4496 8116 4508
rect 8168 4496 8174 4548
rect 2740 4440 6500 4468
rect 2740 4428 2746 4440
rect 6546 4428 6552 4480
rect 6604 4468 6610 4480
rect 6741 4471 6799 4477
rect 6741 4468 6753 4471
rect 6604 4440 6753 4468
rect 6604 4428 6610 4440
rect 6741 4437 6753 4440
rect 6787 4437 6799 4471
rect 8220 4468 8248 4576
rect 8573 4573 8585 4607
rect 8619 4604 8631 4607
rect 10318 4604 10324 4616
rect 8619 4576 10324 4604
rect 8619 4573 8631 4576
rect 8573 4567 8631 4573
rect 10318 4564 10324 4576
rect 10376 4564 10382 4616
rect 8570 4468 8576 4480
rect 8220 4440 8576 4468
rect 6741 4431 6799 4437
rect 8570 4428 8576 4440
rect 8628 4468 8634 4480
rect 9582 4468 9588 4480
rect 8628 4440 9588 4468
rect 8628 4428 8634 4440
rect 9582 4428 9588 4440
rect 9640 4428 9646 4480
rect 3036 4378 10396 4400
rect 3036 4326 7566 4378
rect 7618 4326 7630 4378
rect 7682 4326 7694 4378
rect 7746 4326 7758 4378
rect 7810 4326 7822 4378
rect 7874 4326 10396 4378
rect 3036 4304 10396 4326
rect 5350 4264 5356 4276
rect 5311 4236 5356 4264
rect 5350 4224 5356 4236
rect 5408 4224 5414 4276
rect 5721 4267 5779 4273
rect 5721 4233 5733 4267
rect 5767 4264 5779 4267
rect 5810 4264 5816 4276
rect 5767 4236 5816 4264
rect 5767 4233 5779 4236
rect 5721 4227 5779 4233
rect 5810 4224 5816 4236
rect 5868 4224 5874 4276
rect 5994 4224 6000 4276
rect 6052 4264 6058 4276
rect 6052 4236 7328 4264
rect 6052 4224 6058 4236
rect 6362 4196 6368 4208
rect 5368 4168 6368 4196
rect 3326 4128 3332 4140
rect 3287 4100 3332 4128
rect 3326 4088 3332 4100
rect 3384 4128 3390 4140
rect 3970 4128 3976 4140
rect 3384 4100 3976 4128
rect 3384 4088 3390 4100
rect 3970 4088 3976 4100
rect 4028 4088 4034 4140
rect 4062 4088 4068 4140
rect 4120 4128 4126 4140
rect 5077 4131 5135 4137
rect 4120 4100 4844 4128
rect 4120 4088 4126 4100
rect 4816 4060 4844 4100
rect 5077 4097 5089 4131
rect 5123 4128 5135 4131
rect 5368 4128 5396 4168
rect 6362 4156 6368 4168
rect 6420 4156 6426 4208
rect 7300 4196 7328 4236
rect 8110 4224 8116 4276
rect 8168 4264 8174 4276
rect 8846 4264 8852 4276
rect 8168 4236 8852 4264
rect 8168 4224 8174 4236
rect 8846 4224 8852 4236
rect 8904 4224 8910 4276
rect 9398 4224 9404 4276
rect 9456 4264 9462 4276
rect 16850 4264 16856 4276
rect 9456 4236 16856 4264
rect 9456 4224 9462 4236
rect 16850 4224 16856 4236
rect 16908 4224 16914 4276
rect 8202 4196 8208 4208
rect 7300 4168 8208 4196
rect 8202 4156 8208 4168
rect 8260 4156 8266 4208
rect 5123 4100 5396 4128
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 5442 4088 5448 4140
rect 5500 4128 5506 4140
rect 6914 4128 6920 4140
rect 5500 4100 6408 4128
rect 6875 4100 6920 4128
rect 5500 4088 5506 4100
rect 5350 4069 5356 4072
rect 5169 4063 5227 4069
rect 5169 4060 5181 4063
rect 4816 4032 5181 4060
rect 5169 4029 5181 4032
rect 5215 4029 5227 4063
rect 5169 4023 5227 4029
rect 5323 4063 5356 4069
rect 5323 4029 5335 4063
rect 5323 4023 5356 4029
rect 5350 4020 5356 4023
rect 5408 4020 5414 4072
rect 5626 4020 5632 4072
rect 5684 4060 5690 4072
rect 6273 4063 6331 4069
rect 6273 4060 6285 4063
rect 5684 4032 6285 4060
rect 5684 4020 5690 4032
rect 6273 4029 6285 4032
rect 6319 4029 6331 4063
rect 6380 4060 6408 4100
rect 6914 4088 6920 4100
rect 6972 4088 6978 4140
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4128 7435 4131
rect 7466 4128 7472 4140
rect 7423 4100 7472 4128
rect 7423 4097 7435 4100
rect 7377 4091 7435 4097
rect 7466 4088 7472 4100
rect 7524 4088 7530 4140
rect 13538 4088 13544 4140
rect 13596 4128 13602 4140
rect 17126 4128 17132 4140
rect 13596 4100 17132 4128
rect 13596 4088 13602 4100
rect 17126 4088 17132 4100
rect 17184 4088 17190 4140
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6380 4032 6837 4060
rect 6273 4023 6331 4029
rect 6825 4029 6837 4032
rect 6871 4060 6883 4063
rect 6871 4032 7512 4060
rect 6871 4029 6883 4032
rect 6825 4023 6883 4029
rect 3605 3995 3663 4001
rect 3605 3961 3617 3995
rect 3651 3992 3663 3995
rect 3878 3992 3884 4004
rect 3651 3964 3884 3992
rect 3651 3961 3663 3964
rect 3605 3955 3663 3961
rect 3878 3952 3884 3964
rect 3936 3952 3942 4004
rect 4062 3952 4068 4004
rect 4120 3952 4126 4004
rect 6641 3995 6699 4001
rect 4908 3964 5764 3992
rect 2774 3884 2780 3936
rect 2832 3924 2838 3936
rect 3418 3924 3424 3936
rect 2832 3896 3424 3924
rect 2832 3884 2838 3896
rect 3418 3884 3424 3896
rect 3476 3884 3482 3936
rect 3694 3884 3700 3936
rect 3752 3924 3758 3936
rect 4908 3924 4936 3964
rect 3752 3896 4936 3924
rect 3752 3884 3758 3896
rect 5258 3884 5264 3936
rect 5316 3924 5322 3936
rect 5626 3924 5632 3936
rect 5316 3896 5632 3924
rect 5316 3884 5322 3896
rect 5626 3884 5632 3896
rect 5684 3884 5690 3936
rect 5736 3924 5764 3964
rect 6641 3961 6653 3995
rect 6687 3992 6699 3995
rect 6730 3992 6736 4004
rect 6687 3964 6736 3992
rect 6687 3961 6699 3964
rect 6641 3955 6699 3961
rect 6730 3952 6736 3964
rect 6788 3952 6794 4004
rect 7193 3995 7251 4001
rect 7193 3961 7205 3995
rect 7239 3992 7251 3995
rect 7484 3992 7512 4032
rect 8478 3992 8484 4004
rect 7239 3964 7420 3992
rect 7484 3964 8484 3992
rect 7239 3961 7251 3964
rect 7193 3955 7251 3961
rect 6549 3927 6607 3933
rect 6549 3924 6561 3927
rect 5736 3896 6561 3924
rect 6549 3893 6561 3896
rect 6595 3893 6607 3927
rect 7392 3924 7420 3964
rect 8478 3952 8484 3964
rect 8536 3992 8542 4004
rect 8536 3964 9628 3992
rect 8536 3952 8542 3964
rect 9600 3936 9628 3964
rect 9214 3924 9220 3936
rect 7392 3896 9220 3924
rect 6549 3887 6607 3893
rect 9214 3884 9220 3896
rect 9272 3884 9278 3936
rect 9582 3884 9588 3936
rect 9640 3884 9646 3936
rect 3036 3834 10396 3856
rect 3036 3782 5066 3834
rect 5118 3782 5130 3834
rect 5182 3782 5194 3834
rect 5246 3782 5258 3834
rect 5310 3782 5322 3834
rect 5374 3782 10396 3834
rect 3036 3760 10396 3782
rect 3142 3680 3148 3732
rect 3200 3720 3206 3732
rect 3329 3723 3387 3729
rect 3329 3720 3341 3723
rect 3200 3692 3341 3720
rect 3200 3680 3206 3692
rect 3329 3689 3341 3692
rect 3375 3689 3387 3723
rect 3329 3683 3387 3689
rect 3970 3680 3976 3732
rect 4028 3720 4034 3732
rect 5997 3723 6055 3729
rect 4028 3692 5120 3720
rect 4028 3680 4034 3692
rect 3418 3612 3424 3664
rect 3476 3652 3482 3664
rect 4801 3655 4859 3661
rect 3476 3624 3634 3652
rect 3476 3612 3482 3624
rect 4801 3621 4813 3655
rect 4847 3652 4859 3655
rect 4890 3652 4896 3664
rect 4847 3624 4896 3652
rect 4847 3621 4859 3624
rect 4801 3615 4859 3621
rect 4890 3612 4896 3624
rect 4948 3612 4954 3664
rect 5092 3593 5120 3692
rect 5997 3689 6009 3723
rect 6043 3720 6055 3723
rect 6086 3720 6092 3732
rect 6043 3692 6092 3720
rect 6043 3689 6055 3692
rect 5997 3683 6055 3689
rect 6086 3680 6092 3692
rect 6144 3680 6150 3732
rect 7190 3720 7196 3732
rect 7151 3692 7196 3720
rect 7190 3680 7196 3692
rect 7248 3680 7254 3732
rect 8481 3723 8539 3729
rect 8481 3689 8493 3723
rect 8527 3720 8539 3723
rect 9030 3720 9036 3732
rect 8527 3692 9036 3720
rect 8527 3689 8539 3692
rect 8481 3683 8539 3689
rect 9030 3680 9036 3692
rect 9088 3720 9094 3732
rect 9953 3723 10011 3729
rect 9088 3692 9536 3720
rect 9088 3680 9094 3692
rect 7282 3612 7288 3664
rect 7340 3652 7346 3664
rect 7340 3624 9076 3652
rect 7340 3612 7346 3624
rect 5077 3587 5135 3593
rect 5077 3553 5089 3587
rect 5123 3553 5135 3587
rect 5077 3547 5135 3553
rect 5442 3544 5448 3596
rect 5500 3584 5506 3596
rect 5905 3587 5963 3593
rect 5905 3584 5917 3587
rect 5500 3556 5917 3584
rect 5500 3544 5506 3556
rect 5905 3553 5917 3556
rect 5951 3553 5963 3587
rect 5905 3547 5963 3553
rect 8113 3587 8171 3593
rect 8113 3553 8125 3587
rect 8159 3584 8171 3587
rect 8389 3587 8447 3593
rect 8159 3556 8340 3584
rect 8159 3553 8171 3556
rect 8113 3547 8171 3553
rect 3050 3476 3056 3528
rect 3108 3516 3114 3528
rect 3786 3516 3792 3528
rect 3108 3488 3792 3516
rect 3108 3476 3114 3488
rect 3786 3476 3792 3488
rect 3844 3476 3850 3528
rect 4062 3476 4068 3528
rect 4120 3516 4126 3528
rect 5350 3516 5356 3528
rect 4120 3488 5356 3516
rect 4120 3476 4126 3488
rect 5350 3476 5356 3488
rect 5408 3476 5414 3528
rect 5626 3476 5632 3528
rect 5684 3516 5690 3528
rect 5721 3519 5779 3525
rect 5721 3516 5733 3519
rect 5684 3488 5733 3516
rect 5684 3476 5690 3488
rect 5721 3485 5733 3488
rect 5767 3485 5779 3519
rect 5721 3479 5779 3485
rect 4982 3340 4988 3392
rect 5040 3380 5046 3392
rect 5169 3383 5227 3389
rect 5169 3380 5181 3383
rect 5040 3352 5181 3380
rect 5040 3340 5046 3352
rect 5169 3349 5181 3352
rect 5215 3349 5227 3383
rect 8312 3380 8340 3556
rect 8389 3553 8401 3587
rect 8435 3553 8447 3587
rect 8846 3584 8852 3596
rect 8807 3556 8852 3584
rect 8389 3547 8447 3553
rect 8404 3516 8432 3547
rect 8846 3544 8852 3556
rect 8904 3544 8910 3596
rect 9048 3593 9076 3624
rect 9033 3587 9091 3593
rect 9033 3553 9045 3587
rect 9079 3553 9091 3587
rect 9214 3584 9220 3596
rect 9127 3556 9220 3584
rect 9033 3547 9091 3553
rect 9214 3544 9220 3556
rect 9272 3584 9278 3596
rect 9508 3593 9536 3692
rect 9953 3689 9965 3723
rect 9999 3720 10011 3723
rect 10042 3720 10048 3732
rect 9999 3692 10048 3720
rect 9999 3689 10011 3692
rect 9953 3683 10011 3689
rect 10042 3680 10048 3692
rect 10100 3680 10106 3732
rect 9582 3612 9588 3664
rect 9640 3652 9646 3664
rect 9640 3624 9904 3652
rect 9640 3612 9646 3624
rect 9876 3593 9904 3624
rect 9493 3587 9551 3593
rect 9272 3556 9444 3584
rect 9272 3544 9278 3556
rect 9122 3516 9128 3528
rect 8404 3488 9128 3516
rect 9122 3476 9128 3488
rect 9180 3476 9186 3528
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3485 9367 3519
rect 9416 3516 9444 3556
rect 9493 3553 9505 3587
rect 9539 3553 9551 3587
rect 9493 3547 9551 3553
rect 9861 3587 9919 3593
rect 9861 3553 9873 3587
rect 9907 3553 9919 3587
rect 9861 3547 9919 3553
rect 22094 3516 22100 3528
rect 9416 3488 22100 3516
rect 9309 3479 9367 3485
rect 9214 3408 9220 3460
rect 9272 3448 9278 3460
rect 9324 3448 9352 3479
rect 22094 3476 22100 3488
rect 22152 3476 22158 3528
rect 10410 3448 10416 3460
rect 9272 3420 9352 3448
rect 9416 3420 10416 3448
rect 9272 3408 9278 3420
rect 9416 3380 9444 3420
rect 10410 3408 10416 3420
rect 10468 3408 10474 3460
rect 8312 3352 9444 3380
rect 9677 3383 9735 3389
rect 5169 3343 5227 3349
rect 9677 3349 9689 3383
rect 9723 3380 9735 3383
rect 10502 3380 10508 3392
rect 9723 3352 10508 3380
rect 9723 3349 9735 3352
rect 9677 3343 9735 3349
rect 10502 3340 10508 3352
rect 10560 3340 10566 3392
rect 3036 3290 10396 3312
rect 3036 3238 7566 3290
rect 7618 3238 7630 3290
rect 7682 3238 7694 3290
rect 7746 3238 7758 3290
rect 7810 3238 7822 3290
rect 7874 3238 10396 3290
rect 3036 3216 10396 3238
rect 3234 3136 3240 3188
rect 3292 3176 3298 3188
rect 3329 3179 3387 3185
rect 3329 3176 3341 3179
rect 3292 3148 3341 3176
rect 3292 3136 3298 3148
rect 3329 3145 3341 3148
rect 3375 3145 3387 3179
rect 3329 3139 3387 3145
rect 4430 3136 4436 3188
rect 4488 3176 4494 3188
rect 5261 3179 5319 3185
rect 5261 3176 5273 3179
rect 4488 3148 5273 3176
rect 4488 3136 4494 3148
rect 5261 3145 5273 3148
rect 5307 3145 5319 3179
rect 5261 3139 5319 3145
rect 5350 3136 5356 3188
rect 5408 3176 5414 3188
rect 9674 3176 9680 3188
rect 5408 3148 9680 3176
rect 5408 3136 5414 3148
rect 9674 3136 9680 3148
rect 9732 3136 9738 3188
rect 10045 3179 10103 3185
rect 10045 3145 10057 3179
rect 10091 3176 10103 3179
rect 11054 3176 11060 3188
rect 10091 3148 11060 3176
rect 10091 3145 10103 3148
rect 10045 3139 10103 3145
rect 11054 3136 11060 3148
rect 11112 3136 11118 3188
rect 5721 3111 5779 3117
rect 5721 3077 5733 3111
rect 5767 3108 5779 3111
rect 6638 3108 6644 3120
rect 5767 3080 6644 3108
rect 5767 3077 5779 3080
rect 5721 3071 5779 3077
rect 6638 3068 6644 3080
rect 6696 3068 6702 3120
rect 4062 3000 4068 3052
rect 4120 3040 4126 3052
rect 5077 3043 5135 3049
rect 5077 3040 5089 3043
rect 4120 3012 5089 3040
rect 4120 3000 4126 3012
rect 5077 3009 5089 3012
rect 5123 3009 5135 3043
rect 5077 3003 5135 3009
rect 7377 3043 7435 3049
rect 7377 3009 7389 3043
rect 7423 3040 7435 3043
rect 11146 3040 11152 3052
rect 7423 3012 11152 3040
rect 7423 3009 7435 3012
rect 7377 3003 7435 3009
rect 11146 3000 11152 3012
rect 11204 3000 11210 3052
rect 5902 2972 5908 2984
rect 5863 2944 5908 2972
rect 5902 2932 5908 2944
rect 5960 2932 5966 2984
rect 8018 2972 8024 2984
rect 7979 2944 8024 2972
rect 8018 2932 8024 2944
rect 8076 2932 8082 2984
rect 8481 2975 8539 2981
rect 8481 2941 8493 2975
rect 8527 2972 8539 2975
rect 8938 2972 8944 2984
rect 8527 2944 8944 2972
rect 8527 2941 8539 2944
rect 8481 2935 8539 2941
rect 8938 2932 8944 2944
rect 8996 2932 9002 2984
rect 4246 2864 4252 2916
rect 4304 2864 4310 2916
rect 4801 2907 4859 2913
rect 4801 2873 4813 2907
rect 4847 2873 4859 2907
rect 4801 2867 4859 2873
rect 4816 2836 4844 2867
rect 4890 2864 4896 2916
rect 4948 2904 4954 2916
rect 5353 2907 5411 2913
rect 5353 2904 5365 2907
rect 4948 2876 5365 2904
rect 4948 2864 4954 2876
rect 5353 2873 5365 2876
rect 5399 2873 5411 2907
rect 5353 2867 5411 2873
rect 6454 2836 6460 2848
rect 4816 2808 6460 2836
rect 6454 2796 6460 2808
rect 6512 2796 6518 2848
rect 3036 2746 10396 2768
rect 3036 2694 5066 2746
rect 5118 2694 5130 2746
rect 5182 2694 5194 2746
rect 5246 2694 5258 2746
rect 5310 2694 5322 2746
rect 5374 2694 10396 2746
rect 3036 2672 10396 2694
rect 3970 2632 3976 2644
rect 3804 2604 3976 2632
rect 3050 2524 3056 2576
rect 3108 2564 3114 2576
rect 3804 2573 3832 2604
rect 3970 2592 3976 2604
rect 4028 2592 4034 2644
rect 4249 2635 4307 2641
rect 4249 2601 4261 2635
rect 4295 2601 4307 2635
rect 4249 2595 4307 2601
rect 3789 2567 3847 2573
rect 3108 2536 3740 2564
rect 3108 2524 3114 2536
rect 3712 2508 3740 2536
rect 3789 2533 3801 2567
rect 3835 2533 3847 2567
rect 3789 2527 3847 2533
rect 4157 2567 4215 2573
rect 4157 2533 4169 2567
rect 4203 2533 4215 2567
rect 4264 2564 4292 2595
rect 4338 2592 4344 2644
rect 4396 2632 4402 2644
rect 5261 2635 5319 2641
rect 5261 2632 5273 2635
rect 4396 2604 5273 2632
rect 4396 2592 4402 2604
rect 5261 2601 5273 2604
rect 5307 2601 5319 2635
rect 5534 2632 5540 2644
rect 5495 2604 5540 2632
rect 5261 2595 5319 2601
rect 5534 2592 5540 2604
rect 5592 2592 5598 2644
rect 5626 2592 5632 2644
rect 5684 2592 5690 2644
rect 5718 2592 5724 2644
rect 5776 2632 5782 2644
rect 5997 2635 6055 2641
rect 5997 2632 6009 2635
rect 5776 2604 6009 2632
rect 5776 2592 5782 2604
rect 5997 2601 6009 2604
rect 6043 2601 6055 2635
rect 8386 2632 8392 2644
rect 8347 2604 8392 2632
rect 5997 2595 6055 2601
rect 8386 2592 8392 2604
rect 8444 2592 8450 2644
rect 8662 2632 8668 2644
rect 8623 2604 8668 2632
rect 8662 2592 8668 2604
rect 8720 2592 8726 2644
rect 9401 2635 9459 2641
rect 9401 2601 9413 2635
rect 9447 2632 9459 2635
rect 9490 2632 9496 2644
rect 9447 2604 9496 2632
rect 9447 2601 9459 2604
rect 9401 2595 9459 2601
rect 9490 2592 9496 2604
rect 9548 2592 9554 2644
rect 9674 2592 9680 2644
rect 9732 2632 9738 2644
rect 9769 2635 9827 2641
rect 9769 2632 9781 2635
rect 9732 2604 9781 2632
rect 9732 2592 9738 2604
rect 9769 2601 9781 2604
rect 9815 2632 9827 2635
rect 10778 2632 10784 2644
rect 9815 2604 10784 2632
rect 9815 2601 9827 2604
rect 9769 2595 9827 2601
rect 10778 2592 10784 2604
rect 10836 2592 10842 2644
rect 5644 2564 5672 2592
rect 4264 2536 5672 2564
rect 5813 2567 5871 2573
rect 4157 2527 4215 2533
rect 5813 2533 5825 2567
rect 5859 2564 5871 2567
rect 6638 2564 6644 2576
rect 5859 2536 6644 2564
rect 5859 2533 5871 2536
rect 5813 2527 5871 2533
rect 3418 2496 3424 2508
rect 3379 2468 3424 2496
rect 3418 2456 3424 2468
rect 3476 2456 3482 2508
rect 3694 2496 3700 2508
rect 3607 2468 3700 2496
rect 3694 2456 3700 2468
rect 3752 2486 3758 2508
rect 4172 2496 4200 2527
rect 6638 2524 6644 2536
rect 6696 2524 6702 2576
rect 7374 2524 7380 2576
rect 7432 2564 7438 2576
rect 7432 2536 8892 2564
rect 7432 2524 7438 2536
rect 3804 2486 4200 2496
rect 3752 2468 4200 2486
rect 4617 2499 4675 2505
rect 3752 2458 3832 2468
rect 4617 2465 4629 2499
rect 4663 2465 4675 2499
rect 4890 2496 4896 2508
rect 4851 2468 4896 2496
rect 4617 2459 4675 2465
rect 3752 2456 3758 2458
rect 2866 2388 2872 2440
rect 2924 2428 2930 2440
rect 4433 2431 4491 2437
rect 4433 2428 4445 2431
rect 2924 2400 4445 2428
rect 2924 2388 2930 2400
rect 4433 2397 4445 2400
rect 4479 2397 4491 2431
rect 4433 2391 4491 2397
rect 4632 2360 4660 2459
rect 4890 2456 4896 2468
rect 4948 2456 4954 2508
rect 5350 2496 5356 2508
rect 5311 2468 5356 2496
rect 5350 2456 5356 2468
rect 5408 2496 5414 2508
rect 5629 2499 5687 2505
rect 5629 2496 5641 2499
rect 5408 2468 5641 2496
rect 5408 2456 5414 2468
rect 5629 2465 5641 2468
rect 5675 2496 5687 2499
rect 5905 2499 5963 2505
rect 5905 2496 5917 2499
rect 5675 2468 5917 2496
rect 5675 2465 5687 2468
rect 5629 2459 5687 2465
rect 5905 2465 5917 2468
rect 5951 2465 5963 2499
rect 6546 2496 6552 2508
rect 6507 2468 6552 2496
rect 5905 2459 5963 2465
rect 6546 2456 6552 2468
rect 6604 2456 6610 2508
rect 8478 2496 8484 2508
rect 8439 2468 8484 2496
rect 8478 2456 8484 2468
rect 8536 2456 8542 2508
rect 8570 2456 8576 2508
rect 8628 2496 8634 2508
rect 8754 2496 8760 2508
rect 8628 2468 8760 2496
rect 8628 2456 8634 2468
rect 8754 2456 8760 2468
rect 8812 2456 8818 2508
rect 8864 2496 8892 2536
rect 9030 2524 9036 2576
rect 9088 2564 9094 2576
rect 9125 2567 9183 2573
rect 9125 2564 9137 2567
rect 9088 2536 9137 2564
rect 9088 2524 9094 2536
rect 9125 2533 9137 2536
rect 9171 2533 9183 2567
rect 16666 2564 16672 2576
rect 9125 2527 9183 2533
rect 12406 2536 16672 2564
rect 9493 2499 9551 2505
rect 9493 2496 9505 2499
rect 8864 2468 9505 2496
rect 9493 2465 9505 2468
rect 9539 2496 9551 2499
rect 9861 2499 9919 2505
rect 9861 2496 9873 2499
rect 9539 2468 9873 2496
rect 9539 2465 9551 2468
rect 9493 2459 9551 2465
rect 9861 2465 9873 2468
rect 9907 2465 9919 2499
rect 9861 2459 9919 2465
rect 5718 2388 5724 2440
rect 5776 2428 5782 2440
rect 12406 2428 12434 2536
rect 16666 2524 16672 2536
rect 16724 2524 16730 2576
rect 5776 2400 12434 2428
rect 5776 2388 5782 2400
rect 5994 2360 6000 2372
rect 4632 2332 6000 2360
rect 5994 2320 6000 2332
rect 6052 2320 6058 2372
rect 8113 2363 8171 2369
rect 8113 2329 8125 2363
rect 8159 2360 8171 2363
rect 13814 2360 13820 2372
rect 8159 2332 13820 2360
rect 8159 2329 8171 2332
rect 8113 2323 8171 2329
rect 13814 2320 13820 2332
rect 13872 2320 13878 2372
rect 3418 2252 3424 2304
rect 3476 2292 3482 2304
rect 3513 2295 3571 2301
rect 3513 2292 3525 2295
rect 3476 2264 3525 2292
rect 3476 2252 3482 2264
rect 3513 2261 3525 2264
rect 3559 2261 3571 2295
rect 3878 2292 3884 2304
rect 3839 2264 3884 2292
rect 3513 2255 3571 2261
rect 3878 2252 3884 2264
rect 3936 2252 3942 2304
rect 4982 2292 4988 2304
rect 4943 2264 4988 2292
rect 4982 2252 4988 2264
rect 5040 2252 5046 2304
rect 5074 2252 5080 2304
rect 5132 2292 5138 2304
rect 6822 2292 6828 2304
rect 5132 2264 6828 2292
rect 5132 2252 5138 2264
rect 6822 2252 6828 2264
rect 6880 2252 6886 2304
rect 8662 2252 8668 2304
rect 8720 2292 8726 2304
rect 9033 2295 9091 2301
rect 9033 2292 9045 2295
rect 8720 2264 9045 2292
rect 8720 2252 8726 2264
rect 9033 2261 9045 2264
rect 9079 2261 9091 2295
rect 9033 2255 9091 2261
rect 3036 2202 10396 2224
rect 3036 2150 7566 2202
rect 7618 2150 7630 2202
rect 7682 2150 7694 2202
rect 7746 2150 7758 2202
rect 7810 2150 7822 2202
rect 7874 2150 10396 2202
rect 3036 2128 10396 2150
rect 2682 2048 2688 2100
rect 2740 2088 2746 2100
rect 3881 2091 3939 2097
rect 3881 2088 3893 2091
rect 2740 2060 3893 2088
rect 2740 2048 2746 2060
rect 3881 2057 3893 2060
rect 3927 2057 3939 2091
rect 3881 2051 3939 2057
rect 4249 2091 4307 2097
rect 4249 2057 4261 2091
rect 4295 2088 4307 2091
rect 4430 2088 4436 2100
rect 4295 2060 4436 2088
rect 4295 2057 4307 2060
rect 4249 2051 4307 2057
rect 4430 2048 4436 2060
rect 4488 2048 4494 2100
rect 4798 2088 4804 2100
rect 4759 2060 4804 2088
rect 4798 2048 4804 2060
rect 4856 2048 4862 2100
rect 5353 2091 5411 2097
rect 5353 2057 5365 2091
rect 5399 2088 5411 2091
rect 5442 2088 5448 2100
rect 5399 2060 5448 2088
rect 5399 2057 5411 2060
rect 5353 2051 5411 2057
rect 5442 2048 5448 2060
rect 5500 2048 5506 2100
rect 5813 2091 5871 2097
rect 5813 2057 5825 2091
rect 5859 2088 5871 2091
rect 5902 2088 5908 2100
rect 5859 2060 5908 2088
rect 5859 2057 5871 2060
rect 5813 2051 5871 2057
rect 5902 2048 5908 2060
rect 5960 2048 5966 2100
rect 5994 2048 6000 2100
rect 6052 2088 6058 2100
rect 6052 2060 7144 2088
rect 6052 2048 6058 2060
rect 3510 1980 3516 2032
rect 3568 2020 3574 2032
rect 4525 2023 4583 2029
rect 4525 2020 4537 2023
rect 3568 1992 4537 2020
rect 3568 1980 3574 1992
rect 4525 1989 4537 1992
rect 4571 1989 4583 2023
rect 4525 1983 4583 1989
rect 4706 1980 4712 2032
rect 4764 2020 4770 2032
rect 5077 2023 5135 2029
rect 5077 2020 5089 2023
rect 4764 1992 5089 2020
rect 4764 1980 4770 1992
rect 5077 1989 5089 1992
rect 5123 1989 5135 2023
rect 5460 2020 5488 2048
rect 6086 2020 6092 2032
rect 5460 1992 6092 2020
rect 5077 1983 5135 1989
rect 6086 1980 6092 1992
rect 6144 1980 6150 2032
rect 6917 2023 6975 2029
rect 6917 1989 6929 2023
rect 6963 2020 6975 2023
rect 7006 2020 7012 2032
rect 6963 1992 7012 2020
rect 6963 1989 6975 1992
rect 6917 1983 6975 1989
rect 7006 1980 7012 1992
rect 7064 1980 7070 2032
rect 7116 2020 7144 2060
rect 7466 2048 7472 2100
rect 7524 2088 7530 2100
rect 16758 2088 16764 2100
rect 7524 2060 16764 2088
rect 7524 2048 7530 2060
rect 16758 2048 16764 2060
rect 16816 2048 16822 2100
rect 20622 2020 20628 2032
rect 7116 1992 20628 2020
rect 20622 1980 20628 1992
rect 20680 1980 20686 2032
rect 3878 1912 3884 1964
rect 3936 1952 3942 1964
rect 7098 1952 7104 1964
rect 3936 1924 7104 1952
rect 3936 1912 3942 1924
rect 7098 1912 7104 1924
rect 7156 1912 7162 1964
rect 9401 1955 9459 1961
rect 9401 1921 9413 1955
rect 9447 1952 9459 1955
rect 13630 1952 13636 1964
rect 9447 1924 13636 1952
rect 9447 1921 9459 1924
rect 9401 1915 9459 1921
rect 13630 1912 13636 1924
rect 13688 1912 13694 1964
rect 2682 1844 2688 1896
rect 2740 1884 2746 1896
rect 3789 1887 3847 1893
rect 3789 1884 3801 1887
rect 2740 1856 3801 1884
rect 2740 1844 2746 1856
rect 3789 1853 3801 1856
rect 3835 1853 3847 1887
rect 4062 1884 4068 1896
rect 4023 1856 4068 1884
rect 3789 1847 3847 1853
rect 4062 1844 4068 1856
rect 4120 1844 4126 1896
rect 4614 1884 4620 1896
rect 4575 1856 4620 1884
rect 4614 1844 4620 1856
rect 4672 1884 4678 1896
rect 4893 1887 4951 1893
rect 4893 1884 4905 1887
rect 4672 1856 4905 1884
rect 4672 1844 4678 1856
rect 4893 1853 4905 1856
rect 4939 1884 4951 1887
rect 5169 1887 5227 1893
rect 5169 1884 5181 1887
rect 4939 1856 5181 1884
rect 4939 1853 4951 1856
rect 4893 1847 4951 1853
rect 5169 1853 5181 1856
rect 5215 1884 5227 1887
rect 5350 1884 5356 1896
rect 5215 1856 5356 1884
rect 5215 1853 5227 1856
rect 5169 1847 5227 1853
rect 5350 1844 5356 1856
rect 5408 1844 5414 1896
rect 7926 1884 7932 1896
rect 7887 1856 7932 1884
rect 7926 1844 7932 1856
rect 7984 1844 7990 1896
rect 9766 1884 9772 1896
rect 9727 1856 9772 1884
rect 9766 1844 9772 1856
rect 9824 1844 9830 1896
rect 3234 1776 3240 1828
rect 3292 1816 3298 1828
rect 3421 1819 3479 1825
rect 3421 1816 3433 1819
rect 3292 1788 3433 1816
rect 3292 1776 3298 1788
rect 3421 1785 3433 1788
rect 3467 1785 3479 1819
rect 3421 1779 3479 1785
rect 3602 1776 3608 1828
rect 3660 1816 3666 1828
rect 3660 1788 5580 1816
rect 3660 1776 3666 1788
rect 3513 1751 3571 1757
rect 3513 1717 3525 1751
rect 3559 1748 3571 1751
rect 5074 1748 5080 1760
rect 3559 1720 5080 1748
rect 3559 1717 3571 1720
rect 3513 1711 3571 1717
rect 5074 1708 5080 1720
rect 5132 1708 5138 1760
rect 5552 1748 5580 1788
rect 7374 1776 7380 1828
rect 7432 1816 7438 1828
rect 7432 1788 12434 1816
rect 7432 1776 7438 1788
rect 8294 1748 8300 1760
rect 5552 1720 8300 1748
rect 8294 1708 8300 1720
rect 8352 1708 8358 1760
rect 12406 1748 12434 1788
rect 13446 1748 13452 1760
rect 12406 1720 13452 1748
rect 13446 1708 13452 1720
rect 13504 1708 13510 1760
rect 3036 1658 10396 1680
rect 3036 1606 5066 1658
rect 5118 1606 5130 1658
rect 5182 1606 5194 1658
rect 5246 1606 5258 1658
rect 5310 1606 5322 1658
rect 5374 1606 10396 1658
rect 3036 1584 10396 1606
rect 14 1504 20 1556
rect 72 1544 78 1556
rect 3234 1544 3240 1556
rect 72 1516 3240 1544
rect 72 1504 78 1516
rect 3234 1504 3240 1516
rect 3292 1504 3298 1556
rect 4065 1547 4123 1553
rect 4065 1513 4077 1547
rect 4111 1544 4123 1547
rect 4890 1544 4896 1556
rect 4111 1516 4896 1544
rect 4111 1513 4123 1516
rect 4065 1507 4123 1513
rect 4890 1504 4896 1516
rect 4948 1504 4954 1556
rect 5169 1547 5227 1553
rect 5169 1513 5181 1547
rect 5215 1544 5227 1547
rect 5718 1544 5724 1556
rect 5215 1516 5724 1544
rect 5215 1513 5227 1516
rect 5169 1507 5227 1513
rect 5718 1504 5724 1516
rect 5776 1504 5782 1556
rect 7466 1544 7472 1556
rect 6012 1516 7472 1544
rect 1026 1436 1032 1488
rect 1084 1476 1090 1488
rect 4982 1476 4988 1488
rect 1084 1448 4988 1476
rect 1084 1436 1090 1448
rect 4982 1436 4988 1448
rect 5040 1436 5046 1488
rect 5074 1436 5080 1488
rect 5132 1476 5138 1488
rect 6012 1476 6040 1516
rect 7466 1504 7472 1516
rect 7524 1504 7530 1556
rect 8113 1547 8171 1553
rect 8113 1513 8125 1547
rect 8159 1544 8171 1547
rect 8159 1516 16574 1544
rect 8159 1513 8171 1516
rect 8113 1507 8171 1513
rect 16546 1488 16574 1516
rect 9217 1479 9275 1485
rect 9217 1476 9229 1479
rect 5132 1448 6040 1476
rect 6104 1448 9229 1476
rect 5132 1436 5138 1448
rect 3050 1368 3056 1420
rect 3108 1408 3114 1420
rect 3881 1411 3939 1417
rect 3881 1408 3893 1411
rect 3108 1380 3893 1408
rect 3108 1368 3114 1380
rect 3881 1377 3893 1380
rect 3927 1408 3939 1411
rect 4246 1408 4252 1420
rect 3927 1380 4252 1408
rect 3927 1377 3939 1380
rect 3881 1371 3939 1377
rect 4246 1368 4252 1380
rect 4304 1368 4310 1420
rect 6104 1417 6132 1448
rect 9217 1445 9229 1448
rect 9263 1445 9275 1479
rect 9398 1476 9404 1488
rect 9359 1448 9404 1476
rect 9217 1439 9275 1445
rect 9398 1436 9404 1448
rect 9456 1436 9462 1488
rect 9677 1479 9735 1485
rect 9677 1445 9689 1479
rect 9723 1445 9735 1479
rect 16546 1448 16580 1488
rect 9677 1439 9735 1445
rect 6089 1411 6147 1417
rect 6089 1377 6101 1411
rect 6135 1377 6147 1411
rect 6270 1408 6276 1420
rect 6231 1380 6276 1408
rect 6089 1371 6147 1377
rect 6270 1368 6276 1380
rect 6328 1368 6334 1420
rect 8570 1408 8576 1420
rect 8531 1380 8576 1408
rect 8570 1368 8576 1380
rect 8628 1368 8634 1420
rect 9692 1408 9720 1439
rect 16574 1436 16580 1448
rect 16632 1436 16638 1488
rect 8680 1380 9720 1408
rect 9861 1411 9919 1417
rect 2498 1300 2504 1352
rect 2556 1340 2562 1352
rect 3329 1343 3387 1349
rect 3329 1340 3341 1343
rect 2556 1312 3341 1340
rect 2556 1300 2562 1312
rect 3329 1309 3341 1312
rect 3375 1309 3387 1343
rect 3329 1303 3387 1309
rect 5994 1300 6000 1352
rect 6052 1340 6058 1352
rect 8680 1340 8708 1380
rect 9861 1377 9873 1411
rect 9907 1377 9919 1411
rect 9861 1371 9919 1377
rect 6052 1312 8708 1340
rect 8757 1343 8815 1349
rect 6052 1300 6058 1312
rect 8757 1309 8769 1343
rect 8803 1340 8815 1343
rect 9122 1340 9128 1352
rect 8803 1312 9128 1340
rect 8803 1309 8815 1312
rect 8757 1303 8815 1309
rect 9122 1300 9128 1312
rect 9180 1300 9186 1352
rect 9674 1340 9680 1352
rect 9416 1312 9680 1340
rect 9416 1272 9444 1312
rect 9674 1300 9680 1312
rect 9732 1340 9738 1352
rect 9876 1340 9904 1371
rect 9732 1312 9904 1340
rect 9732 1300 9738 1312
rect 8864 1244 9444 1272
rect 9585 1275 9643 1281
rect 1486 1164 1492 1216
rect 1544 1204 1550 1216
rect 2682 1204 2688 1216
rect 1544 1176 2688 1204
rect 1544 1164 1550 1176
rect 2682 1164 2688 1176
rect 2740 1164 2746 1216
rect 3326 1164 3332 1216
rect 3384 1204 3390 1216
rect 8864 1213 8892 1244
rect 9585 1241 9597 1275
rect 9631 1272 9643 1275
rect 9858 1272 9864 1284
rect 9631 1244 9864 1272
rect 9631 1241 9643 1244
rect 9585 1235 9643 1241
rect 9858 1232 9864 1244
rect 9916 1232 9922 1284
rect 16574 1272 16580 1284
rect 12406 1244 16580 1272
rect 3513 1207 3571 1213
rect 3513 1204 3525 1207
rect 3384 1176 3525 1204
rect 3384 1164 3390 1176
rect 3513 1173 3525 1176
rect 3559 1204 3571 1207
rect 8297 1207 8355 1213
rect 8297 1204 8309 1207
rect 3559 1176 8309 1204
rect 3559 1173 3571 1176
rect 3513 1167 3571 1173
rect 8297 1173 8309 1176
rect 8343 1204 8355 1207
rect 8849 1207 8907 1213
rect 8849 1204 8861 1207
rect 8343 1176 8861 1204
rect 8343 1173 8355 1176
rect 8297 1167 8355 1173
rect 8849 1173 8861 1176
rect 8895 1173 8907 1207
rect 9030 1204 9036 1216
rect 8991 1176 9036 1204
rect 8849 1167 8907 1173
rect 9030 1164 9036 1176
rect 9088 1164 9094 1216
rect 9122 1164 9128 1216
rect 9180 1204 9186 1216
rect 12406 1204 12434 1244
rect 16574 1232 16580 1244
rect 16632 1232 16638 1284
rect 9180 1176 12434 1204
rect 9180 1164 9186 1176
rect 920 1114 10396 1136
rect 920 1062 2566 1114
rect 2618 1062 2630 1114
rect 2682 1062 2694 1114
rect 2746 1062 2758 1114
rect 2810 1062 2822 1114
rect 2874 1062 7566 1114
rect 7618 1062 7630 1114
rect 7682 1062 7694 1114
rect 7746 1062 7758 1114
rect 7810 1062 7822 1114
rect 7874 1062 10396 1114
rect 920 1040 10396 1062
rect 1486 1000 1492 1012
rect 1447 972 1492 1000
rect 1486 960 1492 972
rect 1544 960 1550 1012
rect 2501 1003 2559 1009
rect 2501 969 2513 1003
rect 2547 1000 2559 1003
rect 2869 1003 2927 1009
rect 2547 972 2774 1000
rect 2547 969 2559 972
rect 2501 963 2559 969
rect 1118 892 1124 944
rect 1176 932 1182 944
rect 1673 935 1731 941
rect 1673 932 1685 935
rect 1176 904 1685 932
rect 1176 892 1182 904
rect 1673 901 1685 904
rect 1719 901 1731 935
rect 1673 895 1731 901
rect 2317 935 2375 941
rect 2317 901 2329 935
rect 2363 932 2375 935
rect 2406 932 2412 944
rect 2363 904 2412 932
rect 2363 901 2375 904
rect 2317 895 2375 901
rect 2406 892 2412 904
rect 2464 892 2470 944
rect 2746 932 2774 972
rect 2869 969 2881 1003
rect 2915 1000 2927 1003
rect 2958 1000 2964 1012
rect 2915 972 2964 1000
rect 2915 969 2927 972
rect 2869 963 2927 969
rect 2958 960 2964 972
rect 3016 960 3022 1012
rect 3050 960 3056 1012
rect 3108 1000 3114 1012
rect 3234 1000 3240 1012
rect 3108 972 3153 1000
rect 3195 972 3240 1000
rect 3108 960 3114 972
rect 3234 960 3240 972
rect 3292 960 3298 1012
rect 3694 1000 3700 1012
rect 3655 972 3700 1000
rect 3694 960 3700 972
rect 3752 960 3758 1012
rect 3973 1003 4031 1009
rect 3973 969 3985 1003
rect 4019 1000 4031 1003
rect 4154 1000 4160 1012
rect 4019 972 4160 1000
rect 4019 969 4031 972
rect 3973 963 4031 969
rect 4154 960 4160 972
rect 4212 960 4218 1012
rect 5074 1000 5080 1012
rect 5035 972 5080 1000
rect 5074 960 5080 972
rect 5132 960 5138 1012
rect 5810 960 5816 1012
rect 5868 1000 5874 1012
rect 9217 1003 9275 1009
rect 9217 1000 9229 1003
rect 5868 972 9229 1000
rect 5868 960 5874 972
rect 9217 969 9229 972
rect 9263 1000 9275 1003
rect 9263 972 9444 1000
rect 9263 969 9275 972
rect 9217 963 9275 969
rect 3326 932 3332 944
rect 2746 904 3332 932
rect 3326 892 3332 904
rect 3384 892 3390 944
rect 3421 935 3479 941
rect 3421 901 3433 935
rect 3467 932 3479 935
rect 4522 932 4528 944
rect 3467 904 4528 932
rect 3467 901 3479 904
rect 3421 895 3479 901
rect 4522 892 4528 904
rect 4580 892 4586 944
rect 5644 904 5948 932
rect 5644 864 5672 904
rect 1412 836 5672 864
rect 1412 805 1440 836
rect 1397 799 1455 805
rect 1397 765 1409 799
rect 1443 765 1455 799
rect 1397 759 1455 765
rect 1857 799 1915 805
rect 1857 765 1869 799
rect 1903 796 1915 799
rect 2314 796 2320 808
rect 1903 768 2320 796
rect 1903 765 1915 768
rect 1857 759 1915 765
rect 2314 756 2320 768
rect 2372 756 2378 808
rect 2590 796 2596 808
rect 2551 768 2596 796
rect 2590 756 2596 768
rect 2648 756 2654 808
rect 2133 731 2191 737
rect 2133 697 2145 731
rect 2179 728 2191 731
rect 5810 728 5816 740
rect 2179 700 5816 728
rect 2179 697 2191 700
rect 2133 691 2191 697
rect 5810 688 5816 700
rect 5868 688 5874 740
rect 5920 728 5948 904
rect 6086 892 6092 944
rect 6144 932 6150 944
rect 6181 935 6239 941
rect 6181 932 6193 935
rect 6144 904 6193 932
rect 6144 892 6150 904
rect 6181 901 6193 904
rect 6227 901 6239 935
rect 6181 895 6239 901
rect 7653 935 7711 941
rect 7653 901 7665 935
rect 7699 932 7711 935
rect 9122 932 9128 944
rect 7699 904 9128 932
rect 7699 901 7711 904
rect 7653 895 7711 901
rect 9122 892 9128 904
rect 9180 892 9186 944
rect 9416 932 9444 972
rect 9490 960 9496 1012
rect 9548 1000 9554 1012
rect 9677 1003 9735 1009
rect 9677 1000 9689 1003
rect 9548 972 9689 1000
rect 9548 960 9554 972
rect 9677 969 9689 972
rect 9723 969 9735 1003
rect 17218 1000 17224 1012
rect 9677 963 9735 969
rect 12406 972 17224 1000
rect 12406 932 12434 972
rect 17218 960 17224 972
rect 17276 960 17282 1012
rect 9416 904 12434 932
rect 9030 864 9036 876
rect 6012 836 9036 864
rect 6012 805 6040 836
rect 9030 824 9036 836
rect 9088 824 9094 876
rect 5997 799 6055 805
rect 5997 765 6009 799
rect 6043 765 6055 799
rect 5997 759 6055 765
rect 8573 799 8631 805
rect 8573 765 8585 799
rect 8619 796 8631 799
rect 8662 796 8668 808
rect 8619 768 8668 796
rect 8619 765 8631 768
rect 8573 759 8631 765
rect 8662 756 8668 768
rect 8720 756 8726 808
rect 8754 756 8760 808
rect 8812 796 8818 808
rect 9585 799 9643 805
rect 8812 768 8857 796
rect 8812 756 8818 768
rect 9585 765 9597 799
rect 9631 796 9643 799
rect 9674 796 9680 808
rect 9631 768 9680 796
rect 9631 765 9643 768
rect 9585 759 9643 765
rect 9674 756 9680 768
rect 9732 756 9738 808
rect 9861 731 9919 737
rect 9861 728 9873 731
rect 5920 700 9873 728
rect 9861 697 9873 700
rect 9907 728 9919 731
rect 20714 728 20720 740
rect 9907 700 20720 728
rect 9907 697 9919 700
rect 9861 691 9919 697
rect 20714 688 20720 700
rect 20772 688 20778 740
rect 3326 620 3332 672
rect 3384 660 3390 672
rect 6365 663 6423 669
rect 6365 660 6377 663
rect 3384 632 6377 660
rect 3384 620 3390 632
rect 6365 629 6377 632
rect 6411 660 6423 663
rect 8110 660 8116 672
rect 6411 632 8116 660
rect 6411 629 6423 632
rect 6365 623 6423 629
rect 8110 620 8116 632
rect 8168 660 8174 672
rect 9033 663 9091 669
rect 9033 660 9045 663
rect 8168 632 9045 660
rect 8168 620 8174 632
rect 9033 629 9045 632
rect 9079 629 9091 663
rect 9033 623 9091 629
rect 920 570 10396 592
rect 920 518 5066 570
rect 5118 518 5130 570
rect 5182 518 5194 570
rect 5246 518 5258 570
rect 5310 518 5322 570
rect 5374 518 10396 570
rect 920 496 10396 518
<< via1 >>
rect 1032 12384 1084 12436
rect 8760 12384 8812 12436
rect 2412 12180 2464 12232
rect 6184 12180 6236 12232
rect 3700 12112 3752 12164
rect 7104 12112 7156 12164
rect 5908 12044 5960 12096
rect 10508 12044 10560 12096
rect 2566 11942 2618 11994
rect 2630 11942 2682 11994
rect 2694 11942 2746 11994
rect 2758 11942 2810 11994
rect 2822 11942 2874 11994
rect 7566 11942 7618 11994
rect 7630 11942 7682 11994
rect 7694 11942 7746 11994
rect 7758 11942 7810 11994
rect 7822 11942 7874 11994
rect 9312 11840 9364 11892
rect 5448 11772 5500 11824
rect 5540 11772 5592 11824
rect 7932 11747 7984 11756
rect 1676 11679 1728 11688
rect 1676 11645 1685 11679
rect 1685 11645 1719 11679
rect 1719 11645 1728 11679
rect 1676 11636 1728 11645
rect 3516 11636 3568 11688
rect 1216 11611 1268 11620
rect 1216 11577 1225 11611
rect 1225 11577 1259 11611
rect 1259 11577 1268 11611
rect 1216 11568 1268 11577
rect 1952 11611 2004 11620
rect 1952 11577 1961 11611
rect 1961 11577 1995 11611
rect 1995 11577 2004 11611
rect 1952 11568 2004 11577
rect 2412 11568 2464 11620
rect 3700 11636 3752 11688
rect 4068 11636 4120 11688
rect 5908 11679 5960 11688
rect 1584 11500 1636 11552
rect 3884 11568 3936 11620
rect 4896 11568 4948 11620
rect 4160 11500 4212 11552
rect 5448 11500 5500 11552
rect 5908 11645 5917 11679
rect 5917 11645 5951 11679
rect 5951 11645 5960 11679
rect 5908 11636 5960 11645
rect 6184 11679 6236 11688
rect 6184 11645 6193 11679
rect 6193 11645 6227 11679
rect 6227 11645 6236 11679
rect 6368 11679 6420 11688
rect 6184 11636 6236 11645
rect 6368 11645 6381 11679
rect 6381 11645 6420 11679
rect 6368 11636 6420 11645
rect 7932 11713 7941 11747
rect 7941 11713 7975 11747
rect 7975 11713 7984 11747
rect 7932 11704 7984 11713
rect 8760 11747 8812 11756
rect 8484 11679 8536 11688
rect 8484 11645 8493 11679
rect 8493 11645 8527 11679
rect 8527 11645 8536 11679
rect 8484 11636 8536 11645
rect 8760 11713 8769 11747
rect 8769 11713 8803 11747
rect 8803 11713 8812 11747
rect 8760 11704 8812 11713
rect 9956 11704 10008 11756
rect 9864 11679 9916 11688
rect 8116 11568 8168 11620
rect 9864 11645 9873 11679
rect 9873 11645 9907 11679
rect 9907 11645 9916 11679
rect 9864 11636 9916 11645
rect 10232 11636 10284 11688
rect 9772 11568 9824 11620
rect 6460 11500 6512 11552
rect 6920 11500 6972 11552
rect 7012 11500 7064 11552
rect 9036 11500 9088 11552
rect 9220 11543 9272 11552
rect 9220 11509 9229 11543
rect 9229 11509 9263 11543
rect 9263 11509 9272 11543
rect 9220 11500 9272 11509
rect 5066 11398 5118 11450
rect 5130 11398 5182 11450
rect 5194 11398 5246 11450
rect 5258 11398 5310 11450
rect 5322 11398 5374 11450
rect 1584 11339 1636 11348
rect 1584 11305 1593 11339
rect 1593 11305 1627 11339
rect 1627 11305 1636 11339
rect 1584 11296 1636 11305
rect 4252 11228 4304 11280
rect 7012 11228 7064 11280
rect 7104 11228 7156 11280
rect 9220 11228 9272 11280
rect 1216 11203 1268 11212
rect 1216 11169 1225 11203
rect 1225 11169 1259 11203
rect 1259 11169 1268 11203
rect 1216 11160 1268 11169
rect 1032 11092 1084 11144
rect 1768 11160 1820 11212
rect 2412 11160 2464 11212
rect 3792 11092 3844 11144
rect 4896 11160 4948 11212
rect 6828 11160 6880 11212
rect 4528 11092 4580 11144
rect 6184 11135 6236 11144
rect 6184 11101 6193 11135
rect 6193 11101 6227 11135
rect 6227 11101 6236 11135
rect 6184 11092 6236 11101
rect 6460 11092 6512 11144
rect 7104 11135 7156 11144
rect 7104 11101 7113 11135
rect 7113 11101 7147 11135
rect 7147 11101 7156 11135
rect 7104 11092 7156 11101
rect 9128 11160 9180 11212
rect 8392 11092 8444 11144
rect 1492 10956 1544 11008
rect 3516 10956 3568 11008
rect 5724 11024 5776 11076
rect 10416 11024 10468 11076
rect 16580 11024 16632 11076
rect 4436 10956 4488 11008
rect 4528 10956 4580 11008
rect 4804 10956 4856 11008
rect 7196 10956 7248 11008
rect 2566 10854 2618 10906
rect 2630 10854 2682 10906
rect 2694 10854 2746 10906
rect 2758 10854 2810 10906
rect 2822 10854 2874 10906
rect 7566 10854 7618 10906
rect 7630 10854 7682 10906
rect 7694 10854 7746 10906
rect 7758 10854 7810 10906
rect 7822 10854 7874 10906
rect 4252 10752 4304 10804
rect 4712 10752 4764 10804
rect 5908 10752 5960 10804
rect 6184 10752 6236 10804
rect 6460 10752 6512 10804
rect 9956 10795 10008 10804
rect 9956 10761 9965 10795
rect 9965 10761 9999 10795
rect 9999 10761 10008 10795
rect 9956 10752 10008 10761
rect 7380 10684 7432 10736
rect 6736 10616 6788 10668
rect 9312 10659 9364 10668
rect 9312 10625 9321 10659
rect 9321 10625 9355 10659
rect 9355 10625 9364 10659
rect 9312 10616 9364 10625
rect 1216 10591 1268 10600
rect 1216 10557 1225 10591
rect 1225 10557 1259 10591
rect 1259 10557 1268 10591
rect 1216 10548 1268 10557
rect 1492 10548 1544 10600
rect 1676 10591 1728 10600
rect 1676 10557 1685 10591
rect 1685 10557 1719 10591
rect 1719 10557 1728 10591
rect 1676 10548 1728 10557
rect 2044 10480 2096 10532
rect 1492 10412 1544 10464
rect 2964 10412 3016 10464
rect 3700 10548 3752 10600
rect 3424 10480 3476 10532
rect 4068 10548 4120 10600
rect 5632 10548 5684 10600
rect 6092 10591 6144 10600
rect 6092 10557 6101 10591
rect 6101 10557 6135 10591
rect 6135 10557 6144 10591
rect 6092 10548 6144 10557
rect 6460 10591 6512 10600
rect 6460 10557 6469 10591
rect 6469 10557 6503 10591
rect 6503 10557 6512 10591
rect 6460 10548 6512 10557
rect 4068 10412 4120 10464
rect 4712 10412 4764 10464
rect 6920 10480 6972 10532
rect 9220 10548 9272 10600
rect 9956 10548 10008 10600
rect 7380 10412 7432 10464
rect 7472 10412 7524 10464
rect 9956 10412 10008 10464
rect 5066 10310 5118 10362
rect 5130 10310 5182 10362
rect 5194 10310 5246 10362
rect 5258 10310 5310 10362
rect 5322 10310 5374 10362
rect 2228 10208 2280 10260
rect 1216 10140 1268 10192
rect 2964 10208 3016 10260
rect 4160 10140 4212 10192
rect 1492 10072 1544 10124
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 1952 10047 2004 10056
rect 1952 10013 1961 10047
rect 1961 10013 1995 10047
rect 1995 10013 2004 10047
rect 1952 10004 2004 10013
rect 3884 10047 3936 10056
rect 2136 9868 2188 9920
rect 2320 9868 2372 9920
rect 3240 9868 3292 9920
rect 3884 10013 3893 10047
rect 3893 10013 3927 10047
rect 3927 10013 3936 10047
rect 3884 10004 3936 10013
rect 9680 10208 9732 10260
rect 9772 10208 9824 10260
rect 4528 10004 4580 10056
rect 6368 10072 6420 10124
rect 5540 10004 5592 10056
rect 6920 10004 6972 10056
rect 7196 10072 7248 10124
rect 7288 10004 7340 10056
rect 8024 10004 8076 10056
rect 9956 10115 10008 10124
rect 9956 10081 9965 10115
rect 9965 10081 9999 10115
rect 9999 10081 10008 10115
rect 9956 10072 10008 10081
rect 10784 10072 10836 10124
rect 10232 10004 10284 10056
rect 6552 9936 6604 9988
rect 7104 9936 7156 9988
rect 4252 9868 4304 9920
rect 4528 9868 4580 9920
rect 6184 9868 6236 9920
rect 9772 9936 9824 9988
rect 10140 9868 10192 9920
rect 2566 9766 2618 9818
rect 2630 9766 2682 9818
rect 2694 9766 2746 9818
rect 2758 9766 2810 9818
rect 2822 9766 2874 9818
rect 7566 9766 7618 9818
rect 7630 9766 7682 9818
rect 7694 9766 7746 9818
rect 7758 9766 7810 9818
rect 7822 9766 7874 9818
rect 1952 9664 2004 9716
rect 6552 9664 6604 9716
rect 1676 9460 1728 9512
rect 1860 9528 1912 9580
rect 5448 9596 5500 9648
rect 9680 9639 9732 9648
rect 2136 9528 2188 9580
rect 3700 9528 3752 9580
rect 6368 9528 6420 9580
rect 8484 9528 8536 9580
rect 9312 9528 9364 9580
rect 9680 9605 9689 9639
rect 9689 9605 9723 9639
rect 9723 9605 9732 9639
rect 9680 9596 9732 9605
rect 16856 9596 16908 9648
rect 1584 9324 1636 9376
rect 1768 9324 1820 9376
rect 3516 9460 3568 9512
rect 3884 9503 3936 9512
rect 3884 9469 3893 9503
rect 3893 9469 3927 9503
rect 3927 9469 3936 9503
rect 3884 9460 3936 9469
rect 5724 9503 5776 9512
rect 5724 9469 5733 9503
rect 5733 9469 5767 9503
rect 5767 9469 5776 9503
rect 5724 9460 5776 9469
rect 6552 9503 6604 9512
rect 6552 9469 6561 9503
rect 6561 9469 6595 9503
rect 6595 9469 6604 9503
rect 6552 9460 6604 9469
rect 8852 9460 8904 9512
rect 9128 9503 9180 9512
rect 9128 9469 9137 9503
rect 9137 9469 9171 9503
rect 9171 9469 9180 9503
rect 9128 9460 9180 9469
rect 9864 9503 9916 9512
rect 9864 9469 9873 9503
rect 9873 9469 9907 9503
rect 9907 9469 9916 9503
rect 9864 9460 9916 9469
rect 2872 9392 2924 9444
rect 3148 9435 3200 9444
rect 3148 9401 3157 9435
rect 3157 9401 3191 9435
rect 3191 9401 3200 9435
rect 3148 9392 3200 9401
rect 3792 9392 3844 9444
rect 4712 9392 4764 9444
rect 8208 9392 8260 9444
rect 2320 9324 2372 9376
rect 5448 9324 5500 9376
rect 5724 9324 5776 9376
rect 8300 9324 8352 9376
rect 8760 9367 8812 9376
rect 8760 9333 8769 9367
rect 8769 9333 8803 9367
rect 8803 9333 8812 9367
rect 8760 9324 8812 9333
rect 8852 9324 8904 9376
rect 9312 9324 9364 9376
rect 10600 9324 10652 9376
rect 5066 9222 5118 9274
rect 5130 9222 5182 9274
rect 5194 9222 5246 9274
rect 5258 9222 5310 9274
rect 5322 9222 5374 9274
rect 6552 9120 6604 9172
rect 8944 9120 8996 9172
rect 19800 9392 19852 9444
rect 2044 9052 2096 9104
rect 3700 9052 3752 9104
rect 3884 9052 3936 9104
rect 5540 9052 5592 9104
rect 6184 9052 6236 9104
rect 2964 8984 3016 9036
rect 3332 8984 3384 9036
rect 3792 8984 3844 9036
rect 3976 9027 4028 9036
rect 3976 8993 3985 9027
rect 3985 8993 4019 9027
rect 4019 8993 4028 9027
rect 3976 8984 4028 8993
rect 1584 8959 1636 8968
rect 1584 8925 1593 8959
rect 1593 8925 1627 8959
rect 1627 8925 1636 8959
rect 1584 8916 1636 8925
rect 1768 8916 1820 8968
rect 6552 8984 6604 9036
rect 6736 9027 6788 9036
rect 6736 8993 6745 9027
rect 6745 8993 6779 9027
rect 6779 8993 6788 9027
rect 6736 8984 6788 8993
rect 8484 9052 8536 9104
rect 8760 9052 8812 9104
rect 8208 9027 8260 9036
rect 4252 8916 4304 8968
rect 4712 8916 4764 8968
rect 6184 8916 6236 8968
rect 3792 8848 3844 8900
rect 6644 8916 6696 8968
rect 8208 8993 8217 9027
rect 8217 8993 8251 9027
rect 8251 8993 8260 9027
rect 8208 8984 8260 8993
rect 9772 8984 9824 9036
rect 10324 8984 10376 9036
rect 7288 8959 7340 8968
rect 7288 8925 7297 8959
rect 7297 8925 7331 8959
rect 7331 8925 7340 8959
rect 7288 8916 7340 8925
rect 10048 8959 10100 8968
rect 10048 8925 10057 8959
rect 10057 8925 10091 8959
rect 10091 8925 10100 8959
rect 10048 8916 10100 8925
rect 3332 8780 3384 8832
rect 3884 8780 3936 8832
rect 6736 8780 6788 8832
rect 7012 8780 7064 8832
rect 16672 8780 16724 8832
rect 2566 8678 2618 8730
rect 2630 8678 2682 8730
rect 2694 8678 2746 8730
rect 2758 8678 2810 8730
rect 2822 8678 2874 8730
rect 7566 8678 7618 8730
rect 7630 8678 7682 8730
rect 7694 8678 7746 8730
rect 7758 8678 7810 8730
rect 7822 8678 7874 8730
rect 1768 8576 1820 8628
rect 3148 8576 3200 8628
rect 5356 8576 5408 8628
rect 3240 8508 3292 8560
rect 3976 8440 4028 8492
rect 8484 8508 8536 8560
rect 1124 8372 1176 8424
rect 3148 8372 3200 8424
rect 6000 8440 6052 8492
rect 8668 8440 8720 8492
rect 3240 8304 3292 8356
rect 4252 8304 4304 8356
rect 6184 8372 6236 8424
rect 8576 8415 8628 8424
rect 8576 8381 8585 8415
rect 8585 8381 8619 8415
rect 8619 8381 8628 8415
rect 8576 8372 8628 8381
rect 9128 8508 9180 8560
rect 9496 8508 9548 8560
rect 9680 8508 9732 8560
rect 9220 8415 9272 8424
rect 4896 8304 4948 8356
rect 6644 8304 6696 8356
rect 9220 8381 9229 8415
rect 9229 8381 9263 8415
rect 9263 8381 9272 8415
rect 9220 8372 9272 8381
rect 9312 8415 9364 8424
rect 9312 8381 9322 8415
rect 9322 8381 9356 8415
rect 9356 8381 9364 8415
rect 9312 8372 9364 8381
rect 9680 8415 9732 8424
rect 9680 8381 9689 8415
rect 9689 8381 9723 8415
rect 9723 8381 9732 8415
rect 9680 8372 9732 8381
rect 9956 8372 10008 8424
rect 9128 8347 9180 8356
rect 9128 8313 9137 8347
rect 9137 8313 9171 8347
rect 9171 8313 9180 8347
rect 9128 8304 9180 8313
rect 9588 8347 9640 8356
rect 9588 8313 9597 8347
rect 9597 8313 9631 8347
rect 9631 8313 9640 8347
rect 9588 8304 9640 8313
rect 9772 8304 9824 8356
rect 11244 8372 11296 8424
rect 19616 8372 19668 8424
rect 16764 8304 16816 8356
rect 5724 8236 5776 8288
rect 5908 8236 5960 8288
rect 6552 8236 6604 8288
rect 12348 8236 12400 8288
rect 5066 8134 5118 8186
rect 5130 8134 5182 8186
rect 5194 8134 5246 8186
rect 5258 8134 5310 8186
rect 5322 8134 5374 8186
rect 3424 8032 3476 8084
rect 6828 8075 6880 8084
rect 6828 8041 6837 8075
rect 6837 8041 6871 8075
rect 6871 8041 6880 8075
rect 6828 8032 6880 8041
rect 7288 8032 7340 8084
rect 1768 7964 1820 8016
rect 2412 7964 2464 8016
rect 3516 7964 3568 8016
rect 4252 7964 4304 8016
rect 7932 8032 7984 8084
rect 16948 8032 17000 8084
rect 3424 7896 3476 7948
rect 3700 7896 3752 7948
rect 3884 7939 3936 7948
rect 3884 7905 3893 7939
rect 3893 7905 3927 7939
rect 3927 7905 3936 7939
rect 3884 7896 3936 7905
rect 4896 7896 4948 7948
rect 5448 7896 5500 7948
rect 7104 7896 7156 7948
rect 9128 7896 9180 7948
rect 3516 7871 3568 7880
rect 3516 7837 3525 7871
rect 3525 7837 3559 7871
rect 3559 7837 3568 7871
rect 3516 7828 3568 7837
rect 6368 7828 6420 7880
rect 12348 7896 12400 7948
rect 14096 7896 14148 7948
rect 9496 7871 9548 7880
rect 9496 7837 9505 7871
rect 9505 7837 9539 7871
rect 9539 7837 9548 7871
rect 9496 7828 9548 7837
rect 1492 7692 1544 7744
rect 3240 7692 3292 7744
rect 5908 7735 5960 7744
rect 5908 7701 5925 7735
rect 5925 7701 5959 7735
rect 5959 7701 5960 7735
rect 5908 7692 5960 7701
rect 6276 7692 6328 7744
rect 6828 7692 6880 7744
rect 7288 7692 7340 7744
rect 9588 7760 9640 7812
rect 8760 7692 8812 7744
rect 9956 7735 10008 7744
rect 9956 7701 9965 7735
rect 9965 7701 9999 7735
rect 9999 7701 10008 7735
rect 9956 7692 10008 7701
rect 2566 7590 2618 7642
rect 2630 7590 2682 7642
rect 2694 7590 2746 7642
rect 2758 7590 2810 7642
rect 2822 7590 2874 7642
rect 7566 7590 7618 7642
rect 7630 7590 7682 7642
rect 7694 7590 7746 7642
rect 7758 7590 7810 7642
rect 7822 7590 7874 7642
rect 4252 7488 4304 7540
rect 9128 7488 9180 7540
rect 4068 7420 4120 7472
rect 6000 7420 6052 7472
rect 8576 7420 8628 7472
rect 9588 7420 9640 7472
rect 10232 7420 10284 7472
rect 3240 7352 3292 7404
rect 4252 7352 4304 7404
rect 4528 7352 4580 7404
rect 13544 7420 13596 7472
rect 20168 7352 20220 7404
rect 1492 7327 1544 7336
rect 1492 7293 1500 7327
rect 1500 7293 1534 7327
rect 1534 7293 1544 7327
rect 1492 7284 1544 7293
rect 1584 7327 1636 7336
rect 1584 7293 1593 7327
rect 1593 7293 1627 7327
rect 1627 7293 1636 7327
rect 1584 7284 1636 7293
rect 3332 7284 3384 7336
rect 3700 7284 3752 7336
rect 5448 7284 5500 7336
rect 5632 7284 5684 7336
rect 6276 7284 6328 7336
rect 7012 7284 7064 7336
rect 8576 7327 8628 7336
rect 8576 7293 8585 7327
rect 8585 7293 8619 7327
rect 8619 7293 8628 7327
rect 8576 7284 8628 7293
rect 8668 7284 8720 7336
rect 7104 7216 7156 7268
rect 9496 7327 9548 7336
rect 9496 7293 9505 7327
rect 9505 7293 9539 7327
rect 9539 7293 9548 7327
rect 9496 7284 9548 7293
rect 10232 7284 10284 7336
rect 2136 7191 2188 7200
rect 2136 7157 2145 7191
rect 2145 7157 2179 7191
rect 2179 7157 2188 7191
rect 2136 7148 2188 7157
rect 4160 7148 4212 7200
rect 4620 7148 4672 7200
rect 5632 7191 5684 7200
rect 5632 7157 5641 7191
rect 5641 7157 5675 7191
rect 5675 7157 5684 7191
rect 5632 7148 5684 7157
rect 10600 7216 10652 7268
rect 5066 7046 5118 7098
rect 5130 7046 5182 7098
rect 5194 7046 5246 7098
rect 5258 7046 5310 7098
rect 5322 7046 5374 7098
rect 11060 7080 11112 7132
rect 19892 7080 19944 7132
rect 13636 7012 13688 7064
rect 20260 7012 20312 7064
rect 1584 6944 1636 6996
rect 3700 6944 3752 6996
rect 6276 6944 6328 6996
rect 9312 6944 9364 6996
rect 2412 6876 2464 6928
rect 4528 6876 4580 6928
rect 6000 6876 6052 6928
rect 1676 6851 1728 6860
rect 1676 6817 1685 6851
rect 1685 6817 1719 6851
rect 1719 6817 1728 6851
rect 1676 6808 1728 6817
rect 3424 6851 3476 6860
rect 3424 6817 3433 6851
rect 3433 6817 3467 6851
rect 3467 6817 3476 6851
rect 3424 6808 3476 6817
rect 3884 6783 3936 6792
rect 3884 6749 3893 6783
rect 3893 6749 3927 6783
rect 3927 6749 3936 6783
rect 3884 6740 3936 6749
rect 4896 6808 4948 6860
rect 4160 6740 4212 6792
rect 6184 6783 6236 6792
rect 6184 6749 6193 6783
rect 6193 6749 6227 6783
rect 6227 6749 6236 6783
rect 6184 6740 6236 6749
rect 8116 6876 8168 6928
rect 9220 6876 9272 6928
rect 10232 6876 10284 6928
rect 7104 6851 7156 6860
rect 7104 6817 7113 6851
rect 7113 6817 7147 6851
rect 7147 6817 7156 6851
rect 7104 6808 7156 6817
rect 7380 6808 7432 6860
rect 9772 6808 9824 6860
rect 7196 6740 7248 6792
rect 9496 6740 9548 6792
rect 10232 6740 10284 6792
rect 19340 6808 19392 6860
rect 2044 6604 2096 6656
rect 6276 6604 6328 6656
rect 8576 6604 8628 6656
rect 2566 6502 2618 6554
rect 2630 6502 2682 6554
rect 2694 6502 2746 6554
rect 2758 6502 2810 6554
rect 2822 6502 2874 6554
rect 7566 6502 7618 6554
rect 7630 6502 7682 6554
rect 7694 6502 7746 6554
rect 7758 6502 7810 6554
rect 7822 6502 7874 6554
rect 1676 6400 1728 6452
rect 4252 6400 4304 6452
rect 6184 6400 6236 6452
rect 7840 6332 7892 6384
rect 2964 6264 3016 6316
rect 5816 6307 5868 6316
rect 5816 6273 5825 6307
rect 5825 6273 5859 6307
rect 5859 6273 5868 6307
rect 5816 6264 5868 6273
rect 8668 6264 8720 6316
rect 9036 6332 9088 6384
rect 9956 6307 10008 6316
rect 1584 6196 1636 6248
rect 3608 6239 3660 6248
rect 3608 6205 3617 6239
rect 3617 6205 3651 6239
rect 3651 6205 3660 6239
rect 3608 6196 3660 6205
rect 5724 6196 5776 6248
rect 7288 6239 7340 6248
rect 7288 6205 7297 6239
rect 7297 6205 7331 6239
rect 7331 6205 7340 6239
rect 7288 6196 7340 6205
rect 7748 6196 7800 6248
rect 1492 6103 1544 6112
rect 1492 6069 1501 6103
rect 1501 6069 1535 6103
rect 1535 6069 1544 6103
rect 1492 6060 1544 6069
rect 2964 6128 3016 6180
rect 3976 6128 4028 6180
rect 3424 6103 3476 6112
rect 3424 6069 3433 6103
rect 3433 6069 3467 6103
rect 3467 6069 3476 6103
rect 3424 6060 3476 6069
rect 3700 6060 3752 6112
rect 7012 6128 7064 6180
rect 7840 6103 7892 6112
rect 7840 6069 7857 6103
rect 7857 6069 7891 6103
rect 7891 6069 7892 6103
rect 7840 6060 7892 6069
rect 9404 6196 9456 6248
rect 9956 6273 9965 6307
rect 9965 6273 9999 6307
rect 9999 6273 10008 6307
rect 9956 6264 10008 6273
rect 19708 6264 19760 6316
rect 9220 6128 9272 6180
rect 9588 6128 9640 6180
rect 9404 6060 9456 6112
rect 5066 5958 5118 6010
rect 5130 5958 5182 6010
rect 5194 5958 5246 6010
rect 5258 5958 5310 6010
rect 5322 5958 5374 6010
rect 1400 5899 1452 5908
rect 1400 5865 1409 5899
rect 1409 5865 1443 5899
rect 1443 5865 1452 5899
rect 1400 5856 1452 5865
rect 3884 5856 3936 5908
rect 19432 6060 19484 6112
rect 2964 5788 3016 5840
rect 3332 5788 3384 5840
rect 7288 5788 7340 5840
rect 9864 5788 9916 5840
rect 4068 5720 4120 5772
rect 4896 5720 4948 5772
rect 5356 5720 5408 5772
rect 1676 5695 1728 5704
rect 1676 5661 1685 5695
rect 1685 5661 1719 5695
rect 1719 5661 1728 5695
rect 1676 5652 1728 5661
rect 3700 5652 3752 5704
rect 3976 5695 4028 5704
rect 3976 5661 3985 5695
rect 3985 5661 4019 5695
rect 4019 5661 4028 5695
rect 3976 5652 4028 5661
rect 5080 5652 5132 5704
rect 6000 5695 6052 5704
rect 6000 5661 6009 5695
rect 6009 5661 6043 5695
rect 6043 5661 6052 5695
rect 6000 5652 6052 5661
rect 7104 5720 7156 5772
rect 8760 5720 8812 5772
rect 9036 5720 9088 5772
rect 9496 5720 9548 5772
rect 10416 5720 10468 5772
rect 7288 5652 7340 5704
rect 7380 5652 7432 5704
rect 9404 5695 9456 5704
rect 3056 5584 3108 5636
rect 5356 5584 5408 5636
rect 7748 5584 7800 5636
rect 8668 5584 8720 5636
rect 9404 5661 9413 5695
rect 9413 5661 9447 5695
rect 9447 5661 9456 5695
rect 9404 5652 9456 5661
rect 9588 5652 9640 5704
rect 9772 5652 9824 5704
rect 10140 5652 10192 5704
rect 13820 5652 13872 5704
rect 17040 5652 17092 5704
rect 1676 5516 1728 5568
rect 2136 5516 2188 5568
rect 3332 5516 3384 5568
rect 7288 5516 7340 5568
rect 10232 5584 10284 5636
rect 11152 5584 11204 5636
rect 16672 5584 16724 5636
rect 10140 5516 10192 5568
rect 13452 5516 13504 5568
rect 16948 5516 17000 5568
rect 2566 5414 2618 5466
rect 2630 5414 2682 5466
rect 2694 5414 2746 5466
rect 2758 5414 2810 5466
rect 2822 5414 2874 5466
rect 7566 5414 7618 5466
rect 7630 5414 7682 5466
rect 7694 5414 7746 5466
rect 7758 5414 7810 5466
rect 7822 5414 7874 5466
rect 14096 5380 14148 5432
rect 19524 5380 19576 5432
rect 2044 5312 2096 5364
rect 2780 5312 2832 5364
rect 4528 5312 4580 5364
rect 6644 5312 6696 5364
rect 11244 5312 11296 5364
rect 5632 5244 5684 5296
rect 20076 5312 20128 5364
rect 1768 5176 1820 5228
rect 2504 5176 2556 5228
rect 3608 5176 3660 5228
rect 6000 5176 6052 5228
rect 16580 5176 16632 5228
rect 2964 5108 3016 5160
rect 3700 5108 3752 5160
rect 5908 5108 5960 5160
rect 8300 5151 8352 5160
rect 8300 5117 8309 5151
rect 8309 5117 8343 5151
rect 8343 5117 8352 5151
rect 8300 5108 8352 5117
rect 4528 5040 4580 5092
rect 4896 4972 4948 5024
rect 5080 4972 5132 5024
rect 6552 5040 6604 5092
rect 8576 5040 8628 5092
rect 8760 5040 8812 5092
rect 5632 4972 5684 5024
rect 8300 4972 8352 5024
rect 8852 4972 8904 5024
rect 17316 5040 17368 5092
rect 5066 4870 5118 4922
rect 5130 4870 5182 4922
rect 5194 4870 5246 4922
rect 5258 4870 5310 4922
rect 5322 4870 5374 4922
rect 3884 4768 3936 4820
rect 4160 4811 4212 4820
rect 4160 4777 4169 4811
rect 4169 4777 4203 4811
rect 4203 4777 4212 4811
rect 4160 4768 4212 4777
rect 4252 4768 4304 4820
rect 4528 4768 4580 4820
rect 4988 4768 5040 4820
rect 7012 4768 7064 4820
rect 7380 4768 7432 4820
rect 8116 4811 8168 4820
rect 8116 4777 8125 4811
rect 8125 4777 8159 4811
rect 8159 4777 8168 4811
rect 8116 4768 8168 4777
rect 9404 4768 9456 4820
rect 1308 4700 1360 4752
rect 3608 4700 3660 4752
rect 2228 4632 2280 4684
rect 2872 4632 2924 4684
rect 3424 4675 3476 4684
rect 3424 4641 3433 4675
rect 3433 4641 3467 4675
rect 3467 4641 3476 4675
rect 3424 4632 3476 4641
rect 5356 4700 5408 4752
rect 6000 4700 6052 4752
rect 4620 4632 4672 4684
rect 6552 4632 6604 4684
rect 7104 4675 7156 4684
rect 7104 4641 7143 4675
rect 7143 4641 7156 4675
rect 7104 4632 7156 4641
rect 7288 4675 7340 4684
rect 7288 4641 7297 4675
rect 7297 4641 7331 4675
rect 7331 4641 7340 4675
rect 7288 4632 7340 4641
rect 4344 4607 4396 4616
rect 4344 4573 4353 4607
rect 4353 4573 4387 4607
rect 4387 4573 4396 4607
rect 4344 4564 4396 4573
rect 4896 4564 4948 4616
rect 8116 4632 8168 4684
rect 9588 4700 9640 4752
rect 2688 4428 2740 4480
rect 8116 4496 8168 4548
rect 6552 4428 6604 4480
rect 10324 4564 10376 4616
rect 8576 4428 8628 4480
rect 9588 4428 9640 4480
rect 7566 4326 7618 4378
rect 7630 4326 7682 4378
rect 7694 4326 7746 4378
rect 7758 4326 7810 4378
rect 7822 4326 7874 4378
rect 5356 4267 5408 4276
rect 5356 4233 5365 4267
rect 5365 4233 5399 4267
rect 5399 4233 5408 4267
rect 5356 4224 5408 4233
rect 5816 4224 5868 4276
rect 6000 4224 6052 4276
rect 3332 4131 3384 4140
rect 3332 4097 3341 4131
rect 3341 4097 3375 4131
rect 3375 4097 3384 4131
rect 3332 4088 3384 4097
rect 3976 4088 4028 4140
rect 4068 4088 4120 4140
rect 6368 4156 6420 4208
rect 8116 4224 8168 4276
rect 8852 4224 8904 4276
rect 9404 4224 9456 4276
rect 16856 4224 16908 4276
rect 8208 4156 8260 4208
rect 5448 4088 5500 4140
rect 6920 4131 6972 4140
rect 5356 4063 5408 4072
rect 5356 4029 5369 4063
rect 5369 4029 5408 4063
rect 5356 4020 5408 4029
rect 5632 4020 5684 4072
rect 6920 4097 6929 4131
rect 6929 4097 6963 4131
rect 6963 4097 6972 4131
rect 6920 4088 6972 4097
rect 7472 4088 7524 4140
rect 13544 4088 13596 4140
rect 17132 4088 17184 4140
rect 3884 3952 3936 4004
rect 4068 3952 4120 4004
rect 2780 3884 2832 3936
rect 3424 3884 3476 3936
rect 3700 3884 3752 3936
rect 5264 3884 5316 3936
rect 5632 3884 5684 3936
rect 6736 3952 6788 4004
rect 8484 3952 8536 4004
rect 9220 3884 9272 3936
rect 9588 3884 9640 3936
rect 5066 3782 5118 3834
rect 5130 3782 5182 3834
rect 5194 3782 5246 3834
rect 5258 3782 5310 3834
rect 5322 3782 5374 3834
rect 3148 3680 3200 3732
rect 3976 3680 4028 3732
rect 3424 3612 3476 3664
rect 4896 3612 4948 3664
rect 6092 3680 6144 3732
rect 7196 3723 7248 3732
rect 7196 3689 7205 3723
rect 7205 3689 7239 3723
rect 7239 3689 7248 3723
rect 7196 3680 7248 3689
rect 9036 3680 9088 3732
rect 7288 3612 7340 3664
rect 5448 3544 5500 3596
rect 3056 3476 3108 3528
rect 3792 3476 3844 3528
rect 4068 3476 4120 3528
rect 5356 3476 5408 3528
rect 5632 3476 5684 3528
rect 4988 3340 5040 3392
rect 8852 3587 8904 3596
rect 8852 3553 8861 3587
rect 8861 3553 8895 3587
rect 8895 3553 8904 3587
rect 8852 3544 8904 3553
rect 9220 3587 9272 3596
rect 9220 3553 9229 3587
rect 9229 3553 9263 3587
rect 9263 3553 9272 3587
rect 10048 3680 10100 3732
rect 9588 3612 9640 3664
rect 9220 3544 9272 3553
rect 9128 3476 9180 3528
rect 9220 3408 9272 3460
rect 22100 3476 22152 3528
rect 10416 3408 10468 3460
rect 10508 3340 10560 3392
rect 7566 3238 7618 3290
rect 7630 3238 7682 3290
rect 7694 3238 7746 3290
rect 7758 3238 7810 3290
rect 7822 3238 7874 3290
rect 3240 3136 3292 3188
rect 4436 3136 4488 3188
rect 5356 3136 5408 3188
rect 9680 3136 9732 3188
rect 11060 3136 11112 3188
rect 6644 3068 6696 3120
rect 4068 3000 4120 3052
rect 11152 3000 11204 3052
rect 5908 2975 5960 2984
rect 5908 2941 5917 2975
rect 5917 2941 5951 2975
rect 5951 2941 5960 2975
rect 5908 2932 5960 2941
rect 8024 2975 8076 2984
rect 8024 2941 8033 2975
rect 8033 2941 8067 2975
rect 8067 2941 8076 2975
rect 8024 2932 8076 2941
rect 8944 2932 8996 2984
rect 4252 2864 4304 2916
rect 4896 2864 4948 2916
rect 6460 2796 6512 2848
rect 5066 2694 5118 2746
rect 5130 2694 5182 2746
rect 5194 2694 5246 2746
rect 5258 2694 5310 2746
rect 5322 2694 5374 2746
rect 3056 2524 3108 2576
rect 3976 2592 4028 2644
rect 4344 2592 4396 2644
rect 5540 2635 5592 2644
rect 5540 2601 5549 2635
rect 5549 2601 5583 2635
rect 5583 2601 5592 2635
rect 5540 2592 5592 2601
rect 5632 2592 5684 2644
rect 5724 2592 5776 2644
rect 8392 2635 8444 2644
rect 8392 2601 8401 2635
rect 8401 2601 8435 2635
rect 8435 2601 8444 2635
rect 8392 2592 8444 2601
rect 8668 2635 8720 2644
rect 8668 2601 8677 2635
rect 8677 2601 8711 2635
rect 8711 2601 8720 2635
rect 8668 2592 8720 2601
rect 9496 2592 9548 2644
rect 9680 2592 9732 2644
rect 10784 2592 10836 2644
rect 3424 2499 3476 2508
rect 3424 2465 3433 2499
rect 3433 2465 3467 2499
rect 3467 2465 3476 2499
rect 3424 2456 3476 2465
rect 3700 2456 3752 2508
rect 6644 2524 6696 2576
rect 7380 2524 7432 2576
rect 4896 2499 4948 2508
rect 2872 2388 2924 2440
rect 4896 2465 4905 2499
rect 4905 2465 4939 2499
rect 4939 2465 4948 2499
rect 4896 2456 4948 2465
rect 5356 2499 5408 2508
rect 5356 2465 5365 2499
rect 5365 2465 5399 2499
rect 5399 2465 5408 2499
rect 5356 2456 5408 2465
rect 6552 2499 6604 2508
rect 6552 2465 6561 2499
rect 6561 2465 6595 2499
rect 6595 2465 6604 2499
rect 6552 2456 6604 2465
rect 8484 2499 8536 2508
rect 8484 2465 8493 2499
rect 8493 2465 8527 2499
rect 8527 2465 8536 2499
rect 8484 2456 8536 2465
rect 8576 2456 8628 2508
rect 8760 2499 8812 2508
rect 8760 2465 8769 2499
rect 8769 2465 8803 2499
rect 8803 2465 8812 2499
rect 8760 2456 8812 2465
rect 9036 2524 9088 2576
rect 5724 2388 5776 2440
rect 16672 2524 16724 2576
rect 6000 2320 6052 2372
rect 13820 2320 13872 2372
rect 3424 2252 3476 2304
rect 3884 2295 3936 2304
rect 3884 2261 3893 2295
rect 3893 2261 3927 2295
rect 3927 2261 3936 2295
rect 3884 2252 3936 2261
rect 4988 2295 5040 2304
rect 4988 2261 4997 2295
rect 4997 2261 5031 2295
rect 5031 2261 5040 2295
rect 4988 2252 5040 2261
rect 5080 2252 5132 2304
rect 6828 2252 6880 2304
rect 8668 2252 8720 2304
rect 7566 2150 7618 2202
rect 7630 2150 7682 2202
rect 7694 2150 7746 2202
rect 7758 2150 7810 2202
rect 7822 2150 7874 2202
rect 2688 2048 2740 2100
rect 4436 2048 4488 2100
rect 4804 2091 4856 2100
rect 4804 2057 4813 2091
rect 4813 2057 4847 2091
rect 4847 2057 4856 2091
rect 4804 2048 4856 2057
rect 5448 2091 5500 2100
rect 5448 2057 5457 2091
rect 5457 2057 5491 2091
rect 5491 2057 5500 2091
rect 5448 2048 5500 2057
rect 5908 2048 5960 2100
rect 6000 2091 6052 2100
rect 6000 2057 6009 2091
rect 6009 2057 6043 2091
rect 6043 2057 6052 2091
rect 6000 2048 6052 2057
rect 3516 1980 3568 2032
rect 4712 1980 4764 2032
rect 6092 1980 6144 2032
rect 7012 1980 7064 2032
rect 7472 2048 7524 2100
rect 16764 2048 16816 2100
rect 20628 1980 20680 2032
rect 3884 1912 3936 1964
rect 7104 1912 7156 1964
rect 13636 1912 13688 1964
rect 2688 1844 2740 1896
rect 4068 1887 4120 1896
rect 4068 1853 4077 1887
rect 4077 1853 4111 1887
rect 4111 1853 4120 1887
rect 4068 1844 4120 1853
rect 4620 1887 4672 1896
rect 4620 1853 4629 1887
rect 4629 1853 4663 1887
rect 4663 1853 4672 1887
rect 4620 1844 4672 1853
rect 5356 1844 5408 1896
rect 7932 1887 7984 1896
rect 7932 1853 7941 1887
rect 7941 1853 7975 1887
rect 7975 1853 7984 1887
rect 7932 1844 7984 1853
rect 9772 1887 9824 1896
rect 9772 1853 9781 1887
rect 9781 1853 9815 1887
rect 9815 1853 9824 1887
rect 9772 1844 9824 1853
rect 3240 1776 3292 1828
rect 3608 1776 3660 1828
rect 5080 1708 5132 1760
rect 7380 1776 7432 1828
rect 8300 1708 8352 1760
rect 13452 1708 13504 1760
rect 5066 1606 5118 1658
rect 5130 1606 5182 1658
rect 5194 1606 5246 1658
rect 5258 1606 5310 1658
rect 5322 1606 5374 1658
rect 20 1504 72 1556
rect 3240 1504 3292 1556
rect 4896 1504 4948 1556
rect 5724 1504 5776 1556
rect 1032 1436 1084 1488
rect 4988 1436 5040 1488
rect 5080 1436 5132 1488
rect 7472 1504 7524 1556
rect 3056 1368 3108 1420
rect 4252 1368 4304 1420
rect 9404 1479 9456 1488
rect 9404 1445 9413 1479
rect 9413 1445 9447 1479
rect 9447 1445 9456 1479
rect 9404 1436 9456 1445
rect 6276 1411 6328 1420
rect 6276 1377 6285 1411
rect 6285 1377 6319 1411
rect 6319 1377 6328 1411
rect 6276 1368 6328 1377
rect 8576 1411 8628 1420
rect 8576 1377 8585 1411
rect 8585 1377 8619 1411
rect 8619 1377 8628 1411
rect 8576 1368 8628 1377
rect 16580 1436 16632 1488
rect 2504 1300 2556 1352
rect 6000 1300 6052 1352
rect 9128 1300 9180 1352
rect 9680 1300 9732 1352
rect 1492 1164 1544 1216
rect 2688 1164 2740 1216
rect 3332 1164 3384 1216
rect 9864 1232 9916 1284
rect 9036 1207 9088 1216
rect 9036 1173 9045 1207
rect 9045 1173 9079 1207
rect 9079 1173 9088 1207
rect 9036 1164 9088 1173
rect 9128 1164 9180 1216
rect 16580 1232 16632 1284
rect 2566 1062 2618 1114
rect 2630 1062 2682 1114
rect 2694 1062 2746 1114
rect 2758 1062 2810 1114
rect 2822 1062 2874 1114
rect 7566 1062 7618 1114
rect 7630 1062 7682 1114
rect 7694 1062 7746 1114
rect 7758 1062 7810 1114
rect 7822 1062 7874 1114
rect 1492 1003 1544 1012
rect 1492 969 1501 1003
rect 1501 969 1535 1003
rect 1535 969 1544 1003
rect 1492 960 1544 969
rect 1124 892 1176 944
rect 2412 892 2464 944
rect 2964 960 3016 1012
rect 3056 1003 3108 1012
rect 3056 969 3065 1003
rect 3065 969 3099 1003
rect 3099 969 3108 1003
rect 3240 1003 3292 1012
rect 3056 960 3108 969
rect 3240 969 3249 1003
rect 3249 969 3283 1003
rect 3283 969 3292 1003
rect 3240 960 3292 969
rect 3700 1003 3752 1012
rect 3700 969 3709 1003
rect 3709 969 3743 1003
rect 3743 969 3752 1003
rect 3700 960 3752 969
rect 4160 960 4212 1012
rect 5080 1003 5132 1012
rect 5080 969 5089 1003
rect 5089 969 5123 1003
rect 5123 969 5132 1003
rect 5080 960 5132 969
rect 5816 960 5868 1012
rect 3332 892 3384 944
rect 4528 892 4580 944
rect 2320 756 2372 808
rect 2596 799 2648 808
rect 2596 765 2605 799
rect 2605 765 2639 799
rect 2639 765 2648 799
rect 2596 756 2648 765
rect 5816 688 5868 740
rect 6092 892 6144 944
rect 9128 892 9180 944
rect 9496 960 9548 1012
rect 17224 960 17276 1012
rect 9036 824 9088 876
rect 8668 756 8720 808
rect 8760 799 8812 808
rect 8760 765 8769 799
rect 8769 765 8803 799
rect 8803 765 8812 799
rect 8760 756 8812 765
rect 9680 756 9732 808
rect 20720 688 20772 740
rect 3332 620 3384 672
rect 8116 620 8168 672
rect 5066 518 5118 570
rect 5130 518 5182 570
rect 5194 518 5246 570
rect 5258 518 5310 570
rect 5322 518 5374 570
<< metal2 >>
rect 938 12322 994 13000
rect 1032 12436 1084 12442
rect 1032 12378 1084 12384
rect 32 12294 994 12322
rect 32 1562 60 12294
rect 938 12200 994 12294
rect 1044 11150 1072 12378
rect 1398 12200 1454 13000
rect 1858 12200 1914 13000
rect 2318 12200 2374 13000
rect 2778 12322 2834 13000
rect 3238 12322 3294 13000
rect 3698 12322 3754 13000
rect 2778 12294 3096 12322
rect 2412 12232 2464 12238
rect 1214 11656 1270 11665
rect 1214 11591 1216 11600
rect 1268 11591 1270 11600
rect 1216 11562 1268 11568
rect 1216 11212 1268 11218
rect 1216 11154 1268 11160
rect 1032 11144 1084 11150
rect 1032 11086 1084 11092
rect 20 1556 72 1562
rect 20 1498 72 1504
rect 1044 1494 1072 11086
rect 1228 10606 1256 11154
rect 1216 10600 1268 10606
rect 1216 10542 1268 10548
rect 1228 10198 1256 10542
rect 1216 10192 1268 10198
rect 1216 10134 1268 10140
rect 1412 9674 1440 12200
rect 1676 11688 1728 11694
rect 1676 11630 1728 11636
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1596 11354 1624 11494
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 1492 11008 1544 11014
rect 1492 10950 1544 10956
rect 1504 10606 1532 10950
rect 1688 10606 1716 11630
rect 1768 11212 1820 11218
rect 1768 11154 1820 11160
rect 1492 10600 1544 10606
rect 1492 10542 1544 10548
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1492 10464 1544 10470
rect 1492 10406 1544 10412
rect 1504 10130 1532 10406
rect 1492 10124 1544 10130
rect 1492 10066 1544 10072
rect 1320 9646 1440 9674
rect 1124 8424 1176 8430
rect 1124 8366 1176 8372
rect 1032 1488 1084 1494
rect 1032 1430 1084 1436
rect 1136 950 1164 8366
rect 1320 4758 1348 9646
rect 1504 7834 1532 10066
rect 1688 10062 1716 10542
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1780 9466 1808 11154
rect 1872 9586 1900 12200
rect 1952 11620 2004 11626
rect 1952 11562 2004 11568
rect 1964 10169 1992 11562
rect 2044 10532 2096 10538
rect 2044 10474 2096 10480
rect 1950 10160 2006 10169
rect 1950 10095 2006 10104
rect 1952 10056 2004 10062
rect 1952 9998 2004 10004
rect 1964 9722 1992 9998
rect 1952 9716 2004 9722
rect 1952 9658 2004 9664
rect 1860 9580 1912 9586
rect 1860 9522 1912 9528
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1596 8974 1624 9318
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 1504 7806 1624 7834
rect 1492 7744 1544 7750
rect 1492 7686 1544 7692
rect 1504 7342 1532 7686
rect 1596 7342 1624 7806
rect 1492 7336 1544 7342
rect 1412 7296 1492 7324
rect 1412 5914 1440 7296
rect 1492 7278 1544 7284
rect 1584 7336 1636 7342
rect 1584 7278 1636 7284
rect 1596 7002 1624 7278
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1688 6866 1716 9454
rect 1780 9438 1992 9466
rect 1768 9376 1820 9382
rect 1820 9336 1900 9364
rect 1768 9318 1820 9324
rect 1768 8968 1820 8974
rect 1768 8910 1820 8916
rect 1780 8634 1808 8910
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1768 8016 1820 8022
rect 1768 7958 1820 7964
rect 1676 6860 1728 6866
rect 1676 6802 1728 6808
rect 1688 6458 1716 6802
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1582 6352 1638 6361
rect 1582 6287 1638 6296
rect 1596 6254 1624 6287
rect 1584 6248 1636 6254
rect 1490 6216 1546 6225
rect 1584 6190 1636 6196
rect 1490 6151 1546 6160
rect 1504 6118 1532 6151
rect 1492 6112 1544 6118
rect 1492 6054 1544 6060
rect 1400 5908 1452 5914
rect 1400 5850 1452 5856
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 1688 5574 1716 5646
rect 1676 5568 1728 5574
rect 1676 5510 1728 5516
rect 1780 5234 1808 7958
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 1308 4752 1360 4758
rect 1308 4694 1360 4700
rect 1872 4593 1900 9336
rect 1964 8616 1992 9438
rect 2056 9110 2084 10474
rect 2332 10418 2360 12200
rect 2778 12200 2834 12294
rect 2412 12174 2464 12180
rect 2424 11626 2452 12174
rect 2566 11996 2874 12005
rect 2566 11994 2572 11996
rect 2628 11994 2652 11996
rect 2708 11994 2732 11996
rect 2788 11994 2812 11996
rect 2868 11994 2874 11996
rect 2628 11942 2630 11994
rect 2810 11942 2812 11994
rect 2566 11940 2572 11942
rect 2628 11940 2652 11942
rect 2708 11940 2732 11942
rect 2788 11940 2812 11942
rect 2868 11940 2874 11942
rect 2566 11931 2874 11940
rect 2412 11620 2464 11626
rect 2412 11562 2464 11568
rect 2424 11218 2452 11562
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 2566 10908 2874 10917
rect 2566 10906 2572 10908
rect 2628 10906 2652 10908
rect 2708 10906 2732 10908
rect 2788 10906 2812 10908
rect 2868 10906 2874 10908
rect 2628 10854 2630 10906
rect 2810 10854 2812 10906
rect 2566 10852 2572 10854
rect 2628 10852 2652 10854
rect 2708 10852 2732 10854
rect 2788 10852 2812 10854
rect 2868 10852 2874 10854
rect 2566 10843 2874 10852
rect 2964 10464 3016 10470
rect 2332 10390 2452 10418
rect 2964 10406 3016 10412
rect 2228 10260 2280 10266
rect 2280 10220 2360 10248
rect 2228 10202 2280 10208
rect 2332 9926 2360 10220
rect 2136 9920 2188 9926
rect 2320 9920 2372 9926
rect 2136 9862 2188 9868
rect 2226 9888 2282 9897
rect 2148 9586 2176 9862
rect 2320 9862 2372 9868
rect 2226 9823 2282 9832
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 2044 9104 2096 9110
rect 2044 9046 2096 9052
rect 1964 8588 2084 8616
rect 2056 6662 2084 8588
rect 2148 7206 2176 9522
rect 2136 7200 2188 7206
rect 2136 7142 2188 7148
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 2056 5370 2084 6598
rect 2148 5574 2176 7142
rect 2136 5568 2188 5574
rect 2136 5510 2188 5516
rect 2044 5364 2096 5370
rect 2044 5306 2096 5312
rect 2240 4690 2268 9823
rect 2320 9376 2372 9382
rect 2320 9318 2372 9324
rect 2228 4684 2280 4690
rect 2228 4626 2280 4632
rect 1858 4584 1914 4593
rect 1858 4519 1914 4528
rect 1492 1216 1544 1222
rect 1492 1158 1544 1164
rect 1504 1018 1532 1158
rect 1492 1012 1544 1018
rect 1492 954 1544 960
rect 1124 944 1176 950
rect 1124 886 1176 892
rect 2332 814 2360 9318
rect 2424 8022 2452 10390
rect 2976 10266 3004 10406
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 2566 9820 2874 9829
rect 2566 9818 2572 9820
rect 2628 9818 2652 9820
rect 2708 9818 2732 9820
rect 2788 9818 2812 9820
rect 2868 9818 2874 9820
rect 2628 9766 2630 9818
rect 2810 9766 2812 9818
rect 2566 9764 2572 9766
rect 2628 9764 2652 9766
rect 2708 9764 2732 9766
rect 2788 9764 2812 9766
rect 2868 9764 2874 9766
rect 2566 9755 2874 9764
rect 2976 9489 3004 10202
rect 2962 9480 3018 9489
rect 2872 9444 2924 9450
rect 2924 9424 2962 9432
rect 2924 9415 3018 9424
rect 2924 9404 3004 9415
rect 2872 9386 2924 9392
rect 2976 9355 3004 9404
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 2566 8732 2874 8741
rect 2566 8730 2572 8732
rect 2628 8730 2652 8732
rect 2708 8730 2732 8732
rect 2788 8730 2812 8732
rect 2868 8730 2874 8732
rect 2628 8678 2630 8730
rect 2810 8678 2812 8730
rect 2566 8676 2572 8678
rect 2628 8676 2652 8678
rect 2708 8676 2732 8678
rect 2788 8676 2812 8678
rect 2868 8676 2874 8678
rect 2566 8667 2874 8676
rect 2412 8016 2464 8022
rect 2412 7958 2464 7964
rect 2566 7644 2874 7653
rect 2566 7642 2572 7644
rect 2628 7642 2652 7644
rect 2708 7642 2732 7644
rect 2788 7642 2812 7644
rect 2868 7642 2874 7644
rect 2628 7590 2630 7642
rect 2810 7590 2812 7642
rect 2566 7588 2572 7590
rect 2628 7588 2652 7590
rect 2708 7588 2732 7590
rect 2788 7588 2812 7590
rect 2868 7588 2874 7590
rect 2566 7579 2874 7588
rect 2412 6928 2464 6934
rect 2412 6870 2464 6876
rect 2424 5352 2452 6870
rect 2566 6556 2874 6565
rect 2566 6554 2572 6556
rect 2628 6554 2652 6556
rect 2708 6554 2732 6556
rect 2788 6554 2812 6556
rect 2868 6554 2874 6556
rect 2628 6502 2630 6554
rect 2810 6502 2812 6554
rect 2566 6500 2572 6502
rect 2628 6500 2652 6502
rect 2708 6500 2732 6502
rect 2788 6500 2812 6502
rect 2868 6500 2874 6502
rect 2566 6491 2874 6500
rect 2976 6322 3004 8978
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 2964 6180 3016 6186
rect 2964 6122 3016 6128
rect 2976 6089 3004 6122
rect 2962 6080 3018 6089
rect 2962 6015 3018 6024
rect 2976 5846 3004 6015
rect 2964 5840 3016 5846
rect 2964 5782 3016 5788
rect 2566 5468 2874 5477
rect 2566 5466 2572 5468
rect 2628 5466 2652 5468
rect 2708 5466 2732 5468
rect 2788 5466 2812 5468
rect 2868 5466 2874 5468
rect 2628 5414 2630 5466
rect 2810 5414 2812 5466
rect 2566 5412 2572 5414
rect 2628 5412 2652 5414
rect 2708 5412 2732 5414
rect 2788 5412 2812 5414
rect 2868 5412 2874 5414
rect 2566 5403 2874 5412
rect 2780 5364 2832 5370
rect 2424 5324 2728 5352
rect 2504 5228 2556 5234
rect 2504 5170 2556 5176
rect 2410 4040 2466 4049
rect 2410 3975 2466 3984
rect 2424 950 2452 3975
rect 2516 1358 2544 5170
rect 2700 4486 2728 5324
rect 2780 5306 2832 5312
rect 2688 4480 2740 4486
rect 2688 4422 2740 4428
rect 2700 2106 2728 4422
rect 2792 3942 2820 5306
rect 2976 5166 3004 5782
rect 3068 5642 3096 12294
rect 3238 12294 3372 12322
rect 3238 12200 3294 12294
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3148 9444 3200 9450
rect 3148 9386 3200 9392
rect 3160 8634 3188 9386
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 3252 8566 3280 9862
rect 3344 9042 3372 12294
rect 3620 12294 3754 12322
rect 3516 11688 3568 11694
rect 3516 11630 3568 11636
rect 3528 11014 3556 11630
rect 3516 11008 3568 11014
rect 3516 10950 3568 10956
rect 3424 10532 3476 10538
rect 3424 10474 3476 10480
rect 3332 9036 3384 9042
rect 3332 8978 3384 8984
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 3240 8560 3292 8566
rect 3238 8528 3240 8537
rect 3292 8528 3294 8537
rect 3238 8463 3294 8472
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 3056 5636 3108 5642
rect 3056 5578 3108 5584
rect 2964 5160 3016 5166
rect 2964 5102 3016 5108
rect 2872 4684 2924 4690
rect 2872 4626 2924 4632
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2884 2446 2912 4626
rect 3068 3618 3096 5578
rect 3160 3738 3188 8366
rect 3240 8356 3292 8362
rect 3240 8298 3292 8304
rect 3252 7750 3280 8298
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 2976 3590 3096 3618
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 2688 2100 2740 2106
rect 2688 2042 2740 2048
rect 2688 1896 2740 1902
rect 2688 1838 2740 1844
rect 2504 1352 2556 1358
rect 2504 1294 2556 1300
rect 2700 1222 2728 1838
rect 2688 1216 2740 1222
rect 2688 1158 2740 1164
rect 2566 1116 2874 1125
rect 2566 1114 2572 1116
rect 2628 1114 2652 1116
rect 2708 1114 2732 1116
rect 2788 1114 2812 1116
rect 2868 1114 2874 1116
rect 2628 1062 2630 1114
rect 2810 1062 2812 1114
rect 2566 1060 2572 1062
rect 2628 1060 2652 1062
rect 2708 1060 2732 1062
rect 2788 1060 2812 1062
rect 2868 1060 2874 1062
rect 2566 1051 2874 1060
rect 2976 1018 3004 3590
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 3068 2582 3096 3470
rect 3252 3194 3280 7346
rect 3344 7342 3372 8774
rect 3436 8090 3464 10474
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3528 8022 3556 9454
rect 3620 8514 3648 12294
rect 3698 12200 3754 12294
rect 4158 12322 4214 13000
rect 4158 12294 4384 12322
rect 4158 12200 4214 12294
rect 3700 12164 3752 12170
rect 3700 12106 3752 12112
rect 3712 11694 3740 12106
rect 3700 11688 3752 11694
rect 3700 11630 3752 11636
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 3712 10606 3740 11630
rect 3884 11620 3936 11626
rect 3884 11562 3936 11568
rect 3792 11144 3844 11150
rect 3792 11086 3844 11092
rect 3700 10600 3752 10606
rect 3700 10542 3752 10548
rect 3700 9580 3752 9586
rect 3700 9522 3752 9528
rect 3712 9110 3740 9522
rect 3804 9450 3832 11086
rect 3896 10849 3924 11562
rect 3882 10840 3938 10849
rect 3882 10775 3938 10784
rect 4080 10606 4108 11630
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 3896 9897 3924 9998
rect 3882 9888 3938 9897
rect 3882 9823 3938 9832
rect 4080 9738 4108 10406
rect 4172 10198 4200 11494
rect 4252 11280 4304 11286
rect 4252 11222 4304 11228
rect 4264 10810 4292 11222
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 4160 10192 4212 10198
rect 4160 10134 4212 10140
rect 4252 9920 4304 9926
rect 4158 9888 4214 9897
rect 4252 9862 4304 9868
rect 4158 9823 4214 9832
rect 3896 9710 4108 9738
rect 3896 9674 3924 9710
rect 3896 9646 4016 9674
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 3792 9444 3844 9450
rect 3792 9386 3844 9392
rect 3896 9110 3924 9454
rect 3700 9104 3752 9110
rect 3700 9046 3752 9052
rect 3884 9104 3936 9110
rect 3884 9046 3936 9052
rect 3988 9042 4016 9646
rect 3792 9036 3844 9042
rect 3792 8978 3844 8984
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 3804 8906 3832 8978
rect 3792 8900 3844 8906
rect 3792 8842 3844 8848
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 3988 8786 4016 8978
rect 3620 8486 3832 8514
rect 3698 8256 3754 8265
rect 3698 8191 3754 8200
rect 3516 8016 3568 8022
rect 3568 7976 3648 8004
rect 3516 7958 3568 7964
rect 3424 7948 3476 7954
rect 3424 7890 3476 7896
rect 3332 7336 3384 7342
rect 3332 7278 3384 7284
rect 3344 5846 3372 7278
rect 3436 6866 3464 7890
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3332 5840 3384 5846
rect 3332 5782 3384 5788
rect 3332 5568 3384 5574
rect 3332 5510 3384 5516
rect 3344 4146 3372 5510
rect 3436 4690 3464 6054
rect 3424 4684 3476 4690
rect 3424 4626 3476 4632
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3424 3936 3476 3942
rect 3424 3878 3476 3884
rect 3436 3670 3464 3878
rect 3424 3664 3476 3670
rect 3424 3606 3476 3612
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3436 2774 3464 3606
rect 3344 2746 3464 2774
rect 3056 2576 3108 2582
rect 3056 2518 3108 2524
rect 3240 1828 3292 1834
rect 3240 1770 3292 1776
rect 3252 1562 3280 1770
rect 3240 1556 3292 1562
rect 3240 1498 3292 1504
rect 3056 1420 3108 1426
rect 3056 1362 3108 1368
rect 3068 1018 3096 1362
rect 3252 1018 3280 1498
rect 3344 1222 3372 2746
rect 3422 2680 3478 2689
rect 3422 2615 3478 2624
rect 3436 2514 3464 2615
rect 3424 2508 3476 2514
rect 3424 2450 3476 2456
rect 3424 2304 3476 2310
rect 3424 2246 3476 2252
rect 3436 1850 3464 2246
rect 3528 2038 3556 7822
rect 3620 7324 3648 7976
rect 3712 7954 3740 8191
rect 3700 7948 3752 7954
rect 3700 7890 3752 7896
rect 3700 7336 3752 7342
rect 3620 7296 3700 7324
rect 3700 7278 3752 7284
rect 3700 6996 3752 7002
rect 3700 6938 3752 6944
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3620 5234 3648 6190
rect 3712 6118 3740 6938
rect 3700 6112 3752 6118
rect 3700 6054 3752 6060
rect 3712 5817 3740 6054
rect 3698 5808 3754 5817
rect 3698 5743 3754 5752
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3712 5166 3740 5646
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 3608 4752 3660 4758
rect 3608 4694 3660 4700
rect 3620 2553 3648 4694
rect 3712 3942 3740 5102
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 3804 3534 3832 8486
rect 3896 7954 3924 8774
rect 3988 8758 4108 8786
rect 3974 8528 4030 8537
rect 3974 8463 3976 8472
rect 4028 8463 4030 8472
rect 3976 8434 4028 8440
rect 3884 7948 3936 7954
rect 3884 7890 3936 7896
rect 3896 6882 3924 7890
rect 4080 7478 4108 8758
rect 4068 7472 4120 7478
rect 4068 7414 4120 7420
rect 4172 7206 4200 9823
rect 4264 8974 4292 9862
rect 4252 8968 4304 8974
rect 4252 8910 4304 8916
rect 4252 8356 4304 8362
rect 4252 8298 4304 8304
rect 4264 8265 4292 8298
rect 4250 8256 4306 8265
rect 4250 8191 4306 8200
rect 4252 8016 4304 8022
rect 4252 7958 4304 7964
rect 4264 7546 4292 7958
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 4264 6882 4292 7346
rect 3896 6854 4016 6882
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3896 5914 3924 6734
rect 3988 6186 4016 6854
rect 4080 6854 4292 6882
rect 3976 6180 4028 6186
rect 3976 6122 4028 6128
rect 3974 6080 4030 6089
rect 3974 6015 4030 6024
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3896 4826 3924 5850
rect 3988 5710 4016 6015
rect 4080 5778 4108 6854
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 3988 5137 4016 5646
rect 3974 5128 4030 5137
rect 4030 5086 4108 5114
rect 3974 5063 4030 5072
rect 3884 4820 3936 4826
rect 3884 4762 3936 4768
rect 4080 4146 4108 5086
rect 4172 4826 4200 6734
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4264 4826 4292 6394
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4252 4820 4304 4826
rect 4252 4762 4304 4768
rect 4356 4706 4384 12294
rect 4618 12200 4674 13000
rect 5078 12200 5134 13000
rect 5538 12322 5594 13000
rect 5538 12294 5856 12322
rect 5538 12200 5594 12294
rect 4528 11144 4580 11150
rect 4528 11086 4580 11092
rect 4540 11014 4568 11086
rect 4436 11008 4488 11014
rect 4436 10950 4488 10956
rect 4528 11008 4580 11014
rect 4528 10950 4580 10956
rect 4172 4678 4384 4706
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 3882 4040 3938 4049
rect 3882 3975 3884 3984
rect 3936 3975 3938 3984
rect 3884 3946 3936 3952
rect 3988 3738 4016 4082
rect 4068 4004 4120 4010
rect 4068 3946 4120 3952
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 3988 3074 4016 3674
rect 4080 3534 4108 3946
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 3988 3058 4108 3074
rect 3988 3052 4120 3058
rect 3988 3046 4068 3052
rect 3988 2774 4016 3046
rect 4068 2994 4120 3000
rect 3896 2746 4016 2774
rect 3606 2544 3662 2553
rect 3896 2530 3924 2746
rect 4172 2666 4200 4678
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4250 2952 4306 2961
rect 4250 2887 4252 2896
rect 4304 2887 4306 2896
rect 4252 2858 4304 2864
rect 3988 2650 4200 2666
rect 3976 2644 4200 2650
rect 4028 2638 4200 2644
rect 3976 2586 4028 2592
rect 3606 2479 3662 2488
rect 3700 2508 3752 2514
rect 3896 2502 4108 2530
rect 3700 2450 3752 2456
rect 3516 2032 3568 2038
rect 3516 1974 3568 1980
rect 3436 1834 3648 1850
rect 3436 1828 3660 1834
rect 3436 1822 3608 1828
rect 3608 1770 3660 1776
rect 3332 1216 3384 1222
rect 3332 1158 3384 1164
rect 3712 1018 3740 2450
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 3896 1970 3924 2246
rect 3884 1964 3936 1970
rect 3884 1906 3936 1912
rect 4080 1902 4108 2502
rect 4068 1896 4120 1902
rect 4068 1838 4120 1844
rect 4172 1018 4200 2638
rect 4264 1426 4292 2858
rect 4356 2650 4384 4558
rect 4448 3194 4476 10950
rect 4528 10056 4580 10062
rect 4528 9998 4580 10004
rect 4540 9926 4568 9998
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 4632 8786 4660 12200
rect 4896 11620 4948 11626
rect 5092 11608 5120 12200
rect 5460 11886 5672 11914
rect 5460 11830 5488 11886
rect 5448 11824 5500 11830
rect 5448 11766 5500 11772
rect 5540 11824 5592 11830
rect 5540 11766 5592 11772
rect 4896 11562 4948 11568
rect 5000 11580 5120 11608
rect 4908 11218 4936 11562
rect 4896 11212 4948 11218
rect 4896 11154 4948 11160
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 4710 10840 4766 10849
rect 4710 10775 4712 10784
rect 4764 10775 4766 10784
rect 4712 10746 4764 10752
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4724 9450 4752 10406
rect 4712 9444 4764 9450
rect 4712 9386 4764 9392
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4540 8758 4660 8786
rect 4540 7410 4568 8758
rect 4528 7404 4580 7410
rect 4528 7346 4580 7352
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4528 6928 4580 6934
rect 4528 6870 4580 6876
rect 4540 5370 4568 6870
rect 4528 5364 4580 5370
rect 4528 5306 4580 5312
rect 4526 5128 4582 5137
rect 4526 5063 4528 5072
rect 4580 5063 4582 5072
rect 4528 5034 4580 5040
rect 4632 4865 4660 7142
rect 4618 4856 4674 4865
rect 4528 4820 4580 4826
rect 4618 4791 4674 4800
rect 4528 4762 4580 4768
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4434 2816 4490 2825
rect 4434 2751 4490 2760
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 4448 2106 4476 2751
rect 4540 2689 4568 4762
rect 4620 4684 4672 4690
rect 4620 4626 4672 4632
rect 4526 2680 4582 2689
rect 4526 2615 4582 2624
rect 4436 2100 4488 2106
rect 4436 2042 4488 2048
rect 4252 1420 4304 1426
rect 4252 1362 4304 1368
rect 2964 1012 3016 1018
rect 2964 954 3016 960
rect 3056 1012 3108 1018
rect 3056 954 3108 960
rect 3240 1012 3292 1018
rect 3240 954 3292 960
rect 3700 1012 3752 1018
rect 3700 954 3752 960
rect 4160 1012 4212 1018
rect 4160 954 4212 960
rect 4540 950 4568 2615
rect 4632 1902 4660 4626
rect 4724 2038 4752 8910
rect 4816 2106 4844 10950
rect 4896 8356 4948 8362
rect 4896 8298 4948 8304
rect 4908 7954 4936 8298
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 4908 5778 4936 6802
rect 4896 5772 4948 5778
rect 4896 5714 4948 5720
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4908 4622 4936 4966
rect 5000 4826 5028 11580
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5066 11452 5374 11461
rect 5066 11450 5072 11452
rect 5128 11450 5152 11452
rect 5208 11450 5232 11452
rect 5288 11450 5312 11452
rect 5368 11450 5374 11452
rect 5128 11398 5130 11450
rect 5310 11398 5312 11450
rect 5066 11396 5072 11398
rect 5128 11396 5152 11398
rect 5208 11396 5232 11398
rect 5288 11396 5312 11398
rect 5368 11396 5374 11398
rect 5066 11387 5374 11396
rect 5066 10364 5374 10373
rect 5066 10362 5072 10364
rect 5128 10362 5152 10364
rect 5208 10362 5232 10364
rect 5288 10362 5312 10364
rect 5368 10362 5374 10364
rect 5128 10310 5130 10362
rect 5310 10310 5312 10362
rect 5066 10308 5072 10310
rect 5128 10308 5152 10310
rect 5208 10308 5232 10310
rect 5288 10308 5312 10310
rect 5368 10308 5374 10310
rect 5066 10299 5374 10308
rect 5460 9654 5488 11494
rect 5552 10062 5580 11766
rect 5644 10606 5672 11886
rect 5724 11076 5776 11082
rect 5724 11018 5776 11024
rect 5632 10600 5684 10606
rect 5630 10568 5632 10577
rect 5684 10568 5686 10577
rect 5630 10503 5686 10512
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5448 9648 5500 9654
rect 5448 9590 5500 9596
rect 5736 9518 5764 11018
rect 5724 9512 5776 9518
rect 5630 9480 5686 9489
rect 5724 9454 5776 9460
rect 5630 9415 5686 9424
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5066 9276 5374 9285
rect 5066 9274 5072 9276
rect 5128 9274 5152 9276
rect 5208 9274 5232 9276
rect 5288 9274 5312 9276
rect 5368 9274 5374 9276
rect 5128 9222 5130 9274
rect 5310 9222 5312 9274
rect 5066 9220 5072 9222
rect 5128 9220 5152 9222
rect 5208 9220 5232 9222
rect 5288 9220 5312 9222
rect 5368 9220 5374 9222
rect 5066 9211 5374 9220
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5368 8537 5396 8570
rect 5354 8528 5410 8537
rect 5354 8463 5410 8472
rect 5066 8188 5374 8197
rect 5066 8186 5072 8188
rect 5128 8186 5152 8188
rect 5208 8186 5232 8188
rect 5288 8186 5312 8188
rect 5368 8186 5374 8188
rect 5128 8134 5130 8186
rect 5310 8134 5312 8186
rect 5066 8132 5072 8134
rect 5128 8132 5152 8134
rect 5208 8132 5232 8134
rect 5288 8132 5312 8134
rect 5368 8132 5374 8134
rect 5066 8123 5374 8132
rect 5460 7954 5488 9318
rect 5540 9104 5592 9110
rect 5540 9046 5592 9052
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5066 7100 5374 7109
rect 5066 7098 5072 7100
rect 5128 7098 5152 7100
rect 5208 7098 5232 7100
rect 5288 7098 5312 7100
rect 5368 7098 5374 7100
rect 5128 7046 5130 7098
rect 5310 7046 5312 7098
rect 5066 7044 5072 7046
rect 5128 7044 5152 7046
rect 5208 7044 5232 7046
rect 5288 7044 5312 7046
rect 5368 7044 5374 7046
rect 5066 7035 5374 7044
rect 5066 6012 5374 6021
rect 5066 6010 5072 6012
rect 5128 6010 5152 6012
rect 5208 6010 5232 6012
rect 5288 6010 5312 6012
rect 5368 6010 5374 6012
rect 5128 5958 5130 6010
rect 5310 5958 5312 6010
rect 5066 5956 5072 5958
rect 5128 5956 5152 5958
rect 5208 5956 5232 5958
rect 5288 5956 5312 5958
rect 5368 5956 5374 5958
rect 5066 5947 5374 5956
rect 5354 5808 5410 5817
rect 5354 5743 5356 5752
rect 5408 5743 5410 5752
rect 5356 5714 5408 5720
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 5092 5030 5120 5646
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 5368 5137 5396 5578
rect 5354 5128 5410 5137
rect 5354 5063 5410 5072
rect 5080 5024 5132 5030
rect 5080 4966 5132 4972
rect 5066 4924 5374 4933
rect 5066 4922 5072 4924
rect 5128 4922 5152 4924
rect 5208 4922 5232 4924
rect 5288 4922 5312 4924
rect 5368 4922 5374 4924
rect 5128 4870 5130 4922
rect 5310 4870 5312 4922
rect 5066 4868 5072 4870
rect 5128 4868 5152 4870
rect 5208 4868 5232 4870
rect 5288 4868 5312 4870
rect 5368 4868 5374 4870
rect 5066 4859 5374 4868
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 5356 4752 5408 4758
rect 5262 4720 5318 4729
rect 5356 4694 5408 4700
rect 5262 4655 5318 4664
rect 4896 4616 4948 4622
rect 4948 4576 5028 4604
rect 4896 4558 4948 4564
rect 4896 3664 4948 3670
rect 4894 3632 4896 3641
rect 4948 3632 4950 3641
rect 4894 3567 4950 3576
rect 5000 3398 5028 4576
rect 5276 3942 5304 4655
rect 5368 4282 5396 4694
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5354 4176 5410 4185
rect 5460 4146 5488 7278
rect 5354 4111 5410 4120
rect 5448 4140 5500 4146
rect 5368 4078 5396 4111
rect 5448 4082 5500 4088
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 5066 3836 5374 3845
rect 5066 3834 5072 3836
rect 5128 3834 5152 3836
rect 5208 3834 5232 3836
rect 5288 3834 5312 3836
rect 5368 3834 5374 3836
rect 5128 3782 5130 3834
rect 5310 3782 5312 3834
rect 5066 3780 5072 3782
rect 5128 3780 5152 3782
rect 5208 3780 5232 3782
rect 5288 3780 5312 3782
rect 5368 3780 5374 3782
rect 5066 3771 5374 3780
rect 5460 3602 5488 4082
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 5368 3194 5396 3470
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 5446 2952 5502 2961
rect 4896 2916 4948 2922
rect 5446 2887 5502 2896
rect 4896 2858 4948 2864
rect 4908 2825 4936 2858
rect 4894 2816 4950 2825
rect 4894 2751 4950 2760
rect 5066 2748 5374 2757
rect 5066 2746 5072 2748
rect 5128 2746 5152 2748
rect 5208 2746 5232 2748
rect 5288 2746 5312 2748
rect 5368 2746 5374 2748
rect 5128 2694 5130 2746
rect 5310 2694 5312 2746
rect 5066 2692 5072 2694
rect 5128 2692 5152 2694
rect 5208 2692 5232 2694
rect 5288 2692 5312 2694
rect 5368 2692 5374 2694
rect 5066 2683 5374 2692
rect 4894 2544 4950 2553
rect 4894 2479 4896 2488
rect 4948 2479 4950 2488
rect 5356 2508 5408 2514
rect 4896 2450 4948 2456
rect 5356 2450 5408 2456
rect 4804 2100 4856 2106
rect 4804 2042 4856 2048
rect 4712 2032 4764 2038
rect 4712 1974 4764 1980
rect 4620 1896 4672 1902
rect 4620 1838 4672 1844
rect 4908 1562 4936 2450
rect 4988 2304 5040 2310
rect 4988 2246 5040 2252
rect 5080 2304 5132 2310
rect 5080 2246 5132 2252
rect 4896 1556 4948 1562
rect 4896 1498 4948 1504
rect 5000 1494 5028 2246
rect 5092 1766 5120 2246
rect 5368 1902 5396 2450
rect 5460 2106 5488 2887
rect 5552 2650 5580 9046
rect 5644 7342 5672 9415
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 5736 8401 5764 9318
rect 5722 8392 5778 8401
rect 5722 8327 5778 8336
rect 5736 8294 5764 8327
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5632 7336 5684 7342
rect 5630 7304 5632 7313
rect 5828 7324 5856 12294
rect 5998 12200 6054 13000
rect 6458 12322 6514 13000
rect 22098 12608 22154 12617
rect 22098 12543 22154 12552
rect 8760 12436 8812 12442
rect 8760 12378 8812 12384
rect 6458 12294 6684 12322
rect 6184 12232 6236 12238
rect 5908 12096 5960 12102
rect 5908 12038 5960 12044
rect 5920 11694 5948 12038
rect 5908 11688 5960 11694
rect 5908 11630 5960 11636
rect 5908 10804 5960 10810
rect 5908 10746 5960 10752
rect 5920 8294 5948 10746
rect 6012 8498 6040 12200
rect 6458 12200 6514 12294
rect 6184 12174 6236 12180
rect 6196 11694 6224 12174
rect 6184 11688 6236 11694
rect 6368 11688 6420 11694
rect 6184 11630 6236 11636
rect 6288 11636 6368 11642
rect 6288 11630 6420 11636
rect 6288 11614 6408 11630
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6196 10810 6224 11086
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6092 10600 6144 10606
rect 6092 10542 6144 10548
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 5684 7304 5686 7313
rect 5630 7239 5686 7248
rect 5736 7296 5856 7324
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5644 5302 5672 7142
rect 5736 6361 5764 7296
rect 5722 6352 5778 6361
rect 5722 6287 5778 6296
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 5724 6248 5776 6254
rect 5724 6190 5776 6196
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5644 4078 5672 4966
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5644 3534 5672 3878
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 5736 2650 5764 6190
rect 5828 4282 5856 6258
rect 5920 5166 5948 7686
rect 6000 7472 6052 7478
rect 6000 7414 6052 7420
rect 6012 6934 6040 7414
rect 6000 6928 6052 6934
rect 6000 6870 6052 6876
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 6012 5234 6040 5646
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 6012 4758 6040 5170
rect 6000 4752 6052 4758
rect 6000 4694 6052 4700
rect 5906 4584 5962 4593
rect 5906 4519 5962 4528
rect 5816 4276 5868 4282
rect 5816 4218 5868 4224
rect 5814 4176 5870 4185
rect 5814 4111 5870 4120
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 5644 2530 5672 2586
rect 5828 2530 5856 4111
rect 5920 2990 5948 4519
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 6012 4049 6040 4218
rect 5998 4040 6054 4049
rect 5998 3975 6054 3984
rect 6104 3738 6132 10542
rect 6288 10146 6316 11614
rect 6460 11552 6512 11558
rect 6460 11494 6512 11500
rect 6472 11150 6500 11494
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 6472 10606 6500 10746
rect 6460 10600 6512 10606
rect 6460 10542 6512 10548
rect 6288 10130 6408 10146
rect 6288 10124 6420 10130
rect 6288 10118 6368 10124
rect 6184 9920 6236 9926
rect 6184 9862 6236 9868
rect 6196 9110 6224 9862
rect 6184 9104 6236 9110
rect 6184 9046 6236 9052
rect 6184 8968 6236 8974
rect 6184 8910 6236 8916
rect 6196 8430 6224 8910
rect 6184 8424 6236 8430
rect 6184 8366 6236 8372
rect 6288 7750 6316 10118
rect 6368 10066 6420 10072
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6380 7886 6408 9522
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6276 7336 6328 7342
rect 6276 7278 6328 7284
rect 6288 7002 6316 7278
rect 6276 6996 6328 7002
rect 6276 6938 6328 6944
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 6196 6458 6224 6734
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 5908 2984 5960 2990
rect 5908 2926 5960 2932
rect 5644 2502 5856 2530
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 5448 2100 5500 2106
rect 5448 2042 5500 2048
rect 5356 1896 5408 1902
rect 5356 1838 5408 1844
rect 5080 1760 5132 1766
rect 5080 1702 5132 1708
rect 5066 1660 5374 1669
rect 5066 1658 5072 1660
rect 5128 1658 5152 1660
rect 5208 1658 5232 1660
rect 5288 1658 5312 1660
rect 5368 1658 5374 1660
rect 5128 1606 5130 1658
rect 5310 1606 5312 1658
rect 5066 1604 5072 1606
rect 5128 1604 5152 1606
rect 5208 1604 5232 1606
rect 5288 1604 5312 1606
rect 5368 1604 5374 1606
rect 5066 1595 5374 1604
rect 5736 1562 5764 2382
rect 5920 2106 5948 2926
rect 6000 2372 6052 2378
rect 6000 2314 6052 2320
rect 6012 2106 6040 2314
rect 5908 2100 5960 2106
rect 5908 2042 5960 2048
rect 6000 2100 6052 2106
rect 6000 2042 6052 2048
rect 6092 2032 6144 2038
rect 6092 1974 6144 1980
rect 5724 1556 5776 1562
rect 5724 1498 5776 1504
rect 4988 1488 5040 1494
rect 4988 1430 5040 1436
rect 5080 1488 5132 1494
rect 5080 1430 5132 1436
rect 5092 1018 5120 1430
rect 6000 1352 6052 1358
rect 6104 1340 6132 1974
rect 6288 1426 6316 6598
rect 6380 4214 6408 7822
rect 6368 4208 6420 4214
rect 6368 4150 6420 4156
rect 6472 2854 6500 10542
rect 6552 9988 6604 9994
rect 6552 9930 6604 9936
rect 6564 9722 6592 9930
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 6564 9178 6592 9454
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6656 9081 6684 12294
rect 7104 12164 7156 12170
rect 7104 12106 7156 12112
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6642 9072 6698 9081
rect 6552 9036 6604 9042
rect 6748 9042 6776 10610
rect 6642 9007 6698 9016
rect 6736 9036 6788 9042
rect 6552 8978 6604 8984
rect 6736 8978 6788 8984
rect 6564 8537 6592 8978
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6550 8528 6606 8537
rect 6550 8463 6606 8472
rect 6656 8362 6684 8910
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6564 5250 6592 8230
rect 6656 5370 6684 8298
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6564 5222 6684 5250
rect 6552 5092 6604 5098
rect 6552 5034 6604 5040
rect 6564 4690 6592 5034
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6552 4480 6604 4486
rect 6552 4422 6604 4428
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 6564 2514 6592 4422
rect 6656 3126 6684 5222
rect 6748 4010 6776 8774
rect 6840 8090 6868 11154
rect 6932 10538 6960 11494
rect 7024 11286 7052 11494
rect 7116 11286 7144 12106
rect 7566 11996 7874 12005
rect 7566 11994 7572 11996
rect 7628 11994 7652 11996
rect 7708 11994 7732 11996
rect 7788 11994 7812 11996
rect 7868 11994 7874 11996
rect 7628 11942 7630 11994
rect 7810 11942 7812 11994
rect 7566 11940 7572 11942
rect 7628 11940 7652 11942
rect 7708 11940 7732 11942
rect 7788 11940 7812 11942
rect 7868 11940 7874 11942
rect 7566 11931 7874 11940
rect 8772 11762 8800 12378
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 7012 11280 7064 11286
rect 7012 11222 7064 11228
rect 7104 11280 7156 11286
rect 7104 11222 7156 11228
rect 7116 11150 7144 11222
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 7208 10130 7236 10950
rect 7566 10908 7874 10917
rect 7566 10906 7572 10908
rect 7628 10906 7652 10908
rect 7708 10906 7732 10908
rect 7788 10906 7812 10908
rect 7868 10906 7874 10908
rect 7628 10854 7630 10906
rect 7810 10854 7812 10906
rect 7566 10852 7572 10854
rect 7628 10852 7652 10854
rect 7708 10852 7732 10854
rect 7788 10852 7812 10854
rect 7868 10852 7874 10854
rect 7566 10843 7874 10852
rect 7380 10736 7432 10742
rect 7380 10678 7432 10684
rect 7392 10554 7420 10678
rect 7300 10526 7420 10554
rect 7470 10568 7526 10577
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 7300 10062 7328 10526
rect 7470 10503 7526 10512
rect 7484 10470 7512 10503
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 6828 7744 6880 7750
rect 6828 7686 6880 7692
rect 6736 4004 6788 4010
rect 6736 3946 6788 3952
rect 6644 3120 6696 3126
rect 6644 3062 6696 3068
rect 6748 2774 6776 3946
rect 6656 2746 6776 2774
rect 6656 2582 6684 2746
rect 6644 2576 6696 2582
rect 6644 2518 6696 2524
rect 6552 2508 6604 2514
rect 6552 2450 6604 2456
rect 6840 2310 6868 7686
rect 6932 4146 6960 9998
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 7012 8832 7064 8838
rect 7012 8774 7064 8780
rect 7024 7342 7052 8774
rect 7116 7954 7144 9930
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7300 8090 7328 8910
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 7116 7426 7144 7890
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7116 7398 7236 7426
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 7104 7268 7156 7274
rect 7104 7210 7156 7216
rect 7116 6866 7144 7210
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 7208 6798 7236 7398
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 7300 6338 7328 7686
rect 7392 6866 7420 10406
rect 7566 9820 7874 9829
rect 7566 9818 7572 9820
rect 7628 9818 7652 9820
rect 7708 9818 7732 9820
rect 7788 9818 7812 9820
rect 7868 9818 7874 9820
rect 7628 9766 7630 9818
rect 7810 9766 7812 9818
rect 7566 9764 7572 9766
rect 7628 9764 7652 9766
rect 7708 9764 7732 9766
rect 7788 9764 7812 9766
rect 7868 9764 7874 9766
rect 7566 9755 7874 9764
rect 7566 8732 7874 8741
rect 7566 8730 7572 8732
rect 7628 8730 7652 8732
rect 7708 8730 7732 8732
rect 7788 8730 7812 8732
rect 7868 8730 7874 8732
rect 7628 8678 7630 8730
rect 7810 8678 7812 8730
rect 7566 8676 7572 8678
rect 7628 8676 7652 8678
rect 7708 8676 7732 8678
rect 7788 8676 7812 8678
rect 7868 8676 7874 8678
rect 7566 8667 7874 8676
rect 7470 8392 7526 8401
rect 7470 8327 7526 8336
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 7208 6310 7328 6338
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 7024 4826 7052 6122
rect 7104 5772 7156 5778
rect 7104 5714 7156 5720
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 7116 4690 7144 5714
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 6828 2304 6880 2310
rect 6828 2246 6880 2252
rect 7012 2032 7064 2038
rect 7012 1974 7064 1980
rect 7024 1816 7052 1974
rect 7116 1970 7144 4626
rect 7208 3738 7236 6310
rect 7288 6248 7340 6254
rect 7288 6190 7340 6196
rect 7300 5846 7328 6190
rect 7288 5840 7340 5846
rect 7288 5782 7340 5788
rect 7392 5710 7420 6802
rect 7288 5704 7340 5710
rect 7288 5646 7340 5652
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7300 5574 7328 5646
rect 7288 5568 7340 5574
rect 7484 5556 7512 8327
rect 7944 8090 7972 11698
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 9126 11656 9182 11665
rect 8116 11620 8168 11626
rect 8116 11562 8168 11568
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 7932 8084 7984 8090
rect 7932 8026 7984 8032
rect 7566 7644 7874 7653
rect 7566 7642 7572 7644
rect 7628 7642 7652 7644
rect 7708 7642 7732 7644
rect 7788 7642 7812 7644
rect 7868 7642 7874 7644
rect 7628 7590 7630 7642
rect 7810 7590 7812 7642
rect 7566 7588 7572 7590
rect 7628 7588 7652 7590
rect 7708 7588 7732 7590
rect 7788 7588 7812 7590
rect 7868 7588 7874 7590
rect 7566 7579 7874 7588
rect 8036 7154 8064 9998
rect 8128 7313 8156 11562
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8208 9444 8260 9450
rect 8208 9386 8260 9392
rect 8220 9042 8248 9386
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8114 7304 8170 7313
rect 8114 7239 8170 7248
rect 8036 7126 8248 7154
rect 8116 6928 8168 6934
rect 8116 6870 8168 6876
rect 8022 6624 8078 6633
rect 7566 6556 7874 6565
rect 8022 6559 8078 6568
rect 7566 6554 7572 6556
rect 7628 6554 7652 6556
rect 7708 6554 7732 6556
rect 7788 6554 7812 6556
rect 7868 6554 7874 6556
rect 7628 6502 7630 6554
rect 7810 6502 7812 6554
rect 7566 6500 7572 6502
rect 7628 6500 7652 6502
rect 7708 6500 7732 6502
rect 7788 6500 7812 6502
rect 7868 6500 7874 6502
rect 7566 6491 7874 6500
rect 7840 6384 7892 6390
rect 7838 6352 7840 6361
rect 7892 6352 7894 6361
rect 7838 6287 7894 6296
rect 7748 6248 7800 6254
rect 7748 6190 7800 6196
rect 7760 5642 7788 6190
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7852 5658 7880 6054
rect 7748 5636 7800 5642
rect 7852 5630 7972 5658
rect 7748 5578 7800 5584
rect 7288 5510 7340 5516
rect 7392 5528 7512 5556
rect 7300 4690 7328 5510
rect 7392 4826 7420 5528
rect 7566 5468 7874 5477
rect 7566 5466 7572 5468
rect 7628 5466 7652 5468
rect 7708 5466 7732 5468
rect 7788 5466 7812 5468
rect 7868 5466 7874 5468
rect 7628 5414 7630 5466
rect 7810 5414 7812 5466
rect 7566 5412 7572 5414
rect 7628 5412 7652 5414
rect 7708 5412 7732 5414
rect 7788 5412 7812 5414
rect 7868 5412 7874 5414
rect 7566 5403 7874 5412
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 7300 3670 7328 4626
rect 7288 3664 7340 3670
rect 7288 3606 7340 3612
rect 7392 2582 7420 4762
rect 7470 4584 7526 4593
rect 7470 4519 7526 4528
rect 7484 4146 7512 4519
rect 7566 4380 7874 4389
rect 7566 4378 7572 4380
rect 7628 4378 7652 4380
rect 7708 4378 7732 4380
rect 7788 4378 7812 4380
rect 7868 4378 7874 4380
rect 7628 4326 7630 4378
rect 7810 4326 7812 4378
rect 7566 4324 7572 4326
rect 7628 4324 7652 4326
rect 7708 4324 7732 4326
rect 7788 4324 7812 4326
rect 7868 4324 7874 4326
rect 7566 4315 7874 4324
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7566 3292 7874 3301
rect 7566 3290 7572 3292
rect 7628 3290 7652 3292
rect 7708 3290 7732 3292
rect 7788 3290 7812 3292
rect 7868 3290 7874 3292
rect 7628 3238 7630 3290
rect 7810 3238 7812 3290
rect 7566 3236 7572 3238
rect 7628 3236 7652 3238
rect 7708 3236 7732 3238
rect 7788 3236 7812 3238
rect 7868 3236 7874 3238
rect 7566 3227 7874 3236
rect 7380 2576 7432 2582
rect 7380 2518 7432 2524
rect 7566 2204 7874 2213
rect 7566 2202 7572 2204
rect 7628 2202 7652 2204
rect 7708 2202 7732 2204
rect 7788 2202 7812 2204
rect 7868 2202 7874 2204
rect 7628 2150 7630 2202
rect 7810 2150 7812 2202
rect 7566 2148 7572 2150
rect 7628 2148 7652 2150
rect 7708 2148 7732 2150
rect 7788 2148 7812 2150
rect 7868 2148 7874 2150
rect 7566 2139 7874 2148
rect 7472 2100 7524 2106
rect 7472 2042 7524 2048
rect 7104 1964 7156 1970
rect 7104 1906 7156 1912
rect 7380 1828 7432 1834
rect 7024 1788 7380 1816
rect 7380 1770 7432 1776
rect 7484 1562 7512 2042
rect 7944 1902 7972 5630
rect 8036 2990 8064 6559
rect 8128 4826 8156 6870
rect 8116 4820 8168 4826
rect 8116 4762 8168 4768
rect 8114 4720 8170 4729
rect 8114 4655 8116 4664
rect 8168 4655 8170 4664
rect 8116 4626 8168 4632
rect 8116 4548 8168 4554
rect 8116 4490 8168 4496
rect 8128 4282 8156 4490
rect 8116 4276 8168 4282
rect 8116 4218 8168 4224
rect 8220 4214 8248 7126
rect 8312 5166 8340 9318
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 8206 4040 8262 4049
rect 8206 3975 8262 3984
rect 8024 2984 8076 2990
rect 8024 2926 8076 2932
rect 8220 2774 8248 3975
rect 8128 2746 8248 2774
rect 7932 1896 7984 1902
rect 7932 1838 7984 1844
rect 7472 1556 7524 1562
rect 7472 1498 7524 1504
rect 6276 1420 6328 1426
rect 6276 1362 6328 1368
rect 6052 1312 6132 1340
rect 6000 1294 6052 1300
rect 5080 1012 5132 1018
rect 5080 954 5132 960
rect 5816 1012 5868 1018
rect 5816 954 5868 960
rect 2412 944 2464 950
rect 3332 944 3384 950
rect 2412 886 2464 892
rect 2594 912 2650 921
rect 3332 886 3384 892
rect 4528 944 4580 950
rect 4528 886 4580 892
rect 2594 847 2650 856
rect 2608 814 2636 847
rect 2320 808 2372 814
rect 2320 750 2372 756
rect 2596 808 2648 814
rect 2596 750 2648 756
rect 3344 678 3372 886
rect 5828 746 5856 954
rect 6104 950 6132 1312
rect 7566 1116 7874 1125
rect 7566 1114 7572 1116
rect 7628 1114 7652 1116
rect 7708 1114 7732 1116
rect 7788 1114 7812 1116
rect 7868 1114 7874 1116
rect 7628 1062 7630 1114
rect 7810 1062 7812 1114
rect 7566 1060 7572 1062
rect 7628 1060 7652 1062
rect 7708 1060 7732 1062
rect 7788 1060 7812 1062
rect 7868 1060 7874 1062
rect 7566 1051 7874 1060
rect 6092 944 6144 950
rect 6092 886 6144 892
rect 5816 740 5868 746
rect 5816 682 5868 688
rect 8128 678 8156 2746
rect 8312 1766 8340 4966
rect 8404 2650 8432 11086
rect 8496 9586 8524 11630
rect 9126 11591 9182 11600
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 8852 9512 8904 9518
rect 8852 9454 8904 9460
rect 8864 9382 8892 9454
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8852 9376 8904 9382
rect 8852 9318 8904 9324
rect 8772 9110 8800 9318
rect 8484 9104 8536 9110
rect 8484 9046 8536 9052
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8496 8566 8524 9046
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 8496 4468 8524 8502
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8588 7478 8616 8366
rect 8576 7472 8628 7478
rect 8576 7414 8628 7420
rect 8680 7342 8708 8434
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8576 7336 8628 7342
rect 8574 7304 8576 7313
rect 8668 7336 8720 7342
rect 8628 7304 8630 7313
rect 8668 7278 8720 7284
rect 8574 7239 8630 7248
rect 8576 6656 8628 6662
rect 8574 6624 8576 6633
rect 8772 6633 8800 7686
rect 8628 6624 8630 6633
rect 8574 6559 8630 6568
rect 8758 6624 8814 6633
rect 8758 6559 8814 6568
rect 8758 6352 8814 6361
rect 8668 6316 8720 6322
rect 8588 6276 8668 6304
rect 8588 5098 8616 6276
rect 8758 6287 8814 6296
rect 8668 6258 8720 6264
rect 8772 5778 8800 6287
rect 8760 5772 8812 5778
rect 8760 5714 8812 5720
rect 8668 5636 8720 5642
rect 8668 5578 8720 5584
rect 8576 5092 8628 5098
rect 8576 5034 8628 5040
rect 8576 4480 8628 4486
rect 8496 4440 8576 4468
rect 8576 4422 8628 4428
rect 8484 4004 8536 4010
rect 8484 3946 8536 3952
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 8496 2514 8524 3946
rect 8680 2650 8708 5578
rect 8760 5092 8812 5098
rect 8760 5034 8812 5040
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 8772 2514 8800 5034
rect 8864 5030 8892 9318
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 8956 7449 8984 9114
rect 8942 7440 8998 7449
rect 8942 7375 8998 7384
rect 8942 7304 8998 7313
rect 8942 7239 8998 7248
rect 8956 6372 8984 7239
rect 9048 6497 9076 11494
rect 9140 11218 9168 11591
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 9232 11286 9260 11494
rect 9220 11280 9272 11286
rect 9220 11222 9272 11228
rect 9128 11212 9180 11218
rect 9128 11154 9180 11160
rect 9324 10674 9352 11834
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 9864 11688 9916 11694
rect 9864 11630 9916 11636
rect 9772 11620 9824 11626
rect 9772 11562 9824 11568
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9220 10600 9272 10606
rect 9220 10542 9272 10548
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 9140 8566 9168 9454
rect 9128 8560 9180 8566
rect 9128 8502 9180 8508
rect 9232 8430 9260 10542
rect 9784 10266 9812 11562
rect 9876 10690 9904 11630
rect 9968 10810 9996 11698
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 9876 10662 9996 10690
rect 9968 10606 9996 10662
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 9968 10470 9996 10542
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 9692 9654 9720 10202
rect 9968 10130 9996 10406
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 10244 10062 10272 11630
rect 10416 11076 10468 11082
rect 10416 11018 10468 11024
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9324 9382 9352 9522
rect 9312 9376 9364 9382
rect 9312 9318 9364 9324
rect 9784 9042 9812 9930
rect 10140 9920 10192 9926
rect 10140 9862 10192 9868
rect 9864 9512 9916 9518
rect 9864 9454 9916 9460
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9496 8560 9548 8566
rect 9496 8502 9548 8508
rect 9680 8560 9732 8566
rect 9680 8502 9732 8508
rect 9220 8424 9272 8430
rect 9220 8366 9272 8372
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9128 8356 9180 8362
rect 9128 8298 9180 8304
rect 9140 7954 9168 8298
rect 9128 7948 9180 7954
rect 9128 7890 9180 7896
rect 9126 7576 9182 7585
rect 9126 7511 9128 7520
rect 9180 7511 9182 7520
rect 9128 7482 9180 7488
rect 9126 7440 9182 7449
rect 9126 7375 9182 7384
rect 9034 6488 9090 6497
rect 9034 6423 9090 6432
rect 9036 6384 9088 6390
rect 8956 6344 9036 6372
rect 9036 6326 9088 6332
rect 8942 6216 8998 6225
rect 8942 6151 8998 6160
rect 8852 5024 8904 5030
rect 8852 4966 8904 4972
rect 8852 4276 8904 4282
rect 8852 4218 8904 4224
rect 8864 3602 8892 4218
rect 8852 3596 8904 3602
rect 8852 3538 8904 3544
rect 8956 2990 8984 6151
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 9048 4185 9076 5714
rect 9034 4176 9090 4185
rect 9034 4111 9090 4120
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 9048 2582 9076 3674
rect 9140 3534 9168 7375
rect 9232 6934 9260 8366
rect 9324 7857 9352 8366
rect 9508 7993 9536 8502
rect 9692 8430 9720 8502
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9588 8356 9640 8362
rect 9588 8298 9640 8304
rect 9772 8356 9824 8362
rect 9772 8298 9824 8304
rect 9600 8129 9628 8298
rect 9586 8120 9642 8129
rect 9586 8055 9642 8064
rect 9494 7984 9550 7993
rect 9494 7919 9550 7928
rect 9496 7880 9548 7886
rect 9310 7848 9366 7857
rect 9310 7783 9366 7792
rect 9494 7848 9496 7857
rect 9548 7848 9550 7857
rect 9494 7783 9550 7792
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9600 7585 9628 7754
rect 9310 7576 9366 7585
rect 9586 7576 9642 7585
rect 9366 7520 9536 7528
rect 9310 7511 9536 7520
rect 9586 7511 9642 7520
rect 9325 7500 9536 7511
rect 9508 7460 9536 7500
rect 9588 7472 9640 7478
rect 9508 7432 9588 7460
rect 9588 7414 9640 7420
rect 9496 7336 9548 7342
rect 9310 7304 9366 7313
rect 9496 7278 9548 7284
rect 9586 7304 9642 7313
rect 9310 7239 9366 7248
rect 9324 7002 9352 7239
rect 9312 6996 9364 7002
rect 9312 6938 9364 6944
rect 9220 6928 9272 6934
rect 9508 6905 9536 7278
rect 9586 7239 9642 7248
rect 9220 6870 9272 6876
rect 9494 6896 9550 6905
rect 9232 6186 9260 6870
rect 9494 6831 9550 6840
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9402 6352 9458 6361
rect 9402 6287 9458 6296
rect 9416 6254 9444 6287
rect 9404 6248 9456 6254
rect 9404 6190 9456 6196
rect 9220 6180 9272 6186
rect 9220 6122 9272 6128
rect 9404 6112 9456 6118
rect 9402 6080 9404 6089
rect 9456 6080 9458 6089
rect 9402 6015 9458 6024
rect 9508 5778 9536 6734
rect 9600 6186 9628 7239
rect 9784 6866 9812 8298
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9588 6180 9640 6186
rect 9588 6122 9640 6128
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9600 5710 9628 6122
rect 9876 5846 9904 9454
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 9956 8424 10008 8430
rect 9954 8392 9956 8401
rect 10008 8392 10010 8401
rect 9954 8327 10010 8336
rect 9956 7744 10008 7750
rect 9956 7686 10008 7692
rect 9968 6322 9996 7686
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 9864 5840 9916 5846
rect 9864 5782 9916 5788
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9416 4826 9444 5646
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 9588 4752 9640 4758
rect 9508 4712 9588 4740
rect 9404 4276 9456 4282
rect 9404 4218 9456 4224
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9232 3602 9260 3878
rect 9220 3596 9272 3602
rect 9220 3538 9272 3544
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 9218 3496 9274 3505
rect 9036 2576 9088 2582
rect 9036 2518 9088 2524
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 8576 2508 8628 2514
rect 8576 2450 8628 2456
rect 8760 2508 8812 2514
rect 8760 2450 8812 2456
rect 8300 1760 8352 1766
rect 8300 1702 8352 1708
rect 8588 1426 8616 2450
rect 8668 2304 8720 2310
rect 8668 2246 8720 2252
rect 8576 1420 8628 1426
rect 8576 1362 8628 1368
rect 8680 814 8708 2246
rect 9140 1358 9168 3470
rect 9218 3431 9220 3440
rect 9272 3431 9274 3440
rect 9220 3402 9272 3408
rect 9416 1494 9444 4218
rect 9508 2650 9536 4712
rect 9588 4694 9640 4700
rect 9600 4486 9628 4694
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 9600 3670 9628 3878
rect 9588 3664 9640 3670
rect 9588 3606 9640 3612
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9692 2650 9720 3130
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9784 1902 9812 5646
rect 9772 1896 9824 1902
rect 9772 1838 9824 1844
rect 9404 1488 9456 1494
rect 9404 1430 9456 1436
rect 9128 1352 9180 1358
rect 9128 1294 9180 1300
rect 9036 1216 9088 1222
rect 9036 1158 9088 1164
rect 9128 1216 9180 1222
rect 9128 1158 9180 1164
rect 8758 912 8814 921
rect 9048 882 9076 1158
rect 9140 950 9168 1158
rect 9416 1034 9444 1430
rect 9680 1352 9732 1358
rect 9680 1294 9732 1300
rect 9416 1018 9536 1034
rect 9416 1012 9548 1018
rect 9416 1006 9496 1012
rect 9496 954 9548 960
rect 9128 944 9180 950
rect 9128 886 9180 892
rect 8758 847 8814 856
rect 9036 876 9088 882
rect 8772 814 8800 847
rect 9036 818 9088 824
rect 9692 814 9720 1294
rect 9876 1290 9904 5782
rect 10060 3738 10088 8910
rect 10152 5710 10180 9862
rect 10244 7478 10272 9998
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10232 7472 10284 7478
rect 10232 7414 10284 7420
rect 10232 7336 10284 7342
rect 10232 7278 10284 7284
rect 10244 6934 10272 7278
rect 10232 6928 10284 6934
rect 10232 6870 10284 6876
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 10152 5574 10180 5646
rect 10244 5642 10272 6734
rect 10232 5636 10284 5642
rect 10232 5578 10284 5584
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 10336 4622 10364 8978
rect 10428 5778 10456 11018
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 10324 4616 10376 4622
rect 10324 4558 10376 4564
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 10428 3466 10456 5714
rect 10416 3460 10468 3466
rect 10416 3402 10468 3408
rect 10520 3398 10548 12038
rect 17222 11928 17278 11937
rect 17222 11863 17278 11872
rect 16854 11520 16910 11529
rect 16854 11455 16910 11464
rect 16762 11112 16818 11121
rect 16580 11076 16632 11082
rect 16762 11047 16818 11056
rect 16580 11018 16632 11024
rect 10784 10124 10836 10130
rect 10784 10066 10836 10072
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10612 7274 10640 9318
rect 10600 7268 10652 7274
rect 10600 7210 10652 7216
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 10796 2650 10824 10066
rect 16592 9489 16620 11018
rect 16670 10704 16726 10713
rect 16670 10639 16726 10648
rect 16578 9480 16634 9489
rect 16578 9415 16634 9424
rect 16684 8838 16712 10639
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11060 7132 11112 7138
rect 11060 7074 11112 7080
rect 11072 3194 11100 7074
rect 11152 5636 11204 5642
rect 11152 5578 11204 5584
rect 11060 3188 11112 3194
rect 11060 3130 11112 3136
rect 11164 3058 11192 5578
rect 11256 5370 11284 8366
rect 16776 8362 16804 11047
rect 16868 9654 16896 11455
rect 16946 10296 17002 10305
rect 16946 10231 17002 10240
rect 16856 9648 16908 9654
rect 16856 9590 16908 9596
rect 16764 8356 16816 8362
rect 16764 8298 16816 8304
rect 12348 8288 12400 8294
rect 12348 8230 12400 8236
rect 12360 7954 12388 8230
rect 16960 8090 16988 10231
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 12348 7948 12400 7954
rect 12348 7890 12400 7896
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 13544 7472 13596 7478
rect 13544 7414 13596 7420
rect 13452 5568 13504 5574
rect 13452 5510 13504 5516
rect 11244 5364 11296 5370
rect 11244 5306 11296 5312
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 13464 1766 13492 5510
rect 13556 4146 13584 7414
rect 13636 7064 13688 7070
rect 13636 7006 13688 7012
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13648 1970 13676 7006
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 13832 2378 13860 5646
rect 14108 5438 14136 7890
rect 17130 6624 17186 6633
rect 17130 6559 17186 6568
rect 17040 5704 17092 5710
rect 17040 5646 17092 5652
rect 16672 5636 16724 5642
rect 16672 5578 16724 5584
rect 14096 5432 14148 5438
rect 14096 5374 14148 5380
rect 16578 5400 16634 5409
rect 16578 5335 16634 5344
rect 16592 5234 16620 5335
rect 16580 5228 16632 5234
rect 16580 5170 16632 5176
rect 16684 3777 16712 5578
rect 16948 5568 17000 5574
rect 16948 5510 17000 5516
rect 16856 4276 16908 4282
rect 16856 4218 16908 4224
rect 16670 3768 16726 3777
rect 16670 3703 16726 3712
rect 16672 2576 16724 2582
rect 16578 2544 16634 2553
rect 16672 2518 16724 2524
rect 16578 2479 16634 2488
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 13636 1964 13688 1970
rect 13636 1906 13688 1912
rect 13452 1760 13504 1766
rect 13452 1702 13504 1708
rect 16592 1494 16620 2479
rect 16580 1488 16632 1494
rect 16580 1430 16632 1436
rect 16684 1329 16712 2518
rect 16764 2100 16816 2106
rect 16764 2042 16816 2048
rect 16670 1320 16726 1329
rect 9864 1284 9916 1290
rect 9864 1226 9916 1232
rect 16580 1284 16632 1290
rect 16670 1255 16726 1264
rect 16580 1226 16632 1232
rect 16592 921 16620 1226
rect 16578 912 16634 921
rect 16578 847 16634 856
rect 8668 808 8720 814
rect 8668 750 8720 756
rect 8760 808 8812 814
rect 8760 750 8812 756
rect 9680 808 9732 814
rect 9680 750 9732 756
rect 3332 672 3384 678
rect 3332 614 3384 620
rect 8116 672 8168 678
rect 8116 614 8168 620
rect 5066 572 5374 581
rect 5066 570 5072 572
rect 5128 570 5152 572
rect 5208 570 5232 572
rect 5288 570 5312 572
rect 5368 570 5374 572
rect 5128 518 5130 570
rect 5310 518 5312 570
rect 5066 516 5072 518
rect 5128 516 5152 518
rect 5208 516 5232 518
rect 5288 516 5312 518
rect 5368 516 5374 518
rect 5066 507 5374 516
rect 16776 241 16804 2042
rect 16868 1737 16896 4218
rect 16960 2961 16988 5510
rect 17052 3369 17080 5646
rect 17144 4146 17172 6559
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 17038 3360 17094 3369
rect 17038 3295 17094 3304
rect 16946 2952 17002 2961
rect 16946 2887 17002 2896
rect 16854 1728 16910 1737
rect 16854 1663 16910 1672
rect 17236 1018 17264 11863
rect 20626 9888 20682 9897
rect 20626 9823 20682 9832
rect 19800 9444 19852 9450
rect 19800 9386 19852 9392
rect 19338 9072 19394 9081
rect 19338 9007 19394 9016
rect 19352 6866 19380 9007
rect 19706 8664 19762 8673
rect 19706 8599 19762 8608
rect 19616 8424 19668 8430
rect 19616 8366 19668 8372
rect 19430 7440 19486 7449
rect 19430 7375 19486 7384
rect 19340 6860 19392 6866
rect 19340 6802 19392 6808
rect 19444 6118 19472 7375
rect 19522 7032 19578 7041
rect 19522 6967 19578 6976
rect 19432 6112 19484 6118
rect 19432 6054 19484 6060
rect 19536 5438 19564 6967
rect 19628 6225 19656 8366
rect 19720 6322 19748 8599
rect 19708 6316 19760 6322
rect 19708 6258 19760 6264
rect 19614 6216 19670 6225
rect 19614 6151 19670 6160
rect 19812 5817 19840 9386
rect 20074 7848 20130 7857
rect 20074 7783 20130 7792
rect 19892 7132 19944 7138
rect 19892 7074 19944 7080
rect 19798 5808 19854 5817
rect 19798 5743 19854 5752
rect 19524 5432 19576 5438
rect 19524 5374 19576 5380
rect 17316 5092 17368 5098
rect 17316 5034 17368 5040
rect 17328 2145 17356 5034
rect 19904 5001 19932 7074
rect 20088 5370 20116 7783
rect 20168 7404 20220 7410
rect 20168 7346 20220 7352
rect 20076 5364 20128 5370
rect 20076 5306 20128 5312
rect 19890 4992 19946 5001
rect 19890 4927 19946 4936
rect 20180 4593 20208 7346
rect 20260 7064 20312 7070
rect 20260 7006 20312 7012
rect 20166 4584 20222 4593
rect 20166 4519 20222 4528
rect 20272 4185 20300 7006
rect 20258 4176 20314 4185
rect 20258 4111 20314 4120
rect 17314 2136 17370 2145
rect 17314 2071 17370 2080
rect 20640 2038 20668 9823
rect 20718 8256 20774 8265
rect 20718 8191 20774 8200
rect 20628 2032 20680 2038
rect 20628 1974 20680 1980
rect 17224 1012 17276 1018
rect 17224 954 17276 960
rect 20732 746 20760 8191
rect 22112 3534 22140 12543
rect 22100 3528 22152 3534
rect 22100 3470 22152 3476
rect 20720 740 20772 746
rect 20720 682 20772 688
rect 16762 232 16818 241
rect 16762 167 16818 176
<< via2 >>
rect 1214 11620 1270 11656
rect 1214 11600 1216 11620
rect 1216 11600 1268 11620
rect 1268 11600 1270 11620
rect 1950 10104 2006 10160
rect 1582 6296 1638 6352
rect 1490 6160 1546 6216
rect 2572 11994 2628 11996
rect 2652 11994 2708 11996
rect 2732 11994 2788 11996
rect 2812 11994 2868 11996
rect 2572 11942 2618 11994
rect 2618 11942 2628 11994
rect 2652 11942 2682 11994
rect 2682 11942 2694 11994
rect 2694 11942 2708 11994
rect 2732 11942 2746 11994
rect 2746 11942 2758 11994
rect 2758 11942 2788 11994
rect 2812 11942 2822 11994
rect 2822 11942 2868 11994
rect 2572 11940 2628 11942
rect 2652 11940 2708 11942
rect 2732 11940 2788 11942
rect 2812 11940 2868 11942
rect 2572 10906 2628 10908
rect 2652 10906 2708 10908
rect 2732 10906 2788 10908
rect 2812 10906 2868 10908
rect 2572 10854 2618 10906
rect 2618 10854 2628 10906
rect 2652 10854 2682 10906
rect 2682 10854 2694 10906
rect 2694 10854 2708 10906
rect 2732 10854 2746 10906
rect 2746 10854 2758 10906
rect 2758 10854 2788 10906
rect 2812 10854 2822 10906
rect 2822 10854 2868 10906
rect 2572 10852 2628 10854
rect 2652 10852 2708 10854
rect 2732 10852 2788 10854
rect 2812 10852 2868 10854
rect 2226 9832 2282 9888
rect 1858 4528 1914 4584
rect 2572 9818 2628 9820
rect 2652 9818 2708 9820
rect 2732 9818 2788 9820
rect 2812 9818 2868 9820
rect 2572 9766 2618 9818
rect 2618 9766 2628 9818
rect 2652 9766 2682 9818
rect 2682 9766 2694 9818
rect 2694 9766 2708 9818
rect 2732 9766 2746 9818
rect 2746 9766 2758 9818
rect 2758 9766 2788 9818
rect 2812 9766 2822 9818
rect 2822 9766 2868 9818
rect 2572 9764 2628 9766
rect 2652 9764 2708 9766
rect 2732 9764 2788 9766
rect 2812 9764 2868 9766
rect 2962 9424 3018 9480
rect 2572 8730 2628 8732
rect 2652 8730 2708 8732
rect 2732 8730 2788 8732
rect 2812 8730 2868 8732
rect 2572 8678 2618 8730
rect 2618 8678 2628 8730
rect 2652 8678 2682 8730
rect 2682 8678 2694 8730
rect 2694 8678 2708 8730
rect 2732 8678 2746 8730
rect 2746 8678 2758 8730
rect 2758 8678 2788 8730
rect 2812 8678 2822 8730
rect 2822 8678 2868 8730
rect 2572 8676 2628 8678
rect 2652 8676 2708 8678
rect 2732 8676 2788 8678
rect 2812 8676 2868 8678
rect 2572 7642 2628 7644
rect 2652 7642 2708 7644
rect 2732 7642 2788 7644
rect 2812 7642 2868 7644
rect 2572 7590 2618 7642
rect 2618 7590 2628 7642
rect 2652 7590 2682 7642
rect 2682 7590 2694 7642
rect 2694 7590 2708 7642
rect 2732 7590 2746 7642
rect 2746 7590 2758 7642
rect 2758 7590 2788 7642
rect 2812 7590 2822 7642
rect 2822 7590 2868 7642
rect 2572 7588 2628 7590
rect 2652 7588 2708 7590
rect 2732 7588 2788 7590
rect 2812 7588 2868 7590
rect 2572 6554 2628 6556
rect 2652 6554 2708 6556
rect 2732 6554 2788 6556
rect 2812 6554 2868 6556
rect 2572 6502 2618 6554
rect 2618 6502 2628 6554
rect 2652 6502 2682 6554
rect 2682 6502 2694 6554
rect 2694 6502 2708 6554
rect 2732 6502 2746 6554
rect 2746 6502 2758 6554
rect 2758 6502 2788 6554
rect 2812 6502 2822 6554
rect 2822 6502 2868 6554
rect 2572 6500 2628 6502
rect 2652 6500 2708 6502
rect 2732 6500 2788 6502
rect 2812 6500 2868 6502
rect 2962 6024 3018 6080
rect 2572 5466 2628 5468
rect 2652 5466 2708 5468
rect 2732 5466 2788 5468
rect 2812 5466 2868 5468
rect 2572 5414 2618 5466
rect 2618 5414 2628 5466
rect 2652 5414 2682 5466
rect 2682 5414 2694 5466
rect 2694 5414 2708 5466
rect 2732 5414 2746 5466
rect 2746 5414 2758 5466
rect 2758 5414 2788 5466
rect 2812 5414 2822 5466
rect 2822 5414 2868 5466
rect 2572 5412 2628 5414
rect 2652 5412 2708 5414
rect 2732 5412 2788 5414
rect 2812 5412 2868 5414
rect 2410 3984 2466 4040
rect 3238 8508 3240 8528
rect 3240 8508 3292 8528
rect 3292 8508 3294 8528
rect 3238 8472 3294 8508
rect 2572 1114 2628 1116
rect 2652 1114 2708 1116
rect 2732 1114 2788 1116
rect 2812 1114 2868 1116
rect 2572 1062 2618 1114
rect 2618 1062 2628 1114
rect 2652 1062 2682 1114
rect 2682 1062 2694 1114
rect 2694 1062 2708 1114
rect 2732 1062 2746 1114
rect 2746 1062 2758 1114
rect 2758 1062 2788 1114
rect 2812 1062 2822 1114
rect 2822 1062 2868 1114
rect 2572 1060 2628 1062
rect 2652 1060 2708 1062
rect 2732 1060 2788 1062
rect 2812 1060 2868 1062
rect 3882 10784 3938 10840
rect 3882 9832 3938 9888
rect 4158 9832 4214 9888
rect 3698 8200 3754 8256
rect 3422 2624 3478 2680
rect 3698 5752 3754 5808
rect 3974 8492 4030 8528
rect 3974 8472 3976 8492
rect 3976 8472 4028 8492
rect 4028 8472 4030 8492
rect 4250 8200 4306 8256
rect 3974 6024 4030 6080
rect 3974 5072 4030 5128
rect 3882 4004 3938 4040
rect 3882 3984 3884 4004
rect 3884 3984 3936 4004
rect 3936 3984 3938 4004
rect 3606 2488 3662 2544
rect 4250 2916 4306 2952
rect 4250 2896 4252 2916
rect 4252 2896 4304 2916
rect 4304 2896 4306 2916
rect 4710 10804 4766 10840
rect 4710 10784 4712 10804
rect 4712 10784 4764 10804
rect 4764 10784 4766 10804
rect 4526 5092 4582 5128
rect 4526 5072 4528 5092
rect 4528 5072 4580 5092
rect 4580 5072 4582 5092
rect 4618 4800 4674 4856
rect 4434 2760 4490 2816
rect 4526 2624 4582 2680
rect 5072 11450 5128 11452
rect 5152 11450 5208 11452
rect 5232 11450 5288 11452
rect 5312 11450 5368 11452
rect 5072 11398 5118 11450
rect 5118 11398 5128 11450
rect 5152 11398 5182 11450
rect 5182 11398 5194 11450
rect 5194 11398 5208 11450
rect 5232 11398 5246 11450
rect 5246 11398 5258 11450
rect 5258 11398 5288 11450
rect 5312 11398 5322 11450
rect 5322 11398 5368 11450
rect 5072 11396 5128 11398
rect 5152 11396 5208 11398
rect 5232 11396 5288 11398
rect 5312 11396 5368 11398
rect 5072 10362 5128 10364
rect 5152 10362 5208 10364
rect 5232 10362 5288 10364
rect 5312 10362 5368 10364
rect 5072 10310 5118 10362
rect 5118 10310 5128 10362
rect 5152 10310 5182 10362
rect 5182 10310 5194 10362
rect 5194 10310 5208 10362
rect 5232 10310 5246 10362
rect 5246 10310 5258 10362
rect 5258 10310 5288 10362
rect 5312 10310 5322 10362
rect 5322 10310 5368 10362
rect 5072 10308 5128 10310
rect 5152 10308 5208 10310
rect 5232 10308 5288 10310
rect 5312 10308 5368 10310
rect 5630 10548 5632 10568
rect 5632 10548 5684 10568
rect 5684 10548 5686 10568
rect 5630 10512 5686 10548
rect 5630 9424 5686 9480
rect 5072 9274 5128 9276
rect 5152 9274 5208 9276
rect 5232 9274 5288 9276
rect 5312 9274 5368 9276
rect 5072 9222 5118 9274
rect 5118 9222 5128 9274
rect 5152 9222 5182 9274
rect 5182 9222 5194 9274
rect 5194 9222 5208 9274
rect 5232 9222 5246 9274
rect 5246 9222 5258 9274
rect 5258 9222 5288 9274
rect 5312 9222 5322 9274
rect 5322 9222 5368 9274
rect 5072 9220 5128 9222
rect 5152 9220 5208 9222
rect 5232 9220 5288 9222
rect 5312 9220 5368 9222
rect 5354 8472 5410 8528
rect 5072 8186 5128 8188
rect 5152 8186 5208 8188
rect 5232 8186 5288 8188
rect 5312 8186 5368 8188
rect 5072 8134 5118 8186
rect 5118 8134 5128 8186
rect 5152 8134 5182 8186
rect 5182 8134 5194 8186
rect 5194 8134 5208 8186
rect 5232 8134 5246 8186
rect 5246 8134 5258 8186
rect 5258 8134 5288 8186
rect 5312 8134 5322 8186
rect 5322 8134 5368 8186
rect 5072 8132 5128 8134
rect 5152 8132 5208 8134
rect 5232 8132 5288 8134
rect 5312 8132 5368 8134
rect 5072 7098 5128 7100
rect 5152 7098 5208 7100
rect 5232 7098 5288 7100
rect 5312 7098 5368 7100
rect 5072 7046 5118 7098
rect 5118 7046 5128 7098
rect 5152 7046 5182 7098
rect 5182 7046 5194 7098
rect 5194 7046 5208 7098
rect 5232 7046 5246 7098
rect 5246 7046 5258 7098
rect 5258 7046 5288 7098
rect 5312 7046 5322 7098
rect 5322 7046 5368 7098
rect 5072 7044 5128 7046
rect 5152 7044 5208 7046
rect 5232 7044 5288 7046
rect 5312 7044 5368 7046
rect 5072 6010 5128 6012
rect 5152 6010 5208 6012
rect 5232 6010 5288 6012
rect 5312 6010 5368 6012
rect 5072 5958 5118 6010
rect 5118 5958 5128 6010
rect 5152 5958 5182 6010
rect 5182 5958 5194 6010
rect 5194 5958 5208 6010
rect 5232 5958 5246 6010
rect 5246 5958 5258 6010
rect 5258 5958 5288 6010
rect 5312 5958 5322 6010
rect 5322 5958 5368 6010
rect 5072 5956 5128 5958
rect 5152 5956 5208 5958
rect 5232 5956 5288 5958
rect 5312 5956 5368 5958
rect 5354 5772 5410 5808
rect 5354 5752 5356 5772
rect 5356 5752 5408 5772
rect 5408 5752 5410 5772
rect 5354 5072 5410 5128
rect 5072 4922 5128 4924
rect 5152 4922 5208 4924
rect 5232 4922 5288 4924
rect 5312 4922 5368 4924
rect 5072 4870 5118 4922
rect 5118 4870 5128 4922
rect 5152 4870 5182 4922
rect 5182 4870 5194 4922
rect 5194 4870 5208 4922
rect 5232 4870 5246 4922
rect 5246 4870 5258 4922
rect 5258 4870 5288 4922
rect 5312 4870 5322 4922
rect 5322 4870 5368 4922
rect 5072 4868 5128 4870
rect 5152 4868 5208 4870
rect 5232 4868 5288 4870
rect 5312 4868 5368 4870
rect 5262 4664 5318 4720
rect 4894 3612 4896 3632
rect 4896 3612 4948 3632
rect 4948 3612 4950 3632
rect 4894 3576 4950 3612
rect 5354 4120 5410 4176
rect 5072 3834 5128 3836
rect 5152 3834 5208 3836
rect 5232 3834 5288 3836
rect 5312 3834 5368 3836
rect 5072 3782 5118 3834
rect 5118 3782 5128 3834
rect 5152 3782 5182 3834
rect 5182 3782 5194 3834
rect 5194 3782 5208 3834
rect 5232 3782 5246 3834
rect 5246 3782 5258 3834
rect 5258 3782 5288 3834
rect 5312 3782 5322 3834
rect 5322 3782 5368 3834
rect 5072 3780 5128 3782
rect 5152 3780 5208 3782
rect 5232 3780 5288 3782
rect 5312 3780 5368 3782
rect 5446 2896 5502 2952
rect 4894 2760 4950 2816
rect 5072 2746 5128 2748
rect 5152 2746 5208 2748
rect 5232 2746 5288 2748
rect 5312 2746 5368 2748
rect 5072 2694 5118 2746
rect 5118 2694 5128 2746
rect 5152 2694 5182 2746
rect 5182 2694 5194 2746
rect 5194 2694 5208 2746
rect 5232 2694 5246 2746
rect 5246 2694 5258 2746
rect 5258 2694 5288 2746
rect 5312 2694 5322 2746
rect 5322 2694 5368 2746
rect 5072 2692 5128 2694
rect 5152 2692 5208 2694
rect 5232 2692 5288 2694
rect 5312 2692 5368 2694
rect 4894 2508 4950 2544
rect 4894 2488 4896 2508
rect 4896 2488 4948 2508
rect 4948 2488 4950 2508
rect 5722 8336 5778 8392
rect 22098 12552 22154 12608
rect 5630 7284 5632 7304
rect 5632 7284 5684 7304
rect 5684 7284 5686 7304
rect 5630 7248 5686 7284
rect 5722 6296 5778 6352
rect 5906 4528 5962 4584
rect 5814 4120 5870 4176
rect 5998 3984 6054 4040
rect 5072 1658 5128 1660
rect 5152 1658 5208 1660
rect 5232 1658 5288 1660
rect 5312 1658 5368 1660
rect 5072 1606 5118 1658
rect 5118 1606 5128 1658
rect 5152 1606 5182 1658
rect 5182 1606 5194 1658
rect 5194 1606 5208 1658
rect 5232 1606 5246 1658
rect 5246 1606 5258 1658
rect 5258 1606 5288 1658
rect 5312 1606 5322 1658
rect 5322 1606 5368 1658
rect 5072 1604 5128 1606
rect 5152 1604 5208 1606
rect 5232 1604 5288 1606
rect 5312 1604 5368 1606
rect 6642 9016 6698 9072
rect 6550 8472 6606 8528
rect 7572 11994 7628 11996
rect 7652 11994 7708 11996
rect 7732 11994 7788 11996
rect 7812 11994 7868 11996
rect 7572 11942 7618 11994
rect 7618 11942 7628 11994
rect 7652 11942 7682 11994
rect 7682 11942 7694 11994
rect 7694 11942 7708 11994
rect 7732 11942 7746 11994
rect 7746 11942 7758 11994
rect 7758 11942 7788 11994
rect 7812 11942 7822 11994
rect 7822 11942 7868 11994
rect 7572 11940 7628 11942
rect 7652 11940 7708 11942
rect 7732 11940 7788 11942
rect 7812 11940 7868 11942
rect 7572 10906 7628 10908
rect 7652 10906 7708 10908
rect 7732 10906 7788 10908
rect 7812 10906 7868 10908
rect 7572 10854 7618 10906
rect 7618 10854 7628 10906
rect 7652 10854 7682 10906
rect 7682 10854 7694 10906
rect 7694 10854 7708 10906
rect 7732 10854 7746 10906
rect 7746 10854 7758 10906
rect 7758 10854 7788 10906
rect 7812 10854 7822 10906
rect 7822 10854 7868 10906
rect 7572 10852 7628 10854
rect 7652 10852 7708 10854
rect 7732 10852 7788 10854
rect 7812 10852 7868 10854
rect 7470 10512 7526 10568
rect 7572 9818 7628 9820
rect 7652 9818 7708 9820
rect 7732 9818 7788 9820
rect 7812 9818 7868 9820
rect 7572 9766 7618 9818
rect 7618 9766 7628 9818
rect 7652 9766 7682 9818
rect 7682 9766 7694 9818
rect 7694 9766 7708 9818
rect 7732 9766 7746 9818
rect 7746 9766 7758 9818
rect 7758 9766 7788 9818
rect 7812 9766 7822 9818
rect 7822 9766 7868 9818
rect 7572 9764 7628 9766
rect 7652 9764 7708 9766
rect 7732 9764 7788 9766
rect 7812 9764 7868 9766
rect 7572 8730 7628 8732
rect 7652 8730 7708 8732
rect 7732 8730 7788 8732
rect 7812 8730 7868 8732
rect 7572 8678 7618 8730
rect 7618 8678 7628 8730
rect 7652 8678 7682 8730
rect 7682 8678 7694 8730
rect 7694 8678 7708 8730
rect 7732 8678 7746 8730
rect 7746 8678 7758 8730
rect 7758 8678 7788 8730
rect 7812 8678 7822 8730
rect 7822 8678 7868 8730
rect 7572 8676 7628 8678
rect 7652 8676 7708 8678
rect 7732 8676 7788 8678
rect 7812 8676 7868 8678
rect 7470 8336 7526 8392
rect 7572 7642 7628 7644
rect 7652 7642 7708 7644
rect 7732 7642 7788 7644
rect 7812 7642 7868 7644
rect 7572 7590 7618 7642
rect 7618 7590 7628 7642
rect 7652 7590 7682 7642
rect 7682 7590 7694 7642
rect 7694 7590 7708 7642
rect 7732 7590 7746 7642
rect 7746 7590 7758 7642
rect 7758 7590 7788 7642
rect 7812 7590 7822 7642
rect 7822 7590 7868 7642
rect 7572 7588 7628 7590
rect 7652 7588 7708 7590
rect 7732 7588 7788 7590
rect 7812 7588 7868 7590
rect 8114 7248 8170 7304
rect 8022 6568 8078 6624
rect 7572 6554 7628 6556
rect 7652 6554 7708 6556
rect 7732 6554 7788 6556
rect 7812 6554 7868 6556
rect 7572 6502 7618 6554
rect 7618 6502 7628 6554
rect 7652 6502 7682 6554
rect 7682 6502 7694 6554
rect 7694 6502 7708 6554
rect 7732 6502 7746 6554
rect 7746 6502 7758 6554
rect 7758 6502 7788 6554
rect 7812 6502 7822 6554
rect 7822 6502 7868 6554
rect 7572 6500 7628 6502
rect 7652 6500 7708 6502
rect 7732 6500 7788 6502
rect 7812 6500 7868 6502
rect 7838 6332 7840 6352
rect 7840 6332 7892 6352
rect 7892 6332 7894 6352
rect 7838 6296 7894 6332
rect 7572 5466 7628 5468
rect 7652 5466 7708 5468
rect 7732 5466 7788 5468
rect 7812 5466 7868 5468
rect 7572 5414 7618 5466
rect 7618 5414 7628 5466
rect 7652 5414 7682 5466
rect 7682 5414 7694 5466
rect 7694 5414 7708 5466
rect 7732 5414 7746 5466
rect 7746 5414 7758 5466
rect 7758 5414 7788 5466
rect 7812 5414 7822 5466
rect 7822 5414 7868 5466
rect 7572 5412 7628 5414
rect 7652 5412 7708 5414
rect 7732 5412 7788 5414
rect 7812 5412 7868 5414
rect 7470 4528 7526 4584
rect 7572 4378 7628 4380
rect 7652 4378 7708 4380
rect 7732 4378 7788 4380
rect 7812 4378 7868 4380
rect 7572 4326 7618 4378
rect 7618 4326 7628 4378
rect 7652 4326 7682 4378
rect 7682 4326 7694 4378
rect 7694 4326 7708 4378
rect 7732 4326 7746 4378
rect 7746 4326 7758 4378
rect 7758 4326 7788 4378
rect 7812 4326 7822 4378
rect 7822 4326 7868 4378
rect 7572 4324 7628 4326
rect 7652 4324 7708 4326
rect 7732 4324 7788 4326
rect 7812 4324 7868 4326
rect 7572 3290 7628 3292
rect 7652 3290 7708 3292
rect 7732 3290 7788 3292
rect 7812 3290 7868 3292
rect 7572 3238 7618 3290
rect 7618 3238 7628 3290
rect 7652 3238 7682 3290
rect 7682 3238 7694 3290
rect 7694 3238 7708 3290
rect 7732 3238 7746 3290
rect 7746 3238 7758 3290
rect 7758 3238 7788 3290
rect 7812 3238 7822 3290
rect 7822 3238 7868 3290
rect 7572 3236 7628 3238
rect 7652 3236 7708 3238
rect 7732 3236 7788 3238
rect 7812 3236 7868 3238
rect 7572 2202 7628 2204
rect 7652 2202 7708 2204
rect 7732 2202 7788 2204
rect 7812 2202 7868 2204
rect 7572 2150 7618 2202
rect 7618 2150 7628 2202
rect 7652 2150 7682 2202
rect 7682 2150 7694 2202
rect 7694 2150 7708 2202
rect 7732 2150 7746 2202
rect 7746 2150 7758 2202
rect 7758 2150 7788 2202
rect 7812 2150 7822 2202
rect 7822 2150 7868 2202
rect 7572 2148 7628 2150
rect 7652 2148 7708 2150
rect 7732 2148 7788 2150
rect 7812 2148 7868 2150
rect 8114 4684 8170 4720
rect 8114 4664 8116 4684
rect 8116 4664 8168 4684
rect 8168 4664 8170 4684
rect 8206 3984 8262 4040
rect 2594 856 2650 912
rect 7572 1114 7628 1116
rect 7652 1114 7708 1116
rect 7732 1114 7788 1116
rect 7812 1114 7868 1116
rect 7572 1062 7618 1114
rect 7618 1062 7628 1114
rect 7652 1062 7682 1114
rect 7682 1062 7694 1114
rect 7694 1062 7708 1114
rect 7732 1062 7746 1114
rect 7746 1062 7758 1114
rect 7758 1062 7788 1114
rect 7812 1062 7822 1114
rect 7822 1062 7868 1114
rect 7572 1060 7628 1062
rect 7652 1060 7708 1062
rect 7732 1060 7788 1062
rect 7812 1060 7868 1062
rect 9126 11600 9182 11656
rect 8574 7284 8576 7304
rect 8576 7284 8628 7304
rect 8628 7284 8630 7304
rect 8574 7248 8630 7284
rect 8574 6604 8576 6624
rect 8576 6604 8628 6624
rect 8628 6604 8630 6624
rect 8574 6568 8630 6604
rect 8758 6568 8814 6624
rect 8758 6296 8814 6352
rect 8942 7384 8998 7440
rect 8942 7248 8998 7304
rect 9126 7540 9182 7576
rect 9126 7520 9128 7540
rect 9128 7520 9180 7540
rect 9180 7520 9182 7540
rect 9126 7384 9182 7440
rect 9034 6432 9090 6488
rect 8942 6160 8998 6216
rect 9034 4120 9090 4176
rect 9586 8064 9642 8120
rect 9494 7928 9550 7984
rect 9310 7792 9366 7848
rect 9494 7828 9496 7848
rect 9496 7828 9548 7848
rect 9548 7828 9550 7848
rect 9494 7792 9550 7828
rect 9310 7520 9366 7576
rect 9586 7520 9642 7576
rect 9310 7248 9366 7304
rect 9586 7248 9642 7304
rect 9494 6840 9550 6896
rect 9402 6296 9458 6352
rect 9402 6060 9404 6080
rect 9404 6060 9456 6080
rect 9456 6060 9458 6080
rect 9402 6024 9458 6060
rect 9954 8372 9956 8392
rect 9956 8372 10008 8392
rect 10008 8372 10010 8392
rect 9954 8336 10010 8372
rect 9218 3460 9274 3496
rect 9218 3440 9220 3460
rect 9220 3440 9272 3460
rect 9272 3440 9274 3460
rect 8758 856 8814 912
rect 17222 11872 17278 11928
rect 16854 11464 16910 11520
rect 16762 11056 16818 11112
rect 16670 10648 16726 10704
rect 16578 9424 16634 9480
rect 16946 10240 17002 10296
rect 17130 6568 17186 6624
rect 16578 5344 16634 5400
rect 16670 3712 16726 3768
rect 16578 2488 16634 2544
rect 16670 1264 16726 1320
rect 16578 856 16634 912
rect 5072 570 5128 572
rect 5152 570 5208 572
rect 5232 570 5288 572
rect 5312 570 5368 572
rect 5072 518 5118 570
rect 5118 518 5128 570
rect 5152 518 5182 570
rect 5182 518 5194 570
rect 5194 518 5208 570
rect 5232 518 5246 570
rect 5246 518 5258 570
rect 5258 518 5288 570
rect 5312 518 5322 570
rect 5322 518 5368 570
rect 5072 516 5128 518
rect 5152 516 5208 518
rect 5232 516 5288 518
rect 5312 516 5368 518
rect 17038 3304 17094 3360
rect 16946 2896 17002 2952
rect 16854 1672 16910 1728
rect 20626 9832 20682 9888
rect 19338 9016 19394 9072
rect 19706 8608 19762 8664
rect 19430 7384 19486 7440
rect 19522 6976 19578 7032
rect 19614 6160 19670 6216
rect 20074 7792 20130 7848
rect 19798 5752 19854 5808
rect 19890 4936 19946 4992
rect 20166 4528 20222 4584
rect 20258 4120 20314 4176
rect 17314 2080 17370 2136
rect 20718 8200 20774 8256
rect 16762 176 16818 232
<< metal3 >>
rect 22093 12610 22159 12613
rect 22093 12608 22202 12610
rect 22093 12552 22098 12608
rect 22154 12552 22202 12608
rect 22093 12547 22202 12552
rect 22142 12368 22202 12547
rect 14000 12248 34000 12368
rect 2562 12000 2878 12001
rect 2562 11936 2568 12000
rect 2632 11936 2648 12000
rect 2712 11936 2728 12000
rect 2792 11936 2808 12000
rect 2872 11936 2878 12000
rect 2562 11935 2878 11936
rect 7562 12000 7878 12001
rect 7562 11936 7568 12000
rect 7632 11936 7648 12000
rect 7712 11936 7728 12000
rect 7792 11936 7808 12000
rect 7872 11936 7878 12000
rect 7562 11935 7878 11936
rect 14000 11928 34000 11960
rect 14000 11872 17222 11928
rect 17278 11872 34000 11928
rect 14000 11840 34000 11872
rect 1209 11658 1275 11661
rect 9121 11658 9187 11661
rect 1209 11656 9187 11658
rect 1209 11600 1214 11656
rect 1270 11600 9126 11656
rect 9182 11600 9187 11656
rect 1209 11598 9187 11600
rect 1209 11595 1275 11598
rect 9121 11595 9187 11598
rect 14000 11520 34000 11552
rect 14000 11464 16854 11520
rect 16910 11464 34000 11520
rect 5062 11456 5378 11457
rect 5062 11392 5068 11456
rect 5132 11392 5148 11456
rect 5212 11392 5228 11456
rect 5292 11392 5308 11456
rect 5372 11392 5378 11456
rect 14000 11432 34000 11464
rect 5062 11391 5378 11392
rect 14000 11112 34000 11144
rect 14000 11056 16762 11112
rect 16818 11056 34000 11112
rect 14000 11024 34000 11056
rect 2562 10912 2878 10913
rect 2562 10848 2568 10912
rect 2632 10848 2648 10912
rect 2712 10848 2728 10912
rect 2792 10848 2808 10912
rect 2872 10848 2878 10912
rect 2562 10847 2878 10848
rect 7562 10912 7878 10913
rect 7562 10848 7568 10912
rect 7632 10848 7648 10912
rect 7712 10848 7728 10912
rect 7792 10848 7808 10912
rect 7872 10848 7878 10912
rect 7562 10847 7878 10848
rect 3877 10842 3943 10845
rect 4705 10842 4771 10845
rect 3877 10840 4771 10842
rect 3877 10784 3882 10840
rect 3938 10784 4710 10840
rect 4766 10784 4771 10840
rect 3877 10782 4771 10784
rect 3877 10779 3943 10782
rect 4705 10779 4771 10782
rect 14000 10704 34000 10736
rect 14000 10648 16670 10704
rect 16726 10648 34000 10704
rect 14000 10616 34000 10648
rect 5625 10570 5691 10573
rect 7465 10570 7531 10573
rect 5625 10568 7531 10570
rect 5625 10512 5630 10568
rect 5686 10512 7470 10568
rect 7526 10512 7531 10568
rect 5625 10510 7531 10512
rect 5625 10507 5691 10510
rect 7465 10507 7531 10510
rect 5062 10368 5378 10369
rect 5062 10304 5068 10368
rect 5132 10304 5148 10368
rect 5212 10304 5228 10368
rect 5292 10304 5308 10368
rect 5372 10304 5378 10368
rect 5062 10303 5378 10304
rect 14000 10296 34000 10328
rect 14000 10240 16946 10296
rect 17002 10240 34000 10296
rect 14000 10208 34000 10240
rect 1945 10162 2011 10165
rect 1945 10160 2146 10162
rect 1945 10104 1950 10160
rect 2006 10104 2146 10160
rect 1945 10102 2146 10104
rect 1945 10099 2011 10102
rect 2086 9890 2146 10102
rect 2221 9890 2287 9893
rect 2086 9888 2287 9890
rect 2086 9832 2226 9888
rect 2282 9832 2287 9888
rect 2086 9830 2287 9832
rect 2221 9827 2287 9830
rect 3877 9890 3943 9893
rect 4153 9890 4219 9893
rect 3877 9888 4219 9890
rect 3877 9832 3882 9888
rect 3938 9832 4158 9888
rect 4214 9832 4219 9888
rect 3877 9830 4219 9832
rect 3877 9827 3943 9830
rect 4153 9827 4219 9830
rect 14000 9888 34000 9920
rect 14000 9832 20626 9888
rect 20682 9832 34000 9888
rect 2562 9824 2878 9825
rect 2562 9760 2568 9824
rect 2632 9760 2648 9824
rect 2712 9760 2728 9824
rect 2792 9760 2808 9824
rect 2872 9760 2878 9824
rect 2562 9759 2878 9760
rect 7562 9824 7878 9825
rect 7562 9760 7568 9824
rect 7632 9760 7648 9824
rect 7712 9760 7728 9824
rect 7792 9760 7808 9824
rect 7872 9760 7878 9824
rect 14000 9800 34000 9832
rect 7562 9759 7878 9760
rect 2957 9482 3023 9485
rect 5625 9482 5691 9485
rect 2957 9480 5691 9482
rect 2957 9424 2962 9480
rect 3018 9424 5630 9480
rect 5686 9424 5691 9480
rect 2957 9422 5691 9424
rect 2957 9419 3023 9422
rect 5625 9419 5691 9422
rect 14000 9480 34000 9512
rect 14000 9424 16578 9480
rect 16634 9424 34000 9480
rect 14000 9392 34000 9424
rect 5062 9280 5378 9281
rect 5062 9216 5068 9280
rect 5132 9216 5148 9280
rect 5212 9216 5228 9280
rect 5292 9216 5308 9280
rect 5372 9216 5378 9280
rect 5062 9215 5378 9216
rect 6637 9074 6703 9077
rect 7966 9074 7972 9076
rect 6637 9072 7972 9074
rect 6637 9016 6642 9072
rect 6698 9016 7972 9072
rect 6637 9014 7972 9016
rect 6637 9011 6703 9014
rect 7966 9012 7972 9014
rect 8036 9012 8042 9076
rect 14000 9072 34000 9104
rect 14000 9016 19338 9072
rect 19394 9016 34000 9072
rect 14000 8984 34000 9016
rect 2562 8736 2878 8737
rect 2562 8672 2568 8736
rect 2632 8672 2648 8736
rect 2712 8672 2728 8736
rect 2792 8672 2808 8736
rect 2872 8672 2878 8736
rect 2562 8671 2878 8672
rect 7562 8736 7878 8737
rect 7562 8672 7568 8736
rect 7632 8672 7648 8736
rect 7712 8672 7728 8736
rect 7792 8672 7808 8736
rect 7872 8672 7878 8736
rect 7562 8671 7878 8672
rect 14000 8664 34000 8696
rect 14000 8608 19706 8664
rect 19762 8608 34000 8664
rect 14000 8576 34000 8608
rect 3233 8532 3299 8533
rect 3182 8530 3188 8532
rect 3142 8470 3188 8530
rect 3252 8528 3299 8532
rect 3294 8472 3299 8528
rect 3182 8468 3188 8470
rect 3252 8468 3299 8472
rect 3233 8467 3299 8468
rect 3969 8530 4035 8533
rect 5349 8530 5415 8533
rect 3969 8528 5415 8530
rect 3969 8472 3974 8528
rect 4030 8472 5354 8528
rect 5410 8472 5415 8528
rect 3969 8470 5415 8472
rect 3969 8467 4035 8470
rect 5349 8467 5415 8470
rect 6545 8530 6611 8533
rect 9438 8530 9444 8532
rect 6545 8528 9444 8530
rect 6545 8472 6550 8528
rect 6606 8472 9444 8528
rect 6545 8470 9444 8472
rect 6545 8467 6611 8470
rect 9438 8468 9444 8470
rect 9508 8468 9514 8532
rect 5717 8394 5783 8397
rect 7465 8394 7531 8397
rect 9949 8394 10015 8397
rect 5717 8392 10015 8394
rect 5717 8336 5722 8392
rect 5778 8336 7470 8392
rect 7526 8336 9954 8392
rect 10010 8336 10015 8392
rect 5717 8334 10015 8336
rect 5717 8331 5783 8334
rect 7465 8331 7531 8334
rect 9949 8331 10015 8334
rect 3693 8258 3759 8261
rect 4245 8258 4311 8261
rect 3693 8256 4311 8258
rect 3693 8200 3698 8256
rect 3754 8200 4250 8256
rect 4306 8200 4311 8256
rect 3693 8198 4311 8200
rect 3693 8195 3759 8198
rect 4245 8195 4311 8198
rect 14000 8256 34000 8288
rect 14000 8200 20718 8256
rect 20774 8200 34000 8256
rect 5062 8192 5378 8193
rect 5062 8128 5068 8192
rect 5132 8128 5148 8192
rect 5212 8128 5228 8192
rect 5292 8128 5308 8192
rect 5372 8128 5378 8192
rect 14000 8168 34000 8200
rect 5062 8127 5378 8128
rect 9254 8060 9260 8124
rect 9324 8122 9330 8124
rect 9581 8122 9647 8125
rect 9324 8120 9647 8122
rect 9324 8064 9586 8120
rect 9642 8064 9647 8120
rect 9324 8062 9647 8064
rect 9324 8060 9330 8062
rect 9581 8059 9647 8062
rect 8334 7924 8340 7988
rect 8404 7986 8410 7988
rect 9489 7986 9555 7989
rect 8404 7984 9555 7986
rect 8404 7928 9494 7984
rect 9550 7928 9555 7984
rect 8404 7926 9555 7928
rect 8404 7924 8410 7926
rect 9489 7923 9555 7926
rect 9070 7788 9076 7852
rect 9140 7850 9146 7852
rect 9305 7850 9371 7853
rect 9489 7850 9555 7853
rect 9140 7848 9371 7850
rect 9140 7792 9310 7848
rect 9366 7792 9371 7848
rect 9140 7790 9371 7792
rect 9140 7788 9146 7790
rect 9305 7787 9371 7790
rect 9446 7848 9555 7850
rect 9446 7792 9494 7848
rect 9550 7792 9555 7848
rect 9446 7787 9555 7792
rect 14000 7848 34000 7880
rect 14000 7792 20074 7848
rect 20130 7792 34000 7848
rect 2562 7648 2878 7649
rect 2562 7584 2568 7648
rect 2632 7584 2648 7648
rect 2712 7584 2728 7648
rect 2792 7584 2808 7648
rect 2872 7584 2878 7648
rect 2562 7583 2878 7584
rect 7562 7648 7878 7649
rect 7562 7584 7568 7648
rect 7632 7584 7648 7648
rect 7712 7584 7728 7648
rect 7792 7584 7808 7648
rect 7872 7584 7878 7648
rect 7562 7583 7878 7584
rect 9121 7578 9187 7581
rect 9305 7578 9371 7581
rect 9121 7576 9371 7578
rect 9121 7520 9126 7576
rect 9182 7520 9310 7576
rect 9366 7520 9371 7576
rect 9121 7518 9371 7520
rect 9121 7515 9187 7518
rect 9305 7515 9371 7518
rect 8937 7442 9003 7445
rect 9121 7442 9187 7445
rect 8937 7440 9187 7442
rect 8937 7384 8942 7440
rect 8998 7384 9126 7440
rect 9182 7384 9187 7440
rect 8937 7382 9187 7384
rect 8937 7379 9003 7382
rect 9121 7379 9187 7382
rect 4470 7244 4476 7308
rect 4540 7306 4546 7308
rect 5625 7306 5691 7309
rect 8109 7308 8175 7309
rect 8109 7306 8156 7308
rect 4540 7304 5691 7306
rect 4540 7248 5630 7304
rect 5686 7248 5691 7304
rect 4540 7246 5691 7248
rect 8064 7304 8156 7306
rect 8064 7248 8114 7304
rect 8064 7246 8156 7248
rect 4540 7244 4546 7246
rect 5625 7243 5691 7246
rect 8109 7244 8156 7246
rect 8220 7244 8226 7308
rect 8569 7306 8635 7309
rect 8937 7306 9003 7309
rect 8569 7304 9003 7306
rect 8569 7248 8574 7304
rect 8630 7248 8942 7304
rect 8998 7248 9003 7304
rect 8569 7246 9003 7248
rect 8109 7243 8175 7244
rect 8569 7243 8635 7246
rect 8937 7243 9003 7246
rect 9305 7306 9371 7309
rect 9446 7306 9506 7787
rect 14000 7760 34000 7792
rect 9581 7578 9647 7581
rect 9581 7576 9690 7578
rect 9581 7520 9586 7576
rect 9642 7520 9690 7576
rect 9581 7515 9690 7520
rect 9630 7309 9690 7515
rect 14000 7440 34000 7472
rect 14000 7384 19430 7440
rect 19486 7384 34000 7440
rect 14000 7352 34000 7384
rect 9305 7304 9506 7306
rect 9305 7248 9310 7304
rect 9366 7248 9506 7304
rect 9305 7246 9506 7248
rect 9581 7304 9690 7309
rect 9581 7248 9586 7304
rect 9642 7248 9690 7304
rect 9581 7246 9690 7248
rect 9305 7243 9371 7246
rect 9581 7243 9647 7246
rect 5062 7104 5378 7105
rect 5062 7040 5068 7104
rect 5132 7040 5148 7104
rect 5212 7040 5228 7104
rect 5292 7040 5308 7104
rect 5372 7040 5378 7104
rect 5062 7039 5378 7040
rect 14000 7032 34000 7064
rect 14000 6976 19522 7032
rect 19578 6976 34000 7032
rect 14000 6944 34000 6976
rect 2998 6836 3004 6900
rect 3068 6898 3074 6900
rect 9489 6898 9555 6901
rect 3068 6896 9555 6898
rect 3068 6840 9494 6896
rect 9550 6840 9555 6896
rect 3068 6838 9555 6840
rect 3068 6836 3074 6838
rect 9489 6835 9555 6838
rect 8017 6626 8083 6629
rect 8569 6626 8635 6629
rect 8753 6626 8819 6629
rect 8017 6624 8635 6626
rect 8017 6568 8022 6624
rect 8078 6568 8574 6624
rect 8630 6568 8635 6624
rect 8017 6566 8635 6568
rect 8017 6563 8083 6566
rect 8569 6563 8635 6566
rect 8710 6624 8819 6626
rect 8710 6568 8758 6624
rect 8814 6568 8819 6624
rect 8710 6563 8819 6568
rect 14000 6624 34000 6656
rect 14000 6568 17130 6624
rect 17186 6568 34000 6624
rect 2562 6560 2878 6561
rect 2562 6496 2568 6560
rect 2632 6496 2648 6560
rect 2712 6496 2728 6560
rect 2792 6496 2808 6560
rect 2872 6496 2878 6560
rect 2562 6495 2878 6496
rect 7562 6560 7878 6561
rect 7562 6496 7568 6560
rect 7632 6496 7648 6560
rect 7712 6496 7728 6560
rect 7792 6496 7808 6560
rect 7872 6496 7878 6560
rect 7562 6495 7878 6496
rect 8710 6357 8770 6563
rect 14000 6536 34000 6568
rect 9029 6490 9095 6493
rect 8894 6488 9095 6490
rect 8894 6432 9034 6488
rect 9090 6432 9095 6488
rect 8894 6430 9095 6432
rect 1577 6354 1643 6357
rect 5717 6354 5783 6357
rect 7833 6354 7899 6357
rect 1577 6352 7899 6354
rect 1577 6296 1582 6352
rect 1638 6296 5722 6352
rect 5778 6296 7838 6352
rect 7894 6296 7899 6352
rect 1577 6294 7899 6296
rect 8710 6352 8819 6357
rect 8710 6296 8758 6352
rect 8814 6296 8819 6352
rect 8710 6294 8819 6296
rect 1577 6291 1643 6294
rect 5717 6291 5783 6294
rect 7833 6291 7899 6294
rect 8753 6291 8819 6294
rect 8894 6221 8954 6430
rect 9029 6427 9095 6430
rect 9254 6292 9260 6356
rect 9324 6354 9330 6356
rect 9397 6354 9463 6357
rect 9324 6352 9463 6354
rect 9324 6296 9402 6352
rect 9458 6296 9463 6352
rect 9324 6294 9463 6296
rect 9324 6292 9330 6294
rect 9397 6291 9463 6294
rect 1485 6218 1551 6221
rect 8334 6218 8340 6220
rect 1485 6216 8340 6218
rect 1485 6160 1490 6216
rect 1546 6160 8340 6216
rect 1485 6158 8340 6160
rect 1485 6155 1551 6158
rect 8334 6156 8340 6158
rect 8404 6156 8410 6220
rect 8894 6216 9003 6221
rect 8894 6160 8942 6216
rect 8998 6160 9003 6216
rect 8894 6158 9003 6160
rect 8937 6155 9003 6158
rect 14000 6216 34000 6248
rect 14000 6160 19614 6216
rect 19670 6160 34000 6216
rect 14000 6128 34000 6160
rect 2957 6082 3023 6085
rect 3182 6082 3188 6084
rect 2957 6080 3188 6082
rect 2957 6024 2962 6080
rect 3018 6024 3188 6080
rect 2957 6022 3188 6024
rect 2957 6019 3023 6022
rect 3182 6020 3188 6022
rect 3252 6082 3258 6084
rect 3969 6082 4035 6085
rect 3252 6080 4035 6082
rect 3252 6024 3974 6080
rect 4030 6024 4035 6080
rect 3252 6022 4035 6024
rect 3252 6020 3258 6022
rect 3969 6019 4035 6022
rect 9397 6084 9463 6085
rect 9397 6080 9444 6084
rect 9508 6082 9514 6084
rect 9397 6024 9402 6080
rect 9397 6020 9444 6024
rect 9508 6022 9554 6082
rect 9508 6020 9514 6022
rect 9397 6019 9463 6020
rect 5062 6016 5378 6017
rect 5062 5952 5068 6016
rect 5132 5952 5148 6016
rect 5212 5952 5228 6016
rect 5292 5952 5308 6016
rect 5372 5952 5378 6016
rect 5062 5951 5378 5952
rect 3693 5810 3759 5813
rect 5349 5810 5415 5813
rect 3693 5808 5415 5810
rect 3693 5752 3698 5808
rect 3754 5752 5354 5808
rect 5410 5752 5415 5808
rect 3693 5750 5415 5752
rect 3693 5747 3759 5750
rect 5349 5747 5415 5750
rect 14000 5808 34000 5840
rect 14000 5752 19798 5808
rect 19854 5752 34000 5808
rect 14000 5720 34000 5752
rect 2562 5472 2878 5473
rect 2562 5408 2568 5472
rect 2632 5408 2648 5472
rect 2712 5408 2728 5472
rect 2792 5408 2808 5472
rect 2872 5408 2878 5472
rect 2562 5407 2878 5408
rect 7562 5472 7878 5473
rect 7562 5408 7568 5472
rect 7632 5408 7648 5472
rect 7712 5408 7728 5472
rect 7792 5408 7808 5472
rect 7872 5408 7878 5472
rect 7562 5407 7878 5408
rect 14000 5400 34000 5432
rect 14000 5344 16578 5400
rect 16634 5344 34000 5400
rect 14000 5312 34000 5344
rect 3969 5130 4035 5133
rect 4521 5130 4587 5133
rect 3969 5128 4587 5130
rect 3969 5072 3974 5128
rect 4030 5072 4526 5128
rect 4582 5072 4587 5128
rect 3969 5070 4587 5072
rect 3969 5067 4035 5070
rect 4521 5067 4587 5070
rect 5349 5130 5415 5133
rect 5349 5128 5642 5130
rect 5349 5072 5354 5128
rect 5410 5072 5642 5128
rect 5349 5070 5642 5072
rect 5349 5067 5415 5070
rect 5062 4928 5378 4929
rect 5062 4864 5068 4928
rect 5132 4864 5148 4928
rect 5212 4864 5228 4928
rect 5292 4864 5308 4928
rect 5372 4864 5378 4928
rect 5062 4863 5378 4864
rect 4613 4860 4679 4861
rect 4613 4858 4660 4860
rect 4568 4856 4660 4858
rect 4568 4800 4618 4856
rect 4568 4798 4660 4800
rect 4613 4796 4660 4798
rect 4724 4796 4730 4860
rect 4613 4795 4679 4796
rect 5257 4722 5323 4725
rect 5582 4722 5642 5070
rect 14000 4992 34000 5024
rect 14000 4936 19890 4992
rect 19946 4936 34000 4992
rect 14000 4904 34000 4936
rect 5257 4720 5642 4722
rect 5257 4664 5262 4720
rect 5318 4664 5642 4720
rect 5257 4662 5642 4664
rect 8109 4722 8175 4725
rect 8334 4722 8340 4724
rect 8109 4720 8340 4722
rect 8109 4664 8114 4720
rect 8170 4664 8340 4720
rect 8109 4662 8340 4664
rect 5257 4659 5323 4662
rect 8109 4659 8175 4662
rect 8334 4660 8340 4662
rect 8404 4660 8410 4724
rect 1853 4586 1919 4589
rect 5901 4586 5967 4589
rect 1853 4584 5967 4586
rect 1853 4528 1858 4584
rect 1914 4528 5906 4584
rect 5962 4528 5967 4584
rect 1853 4526 5967 4528
rect 1853 4523 1919 4526
rect 5901 4523 5967 4526
rect 7465 4586 7531 4589
rect 9070 4586 9076 4588
rect 7465 4584 9076 4586
rect 7465 4528 7470 4584
rect 7526 4528 9076 4584
rect 7465 4526 9076 4528
rect 7465 4523 7531 4526
rect 9070 4524 9076 4526
rect 9140 4524 9146 4588
rect 14000 4584 34000 4616
rect 14000 4528 20166 4584
rect 20222 4528 34000 4584
rect 14000 4496 34000 4528
rect 7562 4384 7878 4385
rect 7562 4320 7568 4384
rect 7632 4320 7648 4384
rect 7712 4320 7728 4384
rect 7792 4320 7808 4384
rect 7872 4320 7878 4384
rect 7562 4319 7878 4320
rect 5349 4178 5415 4181
rect 5809 4178 5875 4181
rect 9029 4178 9095 4181
rect 5349 4176 9095 4178
rect 5349 4120 5354 4176
rect 5410 4120 5814 4176
rect 5870 4120 9034 4176
rect 9090 4120 9095 4176
rect 5349 4118 9095 4120
rect 5349 4115 5415 4118
rect 5809 4115 5875 4118
rect 9029 4115 9095 4118
rect 14000 4176 34000 4208
rect 14000 4120 20258 4176
rect 20314 4120 34000 4176
rect 14000 4088 34000 4120
rect 2405 4042 2471 4045
rect 2998 4042 3004 4044
rect 2405 4040 3004 4042
rect 2405 3984 2410 4040
rect 2466 3984 3004 4040
rect 2405 3982 3004 3984
rect 2405 3979 2471 3982
rect 2998 3980 3004 3982
rect 3068 3980 3074 4044
rect 3877 4042 3943 4045
rect 5993 4042 6059 4045
rect 8201 4044 8267 4045
rect 8150 4042 8156 4044
rect 3877 4040 6059 4042
rect 3877 3984 3882 4040
rect 3938 3984 5998 4040
rect 6054 3984 6059 4040
rect 3877 3982 6059 3984
rect 8110 3982 8156 4042
rect 8220 4040 8267 4044
rect 8262 3984 8267 4040
rect 3877 3979 3943 3982
rect 5993 3979 6059 3982
rect 8150 3980 8156 3982
rect 8220 3980 8267 3984
rect 8201 3979 8267 3980
rect 5062 3840 5378 3841
rect 5062 3776 5068 3840
rect 5132 3776 5148 3840
rect 5212 3776 5228 3840
rect 5292 3776 5308 3840
rect 5372 3776 5378 3840
rect 5062 3775 5378 3776
rect 14000 3768 34000 3800
rect 14000 3712 16670 3768
rect 16726 3712 34000 3768
rect 14000 3680 34000 3712
rect 4654 3572 4660 3636
rect 4724 3634 4730 3636
rect 4889 3634 4955 3637
rect 4724 3632 4955 3634
rect 4724 3576 4894 3632
rect 4950 3576 4955 3632
rect 4724 3574 4955 3576
rect 4724 3572 4730 3574
rect 4889 3571 4955 3574
rect 9213 3498 9279 3501
rect 2454 3496 9279 3498
rect 2454 3440 9218 3496
rect 9274 3440 9279 3496
rect 2454 3438 9279 3440
rect 2454 3400 2514 3438
rect 9213 3435 9279 3438
rect 14000 3360 34000 3392
rect 14000 3304 17038 3360
rect 17094 3304 34000 3360
rect 7562 3296 7878 3297
rect 7562 3232 7568 3296
rect 7632 3232 7648 3296
rect 7712 3232 7728 3296
rect 7792 3232 7808 3296
rect 7872 3232 7878 3296
rect 14000 3272 34000 3304
rect 7562 3231 7878 3232
rect 4245 2954 4311 2957
rect 4470 2954 4476 2956
rect 4245 2952 4476 2954
rect 4245 2896 4250 2952
rect 4306 2896 4476 2952
rect 4245 2894 4476 2896
rect 4245 2891 4311 2894
rect 4470 2892 4476 2894
rect 4540 2954 4546 2956
rect 5441 2954 5507 2957
rect 4540 2952 5507 2954
rect 4540 2896 5446 2952
rect 5502 2896 5507 2952
rect 4540 2894 5507 2896
rect 4540 2892 4546 2894
rect 5441 2891 5507 2894
rect 14000 2952 34000 2984
rect 14000 2896 16946 2952
rect 17002 2896 34000 2952
rect 14000 2864 34000 2896
rect 4429 2818 4495 2821
rect 4889 2818 4955 2821
rect 4429 2816 4955 2818
rect 4429 2760 4434 2816
rect 4490 2760 4894 2816
rect 4950 2760 4955 2816
rect 4429 2758 4955 2760
rect 4429 2755 4495 2758
rect 4889 2755 4955 2758
rect 5062 2752 5378 2753
rect 5062 2688 5068 2752
rect 5132 2688 5148 2752
rect 5212 2688 5228 2752
rect 5292 2688 5308 2752
rect 5372 2688 5378 2752
rect 5062 2687 5378 2688
rect 3417 2682 3483 2685
rect 4521 2682 4587 2685
rect 3417 2680 4587 2682
rect 3417 2624 3422 2680
rect 3478 2624 4526 2680
rect 4582 2624 4587 2680
rect 3417 2622 4587 2624
rect 3417 2619 3483 2622
rect 4521 2619 4587 2622
rect 3601 2546 3667 2549
rect 4889 2546 4955 2549
rect 3601 2544 4955 2546
rect 3601 2488 3606 2544
rect 3662 2488 4894 2544
rect 4950 2488 4955 2544
rect 3601 2486 4955 2488
rect 3601 2483 3667 2486
rect 4889 2483 4955 2486
rect 14000 2544 34000 2576
rect 14000 2488 16578 2544
rect 16634 2488 34000 2544
rect 14000 2456 34000 2488
rect 7562 2208 7878 2209
rect 7562 2144 7568 2208
rect 7632 2144 7648 2208
rect 7712 2144 7728 2208
rect 7792 2144 7808 2208
rect 7872 2144 7878 2208
rect 7562 2143 7878 2144
rect 14000 2136 34000 2168
rect 14000 2080 17314 2136
rect 17370 2080 34000 2136
rect 14000 2048 34000 2080
rect 14000 1728 34000 1760
rect 14000 1672 16854 1728
rect 16910 1672 34000 1728
rect 5062 1664 5378 1665
rect 5062 1600 5068 1664
rect 5132 1600 5148 1664
rect 5212 1600 5228 1664
rect 5292 1600 5308 1664
rect 5372 1600 5378 1664
rect 14000 1640 34000 1672
rect 5062 1599 5378 1600
rect 14000 1320 34000 1352
rect 14000 1264 16670 1320
rect 16726 1264 34000 1320
rect 14000 1232 34000 1264
rect 2562 1120 2878 1121
rect 2562 1056 2568 1120
rect 2632 1056 2648 1120
rect 2712 1056 2728 1120
rect 2792 1056 2808 1120
rect 2872 1056 2878 1120
rect 2562 1055 2878 1056
rect 7562 1120 7878 1121
rect 7562 1056 7568 1120
rect 7632 1056 7648 1120
rect 7712 1056 7728 1120
rect 7792 1056 7808 1120
rect 7872 1056 7878 1120
rect 7562 1055 7878 1056
rect 2589 914 2655 917
rect 7966 914 7972 916
rect 2589 912 7972 914
rect 2589 856 2594 912
rect 2650 856 7972 912
rect 2589 854 7972 856
rect 2589 851 2655 854
rect 7966 852 7972 854
rect 8036 914 8042 916
rect 8753 914 8819 917
rect 8036 912 8819 914
rect 8036 856 8758 912
rect 8814 856 8819 912
rect 8036 854 8819 856
rect 8036 852 8042 854
rect 8753 851 8819 854
rect 14000 912 34000 944
rect 14000 856 16578 912
rect 16634 856 34000 912
rect 14000 824 34000 856
rect 5062 576 5378 577
rect 5062 512 5068 576
rect 5132 512 5148 576
rect 5212 512 5228 576
rect 5292 512 5308 576
rect 5372 512 5378 576
rect 5062 511 5378 512
rect 14000 416 34000 536
rect 16806 237 16866 416
rect 16757 232 16866 237
rect 16757 176 16762 232
rect 16818 176 16866 232
rect 16757 174 16866 176
rect 16757 171 16823 174
<< via3 >>
rect 2568 11996 2632 12000
rect 2568 11940 2572 11996
rect 2572 11940 2628 11996
rect 2628 11940 2632 11996
rect 2568 11936 2632 11940
rect 2648 11996 2712 12000
rect 2648 11940 2652 11996
rect 2652 11940 2708 11996
rect 2708 11940 2712 11996
rect 2648 11936 2712 11940
rect 2728 11996 2792 12000
rect 2728 11940 2732 11996
rect 2732 11940 2788 11996
rect 2788 11940 2792 11996
rect 2728 11936 2792 11940
rect 2808 11996 2872 12000
rect 2808 11940 2812 11996
rect 2812 11940 2868 11996
rect 2868 11940 2872 11996
rect 2808 11936 2872 11940
rect 7568 11996 7632 12000
rect 7568 11940 7572 11996
rect 7572 11940 7628 11996
rect 7628 11940 7632 11996
rect 7568 11936 7632 11940
rect 7648 11996 7712 12000
rect 7648 11940 7652 11996
rect 7652 11940 7708 11996
rect 7708 11940 7712 11996
rect 7648 11936 7712 11940
rect 7728 11996 7792 12000
rect 7728 11940 7732 11996
rect 7732 11940 7788 11996
rect 7788 11940 7792 11996
rect 7728 11936 7792 11940
rect 7808 11996 7872 12000
rect 7808 11940 7812 11996
rect 7812 11940 7868 11996
rect 7868 11940 7872 11996
rect 7808 11936 7872 11940
rect 5068 11452 5132 11456
rect 5068 11396 5072 11452
rect 5072 11396 5128 11452
rect 5128 11396 5132 11452
rect 5068 11392 5132 11396
rect 5148 11452 5212 11456
rect 5148 11396 5152 11452
rect 5152 11396 5208 11452
rect 5208 11396 5212 11452
rect 5148 11392 5212 11396
rect 5228 11452 5292 11456
rect 5228 11396 5232 11452
rect 5232 11396 5288 11452
rect 5288 11396 5292 11452
rect 5228 11392 5292 11396
rect 5308 11452 5372 11456
rect 5308 11396 5312 11452
rect 5312 11396 5368 11452
rect 5368 11396 5372 11452
rect 5308 11392 5372 11396
rect 2568 10908 2632 10912
rect 2568 10852 2572 10908
rect 2572 10852 2628 10908
rect 2628 10852 2632 10908
rect 2568 10848 2632 10852
rect 2648 10908 2712 10912
rect 2648 10852 2652 10908
rect 2652 10852 2708 10908
rect 2708 10852 2712 10908
rect 2648 10848 2712 10852
rect 2728 10908 2792 10912
rect 2728 10852 2732 10908
rect 2732 10852 2788 10908
rect 2788 10852 2792 10908
rect 2728 10848 2792 10852
rect 2808 10908 2872 10912
rect 2808 10852 2812 10908
rect 2812 10852 2868 10908
rect 2868 10852 2872 10908
rect 2808 10848 2872 10852
rect 7568 10908 7632 10912
rect 7568 10852 7572 10908
rect 7572 10852 7628 10908
rect 7628 10852 7632 10908
rect 7568 10848 7632 10852
rect 7648 10908 7712 10912
rect 7648 10852 7652 10908
rect 7652 10852 7708 10908
rect 7708 10852 7712 10908
rect 7648 10848 7712 10852
rect 7728 10908 7792 10912
rect 7728 10852 7732 10908
rect 7732 10852 7788 10908
rect 7788 10852 7792 10908
rect 7728 10848 7792 10852
rect 7808 10908 7872 10912
rect 7808 10852 7812 10908
rect 7812 10852 7868 10908
rect 7868 10852 7872 10908
rect 7808 10848 7872 10852
rect 5068 10364 5132 10368
rect 5068 10308 5072 10364
rect 5072 10308 5128 10364
rect 5128 10308 5132 10364
rect 5068 10304 5132 10308
rect 5148 10364 5212 10368
rect 5148 10308 5152 10364
rect 5152 10308 5208 10364
rect 5208 10308 5212 10364
rect 5148 10304 5212 10308
rect 5228 10364 5292 10368
rect 5228 10308 5232 10364
rect 5232 10308 5288 10364
rect 5288 10308 5292 10364
rect 5228 10304 5292 10308
rect 5308 10364 5372 10368
rect 5308 10308 5312 10364
rect 5312 10308 5368 10364
rect 5368 10308 5372 10364
rect 5308 10304 5372 10308
rect 2568 9820 2632 9824
rect 2568 9764 2572 9820
rect 2572 9764 2628 9820
rect 2628 9764 2632 9820
rect 2568 9760 2632 9764
rect 2648 9820 2712 9824
rect 2648 9764 2652 9820
rect 2652 9764 2708 9820
rect 2708 9764 2712 9820
rect 2648 9760 2712 9764
rect 2728 9820 2792 9824
rect 2728 9764 2732 9820
rect 2732 9764 2788 9820
rect 2788 9764 2792 9820
rect 2728 9760 2792 9764
rect 2808 9820 2872 9824
rect 2808 9764 2812 9820
rect 2812 9764 2868 9820
rect 2868 9764 2872 9820
rect 2808 9760 2872 9764
rect 7568 9820 7632 9824
rect 7568 9764 7572 9820
rect 7572 9764 7628 9820
rect 7628 9764 7632 9820
rect 7568 9760 7632 9764
rect 7648 9820 7712 9824
rect 7648 9764 7652 9820
rect 7652 9764 7708 9820
rect 7708 9764 7712 9820
rect 7648 9760 7712 9764
rect 7728 9820 7792 9824
rect 7728 9764 7732 9820
rect 7732 9764 7788 9820
rect 7788 9764 7792 9820
rect 7728 9760 7792 9764
rect 7808 9820 7872 9824
rect 7808 9764 7812 9820
rect 7812 9764 7868 9820
rect 7868 9764 7872 9820
rect 7808 9760 7872 9764
rect 5068 9276 5132 9280
rect 5068 9220 5072 9276
rect 5072 9220 5128 9276
rect 5128 9220 5132 9276
rect 5068 9216 5132 9220
rect 5148 9276 5212 9280
rect 5148 9220 5152 9276
rect 5152 9220 5208 9276
rect 5208 9220 5212 9276
rect 5148 9216 5212 9220
rect 5228 9276 5292 9280
rect 5228 9220 5232 9276
rect 5232 9220 5288 9276
rect 5288 9220 5292 9276
rect 5228 9216 5292 9220
rect 5308 9276 5372 9280
rect 5308 9220 5312 9276
rect 5312 9220 5368 9276
rect 5368 9220 5372 9276
rect 5308 9216 5372 9220
rect 7972 9012 8036 9076
rect 2568 8732 2632 8736
rect 2568 8676 2572 8732
rect 2572 8676 2628 8732
rect 2628 8676 2632 8732
rect 2568 8672 2632 8676
rect 2648 8732 2712 8736
rect 2648 8676 2652 8732
rect 2652 8676 2708 8732
rect 2708 8676 2712 8732
rect 2648 8672 2712 8676
rect 2728 8732 2792 8736
rect 2728 8676 2732 8732
rect 2732 8676 2788 8732
rect 2788 8676 2792 8732
rect 2728 8672 2792 8676
rect 2808 8732 2872 8736
rect 2808 8676 2812 8732
rect 2812 8676 2868 8732
rect 2868 8676 2872 8732
rect 2808 8672 2872 8676
rect 7568 8732 7632 8736
rect 7568 8676 7572 8732
rect 7572 8676 7628 8732
rect 7628 8676 7632 8732
rect 7568 8672 7632 8676
rect 7648 8732 7712 8736
rect 7648 8676 7652 8732
rect 7652 8676 7708 8732
rect 7708 8676 7712 8732
rect 7648 8672 7712 8676
rect 7728 8732 7792 8736
rect 7728 8676 7732 8732
rect 7732 8676 7788 8732
rect 7788 8676 7792 8732
rect 7728 8672 7792 8676
rect 7808 8732 7872 8736
rect 7808 8676 7812 8732
rect 7812 8676 7868 8732
rect 7868 8676 7872 8732
rect 7808 8672 7872 8676
rect 3188 8528 3252 8532
rect 3188 8472 3238 8528
rect 3238 8472 3252 8528
rect 3188 8468 3252 8472
rect 9444 8468 9508 8532
rect 5068 8188 5132 8192
rect 5068 8132 5072 8188
rect 5072 8132 5128 8188
rect 5128 8132 5132 8188
rect 5068 8128 5132 8132
rect 5148 8188 5212 8192
rect 5148 8132 5152 8188
rect 5152 8132 5208 8188
rect 5208 8132 5212 8188
rect 5148 8128 5212 8132
rect 5228 8188 5292 8192
rect 5228 8132 5232 8188
rect 5232 8132 5288 8188
rect 5288 8132 5292 8188
rect 5228 8128 5292 8132
rect 5308 8188 5372 8192
rect 5308 8132 5312 8188
rect 5312 8132 5368 8188
rect 5368 8132 5372 8188
rect 5308 8128 5372 8132
rect 9260 8060 9324 8124
rect 8340 7924 8404 7988
rect 9076 7788 9140 7852
rect 2568 7644 2632 7648
rect 2568 7588 2572 7644
rect 2572 7588 2628 7644
rect 2628 7588 2632 7644
rect 2568 7584 2632 7588
rect 2648 7644 2712 7648
rect 2648 7588 2652 7644
rect 2652 7588 2708 7644
rect 2708 7588 2712 7644
rect 2648 7584 2712 7588
rect 2728 7644 2792 7648
rect 2728 7588 2732 7644
rect 2732 7588 2788 7644
rect 2788 7588 2792 7644
rect 2728 7584 2792 7588
rect 2808 7644 2872 7648
rect 2808 7588 2812 7644
rect 2812 7588 2868 7644
rect 2868 7588 2872 7644
rect 2808 7584 2872 7588
rect 7568 7644 7632 7648
rect 7568 7588 7572 7644
rect 7572 7588 7628 7644
rect 7628 7588 7632 7644
rect 7568 7584 7632 7588
rect 7648 7644 7712 7648
rect 7648 7588 7652 7644
rect 7652 7588 7708 7644
rect 7708 7588 7712 7644
rect 7648 7584 7712 7588
rect 7728 7644 7792 7648
rect 7728 7588 7732 7644
rect 7732 7588 7788 7644
rect 7788 7588 7792 7644
rect 7728 7584 7792 7588
rect 7808 7644 7872 7648
rect 7808 7588 7812 7644
rect 7812 7588 7868 7644
rect 7868 7588 7872 7644
rect 7808 7584 7872 7588
rect 4476 7244 4540 7308
rect 8156 7304 8220 7308
rect 8156 7248 8170 7304
rect 8170 7248 8220 7304
rect 8156 7244 8220 7248
rect 5068 7100 5132 7104
rect 5068 7044 5072 7100
rect 5072 7044 5128 7100
rect 5128 7044 5132 7100
rect 5068 7040 5132 7044
rect 5148 7100 5212 7104
rect 5148 7044 5152 7100
rect 5152 7044 5208 7100
rect 5208 7044 5212 7100
rect 5148 7040 5212 7044
rect 5228 7100 5292 7104
rect 5228 7044 5232 7100
rect 5232 7044 5288 7100
rect 5288 7044 5292 7100
rect 5228 7040 5292 7044
rect 5308 7100 5372 7104
rect 5308 7044 5312 7100
rect 5312 7044 5368 7100
rect 5368 7044 5372 7100
rect 5308 7040 5372 7044
rect 3004 6836 3068 6900
rect 2568 6556 2632 6560
rect 2568 6500 2572 6556
rect 2572 6500 2628 6556
rect 2628 6500 2632 6556
rect 2568 6496 2632 6500
rect 2648 6556 2712 6560
rect 2648 6500 2652 6556
rect 2652 6500 2708 6556
rect 2708 6500 2712 6556
rect 2648 6496 2712 6500
rect 2728 6556 2792 6560
rect 2728 6500 2732 6556
rect 2732 6500 2788 6556
rect 2788 6500 2792 6556
rect 2728 6496 2792 6500
rect 2808 6556 2872 6560
rect 2808 6500 2812 6556
rect 2812 6500 2868 6556
rect 2868 6500 2872 6556
rect 2808 6496 2872 6500
rect 7568 6556 7632 6560
rect 7568 6500 7572 6556
rect 7572 6500 7628 6556
rect 7628 6500 7632 6556
rect 7568 6496 7632 6500
rect 7648 6556 7712 6560
rect 7648 6500 7652 6556
rect 7652 6500 7708 6556
rect 7708 6500 7712 6556
rect 7648 6496 7712 6500
rect 7728 6556 7792 6560
rect 7728 6500 7732 6556
rect 7732 6500 7788 6556
rect 7788 6500 7792 6556
rect 7728 6496 7792 6500
rect 7808 6556 7872 6560
rect 7808 6500 7812 6556
rect 7812 6500 7868 6556
rect 7868 6500 7872 6556
rect 7808 6496 7872 6500
rect 9260 6292 9324 6356
rect 8340 6156 8404 6220
rect 3188 6020 3252 6084
rect 9444 6080 9508 6084
rect 9444 6024 9458 6080
rect 9458 6024 9508 6080
rect 9444 6020 9508 6024
rect 5068 6012 5132 6016
rect 5068 5956 5072 6012
rect 5072 5956 5128 6012
rect 5128 5956 5132 6012
rect 5068 5952 5132 5956
rect 5148 6012 5212 6016
rect 5148 5956 5152 6012
rect 5152 5956 5208 6012
rect 5208 5956 5212 6012
rect 5148 5952 5212 5956
rect 5228 6012 5292 6016
rect 5228 5956 5232 6012
rect 5232 5956 5288 6012
rect 5288 5956 5292 6012
rect 5228 5952 5292 5956
rect 5308 6012 5372 6016
rect 5308 5956 5312 6012
rect 5312 5956 5368 6012
rect 5368 5956 5372 6012
rect 5308 5952 5372 5956
rect 2568 5468 2632 5472
rect 2568 5412 2572 5468
rect 2572 5412 2628 5468
rect 2628 5412 2632 5468
rect 2568 5408 2632 5412
rect 2648 5468 2712 5472
rect 2648 5412 2652 5468
rect 2652 5412 2708 5468
rect 2708 5412 2712 5468
rect 2648 5408 2712 5412
rect 2728 5468 2792 5472
rect 2728 5412 2732 5468
rect 2732 5412 2788 5468
rect 2788 5412 2792 5468
rect 2728 5408 2792 5412
rect 2808 5468 2872 5472
rect 2808 5412 2812 5468
rect 2812 5412 2868 5468
rect 2868 5412 2872 5468
rect 2808 5408 2872 5412
rect 7568 5468 7632 5472
rect 7568 5412 7572 5468
rect 7572 5412 7628 5468
rect 7628 5412 7632 5468
rect 7568 5408 7632 5412
rect 7648 5468 7712 5472
rect 7648 5412 7652 5468
rect 7652 5412 7708 5468
rect 7708 5412 7712 5468
rect 7648 5408 7712 5412
rect 7728 5468 7792 5472
rect 7728 5412 7732 5468
rect 7732 5412 7788 5468
rect 7788 5412 7792 5468
rect 7728 5408 7792 5412
rect 7808 5468 7872 5472
rect 7808 5412 7812 5468
rect 7812 5412 7868 5468
rect 7868 5412 7872 5468
rect 7808 5408 7872 5412
rect 5068 4924 5132 4928
rect 5068 4868 5072 4924
rect 5072 4868 5128 4924
rect 5128 4868 5132 4924
rect 5068 4864 5132 4868
rect 5148 4924 5212 4928
rect 5148 4868 5152 4924
rect 5152 4868 5208 4924
rect 5208 4868 5212 4924
rect 5148 4864 5212 4868
rect 5228 4924 5292 4928
rect 5228 4868 5232 4924
rect 5232 4868 5288 4924
rect 5288 4868 5292 4924
rect 5228 4864 5292 4868
rect 5308 4924 5372 4928
rect 5308 4868 5312 4924
rect 5312 4868 5368 4924
rect 5368 4868 5372 4924
rect 5308 4864 5372 4868
rect 4660 4856 4724 4860
rect 4660 4800 4674 4856
rect 4674 4800 4724 4856
rect 4660 4796 4724 4800
rect 8340 4660 8404 4724
rect 9076 4524 9140 4588
rect 7568 4380 7632 4384
rect 7568 4324 7572 4380
rect 7572 4324 7628 4380
rect 7628 4324 7632 4380
rect 7568 4320 7632 4324
rect 7648 4380 7712 4384
rect 7648 4324 7652 4380
rect 7652 4324 7708 4380
rect 7708 4324 7712 4380
rect 7648 4320 7712 4324
rect 7728 4380 7792 4384
rect 7728 4324 7732 4380
rect 7732 4324 7788 4380
rect 7788 4324 7792 4380
rect 7728 4320 7792 4324
rect 7808 4380 7872 4384
rect 7808 4324 7812 4380
rect 7812 4324 7868 4380
rect 7868 4324 7872 4380
rect 7808 4320 7872 4324
rect 3004 3980 3068 4044
rect 8156 4040 8220 4044
rect 8156 3984 8206 4040
rect 8206 3984 8220 4040
rect 8156 3980 8220 3984
rect 5068 3836 5132 3840
rect 5068 3780 5072 3836
rect 5072 3780 5128 3836
rect 5128 3780 5132 3836
rect 5068 3776 5132 3780
rect 5148 3836 5212 3840
rect 5148 3780 5152 3836
rect 5152 3780 5208 3836
rect 5208 3780 5212 3836
rect 5148 3776 5212 3780
rect 5228 3836 5292 3840
rect 5228 3780 5232 3836
rect 5232 3780 5288 3836
rect 5288 3780 5292 3836
rect 5228 3776 5292 3780
rect 5308 3836 5372 3840
rect 5308 3780 5312 3836
rect 5312 3780 5368 3836
rect 5368 3780 5372 3836
rect 5308 3776 5372 3780
rect 4660 3572 4724 3636
rect 7568 3292 7632 3296
rect 7568 3236 7572 3292
rect 7572 3236 7628 3292
rect 7628 3236 7632 3292
rect 7568 3232 7632 3236
rect 7648 3292 7712 3296
rect 7648 3236 7652 3292
rect 7652 3236 7708 3292
rect 7708 3236 7712 3292
rect 7648 3232 7712 3236
rect 7728 3292 7792 3296
rect 7728 3236 7732 3292
rect 7732 3236 7788 3292
rect 7788 3236 7792 3292
rect 7728 3232 7792 3236
rect 7808 3292 7872 3296
rect 7808 3236 7812 3292
rect 7812 3236 7868 3292
rect 7868 3236 7872 3292
rect 7808 3232 7872 3236
rect 4476 2892 4540 2956
rect 5068 2748 5132 2752
rect 5068 2692 5072 2748
rect 5072 2692 5128 2748
rect 5128 2692 5132 2748
rect 5068 2688 5132 2692
rect 5148 2748 5212 2752
rect 5148 2692 5152 2748
rect 5152 2692 5208 2748
rect 5208 2692 5212 2748
rect 5148 2688 5212 2692
rect 5228 2748 5292 2752
rect 5228 2692 5232 2748
rect 5232 2692 5288 2748
rect 5288 2692 5292 2748
rect 5228 2688 5292 2692
rect 5308 2748 5372 2752
rect 5308 2692 5312 2748
rect 5312 2692 5368 2748
rect 5368 2692 5372 2748
rect 5308 2688 5372 2692
rect 7568 2204 7632 2208
rect 7568 2148 7572 2204
rect 7572 2148 7628 2204
rect 7628 2148 7632 2204
rect 7568 2144 7632 2148
rect 7648 2204 7712 2208
rect 7648 2148 7652 2204
rect 7652 2148 7708 2204
rect 7708 2148 7712 2204
rect 7648 2144 7712 2148
rect 7728 2204 7792 2208
rect 7728 2148 7732 2204
rect 7732 2148 7788 2204
rect 7788 2148 7792 2204
rect 7728 2144 7792 2148
rect 7808 2204 7872 2208
rect 7808 2148 7812 2204
rect 7812 2148 7868 2204
rect 7868 2148 7872 2204
rect 7808 2144 7872 2148
rect 5068 1660 5132 1664
rect 5068 1604 5072 1660
rect 5072 1604 5128 1660
rect 5128 1604 5132 1660
rect 5068 1600 5132 1604
rect 5148 1660 5212 1664
rect 5148 1604 5152 1660
rect 5152 1604 5208 1660
rect 5208 1604 5212 1660
rect 5148 1600 5212 1604
rect 5228 1660 5292 1664
rect 5228 1604 5232 1660
rect 5232 1604 5288 1660
rect 5288 1604 5292 1660
rect 5228 1600 5292 1604
rect 5308 1660 5372 1664
rect 5308 1604 5312 1660
rect 5312 1604 5368 1660
rect 5368 1604 5372 1660
rect 5308 1600 5372 1604
rect 2568 1116 2632 1120
rect 2568 1060 2572 1116
rect 2572 1060 2628 1116
rect 2628 1060 2632 1116
rect 2568 1056 2632 1060
rect 2648 1116 2712 1120
rect 2648 1060 2652 1116
rect 2652 1060 2708 1116
rect 2708 1060 2712 1116
rect 2648 1056 2712 1060
rect 2728 1116 2792 1120
rect 2728 1060 2732 1116
rect 2732 1060 2788 1116
rect 2788 1060 2792 1116
rect 2728 1056 2792 1060
rect 2808 1116 2872 1120
rect 2808 1060 2812 1116
rect 2812 1060 2868 1116
rect 2868 1060 2872 1116
rect 2808 1056 2872 1060
rect 7568 1116 7632 1120
rect 7568 1060 7572 1116
rect 7572 1060 7628 1116
rect 7628 1060 7632 1116
rect 7568 1056 7632 1060
rect 7648 1116 7712 1120
rect 7648 1060 7652 1116
rect 7652 1060 7708 1116
rect 7708 1060 7712 1116
rect 7648 1056 7712 1060
rect 7728 1116 7792 1120
rect 7728 1060 7732 1116
rect 7732 1060 7788 1116
rect 7788 1060 7792 1116
rect 7728 1056 7792 1060
rect 7808 1116 7872 1120
rect 7808 1060 7812 1116
rect 7812 1060 7868 1116
rect 7868 1060 7872 1116
rect 7808 1056 7872 1060
rect 7972 852 8036 916
rect 5068 572 5132 576
rect 5068 516 5072 572
rect 5072 516 5128 572
rect 5128 516 5132 572
rect 5068 512 5132 516
rect 5148 572 5212 576
rect 5148 516 5152 572
rect 5152 516 5208 572
rect 5208 516 5212 572
rect 5148 512 5212 516
rect 5228 572 5292 576
rect 5228 516 5232 572
rect 5232 516 5288 572
rect 5288 516 5292 572
rect 5228 512 5292 516
rect 5308 572 5372 576
rect 5308 516 5312 572
rect 5312 516 5368 572
rect 5368 516 5372 572
rect 5308 512 5372 516
<< metal4 >>
rect 2560 12000 2880 12016
rect 2560 11936 2568 12000
rect 2632 11936 2648 12000
rect 2712 11936 2728 12000
rect 2792 11936 2808 12000
rect 2872 11936 2880 12000
rect 2560 11598 2880 11936
rect 2560 11362 2602 11598
rect 2838 11362 2880 11598
rect 2560 10912 2880 11362
rect 2560 10848 2568 10912
rect 2632 10848 2648 10912
rect 2712 10848 2728 10912
rect 2792 10848 2808 10912
rect 2872 10848 2880 10912
rect 2560 9824 2880 10848
rect 2560 9760 2568 9824
rect 2632 9760 2648 9824
rect 2712 9760 2728 9824
rect 2792 9760 2808 9824
rect 2872 9760 2880 9824
rect 2560 8736 2880 9760
rect 2560 8672 2568 8736
rect 2632 8672 2648 8736
rect 2712 8672 2728 8736
rect 2792 8672 2808 8736
rect 2872 8672 2880 8736
rect 2560 8218 2880 8672
rect 3560 9266 3880 12016
rect 3560 9030 3602 9266
rect 3838 9030 3880 9266
rect 3187 8532 3253 8533
rect 3187 8468 3188 8532
rect 3252 8468 3253 8532
rect 3187 8467 3253 8468
rect 2560 7982 2602 8218
rect 2838 7982 2880 8218
rect 2560 7648 2880 7982
rect 2560 7584 2568 7648
rect 2632 7584 2648 7648
rect 2712 7584 2728 7648
rect 2792 7584 2808 7648
rect 2872 7584 2880 7648
rect 2560 6560 2880 7584
rect 3003 6900 3069 6901
rect 3003 6836 3004 6900
rect 3068 6836 3069 6900
rect 3003 6835 3069 6836
rect 2560 6496 2568 6560
rect 2632 6496 2648 6560
rect 2712 6496 2728 6560
rect 2792 6496 2808 6560
rect 2872 6496 2880 6560
rect 2560 5472 2880 6496
rect 2560 5408 2568 5472
rect 2632 5408 2648 5472
rect 2712 5408 2728 5472
rect 2792 5408 2808 5472
rect 2872 5408 2880 5472
rect 2560 4838 2880 5408
rect 2560 4602 2602 4838
rect 2838 4602 2880 4838
rect 1996 4196 2276 4238
rect 1996 3960 2018 4196
rect 2254 3960 2276 4196
rect 1996 3918 2276 3960
rect 1256 2506 1536 2548
rect 1256 2270 1278 2506
rect 1514 2270 1536 2506
rect 1256 2228 1536 2270
rect 2560 1458 2880 4602
rect 3006 4045 3066 6835
rect 3190 6085 3250 8467
rect 3187 6084 3253 6085
rect 3187 6020 3188 6084
rect 3252 6020 3253 6084
rect 3187 6019 3253 6020
rect 3560 5886 3880 9030
rect 5060 11456 5380 12016
rect 5060 11392 5068 11456
rect 5132 11392 5148 11456
rect 5212 11392 5228 11456
rect 5292 11392 5308 11456
rect 5372 11392 5380 11456
rect 5060 10368 5380 11392
rect 5060 10304 5068 10368
rect 5132 10304 5148 10368
rect 5212 10304 5228 10368
rect 5292 10304 5308 10368
rect 5372 10304 5380 10368
rect 5060 9908 5380 10304
rect 5060 9672 5102 9908
rect 5338 9672 5380 9908
rect 5060 9280 5380 9672
rect 5060 9216 5068 9280
rect 5132 9216 5148 9280
rect 5212 9216 5228 9280
rect 5292 9216 5308 9280
rect 5372 9216 5380 9280
rect 5060 8192 5380 9216
rect 5060 8128 5068 8192
rect 5132 8128 5148 8192
rect 5212 8128 5228 8192
rect 5292 8128 5308 8192
rect 5372 8128 5380 8192
rect 4475 7308 4541 7309
rect 4475 7244 4476 7308
rect 4540 7244 4541 7308
rect 4475 7243 4541 7244
rect 3560 5650 3602 5886
rect 3838 5650 3880 5886
rect 3003 4044 3069 4045
rect 3003 3980 3004 4044
rect 3068 3980 3069 4044
rect 3003 3979 3069 3980
rect 2560 1222 2602 1458
rect 2838 1222 2880 1458
rect 2560 1120 2880 1222
rect 2560 1056 2568 1120
rect 2632 1056 2648 1120
rect 2712 1056 2728 1120
rect 2792 1056 2808 1120
rect 2872 1056 2880 1120
rect 2560 496 2880 1056
rect 3560 2506 3880 5650
rect 4478 2957 4538 7243
rect 5060 7104 5380 8128
rect 5060 7040 5068 7104
rect 5132 7040 5148 7104
rect 5212 7040 5228 7104
rect 5292 7040 5308 7104
rect 5372 7040 5380 7104
rect 5060 6528 5380 7040
rect 5060 6292 5102 6528
rect 5338 6292 5380 6528
rect 5060 6016 5380 6292
rect 5060 5952 5068 6016
rect 5132 5952 5148 6016
rect 5212 5952 5228 6016
rect 5292 5952 5308 6016
rect 5372 5952 5380 6016
rect 5060 4928 5380 5952
rect 5060 4864 5068 4928
rect 5132 4864 5148 4928
rect 5212 4864 5228 4928
rect 5292 4864 5308 4928
rect 5372 4864 5380 4928
rect 4659 4860 4725 4861
rect 4659 4796 4660 4860
rect 4724 4796 4725 4860
rect 4659 4795 4725 4796
rect 4662 3637 4722 4795
rect 5060 3840 5380 4864
rect 5060 3776 5068 3840
rect 5132 3776 5148 3840
rect 5212 3776 5228 3840
rect 5292 3776 5308 3840
rect 5372 3776 5380 3840
rect 4659 3636 4725 3637
rect 4659 3572 4660 3636
rect 4724 3572 4725 3636
rect 4659 3571 4725 3572
rect 5060 3148 5380 3776
rect 4475 2956 4541 2957
rect 4475 2892 4476 2956
rect 4540 2892 4541 2956
rect 4475 2891 4541 2892
rect 5060 2912 5102 3148
rect 5338 2912 5380 3148
rect 3560 2270 3602 2506
rect 3838 2270 3880 2506
rect 3560 496 3880 2270
rect 5060 2752 5380 2912
rect 5060 2688 5068 2752
rect 5132 2688 5148 2752
rect 5212 2688 5228 2752
rect 5292 2688 5308 2752
rect 5372 2688 5380 2752
rect 5060 1664 5380 2688
rect 5060 1600 5068 1664
rect 5132 1600 5148 1664
rect 5212 1600 5228 1664
rect 5292 1600 5308 1664
rect 5372 1600 5380 1664
rect 5060 576 5380 1600
rect 5060 512 5068 576
rect 5132 512 5148 576
rect 5212 512 5228 576
rect 5292 512 5308 576
rect 5372 512 5380 576
rect 5060 496 5380 512
rect 6060 10956 6380 12016
rect 6060 10720 6102 10956
rect 6338 10720 6380 10956
rect 6060 7576 6380 10720
rect 6060 7340 6102 7576
rect 6338 7340 6380 7576
rect 6060 4196 6380 7340
rect 6060 3960 6102 4196
rect 6338 3960 6380 4196
rect 6060 496 6380 3960
rect 7560 12000 7880 12016
rect 7560 11936 7568 12000
rect 7632 11936 7648 12000
rect 7712 11936 7728 12000
rect 7792 11936 7808 12000
rect 7872 11936 7880 12000
rect 7560 11598 7880 11936
rect 7560 11362 7602 11598
rect 7838 11362 7880 11598
rect 7560 10912 7880 11362
rect 7560 10848 7568 10912
rect 7632 10848 7648 10912
rect 7712 10848 7728 10912
rect 7792 10848 7808 10912
rect 7872 10848 7880 10912
rect 7560 9824 7880 10848
rect 7560 9760 7568 9824
rect 7632 9760 7648 9824
rect 7712 9760 7728 9824
rect 7792 9760 7808 9824
rect 7872 9760 7880 9824
rect 7560 8736 7880 9760
rect 8560 9266 8880 12016
rect 7971 9076 8037 9077
rect 7971 9012 7972 9076
rect 8036 9012 8037 9076
rect 7971 9011 8037 9012
rect 8560 9030 8602 9266
rect 8838 9030 8880 9266
rect 7560 8672 7568 8736
rect 7632 8672 7648 8736
rect 7712 8672 7728 8736
rect 7792 8672 7808 8736
rect 7872 8672 7880 8736
rect 7560 8218 7880 8672
rect 7560 7982 7602 8218
rect 7838 7982 7880 8218
rect 7560 7648 7880 7982
rect 7560 7584 7568 7648
rect 7632 7584 7648 7648
rect 7712 7584 7728 7648
rect 7792 7584 7808 7648
rect 7872 7584 7880 7648
rect 7560 6560 7880 7584
rect 7560 6496 7568 6560
rect 7632 6496 7648 6560
rect 7712 6496 7728 6560
rect 7792 6496 7808 6560
rect 7872 6496 7880 6560
rect 7560 5472 7880 6496
rect 7560 5408 7568 5472
rect 7632 5408 7648 5472
rect 7712 5408 7728 5472
rect 7792 5408 7808 5472
rect 7872 5408 7880 5472
rect 7560 4838 7880 5408
rect 7560 4602 7602 4838
rect 7838 4602 7880 4838
rect 7560 4384 7880 4602
rect 7560 4320 7568 4384
rect 7632 4320 7648 4384
rect 7712 4320 7728 4384
rect 7792 4320 7808 4384
rect 7872 4320 7880 4384
rect 7560 3296 7880 4320
rect 7560 3232 7568 3296
rect 7632 3232 7648 3296
rect 7712 3232 7728 3296
rect 7792 3232 7808 3296
rect 7872 3232 7880 3296
rect 7560 2208 7880 3232
rect 7560 2144 7568 2208
rect 7632 2144 7648 2208
rect 7712 2144 7728 2208
rect 7792 2144 7808 2208
rect 7872 2144 7880 2208
rect 7560 1458 7880 2144
rect 7560 1222 7602 1458
rect 7838 1222 7880 1458
rect 7560 1120 7880 1222
rect 7560 1056 7568 1120
rect 7632 1056 7648 1120
rect 7712 1056 7728 1120
rect 7792 1056 7808 1120
rect 7872 1056 7880 1120
rect 7560 496 7880 1056
rect 7974 917 8034 9011
rect 8339 7988 8405 7989
rect 8339 7924 8340 7988
rect 8404 7924 8405 7988
rect 8339 7923 8405 7924
rect 8155 7308 8221 7309
rect 8155 7244 8156 7308
rect 8220 7244 8221 7308
rect 8155 7243 8221 7244
rect 8158 4045 8218 7243
rect 8342 6221 8402 7923
rect 8339 6220 8405 6221
rect 8339 6156 8340 6220
rect 8404 6156 8405 6220
rect 8339 6155 8405 6156
rect 8342 4725 8402 6155
rect 8560 5886 8880 9030
rect 9443 8532 9509 8533
rect 9443 8468 9444 8532
rect 9508 8468 9509 8532
rect 9443 8467 9509 8468
rect 9259 8124 9325 8125
rect 9259 8060 9260 8124
rect 9324 8060 9325 8124
rect 9259 8059 9325 8060
rect 9075 7852 9141 7853
rect 9075 7788 9076 7852
rect 9140 7788 9141 7852
rect 9075 7787 9141 7788
rect 8560 5650 8602 5886
rect 8838 5650 8880 5886
rect 8339 4724 8405 4725
rect 8339 4660 8340 4724
rect 8404 4660 8405 4724
rect 8339 4659 8405 4660
rect 8155 4044 8221 4045
rect 8155 3980 8156 4044
rect 8220 3980 8221 4044
rect 8155 3979 8221 3980
rect 8560 2506 8880 5650
rect 9078 4589 9138 7787
rect 9262 6357 9322 8059
rect 9259 6356 9325 6357
rect 9259 6292 9260 6356
rect 9324 6292 9325 6356
rect 9259 6291 9325 6292
rect 9446 6085 9506 8467
rect 9443 6084 9509 6085
rect 9443 6020 9444 6084
rect 9508 6020 9509 6084
rect 9443 6019 9509 6020
rect 9075 4588 9141 4589
rect 9075 4524 9076 4588
rect 9140 4524 9141 4588
rect 9075 4523 9141 4524
rect 8560 2270 8602 2506
rect 8838 2270 8880 2506
rect 7971 916 8037 917
rect 7971 852 7972 916
rect 8036 852 8037 916
rect 7971 851 8037 852
rect 8560 496 8880 2270
<< via4 >>
rect 2602 11362 2838 11598
rect 3602 9030 3838 9266
rect 2602 7982 2838 8218
rect 2602 4602 2838 4838
rect 2018 3960 2254 4196
rect 1278 2270 1514 2506
rect 5102 9672 5338 9908
rect 3602 5650 3838 5886
rect 2602 1222 2838 1458
rect 5102 6292 5338 6528
rect 5102 2912 5338 3148
rect 3602 2270 3838 2506
rect 6102 10720 6338 10956
rect 6102 7340 6338 7576
rect 6102 3960 6338 4196
rect 7602 11362 7838 11598
rect 8602 9030 8838 9266
rect 7602 7982 7838 8218
rect 7602 4602 7838 4838
rect 7602 1222 7838 1458
rect 8602 5650 8838 5886
rect 8602 2270 8838 2506
<< metal5 >>
rect 872 11598 10000 11640
rect 872 11362 2602 11598
rect 2838 11362 7602 11598
rect 7838 11362 10000 11598
rect 872 11320 10000 11362
rect 872 10956 10000 10998
rect 872 10720 6102 10956
rect 6338 10720 10000 10956
rect 872 10678 10000 10720
rect 872 9908 10000 9950
rect 872 9672 5102 9908
rect 5338 9672 10000 9908
rect 872 9630 10000 9672
rect 872 9266 10000 9308
rect 872 9030 3602 9266
rect 3838 9030 8602 9266
rect 8838 9030 10000 9266
rect 872 8988 10000 9030
rect 872 8218 10000 8260
rect 872 7982 2602 8218
rect 2838 7982 7602 8218
rect 7838 7982 10000 8218
rect 872 7940 10000 7982
rect 872 7576 10000 7618
rect 872 7340 6102 7576
rect 6338 7340 10000 7576
rect 872 7298 10000 7340
rect 872 6528 10000 6570
rect 872 6292 5102 6528
rect 5338 6292 10000 6528
rect 872 6250 10000 6292
rect 872 5886 10000 5928
rect 872 5650 3602 5886
rect 3838 5650 8602 5886
rect 8838 5650 10000 5886
rect 872 5608 10000 5650
rect 872 4838 10000 4880
rect 872 4602 2602 4838
rect 2838 4602 7602 4838
rect 7838 4602 10000 4838
rect 872 4560 10000 4602
rect 872 4196 10000 4238
rect 872 3960 2018 4196
rect 2254 3960 6102 4196
rect 6338 3960 10000 4196
rect 872 3918 10000 3960
rect 872 3148 10000 3190
rect 872 2912 5102 3148
rect 5338 2912 10000 3148
rect 872 2870 10000 2912
rect 872 2506 10000 2548
rect 872 2270 1278 2506
rect 1514 2270 3602 2506
rect 3838 2270 8602 2506
rect 8838 2270 10000 2506
rect 872 2228 10000 2270
rect 872 1458 10000 1500
rect 872 1222 2602 1458
rect 2838 1222 7602 1458
rect 7838 1222 10000 1458
rect 872 1180 10000 1222
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A_N $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 10120 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1666464484
transform 1 0 3772 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A_N
timestamp 1666464484
transform -1 0 3128 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1666464484
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A_N
timestamp 1666464484
transform 1 0 5428 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1666464484
transform 1 0 8832 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A_N
timestamp 1666464484
transform -1 0 6348 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__B
timestamp 1666464484
transform 1 0 6348 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__B
timestamp 1666464484
transform 1 0 9016 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__RESET_B
timestamp 1666464484
transform 1 0 8280 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__RESET_B
timestamp 1666464484
transform 1 0 5244 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__RESET_B
timestamp 1666464484
transform 1 0 3496 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__RESET_B
timestamp 1666464484
transform 1 0 6900 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_serial_clock_A
timestamp 1666464484
transform -1 0 3772 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_serial_load_A
timestamp 1666464484
transform 1 0 7360 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout42_A
timestamp 1666464484
transform -1 0 9660 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1666464484
transform -1 0 3312 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1666464484
transform -1 0 8924 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1666464484
transform -1 0 10120 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1666464484
transform -1 0 8924 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1666464484
transform -1 0 4140 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1666464484
transform -1 0 5888 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1666464484
transform -1 0 3496 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1666464484
transform -1 0 2944 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1666464484
transform -1 0 5888 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1666464484
transform -1 0 3864 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1666464484
transform -1 0 4048 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1666464484
transform -1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1666464484
transform -1 0 3496 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1666464484
transform -1 0 9844 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1666464484
transform -1 0 8648 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1666464484
transform -1 0 8832 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1666464484
transform 1 0 9844 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1666464484
transform -1 0 6072 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1666464484
transform 1 0 9200 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1666464484
transform -1 0 9292 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1196 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29
timestamp 1666464484
transform 1 0 3588 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1666464484
transform 1 0 6532 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87
timestamp 1666464484
transform 1 0 8924 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92
timestamp 1666464484
transform 1 0 9384 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99
timestamp 1666464484
transform 1 0 10028 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_30
timestamp 1666464484
transform 1 0 3680 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_99
timestamp 1666464484
transform 1 0 10028 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_99
timestamp 1666464484
transform 1 0 10028 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_50
timestamp 1666464484
transform 1 0 5520 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_84
timestamp 1666464484
transform 1 0 8648 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1666464484
transform 1 0 1196 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1666464484
transform 1 0 1196 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1666464484
transform 1 0 1196 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1666464484
transform 1 0 1196 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_99
timestamp 1666464484
transform 1 0 10028 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1666464484
transform 1 0 1196 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1666464484
transform 1 0 1196 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_60
timestamp 1666464484
transform 1 0 6440 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1666464484
transform 1 0 1196 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_57
timestamp 1666464484
transform 1 0 6164 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_99
timestamp 1666464484
transform 1 0 10028 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 920 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 10396 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 3036 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 10396 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 3036 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 10396 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 3036 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 10396 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 3036 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 10396 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 3036 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 10396 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 3036 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 10396 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 3036 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 10396 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 3036 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 10396 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 920 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 10396 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 920 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 10396 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 920 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 10396 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 920 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 10396 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 920 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 10396 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 920 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 10396 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 920 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 10396 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 920 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 10396 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 920 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 10396 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 920 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 10396 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 920 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 10396 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 920 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 10396 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3496 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1666464484
transform 1 0 6072 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1666464484
transform 1 0 8648 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1666464484
transform 1 0 8188 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1666464484
transform 1 0 5612 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1666464484
transform 1 0 8188 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1666464484
transform 1 0 5612 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1666464484
transform 1 0 8188 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1666464484
transform 1 0 5612 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1666464484
transform 1 0 8188 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1666464484
transform 1 0 5612 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1666464484
transform 1 0 3496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1666464484
transform 1 0 6072 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1666464484
transform 1 0 8648 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1666464484
transform 1 0 3496 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1666464484
transform 1 0 8648 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1666464484
transform 1 0 6072 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1666464484
transform 1 0 3496 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1666464484
transform 1 0 8648 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1666464484
transform 1 0 6072 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1666464484
transform 1 0 3496 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1666464484
transform 1 0 8648 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1666464484
transform 1 0 6072 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1666464484
transform 1 0 3496 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1666464484
transform 1 0 8648 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1666464484
transform 1 0 6072 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1666464484
transform 1 0 3496 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1666464484
transform 1 0 8648 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1666464484
transform 1 0 6072 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1666464484
transform 1 0 3496 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1666464484
transform 1 0 6072 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1666464484
transform 1 0 8648 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _058__1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5888 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _059__14
timestamp 1666464484
transform -1 0 1472 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _060_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9660 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _061_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9108 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _062_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9200 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _063_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 10120 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _064_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9476 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _065_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 8004 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _066_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 10120 0 1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_2  _067_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9292 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__or2_0  _068_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9476 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _069_
timestamp 1666464484
transform 1 0 6164 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__or2_0  _070_
timestamp 1666464484
transform 1 0 3588 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _071_
timestamp 1666464484
transform 1 0 1196 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__or2_0  _072_
timestamp 1666464484
transform 1 0 8740 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _073_
timestamp 1666464484
transform 1 0 6900 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__or2_0  _074_
timestamp 1666464484
transform 1 0 9200 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _075_
timestamp 1666464484
transform -1 0 9200 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__or2_0  _076_
timestamp 1666464484
transform 1 0 6900 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _077_
timestamp 1666464484
transform 1 0 3772 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__or2_0  _078_
timestamp 1666464484
transform 1 0 4324 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _079_
timestamp 1666464484
transform -1 0 1656 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__or2_0  _080_
timestamp 1666464484
transform 1 0 8740 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _081_
timestamp 1666464484
transform 1 0 1196 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__or2_0  _082_
timestamp 1666464484
transform 1 0 9660 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _083_
timestamp 1666464484
transform 1 0 7728 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__or2_0  _084_
timestamp 1666464484
transform -1 0 10120 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _085_
timestamp 1666464484
transform -1 0 10028 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__or2_0  _086_
timestamp 1666464484
transform -1 0 1656 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _087_
timestamp 1666464484
transform -1 0 9660 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__or2_0  _088_
timestamp 1666464484
transform 1 0 3772 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _089_
timestamp 1666464484
transform 1 0 3312 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__or2_0  _090_
timestamp 1666464484
transform 1 0 9660 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _091_
timestamp 1666464484
transform 1 0 5152 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__or2_0  _092_
timestamp 1666464484
transform 1 0 6164 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _093_
timestamp 1666464484
transform -1 0 7360 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _094__2
timestamp 1666464484
transform -1 0 4968 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _095__3
timestamp 1666464484
transform 1 0 3588 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _096__4
timestamp 1666464484
transform 1 0 9844 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _097__5
timestamp 1666464484
transform -1 0 5704 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _098__6
timestamp 1666464484
transform -1 0 4692 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _099__7
timestamp 1666464484
transform -1 0 5244 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _100__8
timestamp 1666464484
transform 1 0 4324 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _101__9
timestamp 1666464484
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _102__10
timestamp 1666464484
transform -1 0 8556 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _103__11
timestamp 1666464484
transform -1 0 4324 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _104__12
timestamp 1666464484
transform -1 0 5428 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _105__13
timestamp 1666464484
transform 1 0 5888 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_2  _106_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6072 0 1 10336
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _107_
timestamp 1666464484
transform 1 0 3496 0 -1 11424
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _108_
timestamp 1666464484
transform 1 0 6900 0 -1 8160
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _109_
timestamp 1666464484
transform -1 0 10120 0 -1 9248
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _110_
timestamp 1666464484
transform 1 0 3864 0 1 9248
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _111_
timestamp 1666464484
transform 1 0 3496 0 -1 8160
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _112_
timestamp 1666464484
transform 1 0 3496 0 -1 10336
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _113_
timestamp 1666464484
transform 1 0 7084 0 -1 7072
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _114_
timestamp 1666464484
transform 1 0 6992 0 -1 10336
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _115_
timestamp 1666464484
transform 1 0 7544 0 -1 11424
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _116_
timestamp 1666464484
transform 1 0 3496 0 -1 7072
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _117_
timestamp 1666464484
transform 1 0 4324 0 -1 4896
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _118_
timestamp 1666464484
transform 1 0 5428 0 1 5984
box -38 -48 2614 592
use sky130_fd_sc_hd__dfrtp_1  _119_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1656 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _120_
timestamp 1666464484
transform -1 0 5152 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _121_
timestamp 1666464484
transform -1 0 5152 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _122_
timestamp 1666464484
transform -1 0 3496 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _123_
timestamp 1666464484
transform 1 0 1656 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _124_
timestamp 1666464484
transform 1 0 1656 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _125_
timestamp 1666464484
transform 1 0 1656 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _126_
timestamp 1666464484
transform 1 0 3772 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _127_
timestamp 1666464484
transform 1 0 3588 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _128_
timestamp 1666464484
transform 1 0 1656 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _129_
timestamp 1666464484
transform 1 0 8280 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _130_
timestamp 1666464484
transform 1 0 4232 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _131_
timestamp 1666464484
transform 1 0 3312 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _132_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6532 0 1 9248
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_2  _133_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 9292 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1666464484
transform 1 0 1288 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _135_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4048 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _136_
timestamp 1666464484
transform -1 0 1656 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 4048 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_load
timestamp 1666464484
transform -1 0 6624 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_serial_clock
timestamp 1666464484
transform -1 0 3496 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_serial_load
timestamp 1666464484
transform -1 0 3496 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_serial_clock
timestamp 1666464484
transform 1 0 4232 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_serial_load
timestamp 1666464484
transform 1 0 1656 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  const_source $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 9292 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout40
timestamp 1666464484
transform -1 0 1656 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout41
timestamp 1666464484
transform 1 0 8740 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout42
timestamp 1666464484
transform -1 0 10028 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout43
timestamp 1666464484
transform 1 0 1288 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout44
timestamp 1666464484
transform -1 0 9660 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout45
timestamp 1666464484
transform -1 0 10028 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout46
timestamp 1666464484
transform 1 0 7360 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout47
timestamp 1666464484
transform 1 0 3680 0 1 1632
box -38 -48 406 592
use gpio_logic_high  gpio_logic_high
timestamp 0
transform 1 0 1196 0 1 1680
box -38 -48 1418 2768
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 6440 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1666464484
transform 1 0 3312 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1666464484
transform 1 0 1472 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1666464484
transform -1 0 6900 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1666464484
transform -1 0 5888 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1666464484
transform 1 0 3588 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1666464484
transform 1 0 3588 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1666464484
transform 1 0 6164 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1666464484
transform -1 0 9476 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1666464484
transform 1 0 6164 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1666464484
transform -1 0 9476 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1666464484
transform 1 0 6164 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1666464484
transform 1 0 6256 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1666464484
transform 1 0 3312 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1666464484
transform 1 0 1288 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1666464484
transform 1 0 8740 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1666464484
transform -1 0 2760 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1666464484
transform 1 0 4784 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1666464484
transform -1 0 6072 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1666464484
transform 1 0 1288 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1666464484
transform -1 0 1656 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1666464484
transform -1 0 6808 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1666464484
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1666464484
transform 1 0 3680 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1666464484
transform 1 0 5704 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1666464484
transform 1 0 3312 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1666464484
transform 1 0 9292 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1666464484
transform -1 0 8924 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1666464484
transform 1 0 8280 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1666464484
transform 1 0 1288 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1666464484
transform -1 0 4784 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1666464484
transform 1 0 2024 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1666464484
transform 1 0 7084 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_16  one_buffer $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 6164 0 -1 1632
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output21
timestamp 1666464484
transform -1 0 8648 0 1 544
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output22
timestamp 1666464484
transform 1 0 6164 0 -1 1632
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output23
timestamp 1666464484
transform -1 0 8096 0 1 1632
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output24
timestamp 1666464484
transform 1 0 6164 0 -1 2720
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output25
timestamp 1666464484
transform -1 0 8096 0 1 2720
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output26
timestamp 1666464484
transform -1 0 10120 0 1 1632
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output27
timestamp 1666464484
transform -1 0 8188 0 -1 3808
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output28
timestamp 1666464484
transform 1 0 8096 0 1 2720
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output29
timestamp 1666464484
transform 1 0 6072 0 1 4896
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output30
timestamp 1666464484
transform 1 0 8096 0 1 4896
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output31
timestamp 1666464484
transform -1 0 8648 0 1 7072
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output32
timestamp 1666464484
transform -1 0 8648 0 1 8160
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output33
timestamp 1666464484
transform -1 0 8648 0 -1 5984
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output34
timestamp 1666464484
transform -1 0 6624 0 1 7072
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output35
timestamp 1666464484
transform 1 0 4048 0 -1 9248
box -38 -48 2062 592
use sky130_fd_sc_hd__clkbuf_2  output36
timestamp 1666464484
transform -1 0 5520 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_16  output37
timestamp 1666464484
transform -1 0 8648 0 1 11424
box -38 -48 2062 592
use sky130_fd_sc_hd__clkbuf_2  output38
timestamp 1666464484
transform -1 0 2024 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_16  output39
timestamp 1666464484
transform -1 0 6072 0 1 11424
box -38 -48 2062 592
use sky130_fd_sc_hd__clkbuf_16  serial_clock_out_buffer
timestamp 1666464484
transform -1 0 3496 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  serial_load_out_buffer
timestamp 1666464484
transform 1 0 1656 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__macro_sparecell  spare_cell $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7452 0 1 3808
box -38 -48 2706 592
use sky130_fd_sc_hd__buf_16  zero_buffer
timestamp 1666464484
transform -1 0 6072 0 1 544
box -38 -48 2062 592
<< labels >>
flabel metal2 s 938 12200 994 13000 0 FreeSans 224 90 0 0 gpio_defaults[0]
port 0 nsew signal input
flabel metal2 s 5538 12200 5594 13000 0 FreeSans 224 90 0 0 gpio_defaults[10]
port 1 nsew signal input
flabel metal2 s 5998 12200 6054 13000 0 FreeSans 224 90 0 0 gpio_defaults[11]
port 2 nsew signal input
flabel metal2 s 6458 12200 6514 13000 0 FreeSans 224 90 0 0 gpio_defaults[12]
port 3 nsew signal input
flabel metal2 s 1398 12200 1454 13000 0 FreeSans 224 90 0 0 gpio_defaults[1]
port 4 nsew signal input
flabel metal2 s 1858 12200 1914 13000 0 FreeSans 224 90 0 0 gpio_defaults[2]
port 5 nsew signal input
flabel metal2 s 2318 12200 2374 13000 0 FreeSans 224 90 0 0 gpio_defaults[3]
port 6 nsew signal input
flabel metal2 s 2778 12200 2834 13000 0 FreeSans 224 90 0 0 gpio_defaults[4]
port 7 nsew signal input
flabel metal2 s 3238 12200 3294 13000 0 FreeSans 224 90 0 0 gpio_defaults[5]
port 8 nsew signal input
flabel metal2 s 3698 12200 3754 13000 0 FreeSans 224 90 0 0 gpio_defaults[6]
port 9 nsew signal input
flabel metal2 s 4158 12200 4214 13000 0 FreeSans 224 90 0 0 gpio_defaults[7]
port 10 nsew signal input
flabel metal2 s 4618 12200 4674 13000 0 FreeSans 224 90 0 0 gpio_defaults[8]
port 11 nsew signal input
flabel metal2 s 5078 12200 5134 13000 0 FreeSans 224 90 0 0 gpio_defaults[9]
port 12 nsew signal input
flabel metal3 s 14000 824 34000 944 0 FreeSans 480 0 0 0 mgmt_gpio_in
port 13 nsew signal tristate
flabel metal3 s 14000 1640 34000 1760 0 FreeSans 480 0 0 0 mgmt_gpio_oeb
port 14 nsew signal input
flabel metal3 s 14000 2048 34000 2168 0 FreeSans 480 0 0 0 mgmt_gpio_out
port 15 nsew signal input
flabel metal3 s 14000 1232 34000 1352 0 FreeSans 480 0 0 0 one
port 16 nsew signal tristate
flabel metal3 s 14000 2456 34000 2576 0 FreeSans 480 0 0 0 pad_gpio_ana_en
port 17 nsew signal tristate
flabel metal3 s 14000 2864 34000 2984 0 FreeSans 480 0 0 0 pad_gpio_ana_pol
port 18 nsew signal tristate
flabel metal3 s 14000 3272 34000 3392 0 FreeSans 480 0 0 0 pad_gpio_ana_sel
port 19 nsew signal tristate
flabel metal3 s 14000 3680 34000 3800 0 FreeSans 480 0 0 0 pad_gpio_dm[0]
port 20 nsew signal tristate
flabel metal3 s 14000 4088 34000 4208 0 FreeSans 480 0 0 0 pad_gpio_dm[1]
port 21 nsew signal tristate
flabel metal3 s 14000 4496 34000 4616 0 FreeSans 480 0 0 0 pad_gpio_dm[2]
port 22 nsew signal tristate
flabel metal3 s 14000 4904 34000 5024 0 FreeSans 480 0 0 0 pad_gpio_holdover
port 23 nsew signal tristate
flabel metal3 s 14000 5312 34000 5432 0 FreeSans 480 0 0 0 pad_gpio_ib_mode_sel
port 24 nsew signal tristate
flabel metal3 s 14000 5720 34000 5840 0 FreeSans 480 0 0 0 pad_gpio_in
port 25 nsew signal input
flabel metal3 s 14000 6128 34000 6248 0 FreeSans 480 0 0 0 pad_gpio_inenb
port 26 nsew signal tristate
flabel metal3 s 14000 6536 34000 6656 0 FreeSans 480 0 0 0 pad_gpio_out
port 27 nsew signal tristate
flabel metal3 s 14000 6944 34000 7064 0 FreeSans 480 0 0 0 pad_gpio_outenb
port 28 nsew signal tristate
flabel metal3 s 14000 7352 34000 7472 0 FreeSans 480 0 0 0 pad_gpio_slow_sel
port 29 nsew signal tristate
flabel metal3 s 14000 7760 34000 7880 0 FreeSans 480 0 0 0 pad_gpio_vtrip_sel
port 30 nsew signal tristate
flabel metal3 s 14000 8168 34000 8288 0 FreeSans 480 0 0 0 resetn
port 31 nsew signal input
flabel metal3 s 14000 8576 34000 8696 0 FreeSans 480 0 0 0 resetn_out
port 32 nsew signal tristate
flabel metal3 s 14000 8984 34000 9104 0 FreeSans 480 0 0 0 serial_clock
port 33 nsew signal input
flabel metal3 s 14000 9392 34000 9512 0 FreeSans 480 0 0 0 serial_clock_out
port 34 nsew signal tristate
flabel metal3 s 14000 9800 34000 9920 0 FreeSans 480 0 0 0 serial_data_in
port 35 nsew signal input
flabel metal3 s 14000 10208 34000 10328 0 FreeSans 480 0 0 0 serial_data_out
port 36 nsew signal tristate
flabel metal3 s 14000 10616 34000 10736 0 FreeSans 480 0 0 0 serial_load
port 37 nsew signal input
flabel metal3 s 14000 11024 34000 11144 0 FreeSans 480 0 0 0 serial_load_out
port 38 nsew signal tristate
flabel metal3 s 14000 11432 34000 11552 0 FreeSans 480 0 0 0 user_gpio_in
port 39 nsew signal tristate
flabel metal3 s 14000 11840 34000 11960 0 FreeSans 480 0 0 0 user_gpio_oeb
port 40 nsew signal input
flabel metal3 s 14000 12248 34000 12368 0 FreeSans 480 0 0 0 user_gpio_out
port 41 nsew signal input
flabel metal4 s 2560 496 2880 12016 0 FreeSans 1920 90 0 0 vccd
port 42 nsew power bidirectional
flabel metal4 s 7560 496 7880 12016 0 FreeSans 1920 90 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 1180 10000 1500 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 4560 10000 4880 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 7940 10000 8260 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 11320 10000 11640 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal4 s 3560 496 3880 12016 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 8560 496 8880 12016 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 872 2228 10000 2548 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 872 5608 10000 5928 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 872 8988 10000 9308 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 5060 496 5380 12016 0 FreeSans 1920 90 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 2870 10000 3190 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 6250 10000 6570 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 9630 10000 9950 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal4 s 6060 496 6380 12016 0 FreeSans 1920 90 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal5 s 872 3918 10000 4238 0 FreeSans 2560 0 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal5 s 872 7298 10000 7618 0 FreeSans 2560 0 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal5 s 872 10678 10000 10998 0 FreeSans 2560 0 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal3 s 14000 416 34000 536 0 FreeSans 480 0 0 0 zero
port 46 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 34000 13000
<< end >>
