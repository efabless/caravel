* NGSPICE file created from housekeeping.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtn_1 abstract view
.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_2 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_2 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4bb_1 abstract view
.subckt sky130_fd_sc_hd__nand4bb_1 A_N B_N C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_2 abstract view
.subckt sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

.subckt housekeeping VGND VPWR debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oeb
+ pad_flash_csb pad_flash_csb_oeb pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ieb
+ pad_flash_io0_oeb pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ieb pad_flash_io1_oeb
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out[0] pwr_ctrl_out[1]
+ pwr_ctrl_out[2] pwr_ctrl_out[3] qspi_enabled reset ser_rx ser_tx serial_clock serial_data_1
+ serial_data_2 serial_load serial_resetn spi_csb spi_enabled spi_sck spi_sdi spi_sdo
+ spi_sdoenb spimemio_flash_clk spimemio_flash_csb spimemio_flash_io0_di spimemio_flash_io0_do
+ spimemio_flash_io0_oeb spimemio_flash_io1_di spimemio_flash_io1_do spimemio_flash_io1_oeb
+ spimemio_flash_io2_di spimemio_flash_io2_do spimemio_flash_io2_oeb spimemio_flash_io3_di
+ spimemio_flash_io3_do spimemio_flash_io3_oeb trap uart_enabled user_clock usr1_vcc_pwrgood
+ usr1_vdd_pwrgood usr2_vcc_pwrgood usr2_vdd_pwrgood wb_ack_o wb_adr_i[0] wb_adr_i[10]
+ wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17]
+ wb_adr_i[18] wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23]
+ wb_adr_i[24] wb_adr_i[25] wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2]
+ wb_adr_i[30] wb_adr_i[31] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7]
+ wb_adr_i[8] wb_adr_i[9] wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11]
+ wb_dat_i[12] wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18]
+ wb_dat_i[19] wb_dat_i[1] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24]
+ wb_dat_i[25] wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30]
+ wb_dat_i[31] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8]
+ wb_dat_i[9] wb_dat_o[0] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14]
+ wb_dat_o[15] wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20]
+ wb_dat_o[21] wb_dat_o[22] wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27]
+ wb_dat_o[28] wb_dat_o[29] wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4]
+ wb_dat_o[5] wb_dat_o[6] wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0]
+ wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] wb_stb_i wb_we_i
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6914_ _7125_/CLK _6914_/D fanout454/X VGND VGND VPWR VPWR _6914_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6845_ _7018_/CLK _6845_/D fanout460/X VGND VGND VPWR VPWR _6845_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_52_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6776_ _6658_/CLK _6776_/D _6428_/X VGND VGND VPWR VPWR _6776_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_168_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3988_ _3988_/A _5220_/C VGND VGND VPWR VPWR _3999_/S sky130_fd_sc_hd__and2_4
X_5727_ _5727_/A _5727_/B _5727_/C _5727_/D VGND VGND VPWR VPWR _5727_/Y sky130_fd_sc_hd__nor4_2
XFILLER_182_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5658_ _5689_/A _5686_/B _5689_/C VGND VGND VPWR VPWR _5658_/X sky130_fd_sc_hd__and3b_4
XFILLER_164_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4609_ _5100_/C _4609_/B _4609_/C _4609_/D VGND VGND VPWR VPWR _4614_/B sky130_fd_sc_hd__and4_1
XFILLER_190_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5589_ _6490_/Q _6492_/Q VGND VGND VPWR VPWR _5589_/Y sky130_fd_sc_hd__nor2_1
Xhold340 hold340/A VGND VGND VPWR VPWR hold340/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold351 hold961/X VGND VGND VPWR VPWR hold962/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold362 hold362/A VGND VGND VPWR VPWR hold362/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold373 _5244_/X VGND VGND VPWR VPWR _6836_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold384 hold384/A VGND VGND VPWR VPWR _6515_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold395 hold395/A VGND VGND VPWR VPWR hold395/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1040 hold24/X VGND VGND VPWR VPWR _3302_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1051 _7123_/Q VGND VGND VPWR VPWR hold396/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1062 _3302_/X VGND VGND VPWR VPWR hold25/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1073 _5261_/X VGND VGND VPWR VPWR _6851_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1084 _5423_/X VGND VGND VPWR VPWR _6995_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_172_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_202 _5985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1095 hold403/X VGND VGND VPWR VPWR _5585_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4960_ _4552_/B _5033_/B _4782_/X VGND VGND VPWR VPWR _4961_/D sky130_fd_sc_hd__a21oi_2
XFILLER_52_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3911_ _5643_/A _3911_/B VGND VGND VPWR VPWR _3912_/B sky130_fd_sc_hd__and2b_1
X_4891_ _5114_/A _5102_/A _5130_/A _5103_/A VGND VGND VPWR VPWR _4892_/D sky130_fd_sc_hd__and4_1
X_6630_ _6749_/CLK _6630_/D fanout439/X VGND VGND VPWR VPWR _6630_/Q sky130_fd_sc_hd__dfrtp_4
X_3842_ _3182_/Y _3846_/S _3840_/B _6461_/Q VGND VGND VPWR VPWR _3842_/X sky130_fd_sc_hd__o211a_1
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6561_ _6568_/CLK _6561_/D VGND VGND VPWR VPWR _6561_/Q sky130_fd_sc_hd__dfxtp_1
X_3773_ input93/X _5226_/A _3303_/X hold40/A _6845_/Q VGND VGND VPWR VPWR _3773_/X
+ sky130_fd_sc_hd__a32o_1
X_5512_ _5512_/A0 _5575_/A1 _5514_/S VGND VGND VPWR VPWR _7074_/D sky130_fd_sc_hd__mux2_1
X_6492_ _7203_/CLK _6492_/D _6399_/A VGND VGND VPWR VPWR _6492_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_8_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5443_ _5443_/A _5551_/B VGND VGND VPWR VPWR _5451_/S sky130_fd_sc_hd__and2_4
XFILLER_172_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5374_ _5374_/A0 _5572_/A1 _5379_/S VGND VGND VPWR VPWR _6951_/D sky130_fd_sc_hd__mux2_1
X_7113_ _7113_/CLK _7113_/D fanout472/X VGND VGND VPWR VPWR _7113_/Q sky130_fd_sc_hd__dfrtp_4
X_4325_ _4325_/A0 _5187_/A1 _4327_/S VGND VGND VPWR VPWR _4325_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7044_ _7131_/CLK hold57/X fanout469/X VGND VGND VPWR VPWR _7044_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_141_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4256_ _4256_/A _5229_/C VGND VGND VPWR VPWR _4261_/S sky130_fd_sc_hd__and2_4
XFILLER_86_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3207_ _7096_/Q VGND VGND VPWR VPWR _3207_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4187_ _4187_/A0 _5196_/A1 _4187_/S VGND VGND VPWR VPWR _4187_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6828_ _7097_/CLK hold92/X fanout468/X VGND VGND VPWR VPWR _6828_/Q sky130_fd_sc_hd__dfrtp_2
X_6759_ _6759_/CLK _6759_/D _6426_/A VGND VGND VPWR VPWR _6759_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_183_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold170 _7198_/Q VGND VGND VPWR VPWR hold170/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold181 hold181/A VGND VGND VPWR VPWR hold181/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold192 hold192/A VGND VGND VPWR VPWR wb_dat_o[24] sky130_fd_sc_hd__buf_12
XFILLER_105_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4110_ _3675_/Y hold869/A _4115_/S VGND VGND VPWR VPWR _6563_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5090_ _4950_/X _4769_/Y _5090_/C _5090_/D VGND VGND VPWR VPWR _5137_/B sky130_fd_sc_hd__and4bb_1
Xhold1809 _4178_/X VGND VGND VPWR VPWR _6620_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4041_ hold941/X hold20/X _4056_/C VGND VGND VPWR VPWR _4041_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5992_ _6014_/A _6017_/B _6007_/C VGND VGND VPWR VPWR _5992_/X sky130_fd_sc_hd__and3_4
X_4943_ _4462_/Y _4938_/X _4791_/C VGND VGND VPWR VPWR _5151_/C sky130_fd_sc_hd__o21a_1
XFILLER_91_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4874_ _4500_/Y _4652_/Y _4873_/Y VGND VGND VPWR VPWR _4875_/D sky130_fd_sc_hd__o21a_1
X_6613_ _6760_/CLK _6613_/D _6433_/A VGND VGND VPWR VPWR _6613_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3825_ _3253_/A _3824_/X _3835_/S VGND VGND VPWR VPWR _6467_/D sky130_fd_sc_hd__mux2_1
XFILLER_137_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6544_ _7194_/CLK _6544_/D VGND VGND VPWR VPWR _6544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3756_ _6973_/Q _5398_/A _3347_/Y _7005_/Q _3755_/X VGND VGND VPWR VPWR _3759_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_5_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_5_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_118_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6475_ _6792_/CLK _6475_/D fanout442/X VGND VGND VPWR VPWR _6475_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_146_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3687_ _7134_/Q hold33/A _5175_/A _6783_/Q _3685_/X VGND VGND VPWR VPWR _3694_/A
+ sky130_fd_sc_hd__a221o_1
X_5426_ hold797/X _5570_/A1 _5433_/S VGND VGND VPWR VPWR _5426_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput220 _7216_/X VGND VGND VPWR VPWR mgmt_gpio_out[18] sky130_fd_sc_hd__buf_12
Xoutput231 _7226_/X VGND VGND VPWR VPWR mgmt_gpio_out[28] sky130_fd_sc_hd__buf_12
Xoutput242 _7208_/X VGND VGND VPWR VPWR mgmt_gpio_out[3] sky130_fd_sc_hd__buf_12
Xoutput253 _3961_/Y VGND VGND VPWR VPWR pad_flash_io0_oeb sky130_fd_sc_hd__buf_12
Xoutput264 _6786_/Q VGND VGND VPWR VPWR pll_div[2] sky130_fd_sc_hd__buf_12
XFILLER_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5357_ _5357_/A0 _5555_/A1 _5361_/S VGND VGND VPWR VPWR _5357_/X sky130_fd_sc_hd__mux2_1
Xoutput275 _6476_/Q VGND VGND VPWR VPWR pll_trim[13] sky130_fd_sc_hd__buf_12
Xoutput286 _6802_/Q VGND VGND VPWR VPWR pll_trim[23] sky130_fd_sc_hd__buf_12
Xoutput297 _6804_/Q VGND VGND VPWR VPWR pwr_ctrl_out[0] sky130_fd_sc_hd__buf_12
X_4308_ _4308_/A0 _5195_/A1 _4309_/S VGND VGND VPWR VPWR _6735_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5288_ _5288_/A0 _5576_/A1 _5289_/S VGND VGND VPWR VPWR _5288_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7027_ _7139_/CLK _7027_/D fanout478/X VGND VGND VPWR VPWR _7027_/Q sky130_fd_sc_hd__dfrtp_4
X_4239_ _5244_/A0 _5559_/A1 _4239_/S VGND VGND VPWR VPWR _4239_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire347 _3636_/Y VGND VGND VPWR VPWR _3675_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout480 fanout481/X VGND VGND VPWR VPWR fanout480/X sky130_fd_sc_hd__buf_12
XFILLER_47_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3610_ _7024_/Q _5452_/A _5398_/A _6976_/Q _3609_/X VGND VGND VPWR VPWR _3614_/C
+ sky130_fd_sc_hd__a221o_1
X_4590_ _4638_/A _4590_/B VGND VGND VPWR VPWR _4590_/Y sky130_fd_sc_hd__nand2_8
XFILLER_190_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3541_ _6799_/Q _3319_/Y _4140_/A _6593_/Q VGND VGND VPWR VPWR _3541_/X sky130_fd_sc_hd__a22o_1
XFILLER_183_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold906 _3391_/Y VGND VGND VPWR VPWR _5218_/S sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold917 hold58/X VGND VGND VPWR VPWR hold917/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_128_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold928 hold928/A VGND VGND VPWR VPWR hold928/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_143_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6260_ _6723_/Q _5978_/X _5995_/X _6600_/Q _6259_/X VGND VGND VPWR VPWR _6263_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_50_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold939 _5476_/X VGND VGND VPWR VPWR hold70/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_3472_ _6985_/Q _5407_/A _4292_/A _6726_/Q _3471_/X VGND VGND VPWR VPWR _3481_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5211_ _5218_/S _5551_/B VGND VGND VPWR VPWR _5217_/S sky130_fd_sc_hd__and2_4
XFILLER_88_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6191_ _6490_/Q _6191_/A2 _5649_/Y VGND VGND VPWR VPWR _6191_/X sky130_fd_sc_hd__a21o_1
XFILLER_130_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2307 hold811/X VGND VGND VPWR VPWR _4034_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5142_ _4688_/A _4995_/B _5023_/C _5141_/X _4815_/X VGND VGND VPWR VPWR _5143_/B
+ sky130_fd_sc_hd__o2111a_1
Xhold2318 _6630_/Q VGND VGND VPWR VPWR hold772/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2329 _6641_/Q VGND VGND VPWR VPWR hold583/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1606 hold680/X VGND VGND VPWR VPWR _4136_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1617 _6768_/Q VGND VGND VPWR VPWR hold110/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1628 hold685/X VGND VGND VPWR VPWR _4257_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5073_ _4776_/A _5073_/B _5073_/C _5100_/B VGND VGND VPWR VPWR _5156_/A sky130_fd_sc_hd__and4b_1
Xhold1639 _4161_/X VGND VGND VPWR VPWR _6606_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_4024_ hold925/X hold20/X _4047_/C VGND VGND VPWR VPWR _4024_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5975_ _6017_/A _6019_/B _6019_/C VGND VGND VPWR VPWR _5976_/B sky130_fd_sc_hd__and3_4
X_4926_ _4633_/B _4698_/Y _4702_/Y _4616_/B _4616_/A VGND VGND VPWR VPWR _4931_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_178_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4857_ _4917_/D _4857_/B _4857_/C VGND VGND VPWR VPWR _4857_/Y sky130_fd_sc_hd__nand3_1
XFILLER_193_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3808_ _3814_/B _6468_/Q _6469_/Q VGND VGND VPWR VPWR _3811_/B sky130_fd_sc_hd__and3b_1
XFILLER_165_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4788_ _4947_/A _4698_/Y _4531_/B VGND VGND VPWR VPWR _4788_/X sky130_fd_sc_hd__o21a_1
XFILLER_181_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6527_ _6711_/CLK _6527_/D _6433_/A VGND VGND VPWR VPWR _6527_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3739_ _3738_/X _3739_/A1 _3739_/S VGND VGND VPWR VPWR _3739_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6458_ _6658_/CLK _6458_/D _6408_/X VGND VGND VPWR VPWR _6458_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_133_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5409_ hold636/X _5580_/A1 _5415_/S VGND VGND VPWR VPWR _6982_/D sky130_fd_sc_hd__mux2_1
XFILLER_134_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6389_ _4222_/B _3189_/Y _4220_/B _6388_/X _6387_/X VGND VGND VPWR VPWR _7204_/D
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_851 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5760_ _5760_/A _5760_/B _5760_/C VGND VGND VPWR VPWR _5760_/Y sky130_fd_sc_hd__nor3_1
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4711_ _4826_/A _4730_/B VGND VGND VPWR VPWR _4924_/B sky130_fd_sc_hd__nand2_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5691_ _7077_/Q _5689_/X _5690_/X _5683_/X VGND VGND VPWR VPWR _5691_/X sky130_fd_sc_hd__a211o_1
XFILLER_148_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4642_ _4640_/Y _4857_/B VGND VGND VPWR VPWR _4642_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_175_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4573_ _4811_/B _4607_/B VGND VGND VPWR VPWR _4757_/A sky130_fd_sc_hd__nand2_1
XFILLER_116_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold703 hold703/A VGND VGND VPWR VPWR hold703/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap422 _4738_/B VGND VGND VPWR VPWR _4666_/A sky130_fd_sc_hd__clkbuf_2
X_6312_ _6587_/Q _5989_/X _6309_/X _6311_/X VGND VGND VPWR VPWR _6313_/C sky130_fd_sc_hd__a211oi_1
Xhold714 hold714/A VGND VGND VPWR VPWR hold714/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3524_ _7089_/Q _5524_/A _4262_/A _6701_/Q VGND VGND VPWR VPWR _3524_/X sky130_fd_sc_hd__a22o_1
Xmax_cap433 _4584_/A VGND VGND VPWR VPWR _4582_/A sky130_fd_sc_hd__clkbuf_2
Xhold725 hold725/A VGND VGND VPWR VPWR hold725/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold736 hold736/A VGND VGND VPWR VPWR hold736/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold747 hold747/A VGND VGND VPWR VPWR hold747/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold758 hold758/A VGND VGND VPWR VPWR hold758/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6243_ _6595_/Q _5991_/X _6018_/X _6718_/Q VGND VGND VPWR VPWR _6243_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold769 hold769/A VGND VGND VPWR VPWR hold769/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3455_ _7074_/Q _5506_/A _3347_/Y _7010_/Q VGND VGND VPWR VPWR _3455_/X sky130_fd_sc_hd__a22o_1
XFILLER_89_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6174_ _7059_/Q _5990_/X _5998_/X _6891_/Q _6173_/X VGND VGND VPWR VPWR _6179_/B
+ sky130_fd_sc_hd__a221o_1
Xhold2104 hold632/X VGND VGND VPWR VPWR _5554_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_3386_ _6448_/Q _6656_/Q VGND VGND VPWR VPWR _3739_/S sky130_fd_sc_hd__nand2_8
Xhold2115 _6878_/Q VGND VGND VPWR VPWR hold765/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2126 _6803_/Q VGND VGND VPWR VPWR hold686/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2137 _4323_/X VGND VGND VPWR VPWR _6747_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5125_ _5139_/B _5125_/B _5125_/C VGND VGND VPWR VPWR _5127_/C sky130_fd_sc_hd__and3_1
Xhold2148 hold715/X VGND VGND VPWR VPWR _4124_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1403 _4210_/X VGND VGND VPWR VPWR _6647_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2159 _6471_/Q VGND VGND VPWR VPWR hold595/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1414 _6538_/Q VGND VGND VPWR VPWR hold328/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1425 _5242_/X VGND VGND VPWR VPWR hold416/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1436 hold137/X VGND VGND VPWR VPWR _4312_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1447 _5579_/X VGND VGND VPWR VPWR hold293/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5056_ _4610_/A _4693_/B _4508_/B VGND VGND VPWR VPWR _5114_/C sky130_fd_sc_hd__o21ai_2
Xhold1458 _7028_/Q VGND VGND VPWR VPWR hold419/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1469 hold616/X VGND VGND VPWR VPWR _4027_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4007_ hold104/X hold78/X _4008_/S VGND VGND VPWR VPWR _4007_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5958_ _6756_/Q _5681_/X _5956_/X _5957_/X VGND VGND VPWR VPWR _5958_/X sky130_fd_sc_hd__a211o_1
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4909_ _4633_/B _4688_/A _4872_/A _4889_/B VGND VGND VPWR VPWR _5123_/A sky130_fd_sc_hd__o211a_1
XFILLER_187_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5889_ _6693_/Q _5658_/X _5664_/X _6758_/Q VGND VGND VPWR VPWR _5889_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold30 hold30/A VGND VGND VPWR VPWR hold30/X sky130_fd_sc_hd__clkbuf_2
Xhold41 hold41/A VGND VGND VPWR VPWR hold41/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold52 hold52/A VGND VGND VPWR VPWR hold52/X sky130_fd_sc_hd__buf_8
Xhold63 hold63/A VGND VGND VPWR VPWR hold63/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold74 hold74/A VGND VGND VPWR VPWR hold74/X sky130_fd_sc_hd__clkdlybuf4s25_2
XFILLER_75_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold85 hold85/A VGND VGND VPWR VPWR hold85/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold96 hold96/A VGND VGND VPWR VPWR hold96/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1970 _6697_/Q VGND VGND VPWR VPWR hold661/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1981 _6817_/Q VGND VGND VPWR VPWR hold634/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1992 _7030_/Q VGND VGND VPWR VPWR hold604/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_7__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7204_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_43_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_5 _5515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6930_ _7130_/CLK _6930_/D fanout458/X VGND VGND VPWR VPWR _6930_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_82_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6861_ _7109_/CLK _6861_/D fanout457/X VGND VGND VPWR VPWR _6861_/Q sky130_fd_sc_hd__dfstp_2
Xclkbuf_leaf_6_csclk _6727_/CLK VGND VGND VPWR VPWR _6648_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_50_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5812_ _6914_/Q _5670_/X _5685_/X _7074_/Q VGND VGND VPWR VPWR _5812_/X sky130_fd_sc_hd__a22o_1
XFILLER_35_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6792_ _6792_/CLK _6792_/D fanout442/X VGND VGND VPWR VPWR _6792_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5743_ _6855_/Q _5651_/X _5842_/A2 _6847_/Q VGND VGND VPWR VPWR _5743_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5674_ _5686_/A _5679_/B _5688_/C VGND VGND VPWR VPWR _5674_/X sky130_fd_sc_hd__and3b_4
XFILLER_148_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4625_ _4625_/A _4625_/B VGND VGND VPWR VPWR _4625_/Y sky130_fd_sc_hd__nand2_1
XFILLER_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold500 hold500/A VGND VGND VPWR VPWR _6854_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4556_ _4921_/A _4554_/X _4556_/C _5136_/A VGND VGND VPWR VPWR _4556_/X sky130_fd_sc_hd__and4bb_1
Xhold511 hold511/A VGND VGND VPWR VPWR hold511/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold522 hold522/A VGND VGND VPWR VPWR hold522/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold533 hold533/A VGND VGND VPWR VPWR hold533/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold544 hold544/A VGND VGND VPWR VPWR hold544/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3507_ _3530_/B _3523_/B VGND VGND VPWR VPWR _4182_/A sky130_fd_sc_hd__nor2_8
XFILLER_89_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold555 hold555/A VGND VGND VPWR VPWR hold555/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold566 hold566/A VGND VGND VPWR VPWR hold566/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4487_ _4595_/B _4488_/B VGND VGND VPWR VPWR _4972_/A sky130_fd_sc_hd__and2_4
Xhold577 _6586_/Q VGND VGND VPWR VPWR hold577/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold588 hold588/A VGND VGND VPWR VPWR hold588/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6226_ _6535_/Q _5983_/X _6005_/X _6692_/Q VGND VGND VPWR VPWR _6226_/X sky130_fd_sc_hd__a22o_1
Xhold599 hold599/A VGND VGND VPWR VPWR hold599/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3438_ input49/X _4047_/C hold67/A _7122_/Q VGND VGND VPWR VPWR _3438_/X sky130_fd_sc_hd__a22o_2
XFILLER_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _7122_/Q _5978_/X _5995_/X _6922_/Q _6156_/X VGND VGND VPWR VPWR _6163_/A
+ sky130_fd_sc_hd__a221o_1
X_3369_ _7004_/Q _5425_/A _3310_/Y input19/X _3358_/X VGND VGND VPWR VPWR _3369_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1200 _5359_/X VGND VGND VPWR VPWR _6938_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1211 _4067_/X VGND VGND VPWR VPWR _6526_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1222 _4163_/X VGND VGND VPWR VPWR _6608_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5108_ _5108_/A _5108_/B _5108_/C VGND VGND VPWR VPWR _5125_/B sky130_fd_sc_hd__and3_1
Xhold1233 hold123/X VGND VGND VPWR VPWR _5448_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1244 _6888_/Q VGND VGND VPWR VPWR hold175/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6088_ _6088_/A _6088_/B _6088_/C _6088_/D VGND VGND VPWR VPWR _6089_/D sky130_fd_sc_hd__nor4_1
Xhold1255 _4162_/X VGND VGND VPWR VPWR _6607_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1266 hold869/X VGND VGND VPWR VPWR hold232/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1277 _4332_/X VGND VGND VPWR VPWR _6755_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5039_ _5026_/B _4719_/B _4771_/X VGND VGND VPWR VPWR _5039_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_38_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1288 _4285_/X VGND VGND VPWR VPWR _6716_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_26_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1299 hold221/X VGND VGND VPWR VPWR _5233_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput120 wb_adr_i[29] VGND VGND VPWR VPWR _3894_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput131 wb_cyc_i VGND VGND VPWR VPWR _3893_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput142 wb_dat_i[19] VGND VGND VPWR VPWR _6371_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput153 wb_dat_i[29] VGND VGND VPWR VPWR _6377_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput164 wb_rstn_i VGND VGND VPWR VPWR input164/X sky130_fd_sc_hd__buf_8
XFILLER_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2490 _7145_/Q VGND VGND VPWR VPWR _3193_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4410_ _4719_/A _4590_/B VGND VGND VPWR VPWR _4812_/A sky130_fd_sc_hd__and2_4
XFILLER_145_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5390_ hold810/X _5552_/A1 _5397_/S VGND VGND VPWR VPWR _6965_/D sky130_fd_sc_hd__mux2_1
X_4341_ _3890_/Y _4340_/Y _4395_/A VGND VGND VPWR VPWR _4341_/X sky130_fd_sc_hd__o21a_2
XFILLER_126_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7060_ _7116_/CLK _7060_/D fanout455/X VGND VGND VPWR VPWR _7060_/Q sky130_fd_sc_hd__dfrtp_4
X_4272_ _4272_/A0 _5303_/A1 _4273_/S VGND VGND VPWR VPWR _4272_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6011_ _6002_/X _6011_/B VGND VGND VPWR VPWR _6011_/Y sky130_fd_sc_hd__nand2b_4
XFILLER_141_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3223_ _6968_/Q VGND VGND VPWR VPWR _5763_/A sky130_fd_sc_hd__clkinv_2
XFILLER_95_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6913_ _7134_/CLK _6913_/D fanout476/X VGND VGND VPWR VPWR _6913_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_63_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6844_ _7008_/CLK hold28/X fanout474/X VGND VGND VPWR VPWR _6844_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_808 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3987_ _3987_/A0 _5196_/A1 _3987_/S VGND VGND VPWR VPWR _6454_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6775_ _3958_/A1 _6775_/D _6427_/X VGND VGND VPWR VPWR _6775_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_176_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5726_ _6990_/Q _5929_/B _5688_/X _6886_/Q _5725_/X VGND VGND VPWR VPWR _5727_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5657_ _7149_/Q _7148_/Q VGND VGND VPWR VPWR _5689_/C sky130_fd_sc_hd__and2_4
XFILLER_163_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4608_ _4570_/A _4564_/Y _4575_/C _4495_/B VGND VGND VPWR VPWR _4609_/D sky130_fd_sc_hd__a211o_1
X_5588_ _6816_/Q _5611_/A _3197_/Y _5588_/B1 _5587_/X VGND VGND VPWR VPWR _7141_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_123_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold330 hold330/A VGND VGND VPWR VPWR hold330/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold341 hold341/A VGND VGND VPWR VPWR hold341/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4539_ _4621_/A _4972_/A VGND VGND VPWR VPWR _4539_/Y sky130_fd_sc_hd__nand2_2
Xhold352 hold964/X VGND VGND VPWR VPWR hold965/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold363 hold363/A VGND VGND VPWR VPWR hold363/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold374 hold374/A VGND VGND VPWR VPWR hold374/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold385 hold385/A VGND VGND VPWR VPWR hold385/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold396 hold396/A VGND VGND VPWR VPWR hold396/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6209_ _6956_/Q _5997_/X _6012_/X _7004_/Q VGND VGND VPWR VPWR _6209_/X sky130_fd_sc_hd__a22o_1
X_7189_ _7194_/CLK _7189_/D VGND VGND VPWR VPWR _7189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1030 hold171/X VGND VGND VPWR VPWR hold9/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1041 _3260_/X VGND VGND VPWR VPWR _3261_/B sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1052 hold396/X VGND VGND VPWR VPWR _5567_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1063 _3303_/X VGND VGND VPWR VPWR _5207_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1074 _7059_/Q VGND VGND VPWR VPWR hold409/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1085 _6963_/Q VGND VGND VPWR VPWR hold412/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_203 _5986_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1096 _5585_/X VGND VGND VPWR VPWR _7139_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_71_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6691_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_17_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3910_ _7142_/Q _7143_/Q _7144_/Q _7145_/Q VGND VGND VPWR VPWR _3911_/B sky130_fd_sc_hd__and4bb_1
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4890_ _4464_/Y _4601_/A _4601_/B _4581_/X VGND VGND VPWR VPWR _5103_/A sky130_fd_sc_hd__a211o_1
X_3841_ _3841_/A _3841_/B VGND VGND VPWR VPWR _6462_/D sky130_fd_sc_hd__xnor2_1
XFILLER_149_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3772_ _6579_/Q _4128_/A _4212_/A _6649_/Q _3771_/X VGND VGND VPWR VPWR _3772_/X
+ sky130_fd_sc_hd__a221o_2
X_6560_ _6568_/CLK _6560_/D VGND VGND VPWR VPWR _6560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5511_ _5511_/A0 _5583_/A1 _5514_/S VGND VGND VPWR VPWR _7073_/D sky130_fd_sc_hd__mux2_1
X_6491_ _7152_/CLK _6491_/D _6399_/A VGND VGND VPWR VPWR _6491_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_158_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5442_ _5442_/A0 _5577_/A1 _5442_/S VGND VGND VPWR VPWR _7012_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5373_ hold684/X _5580_/A1 _5379_/S VGND VGND VPWR VPWR _6950_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_24_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7136_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_114_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4324_ _4324_/A0 _5193_/A1 _4327_/S VGND VGND VPWR VPWR _4324_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7112_ _7138_/CLK _7112_/D fanout480/X VGND VGND VPWR VPWR _7112_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7043_ _7138_/CLK _7043_/D fanout477/X VGND VGND VPWR VPWR _7043_/Q sky130_fd_sc_hd__dfrtp_4
X_4255_ _4255_/A0 _5196_/A1 _4255_/S VGND VGND VPWR VPWR _4255_/X sky130_fd_sc_hd__mux2_1
X_3206_ _7104_/Q VGND VGND VPWR VPWR _3206_/Y sky130_fd_sc_hd__inv_2
X_4186_ _4186_/A0 _5195_/A1 _4187_/S VGND VGND VPWR VPWR _6627_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_39_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7133_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_83_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_1_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR _6727_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_82_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6827_ _7097_/CLK _6827_/D fanout468/X VGND VGND VPWR VPWR _6827_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6758_ _6759_/CLK _6758_/D _6426_/A VGND VGND VPWR VPWR _6758_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_149_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5709_ _5709_/A1 _5649_/Y _5707_/Y _5708_/X VGND VGND VPWR VPWR _7160_/D sky130_fd_sc_hd__a22o_1
X_6689_ _6817_/CLK _6689_/D fanout445/X VGND VGND VPWR VPWR _6689_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_109_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold160 hold160/A VGND VGND VPWR VPWR hold160/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold171 hold171/A VGND VGND VPWR VPWR hold171/X sky130_fd_sc_hd__clkbuf_2
XFILLER_78_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold182 hold182/A VGND VGND VPWR VPWR hold182/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold193 hold193/A VGND VGND VPWR VPWR hold193/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4040_ _4040_/A0 _4039_/X _4046_/S VGND VGND VPWR VPWR _4040_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5991_ _6017_/A _6007_/C _6016_/C VGND VGND VPWR VPWR _5991_/X sky130_fd_sc_hd__and3_4
XFILLER_52_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4942_ _5026_/B _5033_/A VGND VGND VPWR VPWR _5032_/B sky130_fd_sc_hd__nand2_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4873_ _4988_/A _4607_/B _4526_/X VGND VGND VPWR VPWR _4873_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_178_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6612_ _6760_/CLK _6612_/D _6433_/A VGND VGND VPWR VPWR _6612_/Q sky130_fd_sc_hd__dfrtp_4
X_3824_ _3254_/X _3253_/Y _3827_/B VGND VGND VPWR VPWR _3824_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3755_ _6861_/Q _5272_/A _4077_/A _6535_/Q VGND VGND VPWR VPWR _3755_/X sky130_fd_sc_hd__a22o_1
X_6543_ _7194_/CLK _6543_/D VGND VGND VPWR VPWR _6543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3686_ hold32/X _3686_/B VGND VGND VPWR VPWR _5175_/A sky130_fd_sc_hd__nor2_2
X_6474_ _6792_/CLK _6474_/D fanout442/X VGND VGND VPWR VPWR _6474_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_146_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput210 _3233_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[7] sky130_fd_sc_hd__buf_12
X_5425_ _5425_/A _5569_/B VGND VGND VPWR VPWR _5433_/S sky130_fd_sc_hd__and2_4
Xoutput221 _7217_/X VGND VGND VPWR VPWR mgmt_gpio_out[19] sky130_fd_sc_hd__buf_12
XFILLER_160_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput232 _7227_/X VGND VGND VPWR VPWR mgmt_gpio_out[29] sky130_fd_sc_hd__buf_12
Xoutput243 _7209_/X VGND VGND VPWR VPWR mgmt_gpio_out[4] sky130_fd_sc_hd__buf_12
Xoutput254 _7231_/X VGND VGND VPWR VPWR pad_flash_io1_do sky130_fd_sc_hd__buf_12
X_5356_ _5356_/A0 _5518_/A1 _5361_/S VGND VGND VPWR VPWR _5356_/X sky130_fd_sc_hd__mux2_1
Xoutput265 _6787_/Q VGND VGND VPWR VPWR pll_div[3] sky130_fd_sc_hd__buf_12
XFILLER_160_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput276 _6477_/Q VGND VGND VPWR VPWR pll_trim[14] sky130_fd_sc_hd__buf_12
XFILLER_58_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput287 _6487_/Q VGND VGND VPWR VPWR pll_trim[24] sky130_fd_sc_hd__buf_12
X_4307_ hold558/X _5187_/A1 _4309_/S VGND VGND VPWR VPWR _6734_/D sky130_fd_sc_hd__mux2_1
Xoutput298 _6805_/Q VGND VGND VPWR VPWR pwr_ctrl_out[1] sky130_fd_sc_hd__buf_12
X_5287_ hold989/X _5575_/A1 _5289_/S VGND VGND VPWR VPWR _5287_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7026_ _7035_/CLK _7026_/D fanout456/X VGND VGND VPWR VPWR _7026_/Q sky130_fd_sc_hd__dfrtp_4
X_4238_ _4238_/A0 _4237_/X _4240_/S VGND VGND VPWR VPWR _4238_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4169_ _4169_/A0 _5538_/A1 _4169_/S VGND VGND VPWR VPWR _4169_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire348 _3444_/Y VGND VGND VPWR VPWR _3462_/A sky130_fd_sc_hd__buf_2
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout470 fanout481/X VGND VGND VPWR VPWR fanout470/X sky130_fd_sc_hd__buf_8
XFILLER_120_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout481 fanout482/X VGND VGND VPWR VPWR fanout481/X sky130_fd_sc_hd__buf_12
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3540_ _3540_/A _3550_/B VGND VGND VPWR VPWR _4140_/A sky130_fd_sc_hd__nor2_8
XFILLER_190_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold907 _5216_/X VGND VGND VPWR VPWR _6814_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold918 _5557_/X VGND VGND VPWR VPWR hold59/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_115_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold929 _5243_/X VGND VGND VPWR VPWR _6835_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_3471_ _6841_/Q hold27/A _5178_/A _6788_/Q VGND VGND VPWR VPWR _3471_/X sky130_fd_sc_hd__a22o_1
XFILLER_170_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5210_ _5220_/C _5210_/B VGND VGND VPWR VPWR _6809_/D sky130_fd_sc_hd__and2_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6190_ _6843_/Q _6011_/Y _6189_/Y _6341_/S VGND VGND VPWR VPWR _6190_/X sky130_fd_sc_hd__o211a_1
XFILLER_97_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5141_ _5011_/A _4590_/Y _4676_/Y VGND VGND VPWR VPWR _5141_/X sky130_fd_sc_hd__a21o_1
Xhold2308 _4034_/X VGND VGND VPWR VPWR _6502_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2319 hold772/X VGND VGND VPWR VPWR _4190_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1607 _4136_/X VGND VGND VPWR VPWR _6585_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5072_ _5135_/A _5102_/C _5072_/C _5135_/C VGND VGND VPWR VPWR _5074_/C sky130_fd_sc_hd__and4_1
XFILLER_96_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1618 hold110/X VGND VGND VPWR VPWR _3257_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1629 _4257_/X VGND VGND VPWR VPWR _6692_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4023_ _4023_/A0 _4022_/X _4029_/S VGND VGND VPWR VPWR _4023_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5974_ _7154_/Q _7153_/Q VGND VGND VPWR VPWR _6019_/C sky130_fd_sc_hd__nor2_8
XFILLER_80_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4925_ _4925_/A _5052_/B _4925_/C VGND VGND VPWR VPWR _4925_/X sky130_fd_sc_hd__and3_1
XFILLER_100_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4856_ _4638_/Y _4662_/Y _5073_/B VGND VGND VPWR VPWR _4856_/X sky130_fd_sc_hd__o21a_1
XFILLER_138_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3807_ _3903_/A _3807_/B VGND VGND VPWR VPWR _3814_/B sky130_fd_sc_hd__and2_2
X_4787_ _4411_/Y _4683_/A _4664_/Y _4509_/Y VGND VGND VPWR VPWR _5034_/B sky130_fd_sc_hd__o31a_1
XFILLER_146_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6526_ _6816_/CLK _6526_/D _6414_/A VGND VGND VPWR VPWR _6526_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3738_ _6774_/Q _3737_/Y _3738_/S VGND VGND VPWR VPWR _3738_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6457_ _3958_/A1 _6457_/D _6407_/X VGND VGND VPWR VPWR _6457_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_161_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3669_ _7111_/Q _5551_/A _4116_/A _6571_/Q VGND VGND VPWR VPWR _3669_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5408_ hold664/X _5552_/A1 _5415_/S VGND VGND VPWR VPWR _6981_/D sky130_fd_sc_hd__mux2_1
XFILLER_192_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6388_ _6682_/Q hold11/A _6355_/Y VGND VGND VPWR VPWR _6388_/X sky130_fd_sc_hd__o21ba_1
XFILLER_88_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5339_ _5339_/A0 _5555_/A1 _5343_/S VGND VGND VPWR VPWR _6920_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7009_ _7111_/CLK _7009_/D fanout472/X VGND VGND VPWR VPWR _7009_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_6__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _3950_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_28_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4710_ _4710_/A _5150_/C VGND VGND VPWR VPWR _4832_/C sky130_fd_sc_hd__nand2_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5690_ _6989_/Q _5929_/B _5670_/X _6909_/Q VGND VGND VPWR VPWR _5690_/X sky130_fd_sc_hd__a22o_1
XFILLER_187_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4641_ _4498_/X _4499_/Y _4500_/Y _4501_/X VGND VGND VPWR VPWR _4857_/B sky130_fd_sc_hd__o211a_1
X_4572_ _4637_/B _4823_/A VGND VGND VPWR VPWR _4572_/Y sky130_fd_sc_hd__nor2_1
XFILLER_116_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6311_ _6652_/Q _5996_/X _6012_/X _6750_/Q _6310_/X VGND VGND VPWR VPWR _6311_/X
+ sky130_fd_sc_hd__a221o_1
Xhold704 hold704/A VGND VGND VPWR VPWR hold704/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap423 _4713_/C VGND VGND VPWR VPWR _4738_/B sky130_fd_sc_hd__clkbuf_2
Xhold715 hold715/A VGND VGND VPWR VPWR hold715/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3523_ _3550_/A _3523_/B VGND VGND VPWR VPWR _4262_/A sky130_fd_sc_hd__nor2_4
Xhold726 hold726/A VGND VGND VPWR VPWR hold726/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold737 hold737/A VGND VGND VPWR VPWR hold737/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold748 hold748/A VGND VGND VPWR VPWR hold748/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3454_ _7050_/Q _5479_/A hold27/A _6842_/Q _3436_/X VGND VGND VPWR VPWR _3460_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_116_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6242_ _6242_/A0 _6241_/X _6342_/S VGND VGND VPWR VPWR _6242_/X sky130_fd_sc_hd__mux2_1
Xhold759 hold759/A VGND VGND VPWR VPWR hold759/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_170_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3385_ _3385_/A _3385_/B VGND VGND VPWR VPWR _3385_/Y sky130_fd_sc_hd__nand2_8
X_6173_ _6907_/Q _5985_/X _6018_/X _6971_/Q VGND VGND VPWR VPWR _6173_/X sky130_fd_sc_hd__a22o_1
Xhold2105 _6949_/Q VGND VGND VPWR VPWR hold679/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2116 _6790_/Q VGND VGND VPWR VPWR hold731/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2127 _5201_/X VGND VGND VPWR VPWR hold687/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2138 _6521_/Q VGND VGND VPWR VPWR hold399/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5124_ _4636_/X _5124_/B _5124_/C _5136_/A VGND VGND VPWR VPWR _5125_/C sky130_fd_sc_hd__and4b_1
Xhold2149 _4124_/X VGND VGND VPWR VPWR _6575_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1404 _6859_/Q VGND VGND VPWR VPWR hold356/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1415 _4081_/X VGND VGND VPWR VPWR hold329/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1426 _6539_/Q VGND VGND VPWR VPWR hold516/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_747 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1437 _4312_/X VGND VGND VPWR VPWR _6738_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5055_ _4570_/D _4523_/Y _4931_/B _5054_/X VGND VGND VPWR VPWR _5058_/C sky130_fd_sc_hd__o211a_1
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1448 _6860_/Q VGND VGND VPWR VPWR hold469/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1459 hold419/X VGND VGND VPWR VPWR _5460_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4006_ hold431/X _5503_/A1 _4008_/S VGND VGND VPWR VPWR _6484_/D sky130_fd_sc_hd__mux2_1
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5957_ _6613_/Q _5660_/X _5669_/X _6653_/Q VGND VGND VPWR VPWR _5957_/X sky130_fd_sc_hd__a22o_1
X_4908_ _4636_/X _5127_/B _5127_/A VGND VGND VPWR VPWR _5115_/A sky130_fd_sc_hd__and3b_1
X_5888_ _6595_/Q _5670_/X _5685_/X _6770_/Q VGND VGND VPWR VPWR _5888_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4839_ _4917_/A _4643_/C _4504_/X VGND VGND VPWR VPWR _4839_/X sky130_fd_sc_hd__a21o_1
XFILLER_166_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6509_ _7138_/CLK _6509_/D fanout480/X VGND VGND VPWR VPWR _6509_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold20 hold20/A VGND VGND VPWR VPWR hold20/X sky130_fd_sc_hd__buf_12
XFILLER_102_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold31 hold31/A VGND VGND VPWR VPWR hold31/X sky130_fd_sc_hd__buf_8
XFILLER_102_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold42 hold42/A VGND VGND VPWR VPWR hold42/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold53 hold53/A VGND VGND VPWR VPWR hold53/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold64 hold64/A VGND VGND VPWR VPWR hold64/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold75 hold75/A VGND VGND VPWR VPWR hold75/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1960 _4015_/X VGND VGND VPWR VPWR hold440/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold86 hold86/A VGND VGND VPWR VPWR hold86/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold97 hold97/A VGND VGND VPWR VPWR hold97/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1971 hold661/X VGND VGND VPWR VPWR _4263_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1982 hold634/X VGND VGND VPWR VPWR _5221_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1993 _7054_/Q VGND VGND VPWR VPWR hold683/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_71_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_6 _5326_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6860_ _7124_/CLK _6860_/D fanout458/X VGND VGND VPWR VPWR _6860_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_179_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5811_ _6954_/Q _5672_/X _5679_/X _6906_/Q _5810_/X VGND VGND VPWR VPWR _5811_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6791_ _6793_/CLK _6791_/D fanout442/X VGND VGND VPWR VPWR _6791_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5742_ _6879_/Q _5667_/X _5682_/X _7039_/Q VGND VGND VPWR VPWR _5742_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5673_ _5689_/A _5684_/B _5676_/B VGND VGND VPWR VPWR _5673_/X sky130_fd_sc_hd__and3b_4
XFILLER_191_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4624_ _4569_/C _4655_/A _4901_/B _4622_/X _5098_/A VGND VGND VPWR VPWR _4624_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_163_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold501 hold501/A VGND VGND VPWR VPWR hold501/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4555_ _5026_/B _4948_/A _4392_/X VGND VGND VPWR VPWR _4556_/C sky130_fd_sc_hd__a21oi_1
Xhold512 hold512/A VGND VGND VPWR VPWR hold512/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold523 hold523/A VGND VGND VPWR VPWR hold523/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold534 hold534/A VGND VGND VPWR VPWR hold534/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3506_ _6598_/Q _4146_/A _4122_/A _6578_/Q VGND VGND VPWR VPWR _3506_/X sky130_fd_sc_hd__a22o_1
Xhold545 hold545/A VGND VGND VPWR VPWR hold545/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold556 hold556/A VGND VGND VPWR VPWR hold556/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4486_ _4486_/A _4486_/B VGND VGND VPWR VPWR _4569_/C sky130_fd_sc_hd__nand2_4
Xhold567 hold567/A VGND VGND VPWR VPWR hold567/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold578 hold578/A VGND VGND VPWR VPWR hold578/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6225_ _6742_/Q _6014_/X _6219_/X _6224_/X VGND VGND VPWR VPWR _6230_/A sky130_fd_sc_hd__a211o_1
Xhold589 hold589/A VGND VGND VPWR VPWR hold589/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3437_ input31/X _3307_/Y _3339_/Y _6476_/Q VGND VGND VPWR VPWR _3437_/X sky130_fd_sc_hd__a22o_1
XFILLER_98_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ _3368_/A _3368_/B _3368_/C _3368_/D VGND VGND VPWR VPWR _3368_/Y sky130_fd_sc_hd__nor4_2
X_6156_ hold49/A _6008_/X _6016_/X _7042_/Q VGND VGND VPWR VPWR _6156_/X sky130_fd_sc_hd__a22o_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1201 _6843_/Q VGND VGND VPWR VPWR hold496/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1212 _6994_/Q VGND VGND VPWR VPWR hold476/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1223 _6715_/Q VGND VGND VPWR VPWR hold174/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5107_ _5107_/A _5107_/B _5107_/C VGND VGND VPWR VPWR _5123_/C sky130_fd_sc_hd__and3_1
Xhold1234 _5448_/X VGND VGND VPWR VPWR _7017_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_3299_ _3333_/A _3726_/A VGND VGND VPWR VPWR hold40/A sky130_fd_sc_hd__nor2_8
XFILLER_58_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6087_ _7135_/Q _5977_/X _5984_/X _7095_/Q _6086_/X VGND VGND VPWR VPWR _6088_/D
+ sky130_fd_sc_hd__a221o_1
Xhold1245 hold175/X VGND VGND VPWR VPWR _5303_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1256 _6932_/Q VGND VGND VPWR VPWR hold362/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1267 hold232/X VGND VGND VPWR VPWR hold1267/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1278 _6827_/Q VGND VGND VPWR VPWR hold132/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5038_ _4769_/Y _5038_/B _5038_/C VGND VGND VPWR VPWR _5043_/A sky130_fd_sc_hd__and3b_1
XFILLER_26_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1289 _6561_/Q VGND VGND VPWR VPWR hold868/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6989_ _7077_/CLK _6989_/D fanout456/X VGND VGND VPWR VPWR _6989_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_15_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput110 wb_adr_i[1] VGND VGND VPWR VPWR _4637_/A sky130_fd_sc_hd__clkbuf_16
Xinput121 wb_adr_i[2] VGND VGND VPWR VPWR _4637_/D sky130_fd_sc_hd__buf_12
XFILLER_103_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput132 wb_dat_i[0] VGND VGND VPWR VPWR _6362_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput143 wb_dat_i[1] VGND VGND VPWR VPWR _6364_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput154 wb_dat_i[2] VGND VGND VPWR VPWR _6368_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput165 wb_sel_i[0] VGND VGND VPWR VPWR _6355_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2480 _7177_/Q VGND VGND VPWR VPWR _6142_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_36_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2491 _7180_/Q VGND VGND VPWR VPWR _6217_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1790 hold298/X VGND VGND VPWR VPWR _4197_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_63_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4340_ _4649_/C _4649_/D VGND VGND VPWR VPWR _4340_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4271_ _4271_/A0 _5187_/A1 _4273_/S VGND VGND VPWR VPWR _4271_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6010_ _6010_/A _6010_/B _6010_/C VGND VGND VPWR VPWR _6011_/B sky130_fd_sc_hd__nor3_2
X_3222_ _6976_/Q VGND VGND VPWR VPWR _3222_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6912_ _7091_/CLK _6912_/D fanout471/X VGND VGND VPWR VPWR _6912_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6843_ _7136_/CLK _6843_/D fanout475/X VGND VGND VPWR VPWR _6843_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6774_ _3958_/A1 _6774_/D _6426_/X VGND VGND VPWR VPWR _6774_/Q sky130_fd_sc_hd__dfrtn_1
X_3986_ _3986_/A0 hold106/X _3996_/S VGND VGND VPWR VPWR _3986_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5725_ _6854_/Q _5651_/X _5684_/X _6926_/Q VGND VGND VPWR VPWR _5725_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5656_ _5689_/A _5676_/B _5689_/B VGND VGND VPWR VPWR _5656_/X sky130_fd_sc_hd__and3_4
XFILLER_136_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4607_ _4988_/A _4607_/B VGND VGND VPWR VPWR _4754_/D sky130_fd_sc_hd__nand2_1
XFILLER_191_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5587_ _5610_/A _3915_/Y _6492_/Q VGND VGND VPWR VPWR _5587_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold320 hold320/A VGND VGND VPWR VPWR _6712_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold331 hold331/A VGND VGND VPWR VPWR _6823_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4538_ _4724_/C _4621_/A VGND VGND VPWR VPWR _4894_/A sky130_fd_sc_hd__nand2_1
Xhold342 hold342/A VGND VGND VPWR VPWR hold342/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold353 hold353/A VGND VGND VPWR VPWR hold353/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold364 hold364/A VGND VGND VPWR VPWR hold364/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold375 _5405_/X VGND VGND VPWR VPWR _6979_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold386 hold386/A VGND VGND VPWR VPWR hold386/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4469_ _4917_/A _4469_/B VGND VGND VPWR VPWR _4568_/A sky130_fd_sc_hd__nor2_2
Xhold397 hold397/A VGND VGND VPWR VPWR hold397/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6208_ _7092_/Q _5638_/X _5992_/X _6964_/Q _6207_/X VGND VGND VPWR VPWR _6208_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7188_ _7194_/CLK _7188_/D VGND VGND VPWR VPWR _7188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6139_ _6120_/X _6139_/B _6139_/C VGND VGND VPWR VPWR _6139_/Y sky130_fd_sc_hd__nand3b_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1020 _5477_/X VGND VGND VPWR VPWR _7043_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1031 hold9/X VGND VGND VPWR VPWR _5267_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1042 _3347_/Y VGND VGND VPWR VPWR _5434_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1053 _5567_/X VGND VGND VPWR VPWR _7123_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1064 _5198_/S VGND VGND VPWR VPWR _5199_/S sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1075 hold409/X VGND VGND VPWR VPWR _5495_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1086 hold412/X VGND VGND VPWR VPWR _5387_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_204 _5992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1097 _7075_/Q VGND VGND VPWR VPWR hold408/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_5_csclk _6727_/CLK VGND VGND VPWR VPWR _6761_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_107_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3840_ _3840_/A _3840_/B VGND VGND VPWR VPWR _3841_/B sky130_fd_sc_hd__nand2_1
XFILLER_149_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3771_ _6644_/Q _4206_/A _4328_/A _6752_/Q VGND VGND VPWR VPWR _3771_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5510_ _5510_/A0 _5582_/A1 _5514_/S VGND VGND VPWR VPWR _5510_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6490_ _7152_/CLK _6490_/D _6399_/A VGND VGND VPWR VPWR _6490_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_9_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5441_ hold360/X _5576_/A1 _5442_/S VGND VGND VPWR VPWR _5441_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5372_ hold679/X _5561_/A1 _5379_/S VGND VGND VPWR VPWR _6949_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7111_ _7111_/CLK _7111_/D fanout472/X VGND VGND VPWR VPWR _7111_/Q sky130_fd_sc_hd__dfrtp_4
X_4323_ _4323_/A0 _5208_/A1 _4327_/S VGND VGND VPWR VPWR _4323_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7042_ _7091_/CLK hold70/X fanout471/X VGND VGND VPWR VPWR _7042_/Q sky130_fd_sc_hd__dfrtp_4
X_4254_ _4254_/A0 _5195_/A1 _4255_/S VGND VGND VPWR VPWR _4254_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3205_ _7112_/Q VGND VGND VPWR VPWR _3205_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4185_ hold305/X _4337_/A1 _4187_/S VGND VGND VPWR VPWR _4185_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6826_ _6826_/CLK _6826_/D _6414_/A VGND VGND VPWR VPWR _6826_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6757_ _6757_/CLK _6757_/D fanout447/X VGND VGND VPWR VPWR _6757_/Q sky130_fd_sc_hd__dfrtp_4
X_3969_ _3969_/A _3969_/B VGND VGND VPWR VPWR _6678_/D sky130_fd_sc_hd__nor2_1
X_5708_ _5692_/X _5697_/X _5706_/X _5647_/Y VGND VGND VPWR VPWR _5708_/X sky130_fd_sc_hd__o31a_2
XFILLER_109_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6688_ _6691_/CLK _6688_/D fanout443/X VGND VGND VPWR VPWR _6688_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_176_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5639_ _5639_/A _5639_/B VGND VGND VPWR VPWR _5639_/Y sky130_fd_sc_hd__nor2_1
XFILLER_128_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold150 hold150/A VGND VGND VPWR VPWR _6650_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold161 hold161/A VGND VGND VPWR VPWR _6500_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold172 hold172/A VGND VGND VPWR VPWR _6864_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold183 hold183/A VGND VGND VPWR VPWR hold183/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold194 hold194/A VGND VGND VPWR VPWR hold194/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5990_ _6014_/A _6019_/B _6016_/C VGND VGND VPWR VPWR _5990_/X sky130_fd_sc_hd__and3_4
X_4941_ _4729_/A _4691_/Y _4935_/X _4477_/Y _4534_/Y VGND VGND VPWR VPWR _4963_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_32_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4872_ _4872_/A _5046_/A _4872_/C _4872_/D VGND VGND VPWR VPWR _4875_/C sky130_fd_sc_hd__and4_1
X_6611_ _6648_/CLK _6611_/D fanout449/X VGND VGND VPWR VPWR _6611_/Q sky130_fd_sc_hd__dfstp_4
X_3823_ hold86/A _3826_/B VGND VGND VPWR VPWR _3827_/B sky130_fd_sc_hd__and2_1
XFILLER_119_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6542_ _7194_/CLK _6542_/D VGND VGND VPWR VPWR _6542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3754_ _6989_/Q _5416_/A _5479_/A _7045_/Q _3753_/X VGND VGND VPWR VPWR _3759_/B
+ sky130_fd_sc_hd__a221o_1
X_6473_ _6794_/CLK _6473_/D fanout444/X VGND VGND VPWR VPWR _6473_/Q sky130_fd_sc_hd__dfstp_2
X_3685_ _6758_/Q _4334_/A _4176_/A _6620_/Q VGND VGND VPWR VPWR _3685_/X sky130_fd_sc_hd__a22o_1
X_5424_ _5424_/A0 _5559_/A1 _5424_/S VGND VGND VPWR VPWR _5424_/X sky130_fd_sc_hd__mux2_1
Xoutput200 _3207_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[32] sky130_fd_sc_hd__buf_12
Xoutput211 _3232_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[8] sky130_fd_sc_hd__buf_12
Xoutput222 _3945_/X VGND VGND VPWR VPWR mgmt_gpio_out[1] sky130_fd_sc_hd__buf_12
Xoutput233 _7207_/X VGND VGND VPWR VPWR mgmt_gpio_out[2] sky130_fd_sc_hd__buf_12
XFILLER_160_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput244 _7210_/X VGND VGND VPWR VPWR mgmt_gpio_out[5] sky130_fd_sc_hd__buf_12
X_5355_ hold508/X _5499_/A1 _5361_/S VGND VGND VPWR VPWR _5355_/X sky130_fd_sc_hd__mux2_1
Xoutput255 _3963_/A VGND VGND VPWR VPWR pad_flash_io1_ieb sky130_fd_sc_hd__buf_12
Xoutput266 _6788_/Q VGND VGND VPWR VPWR pll_div[4] sky130_fd_sc_hd__buf_12
Xoutput277 _6478_/Q VGND VGND VPWR VPWR pll_trim[15] sky130_fd_sc_hd__buf_12
X_4306_ _4306_/A0 _5186_/A1 _4309_/S VGND VGND VPWR VPWR _6733_/D sky130_fd_sc_hd__mux2_1
Xoutput288 _6488_/Q VGND VGND VPWR VPWR pll_trim[25] sky130_fd_sc_hd__buf_12
Xoutput299 _6806_/Q VGND VGND VPWR VPWR pwr_ctrl_out[2] sky130_fd_sc_hd__buf_12
X_5286_ _5286_/A0 _5556_/A1 _5289_/S VGND VGND VPWR VPWR _5286_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7025_ _7105_/CLK _7025_/D fanout473/X VGND VGND VPWR VPWR _7025_/Q sky130_fd_sc_hd__dfrtp_4
X_4237_ hold928/X hold78/X _4239_/S VGND VGND VPWR VPWR _4237_/X sky130_fd_sc_hd__mux2_1
X_4168_ _4168_/A0 _5249_/A1 _4169_/S VGND VGND VPWR VPWR _4168_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_5__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7152_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4099_ _3803_/Y hold840/A _4106_/S VGND VGND VPWR VPWR _6553_/D sky130_fd_sc_hd__mux2_1
XFILLER_15_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6809_ _6809_/CLK _6809_/D fanout444/X VGND VGND VPWR VPWR _7206_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_23_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire349 _3368_/Y VGND VGND VPWR VPWR _3385_/A sky130_fd_sc_hd__buf_2
XFILLER_183_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_70_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6792_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_152_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout460 fanout482/X VGND VGND VPWR VPWR fanout460/X sky130_fd_sc_hd__buf_12
XFILLER_171_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout471 fanout481/X VGND VGND VPWR VPWR fanout471/X sky130_fd_sc_hd__buf_12
Xfanout482 input75/X VGND VGND VPWR VPWR fanout482/X sky130_fd_sc_hd__buf_12
XFILLER_48_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_23_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7137_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_38_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7079_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold908 _6763_/Q VGND VGND VPWR VPWR hold908/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_143_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold919 _6882_/Q VGND VGND VPWR VPWR hold919/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_3470_ _3470_/A hold26/X VGND VGND VPWR VPWR _5178_/A sky130_fd_sc_hd__nor2_8
XFILLER_142_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5140_ _5140_/A _5140_/B _5140_/C VGND VGND VPWR VPWR _5140_/X sky130_fd_sc_hd__and3_1
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2309 _6473_/Q VGND VGND VPWR VPWR hold574/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1608 _6972_/Q VGND VGND VPWR VPWR hold512/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5071_ _5135_/C VGND VGND VPWR VPWR _5071_/Y sky130_fd_sc_hd__inv_2
Xhold1619 _3257_/X VGND VGND VPWR VPWR _3259_/B sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4022_ _4052_/A0 _5556_/A1 _4047_/C VGND VGND VPWR VPWR _4022_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5973_ _6015_/B _6008_/A _6018_/B VGND VGND VPWR VPWR _5973_/X sky130_fd_sc_hd__and3_4
XFILLER_80_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4924_ _4924_/A _4924_/B _4924_/C _5046_/B VGND VGND VPWR VPWR _4925_/C sky130_fd_sc_hd__and4_1
XFILLER_33_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4855_ _4570_/D _4655_/A _4590_/Y _4674_/Y VGND VGND VPWR VPWR _4922_/C sky130_fd_sc_hd__o22a_1
XFILLER_193_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3806_ _6657_/Q _6656_/Q VGND VGND VPWR VPWR _3807_/B sky130_fd_sc_hd__nor2_2
XFILLER_119_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4786_ _4729_/A _4698_/Y _5095_/A VGND VGND VPWR VPWR _4786_/X sky130_fd_sc_hd__o21a_1
X_6525_ _6711_/CLK _6525_/D fanout465/X VGND VGND VPWR VPWR _6525_/Q sky130_fd_sc_hd__dfrtp_4
X_3737_ _3737_/A _3737_/B VGND VGND VPWR VPWR _3737_/Y sky130_fd_sc_hd__nand2_4
XFILLER_146_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6456_ _3958_/A1 _6456_/D _6406_/X VGND VGND VPWR VPWR _6456_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_174_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3668_ _6473_/Q _3339_/Y _4262_/A _6699_/Q _3667_/X VGND VGND VPWR VPWR _3673_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5407_ _5407_/A _5407_/B VGND VGND VPWR VPWR _5415_/S sky130_fd_sc_hd__and2_4
X_6387_ _6686_/Q _6357_/A _6358_/A _6386_/Y VGND VGND VPWR VPWR _6387_/X sky130_fd_sc_hd__a31o_1
XFILLER_115_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3599_ _7072_/Q _5506_/A _4065_/A _6528_/Q _3598_/X VGND VGND VPWR VPWR _3604_/B
+ sky130_fd_sc_hd__a221o_1
X_5338_ _5338_/A0 _5518_/A1 _5343_/S VGND VGND VPWR VPWR _6919_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5269_ _5269_/A0 _5575_/A1 _5271_/S VGND VGND VPWR VPWR _5269_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7008_ _7008_/CLK _7008_/D fanout474/X VGND VGND VPWR VPWR _7008_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4640_ _4341_/X _4640_/B VGND VGND VPWR VPWR _4640_/Y sky130_fd_sc_hd__nand2b_4
XFILLER_30_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4571_ _4988_/A _4808_/B VGND VGND VPWR VPWR _4823_/A sky130_fd_sc_hd__nand2_1
X_6310_ _6637_/Q _5994_/X _6018_/X _6720_/Q VGND VGND VPWR VPWR _6310_/X sky130_fd_sc_hd__a22o_1
X_3522_ _6945_/Q _5362_/A _4077_/A _6539_/Q _3520_/X VGND VGND VPWR VPWR _3529_/B
+ sky130_fd_sc_hd__a221o_1
Xhold705 _4060_/X VGND VGND VPWR VPWR _6520_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap424 _4712_/C VGND VGND VPWR VPWR _4713_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold716 hold716/A VGND VGND VPWR VPWR hold716/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold727 hold727/A VGND VGND VPWR VPWR hold727/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold738 hold738/A VGND VGND VPWR VPWR hold738/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6241_ _7180_/Q _6240_/X _6341_/S VGND VGND VPWR VPWR _6241_/X sky130_fd_sc_hd__mux2_1
Xhold749 hold749/A VGND VGND VPWR VPWR hold749/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3453_ _6930_/Q _5344_/A _5515_/A _7082_/Q _3452_/X VGND VGND VPWR VPWR _3461_/B
+ sky130_fd_sc_hd__a221oi_2
XFILLER_131_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6172_ _6915_/Q _5991_/X _5996_/X _7051_/Q _6171_/X VGND VGND VPWR VPWR _6179_/A
+ sky130_fd_sc_hd__a221o_1
X_3384_ _3384_/A _3384_/B _3383_/Y VGND VGND VPWR VPWR _3385_/B sky130_fd_sc_hd__nor3b_4
Xhold2106 _6793_/Q VGND VGND VPWR VPWR hold457/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2117 hold731/X VGND VGND VPWR VPWR _5186_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5123_ _5123_/A _5123_/B _5123_/C _5123_/D VGND VGND VPWR VPWR _5123_/X sky130_fd_sc_hd__and4_1
Xhold2128 _6879_/Q VGND VGND VPWR VPWR hold640/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2139 hold399/X VGND VGND VPWR VPWR _4061_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1405 _5270_/X VGND VGND VPWR VPWR hold357/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1416 _6478_/Q VGND VGND VPWR VPWR hold394/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1427 _4082_/X VGND VGND VPWR VPWR hold517/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1438 _6703_/Q VGND VGND VPWR VPWR hold140/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5054_ _4638_/Y _4698_/Y _4689_/Y _5063_/B VGND VGND VPWR VPWR _5054_/X sky130_fd_sc_hd__o211a_1
XFILLER_85_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1449 hold469/X VGND VGND VPWR VPWR _5271_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4005_ hold473/X _5196_/A1 _4008_/S VGND VGND VPWR VPWR _6483_/D sky130_fd_sc_hd__mux2_1
XFILLER_52_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5956_ _6573_/Q _5674_/X _5680_/X _6711_/Q VGND VGND VPWR VPWR _5956_/X sky130_fd_sc_hd__a22o_1
XFILLER_40_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4907_ hold908/X _5139_/A _4906_/X VGND VGND VPWR VPWR _6763_/D sky130_fd_sc_hd__o21ba_1
X_5887_ _6635_/Q _5671_/X _5886_/X VGND VGND VPWR VPWR _5887_/X sky130_fd_sc_hd__a21o_1
XFILLER_21_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4838_ _4917_/C _4838_/B VGND VGND VPWR VPWR _4857_/C sky130_fd_sc_hd__nor2_1
XFILLER_178_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4769_ _5011_/A _4729_/A _4514_/B VGND VGND VPWR VPWR _4769_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_193_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6508_ _7136_/CLK _6508_/D fanout475/X VGND VGND VPWR VPWR _6508_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_134_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6439_ _3940_/A1 _6439_/D _6394_/X VGND VGND VPWR VPWR _6439_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold10 hold10/A VGND VGND VPWR VPWR hold10/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold21 hold21/A VGND VGND VPWR VPWR hold21/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold32 hold32/A VGND VGND VPWR VPWR hold32/X sky130_fd_sc_hd__buf_12
XFILLER_75_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold43 hold43/A VGND VGND VPWR VPWR hold43/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold54 hold54/A VGND VGND VPWR VPWR hold54/X sky130_fd_sc_hd__buf_12
XFILLER_75_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold65 hold65/A VGND VGND VPWR VPWR hold65/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_188_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold76 hold76/A VGND VGND VPWR VPWR hold76/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1950 _6580_/Q VGND VGND VPWR VPWR hold732/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold87 hold87/A VGND VGND VPWR VPWR hold87/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1961 hold440/X VGND VGND VPWR VPWR _6493_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_63_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold98 hold98/A VGND VGND VPWR VPWR hold98/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1972 _6623_/Q VGND VGND VPWR VPWR hold571/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1983 _5221_/X VGND VGND VPWR VPWR _6817_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1994 _5490_/X VGND VGND VPWR VPWR _7054_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3240__1 _6656_/CLK VGND VGND VPWR VPWR _6436_/CLK sky130_fd_sc_hd__inv_2
XFILLER_189_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_7 _5326_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5810_ _6938_/Q _5659_/X _5687_/X _6922_/Q VGND VGND VPWR VPWR _5810_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6790_ _6793_/CLK _6790_/D _3959_/B VGND VGND VPWR VPWR _6790_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5741_ _6911_/Q _5670_/X _5685_/X _7071_/Q VGND VGND VPWR VPWR _5741_/X sky130_fd_sc_hd__a22o_1
XFILLER_15_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5672_ _5689_/A _5689_/B _5689_/C VGND VGND VPWR VPWR _5672_/X sky130_fd_sc_hd__and3b_4
XFILLER_30_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4623_ _4625_/A _4971_/A VGND VGND VPWR VPWR _5098_/A sky130_fd_sc_hd__nand2_1
XFILLER_136_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4554_ _4637_/B _4590_/B _5033_/A _4959_/A _4553_/Y VGND VGND VPWR VPWR _4554_/X
+ sky130_fd_sc_hd__a311o_1
Xhold502 hold502/A VGND VGND VPWR VPWR hold502/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold513 hold513/A VGND VGND VPWR VPWR hold513/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold524 hold524/A VGND VGND VPWR VPWR hold524/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3505_ _3540_/A _3553_/B VGND VGND VPWR VPWR _4122_/A sky130_fd_sc_hd__nor2_8
Xhold535 hold535/A VGND VGND VPWR VPWR hold535/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold546 hold546/A VGND VGND VPWR VPWR hold546/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4485_ _4486_/A _4485_/B _4568_/A VGND VGND VPWR VPWR _4621_/A sky130_fd_sc_hd__and3_4
XFILLER_143_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold557 hold557/A VGND VGND VPWR VPWR hold557/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold568 hold568/A VGND VGND VPWR VPWR hold568/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6224_ _6589_/Q _5985_/X _5994_/X _6634_/Q _6218_/X VGND VGND VPWR VPWR _6224_/X
+ sky130_fd_sc_hd__a221o_1
Xhold579 hold579/A VGND VGND VPWR VPWR hold579/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3436_ _6850_/Q hold40/A _3431_/Y _7233_/A VGND VGND VPWR VPWR _3436_/X sky130_fd_sc_hd__a22o_1
XFILLER_106_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ _7130_/Q _5973_/X _5988_/X _6874_/Q _6154_/X VGND VGND VPWR VPWR _6155_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _6972_/Q _5389_/A _5308_/A _6900_/Q _3366_/X VGND VGND VPWR VPWR _3368_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1202 hold496/X VGND VGND VPWR VPWR _5252_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5106_ _4569_/A _4523_/Y _4583_/B _4688_/C _4871_/A VGND VGND VPWR VPWR _5107_/C
+ sky130_fd_sc_hd__o221a_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1213 hold476/X VGND VGND VPWR VPWR _5422_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1224 hold174/X VGND VGND VPWR VPWR _4284_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6086_ _6927_/Q _5982_/X _5987_/X _7111_/Q VGND VGND VPWR VPWR _6086_/X sky130_fd_sc_hd__a22o_1
X_3298_ hold31/X _3425_/A VGND VGND VPWR VPWR _3298_/Y sky130_fd_sc_hd__nand2_8
Xhold1235 _6978_/Q VGND VGND VPWR VPWR hold521/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1246 _5303_/X VGND VGND VPWR VPWR _6888_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1257 hold362/X VGND VGND VPWR VPWR _5352_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5037_ _5117_/C _5151_/B _5037_/C VGND VGND VPWR VPWR _5038_/C sky130_fd_sc_hd__and3_1
XFILLER_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1268 _7192_/Q VGND VGND VPWR VPWR hold865/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1279 hold132/X VGND VGND VPWR VPWR _5234_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6988_ _7116_/CLK _6988_/D fanout455/X VGND VGND VPWR VPWR _6988_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_25_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5939_ _6551_/Q _5673_/X _5937_/X _5938_/X VGND VGND VPWR VPWR _5939_/X sky130_fd_sc_hd__a211o_1
XFILLER_139_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput100 wb_adr_i[10] VGND VGND VPWR VPWR _4345_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput111 wb_adr_i[20] VGND VGND VPWR VPWR _4649_/B sky130_fd_sc_hd__buf_12
XFILLER_76_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput122 wb_adr_i[30] VGND VGND VPWR VPWR input122/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput133 wb_dat_i[10] VGND VGND VPWR VPWR _6367_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput144 wb_dat_i[20] VGND VGND VPWR VPWR _6373_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput155 wb_dat_i[30] VGND VGND VPWR VPWR _6380_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput166 wb_sel_i[1] VGND VGND VPWR VPWR _6356_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2470 _7162_/Q VGND VGND VPWR VPWR _5751_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2481 _6470_/Q VGND VGND VPWR VPWR _3811_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2492 _6217_/X VGND VGND VPWR VPWR _7180_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1780 _6453_/Q VGND VGND VPWR VPWR hold617/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1791 _4197_/X VGND VGND VPWR VPWR _6636_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4270_ _4270_/A0 hold135/X _4273_/S VGND VGND VPWR VPWR _4270_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3221_ _6984_/Q VGND VGND VPWR VPWR _3221_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6911_ _7065_/CLK _6911_/D fanout460/X VGND VGND VPWR VPWR _6911_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6842_ _7008_/CLK _6842_/D fanout474/X VGND VGND VPWR VPWR _6842_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6773_ _6794_/CLK _6773_/D fanout445/X VGND VGND VPWR VPWR _6773_/Q sky130_fd_sc_hd__dfrtp_4
X_3985_ _3985_/A0 _5195_/A1 _3987_/S VGND VGND VPWR VPWR _6453_/D sky130_fd_sc_hd__mux2_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5724_ _7046_/Q _5669_/X _5680_/X _6958_/Q _5723_/X VGND VGND VPWR VPWR _5727_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5655_ _5686_/A _5679_/B _5687_/C VGND VGND VPWR VPWR _5655_/X sky130_fd_sc_hd__and3_4
XFILLER_175_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4606_ _4625_/A _4611_/A VGND VGND VPWR VPWR _5073_/B sky130_fd_sc_hd__nand2_2
XFILLER_175_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5586_ hold976/X hold6/X _5586_/S VGND VGND VPWR VPWR _5586_/X sky130_fd_sc_hd__mux2_1
Xhold310 hold310/A VGND VGND VPWR VPWR hold310/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold321 hold321/A VGND VGND VPWR VPWR hold321/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4537_ _4601_/A _4570_/C _4535_/X _4536_/Y VGND VGND VPWR VPWR _4537_/X sky130_fd_sc_hd__o211a_1
Xhold332 hold332/A VGND VGND VPWR VPWR hold332/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold343 hold343/A VGND VGND VPWR VPWR hold343/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold354 hold354/A VGND VGND VPWR VPWR hold354/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold365 hold978/X VGND VGND VPWR VPWR hold979/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold376 hold376/A VGND VGND VPWR VPWR hold376/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4468_ _4638_/B _4488_/B VGND VGND VPWR VPWR _4601_/A sky130_fd_sc_hd__nand2_8
Xhold387 hold983/X VGND VGND VPWR VPWR hold984/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold398 hold398/A VGND VGND VPWR VPWR _6523_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6207_ _7100_/Q _5984_/X _6015_/X _7020_/Q VGND VGND VPWR VPWR _6207_/X sky130_fd_sc_hd__a22o_1
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3419_ _7003_/Q _5425_/A _5506_/A _7075_/Q VGND VGND VPWR VPWR _3419_/X sky130_fd_sc_hd__a22o_1
X_7187_ _7194_/CLK _7187_/D VGND VGND VPWR VPWR _7187_/Q sky130_fd_sc_hd__dfxtp_1
X_4399_ _4637_/D _4575_/C VGND VGND VPWR VPWR _4590_/B sky130_fd_sc_hd__and2b_4
XFILLER_58_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6138_ _6131_/X _6133_/X _6138_/C _6339_/B VGND VGND VPWR VPWR _6139_/C sky130_fd_sc_hd__and4bb_1
Xhold1010 _7229_/A VGND VGND VPWR VPWR hold16/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1021 _7100_/Q VGND VGND VPWR VPWR hold71/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1032 _5267_/X VGND VGND VPWR VPWR hold10/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_133_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1043 _5441_/X VGND VGND VPWR VPWR _7011_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6069_ _6911_/Q _5991_/X _6018_/X _6967_/Q VGND VGND VPWR VPWR _6069_/X sky130_fd_sc_hd__a22o_1
Xhold1054 _7115_/Q VGND VGND VPWR VPWR hold364/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_133_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1065 _5197_/X VGND VGND VPWR VPWR _6800_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_133_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1076 _5495_/X VGND VGND VPWR VPWR _7059_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1087 _5387_/X VGND VGND VPWR VPWR _6963_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_205 _6818_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1098 hold408/X VGND VGND VPWR VPWR _5513_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_26_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3770_ _3770_/A _3770_/B _3770_/C VGND VGND VPWR VPWR _3803_/A sky130_fd_sc_hd__and3_2
XFILLER_32_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5440_ _5440_/A0 _5575_/A1 _5442_/S VGND VGND VPWR VPWR _7010_/D sky130_fd_sc_hd__mux2_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5371_ _5371_/A _5569_/B VGND VGND VPWR VPWR _5379_/S sky130_fd_sc_hd__and2_4
XFILLER_114_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7110_ _7127_/CLK _7110_/D fanout474/X VGND VGND VPWR VPWR _7110_/Q sky130_fd_sc_hd__dfstp_1
X_4322_ _4322_/A _5220_/C VGND VGND VPWR VPWR _4327_/S sky130_fd_sc_hd__and2_4
XFILLER_99_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7041_ _7121_/CLK _7041_/D fanout473/X VGND VGND VPWR VPWR _7041_/Q sky130_fd_sc_hd__dfrtp_4
X_4253_ _4253_/A0 _4337_/A1 _4255_/S VGND VGND VPWR VPWR _4253_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3204_ _7120_/Q VGND VGND VPWR VPWR _3204_/Y sky130_fd_sc_hd__inv_2
X_4184_ _4184_/A0 _5193_/A1 _4187_/S VGND VGND VPWR VPWR _4184_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_4__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7203_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_83_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6825_ _7136_/CLK _6825_/D fanout476/X VGND VGND VPWR VPWR _7230_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6756_ _6760_/CLK _6756_/D _6433_/A VGND VGND VPWR VPWR _6756_/Q sky130_fd_sc_hd__dfrtp_4
X_3968_ _3968_/A _3975_/B VGND VGND VPWR VPWR _6679_/D sky130_fd_sc_hd__and2_1
XFILLER_149_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5707_ _6837_/Q _5707_/B VGND VGND VPWR VPWR _5707_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6687_ _6794_/CLK _6687_/D fanout443/X VGND VGND VPWR VPWR _6687_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3899_ _4345_/A _4345_/B _3899_/C _3899_/D VGND VGND VPWR VPWR _3900_/D sky130_fd_sc_hd__and4bb_2
XFILLER_137_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_494 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5638_ _6014_/A _6017_/B _6019_/B VGND VGND VPWR VPWR _5638_/X sky130_fd_sc_hd__and3_4
XFILLER_164_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5569_ _5569_/A _5569_/B VGND VGND VPWR VPWR _5577_/S sky130_fd_sc_hd__and2_4
XFILLER_117_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold140 hold140/A VGND VGND VPWR VPWR hold140/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold151 hold151/A VGND VGND VPWR VPWR hold151/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold162 hold162/A VGND VGND VPWR VPWR hold162/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold173 hold173/A VGND VGND VPWR VPWR hold173/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold184 hold184/A VGND VGND VPWR VPWR hold184/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold195 hold195/A VGND VGND VPWR VPWR hold195/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4940_ _4462_/Y _4935_/X _4796_/A VGND VGND VPWR VPWR _5162_/A sky130_fd_sc_hd__o21a_1
XFILLER_92_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4871_ _4871_/A _4871_/B _4871_/C _4871_/D VGND VGND VPWR VPWR _4872_/D sky130_fd_sc_hd__and4_1
XFILLER_178_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_551 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6610_ _6759_/CLK _6610_/D fanout449/X VGND VGND VPWR VPWR _6610_/Q sky130_fd_sc_hd__dfrtp_4
X_3822_ _6465_/Q _6464_/Q _3834_/S VGND VGND VPWR VPWR _3826_/B sky130_fd_sc_hd__and3_1
X_6541_ _6568_/CLK _6541_/D VGND VGND VPWR VPWR _6541_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3753_ _6821_/Q _5226_/A _5226_/B _3315_/Y input34/X VGND VGND VPWR VPWR _3753_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_186_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6472_ _6809_/CLK _6472_/D fanout444/X VGND VGND VPWR VPWR _6472_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_146_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3684_ _3684_/A _3684_/B _3684_/C VGND VGND VPWR VPWR _3704_/A sky130_fd_sc_hd__nor3_1
XFILLER_173_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5423_ _5423_/A0 _5576_/A1 _5424_/S VGND VGND VPWR VPWR _5423_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput201 _3206_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[33] sky130_fd_sc_hd__buf_12
Xoutput212 _3231_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[9] sky130_fd_sc_hd__buf_12
XFILLER_160_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput223 _7218_/X VGND VGND VPWR VPWR mgmt_gpio_out[20] sky130_fd_sc_hd__buf_12
Xoutput234 _7228_/X VGND VGND VPWR VPWR mgmt_gpio_out[30] sky130_fd_sc_hd__buf_12
X_5354_ hold784/X _5570_/A1 _5361_/S VGND VGND VPWR VPWR _5354_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput245 _3942_/X VGND VGND VPWR VPWR mgmt_gpio_out[6] sky130_fd_sc_hd__buf_12
XFILLER_114_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput256 _3963_/Y VGND VGND VPWR VPWR pad_flash_io1_oeb sky130_fd_sc_hd__buf_12
Xoutput267 _6782_/Q VGND VGND VPWR VPWR pll_ena sky130_fd_sc_hd__buf_12
XFILLER_142_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4305_ _4305_/A0 _5208_/A1 _4309_/S VGND VGND VPWR VPWR _6732_/D sky130_fd_sc_hd__mux2_1
Xoutput278 _6795_/Q VGND VGND VPWR VPWR pll_trim[16] sky130_fd_sc_hd__buf_12
Xoutput289 _6481_/Q VGND VGND VPWR VPWR pll_trim[2] sky130_fd_sc_hd__buf_12
X_5285_ _5285_/A0 _5555_/A1 _5289_/S VGND VGND VPWR VPWR _5285_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7024_ _7126_/CLK _7024_/D fanout480/X VGND VGND VPWR VPWR _7024_/Q sky130_fd_sc_hd__dfrtp_4
X_4236_ _4236_/A0 _4235_/X _4240_/S VGND VGND VPWR VPWR _6665_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4167_ hold334/X _4337_/A1 _4169_/S VGND VGND VPWR VPWR _6611_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4098_ _6678_/Q _6346_/B VGND VGND VPWR VPWR _4106_/S sky130_fd_sc_hd__nand2_8
XFILLER_71_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_4_csclk _6727_/CLK VGND VGND VPWR VPWR _6759_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6808_ _6808_/CLK _6808_/D fanout440/X VGND VGND VPWR VPWR _6808_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6739_ _6822_/CLK _6739_/D fanout451/X VGND VGND VPWR VPWR _6739_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_136_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout450 fanout482/X VGND VGND VPWR VPWR fanout450/X sky130_fd_sc_hd__clkbuf_16
XFILLER_120_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout461 _6432_/A VGND VGND VPWR VPWR _6433_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_171_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout472 fanout481/X VGND VGND VPWR VPWR fanout472/X sky130_fd_sc_hd__buf_12
XFILLER_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout483 input164/X VGND VGND VPWR VPWR _6346_/B sky130_fd_sc_hd__buf_12
XFILLER_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold909 hold909/A VGND VGND VPWR VPWR hold909/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_6_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5070_ _4476_/X _4568_/Y _4920_/B _4972_/Y VGND VGND VPWR VPWR _5135_/C sky130_fd_sc_hd__o211a_1
XFILLER_150_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1609 hold512/X VGND VGND VPWR VPWR _5397_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4021_ _4021_/A0 _4020_/X _4029_/S VGND VGND VPWR VPWR _4021_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5972_ _7152_/Q _7151_/Q VGND VGND VPWR VPWR _6018_/B sky130_fd_sc_hd__nor2_8
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4923_ _4633_/B _4691_/Y _4846_/X _4894_/B VGND VGND VPWR VPWR _5052_/B sky130_fd_sc_hd__o211a_1
XFILLER_33_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4854_ _4569_/A _4655_/A _4590_/Y _4688_/C VGND VGND VPWR VPWR _4871_/B sky130_fd_sc_hd__o22a_1
XFILLER_178_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3805_ _3805_/A1 _3739_/S _3803_/Y _3804_/X VGND VGND VPWR VPWR _6774_/D sky130_fd_sc_hd__a22o_1
X_4785_ _4718_/A _4463_/B _4570_/D _4691_/Y _4947_/A VGND VGND VPWR VPWR _4785_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_165_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3736_ _3707_/X _3736_/B _3736_/C _3736_/D VGND VGND VPWR VPWR _3737_/B sky130_fd_sc_hd__and4b_2
X_6524_ _7138_/CLK _6524_/D fanout480/X VGND VGND VPWR VPWR _6524_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3667_ _6855_/Q _5263_/A _4334_/A _6759_/Q VGND VGND VPWR VPWR _3667_/X sky130_fd_sc_hd__a22o_1
X_6455_ _6656_/CLK _6455_/D _6405_/X VGND VGND VPWR VPWR _6455_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_173_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5406_ _5406_/A0 _5559_/A1 _5406_/S VGND VGND VPWR VPWR _6980_/D sky130_fd_sc_hd__mux2_1
X_6386_ _3969_/A _6356_/Y _6358_/Y _3967_/A VGND VGND VPWR VPWR _6386_/Y sky130_fd_sc_hd__o22ai_1
X_3598_ _7048_/Q _5479_/A _5169_/A _6772_/Q VGND VGND VPWR VPWR _3598_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5337_ hold766/X _5580_/A1 _5343_/S VGND VGND VPWR VPWR _6918_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5268_ hold99/X hold95/X _5271_/S VGND VGND VPWR VPWR _5268_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7007_ _7079_/CLK _7007_/D fanout470/X VGND VGND VPWR VPWR _7007_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_102_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4219_ _6682_/Q _4220_/B VGND VGND VPWR VPWR _4836_/A sky130_fd_sc_hd__and2b_4
X_5199_ hold376/X _5559_/A1 _5199_/S VGND VGND VPWR VPWR _6802_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4570_ _4570_/A _4570_/B _4570_/C _4570_/D VGND VGND VPWR VPWR _4570_/X sky130_fd_sc_hd__and4_1
X_3521_ _3540_/A _3533_/B VGND VGND VPWR VPWR _4077_/A sky130_fd_sc_hd__nor2_8
Xhold706 hold706/A VGND VGND VPWR VPWR hold706/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap425 _4712_/C VGND VGND VPWR VPWR _4751_/C sky130_fd_sc_hd__buf_2
Xhold717 hold717/A VGND VGND VPWR VPWR hold717/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold728 hold728/A VGND VGND VPWR VPWR hold728/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6240_ _6525_/Q _6339_/B _6239_/X VGND VGND VPWR VPWR _6240_/X sky130_fd_sc_hd__o21ba_1
X_3452_ _6866_/Q _5272_/A _5389_/A _6970_/Q _3451_/X VGND VGND VPWR VPWR _3452_/X
+ sky130_fd_sc_hd__a221o_1
Xhold739 hold739/A VGND VGND VPWR VPWR hold739/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_170_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6171_ _7027_/Q _5971_/X _6014_/X _6995_/Q VGND VGND VPWR VPWR _6171_/X sky130_fd_sc_hd__a22o_1
X_3383_ _3383_/A _3383_/B _3383_/C _3383_/D VGND VGND VPWR VPWR _3383_/Y sky130_fd_sc_hd__nor4_1
XFILLER_130_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2107 _5189_/X VGND VGND VPWR VPWR _6793_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5122_ _4491_/Y _4523_/Y _4583_/B _4676_/Y _4872_/C VGND VGND VPWR VPWR _5123_/D
+ sky130_fd_sc_hd__o221a_1
Xhold2118 _5186_/X VGND VGND VPWR VPWR _6790_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2129 hold640/X VGND VGND VPWR VPWR _5293_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1406 _6745_/Q VGND VGND VPWR VPWR hold327/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1417 _6720_/Q VGND VGND VPWR VPWR hold326/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5053_ _5112_/B _5121_/C _5112_/C _5107_/B VGND VGND VPWR VPWR _5059_/B sky130_fd_sc_hd__and4_1
Xhold1428 _7206_/A VGND VGND VPWR VPWR hold649/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1439 hold140/X VGND VGND VPWR VPWR _4270_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4004_ hold618/X _5195_/A1 _4008_/S VGND VGND VPWR VPWR _6482_/D sky130_fd_sc_hd__mux2_1
XFILLER_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5955_ _6696_/Q _5658_/X _5664_/X _6761_/Q VGND VGND VPWR VPWR _5955_/X sky130_fd_sc_hd__a22o_1
X_4906_ _4906_/A _4906_/B _4906_/C _4906_/D VGND VGND VPWR VPWR _4906_/X sky130_fd_sc_hd__and4_1
X_5886_ _6748_/Q _5666_/X _5689_/X _6625_/Q VGND VGND VPWR VPWR _5886_/X sky130_fd_sc_hd__a22o_1
XFILLER_138_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4837_ _5114_/A _4837_/B VGND VGND VPWR VPWR _5044_/B sky130_fd_sc_hd__and2_1
XFILLER_193_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4768_ _5033_/A _4955_/D VGND VGND VPWR VPWR _5089_/A sky130_fd_sc_hd__nand2_1
XFILLER_107_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6507_ _7138_/CLK _6507_/D fanout478/X VGND VGND VPWR VPWR _6507_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3719_ _6902_/Q _5317_/A _5281_/A _6870_/Q VGND VGND VPWR VPWR _3719_/X sky130_fd_sc_hd__a22o_1
X_4699_ _4710_/A _4702_/B VGND VGND VPWR VPWR _4699_/Y sky130_fd_sc_hd__nand2_1
XFILLER_106_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6438_ _3940_/A1 _6438_/D _6393_/X VGND VGND VPWR VPWR _6438_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6369_ _6368_/X _6369_/A1 _6384_/S VGND VGND VPWR VPWR _7197_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_22_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7105_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold11 hold11/A VGND VGND VPWR VPWR hold11/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold22 hold22/A VGND VGND VPWR VPWR hold22/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold33 hold33/A VGND VGND VPWR VPWR hold33/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold44 hold44/A VGND VGND VPWR VPWR hold44/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold55 hold55/A VGND VGND VPWR VPWR hold55/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1940 _5356_/X VGND VGND VPWR VPWR _6935_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold66 hold66/A VGND VGND VPWR VPWR hold66/X sky130_fd_sc_hd__buf_4
Xhold1951 hold732/X VGND VGND VPWR VPWR _4130_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold77 hold77/A VGND VGND VPWR VPWR hold77/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold88 hold88/A VGND VGND VPWR VPWR hold88/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1962 _6698_/Q VGND VGND VPWR VPWR hold746/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold99 hold99/A VGND VGND VPWR VPWR hold99/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1973 hold571/X VGND VGND VPWR VPWR _4181_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xclkbuf_leaf_37_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7131_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_90_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1984 _7078_/Q VGND VGND VPWR VPWR hold694/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1995 _7064_/Q VGND VGND VPWR VPWR hold708/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] VGND VGND VPWR VPWR clkbuf_0_mgmt_gpio_in[4]/X
+ sky130_fd_sc_hd__clkbuf_16
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_8 hold67/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5740_ _7063_/Q _5671_/X _5733_/X _5735_/X _5739_/X VGND VGND VPWR VPWR _5740_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5671_ _5689_/A _5679_/B _5689_/C VGND VGND VPWR VPWR _5671_/X sky130_fd_sc_hd__and3_4
XFILLER_187_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4622_ _4894_/B _4622_/B _4622_/C _5052_/A VGND VGND VPWR VPWR _4622_/X sky130_fd_sc_hd__and4_1
XFILLER_175_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4553_ _4514_/Y _4526_/X _4553_/C _5090_/C VGND VGND VPWR VPWR _4553_/Y sky130_fd_sc_hd__nand4bb_1
Xhold503 hold503/A VGND VGND VPWR VPWR hold503/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold514 hold514/A VGND VGND VPWR VPWR hold514/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3504_ _3540_/A _3549_/B VGND VGND VPWR VPWR _4146_/A sky130_fd_sc_hd__nor2_4
Xhold525 hold525/A VGND VGND VPWR VPWR hold525/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold536 hold536/A VGND VGND VPWR VPWR hold536/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4484_ _4607_/B _4611_/A VGND VGND VPWR VPWR _4531_/B sky130_fd_sc_hd__nand2_2
Xhold547 hold547/A VGND VGND VPWR VPWR hold547/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold558 hold558/A VGND VGND VPWR VPWR hold558/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6223_ _6702_/Q _5977_/X _5984_/X _6614_/Q _6222_/X VGND VGND VPWR VPWR _6238_/B
+ sky130_fd_sc_hd__a221o_1
X_3435_ input17/X _3310_/Y _3357_/Y _6484_/Q VGND VGND VPWR VPWR _3435_/X sky130_fd_sc_hd__a22o_1
Xhold569 hold569/A VGND VGND VPWR VPWR hold569/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6154_ _6962_/Q _5992_/X _6012_/X _7002_/Q _6153_/X VGND VGND VPWR VPWR _6154_/X
+ sky130_fd_sc_hd__a221o_1
X_3366_ _7140_/Q hold33/A _5335_/A _6924_/Q VGND VGND VPWR VPWR _3366_/X sky130_fd_sc_hd__a22o_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1203 _7094_/Q VGND VGND VPWR VPWR hold222/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_112_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5105_ _5101_/X _5135_/D _5062_/A _5071_/Y VGND VGND VPWR VPWR _5119_/B sky130_fd_sc_hd__a211o_1
Xhold1214 _5422_/X VGND VGND VPWR VPWR _6994_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6085_ _6863_/Q _5999_/X _6019_/X _6983_/Q _6084_/X VGND VGND VPWR VPWR _6088_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_100_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3297_ hold38/X hold66/A VGND VGND VPWR VPWR _3297_/Y sky130_fd_sc_hd__nor2_2
Xhold1225 _4284_/X VGND VGND VPWR VPWR _6715_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1236 hold521/X VGND VGND VPWR VPWR _5404_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1247 _6613_/Q VGND VGND VPWR VPWR hold117/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5036_ _4812_/A _4724_/C _5033_/A VGND VGND VPWR VPWR _5037_/C sky130_fd_sc_hd__o21ai_1
Xhold1258 _5352_/X VGND VGND VPWR VPWR _6932_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1269 hold865/X VGND VGND VPWR VPWR hold211/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6987_ _7123_/CLK _6987_/D fanout479/X VGND VGND VPWR VPWR _6987_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_40_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5938_ _6612_/Q _5660_/X _5669_/X _6652_/Q VGND VGND VPWR VPWR _5938_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5869_ _5869_/A _5869_/B _5869_/C VGND VGND VPWR VPWR _5869_/Y sky130_fd_sc_hd__nor3_1
XFILLER_178_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput101 wb_adr_i[11] VGND VGND VPWR VPWR _4345_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput112 wb_adr_i[21] VGND VGND VPWR VPWR _4720_/C sky130_fd_sc_hd__buf_6
XFILLER_103_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput123 wb_adr_i[31] VGND VGND VPWR VPWR input123/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput134 wb_dat_i[11] VGND VGND VPWR VPWR _6370_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput145 wb_dat_i[21] VGND VGND VPWR VPWR _6376_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2460 _7164_/Q VGND VGND VPWR VPWR _5816_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput156 wb_dat_i[31] VGND VGND VPWR VPWR _6382_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput167 wb_sel_i[2] VGND VGND VPWR VPWR _6358_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2471 _7171_/Q VGND VGND VPWR VPWR _5969_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2482 _7169_/Q VGND VGND VPWR VPWR _5904_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2493 _7160_/Q VGND VGND VPWR VPWR _5709_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1770 hold524/X VGND VGND VPWR VPWR _3981_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1781 hold617/X VGND VGND VPWR VPWR _3985_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1792 _6454_/Q VGND VGND VPWR VPWR hold470/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3220_ _6992_/Q VGND VGND VPWR VPWR _3220_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_140_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_3__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7183_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_121_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6910_ _7126_/CLK _6910_/D fanout475/X VGND VGND VPWR VPWR _6910_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_47_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6841_ _6945_/CLK _6841_/D _6399_/A VGND VGND VPWR VPWR _6841_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6772_ _6794_/CLK _6772_/D fanout445/X VGND VGND VPWR VPWR _6772_/Q sky130_fd_sc_hd__dfrtp_4
X_3984_ _3984_/A0 hold170/X _3996_/S VGND VGND VPWR VPWR _3984_/X sky130_fd_sc_hd__mux2_2
X_5723_ _7014_/Q _5664_/X _5668_/X _7054_/Q VGND VGND VPWR VPWR _5723_/X sky130_fd_sc_hd__a22o_1
X_5654_ _7148_/Q _7149_/Q VGND VGND VPWR VPWR _5687_/C sky130_fd_sc_hd__and2b_4
XFILLER_176_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4605_ _4580_/Y _4969_/B _4584_/Y _4604_/X VGND VGND VPWR VPWR _4609_/C sky130_fd_sc_hd__a31o_1
XFILLER_191_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5585_ _5585_/A0 _5585_/A1 _5586_/S VGND VGND VPWR VPWR _5585_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold300 _5240_/X VGND VGND VPWR VPWR _6832_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold311 hold311/A VGND VGND VPWR VPWR hold311/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4536_ _4607_/B _4562_/A VGND VGND VPWR VPWR _4536_/Y sky130_fd_sc_hd__nand2_1
Xhold322 hold322/A VGND VGND VPWR VPWR hold322/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold333 hold333/A VGND VGND VPWR VPWR hold333/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold344 hold344/A VGND VGND VPWR VPWR hold344/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold355 _4052_/X VGND VGND VPWR VPWR _6513_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold366 hold366/A VGND VGND VPWR VPWR hold366/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4467_ _4638_/B _4488_/B VGND VGND VPWR VPWR _4934_/B sky130_fd_sc_hd__and2_4
Xhold377 hold377/A VGND VGND VPWR VPWR hold377/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold388 hold388/A VGND VGND VPWR VPWR hold388/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6206_ _7052_/Q _5996_/X _6005_/X _6948_/Q _6205_/X VGND VGND VPWR VPWR _6206_/X
+ sky130_fd_sc_hd__a221o_1
Xhold399 hold399/A VGND VGND VPWR VPWR hold399/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3418_ _6923_/Q _5335_/A _5353_/A _6939_/Q _3417_/X VGND VGND VPWR VPWR _3421_/C
+ sky130_fd_sc_hd__a221o_2
X_7186_ _7186_/CLK _7186_/D _6346_/B VGND VGND VPWR VPWR _7186_/Q sky130_fd_sc_hd__dfrtp_4
X_4398_ _4637_/A _4637_/B VGND VGND VPWR VPWR _4495_/B sky130_fd_sc_hd__nand2_8
XFILLER_86_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3349_ _3349_/A _3470_/A VGND VGND VPWR VPWR _5407_/A sky130_fd_sc_hd__nor2_8
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1000 hold381/X VGND VGND VPWR VPWR _5431_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6137_ _7041_/Q _6016_/X _6134_/X _6136_/X VGND VGND VPWR VPWR _6138_/C sky130_fd_sc_hd__a211oi_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1011 hold16/X VGND VGND VPWR VPWR _4249_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1022 hold71/X VGND VGND VPWR VPWR _5541_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_58_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1033 hold10/X VGND VGND VPWR VPWR _6856_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1044 _7027_/Q VGND VGND VPWR VPWR hold389/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6068_ _6855_/Q _5983_/X _6005_/X _6943_/Q VGND VGND VPWR VPWR _6068_/X sky130_fd_sc_hd__a22o_1
Xhold1055 hold364/X VGND VGND VPWR VPWR _5558_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1066 _7058_/Q VGND VGND VPWR VPWR hold429/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_100_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1077 _6986_/Q VGND VGND VPWR VPWR hold433/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_100_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1088 _7228_/A VGND VGND VPWR VPWR hold386/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5019_ _4826_/B _4990_/Y _5018_/X _4683_/A VGND VGND VPWR VPWR _5022_/C sky130_fd_sc_hd__o2bb2a_1
XFILLER_73_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1099 _5513_/X VGND VGND VPWR VPWR _7075_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_206 _3881_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2290 hold803/X VGND VGND VPWR VPWR _4287_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_64_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5370_ _5370_/A0 hold6/X _5370_/S VGND VGND VPWR VPWR _5370_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4321_ _4321_/A0 _4339_/A1 _4321_/S VGND VGND VPWR VPWR _6746_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4252_ _4252_/A0 _5186_/A1 _4255_/S VGND VGND VPWR VPWR _4252_/X sky130_fd_sc_hd__mux2_1
X_7040_ _7126_/CLK _7040_/D fanout475/X VGND VGND VPWR VPWR _7040_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_113_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3203_ _7128_/Q VGND VGND VPWR VPWR _3203_/Y sky130_fd_sc_hd__inv_2
X_4183_ _4183_/A0 _5221_/A1 _4187_/S VGND VGND VPWR VPWR _4183_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6824_ _6826_/CLK _6824_/D _6414_/A VGND VGND VPWR VPWR _6824_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6755_ _6760_/CLK _6755_/D _6432_/A VGND VGND VPWR VPWR _6755_/Q sky130_fd_sc_hd__dfrtp_4
X_3967_ _3967_/A _3969_/B VGND VGND VPWR VPWR _6681_/D sky130_fd_sc_hd__nor2_1
X_5706_ _6973_/Q _5660_/X _5699_/X _5701_/X _5705_/X VGND VGND VPWR VPWR _5706_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_50_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6686_ _7152_/CLK _6686_/D fanout484/X VGND VGND VPWR VPWR _6686_/Q sky130_fd_sc_hd__dfrtp_4
X_3898_ _3898_/A _3898_/B _3898_/C VGND VGND VPWR VPWR _3899_/D sky130_fd_sc_hd__and3_1
XFILLER_12_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5637_ _5637_/A _7156_/Q VGND VGND VPWR VPWR _6019_/B sky130_fd_sc_hd__nor2_8
XFILLER_148_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5568_ _5568_/A0 _5577_/A1 _5568_/S VGND VGND VPWR VPWR _5568_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold130 hold130/A VGND VGND VPWR VPWR hold130/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold141 hold141/A VGND VGND VPWR VPWR hold141/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4519_ _4637_/D _4522_/B VGND VGND VPWR VPWR _4917_/D sky130_fd_sc_hd__nor2_4
Xhold152 hold152/A VGND VGND VPWR VPWR hold152/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold163 hold163/A VGND VGND VPWR VPWR _6668_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5499_ _5499_/A0 _5499_/A1 _5505_/S VGND VGND VPWR VPWR _5499_/X sky130_fd_sc_hd__mux2_1
Xhold174 hold174/A VGND VGND VPWR VPWR hold174/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold185 hold185/A VGND VGND VPWR VPWR hold185/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold196 hold196/A VGND VGND VPWR VPWR hold853/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7169_ _7186_/CLK _7169_/D fanout466/X VGND VGND VPWR VPWR _7169_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4870_ _4870_/A _4870_/B _4870_/C _4870_/D VGND VGND VPWR VPWR _4871_/D sky130_fd_sc_hd__and4_1
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3821_ _6463_/Q _6462_/Q _6461_/Q _6460_/Q VGND VGND VPWR VPWR _3834_/S sky130_fd_sc_hd__and4_1
XFILLER_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6540_ _6568_/CLK _6540_/D VGND VGND VPWR VPWR _6540_/Q sky130_fd_sc_hd__dfxtp_1
X_3752_ _6909_/Q _5326_/A _4316_/A _6742_/Q _3751_/X VGND VGND VPWR VPWR _3759_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6471_ _6809_/CLK _6471_/D fanout444/X VGND VGND VPWR VPWR _6471_/Q sky130_fd_sc_hd__dfstp_2
X_3683_ input12/X _3310_/Y _5169_/A _6770_/Q _3682_/X VGND VGND VPWR VPWR _3684_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_173_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5422_ _5422_/A0 _5575_/A1 _5424_/S VGND VGND VPWR VPWR _5422_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput202 _3205_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[34] sky130_fd_sc_hd__buf_12
Xoutput213 _3946_/X VGND VGND VPWR VPWR mgmt_gpio_out[0] sky130_fd_sc_hd__buf_12
Xoutput224 _7219_/X VGND VGND VPWR VPWR mgmt_gpio_out[21] sky130_fd_sc_hd__buf_12
XFILLER_99_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput235 _7229_/X VGND VGND VPWR VPWR mgmt_gpio_out[31] sky130_fd_sc_hd__buf_12
X_5353_ _5353_/A _5551_/B VGND VGND VPWR VPWR _5361_/S sky130_fd_sc_hd__and2_4
Xoutput246 _7211_/X VGND VGND VPWR VPWR mgmt_gpio_out[7] sky130_fd_sc_hd__buf_12
Xoutput257 _6792_/Q VGND VGND VPWR VPWR pll90_sel[0] sky130_fd_sc_hd__buf_12
X_4304_ _4304_/A _5220_/C VGND VGND VPWR VPWR _4309_/S sky130_fd_sc_hd__and2_4
Xoutput268 _6789_/Q VGND VGND VPWR VPWR pll_sel[0] sky130_fd_sc_hd__buf_12
Xoutput279 _6796_/Q VGND VGND VPWR VPWR pll_trim[17] sky130_fd_sc_hd__buf_12
XFILLER_87_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5284_ _5284_/A0 _5572_/A1 _5289_/S VGND VGND VPWR VPWR _5284_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7023_ _7139_/CLK _7023_/D fanout478/X VGND VGND VPWR VPWR _7023_/Q sky130_fd_sc_hd__dfrtp_4
X_4235_ _5242_/A0 _5503_/A1 _4239_/S VGND VGND VPWR VPWR _4235_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4166_ _4166_/A0 _5193_/A1 _4169_/S VGND VGND VPWR VPWR _6610_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4097_ _4097_/A0 _5196_/A1 _4097_/S VGND VGND VPWR VPWR _6552_/D sky130_fd_sc_hd__mux2_1
XFILLER_70_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6807_ _6833_/CLK _6807_/D fanout454/X VGND VGND VPWR VPWR _6807_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_24_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4999_ _5010_/B _4999_/B _5139_/B _4999_/D VGND VGND VPWR VPWR _5000_/B sky130_fd_sc_hd__and4_1
XFILLER_139_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6738_ _6822_/CLK _6738_/D fanout451/X VGND VGND VPWR VPWR _6738_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6669_ _7016_/CLK _6669_/D fanout476/X VGND VGND VPWR VPWR _7223_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout440 _3959_/B VGND VGND VPWR VPWR fanout440/X sky130_fd_sc_hd__buf_8
Xfanout451 fanout453/X VGND VGND VPWR VPWR fanout451/X sky130_fd_sc_hd__buf_12
Xfanout462 fanout466/X VGND VGND VPWR VPWR _6432_/A sky130_fd_sc_hd__buf_6
Xfanout473 fanout481/X VGND VGND VPWR VPWR fanout473/X sky130_fd_sc_hd__buf_12
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout484 input164/X VGND VGND VPWR VPWR fanout484/X sky130_fd_sc_hd__buf_8
XFILLER_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4020_ _4051_/A0 _5555_/A1 _4047_/C VGND VGND VPWR VPWR _4020_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5971_ _6015_/B _6014_/A _6019_/B VGND VGND VPWR VPWR _5971_/X sky130_fd_sc_hd__and3_4
X_4922_ _4922_/A _4922_/B _4922_/C VGND VGND VPWR VPWR _4925_/A sky130_fd_sc_hd__and3_1
XFILLER_80_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4853_ _4510_/A _4655_/A _4590_/Y _4995_/A VGND VGND VPWR VPWR _4924_/C sky130_fd_sc_hd__o22a_1
XFILLER_178_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3804_ _6448_/Q _6656_/Q _3857_/B VGND VGND VPWR VPWR _3804_/X sky130_fd_sc_hd__and3_1
X_4784_ _4466_/A _4477_/Y _4510_/B _4736_/Y _4407_/Y VGND VGND VPWR VPWR _4784_/X
+ sky130_fd_sc_hd__o32a_1
X_6523_ _6523_/CLK _6523_/D fanout481/X VGND VGND VPWR VPWR _6523_/Q sky130_fd_sc_hd__dfrtp_1
X_3735_ _3735_/A _3735_/B _3735_/C _3735_/D VGND VGND VPWR VPWR _3735_/Y sky130_fd_sc_hd__nor4_1
XFILLER_146_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6454_ _6792_/CLK _6454_/D fanout442/X VGND VGND VPWR VPWR _6454_/Q sky130_fd_sc_hd__dfrtp_4
X_3666_ _7127_/Q _5569_/A _5344_/A _6927_/Q _3665_/X VGND VGND VPWR VPWR _3673_/A
+ sky130_fd_sc_hd__a221o_1
X_5405_ hold374/X _5576_/A1 _5406_/S VGND VGND VPWR VPWR _5405_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6385_ _3184_/Y _3189_/Y _6385_/A3 _4836_/A _4222_/Y VGND VGND VPWR VPWR _7203_/D
+ sky130_fd_sc_hd__a41o_2
XFILLER_161_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3597_ _6474_/Q _3339_/Y _4322_/A _6750_/Q _3596_/X VGND VGND VPWR VPWR _3604_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5336_ hold678/X _5561_/A1 _5343_/S VGND VGND VPWR VPWR _6917_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5267_ _6856_/Q _5267_/A1 _5271_/S VGND VGND VPWR VPWR _5267_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7006_ _7103_/CLK _7006_/D fanout472/X VGND VGND VPWR VPWR _7006_/Q sky130_fd_sc_hd__dfstp_4
X_4218_ _6684_/Q _6685_/Q _6686_/Q VGND VGND VPWR VPWR _4218_/Y sky130_fd_sc_hd__nor3_4
X_5198_ hold105/X hold78/X _5198_/S VGND VGND VPWR VPWR _5198_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4149_ hold572/X _5187_/A1 _4151_/S VGND VGND VPWR VPWR _6596_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_747 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3520_ _7137_/Q hold33/A _5290_/A _6881_/Q VGND VGND VPWR VPWR _3520_/X sky130_fd_sc_hd__a22o_1
Xhold707 hold707/A VGND VGND VPWR VPWR hold707/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap426 _4672_/B VGND VGND VPWR VPWR _4712_/C sky130_fd_sc_hd__clkbuf_2
Xhold718 hold718/A VGND VGND VPWR VPWR hold718/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold729 _5208_/X VGND VGND VPWR VPWR _6808_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3451_ _6978_/Q _5398_/A _5524_/A _7090_/Q _3450_/X VGND VGND VPWR VPWR _3451_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3382_ _6932_/Q _5344_/A _5263_/A _6860_/Q _3381_/X VGND VGND VPWR VPWR _3383_/D
+ sky130_fd_sc_hd__a221o_1
X_6170_ _7099_/Q _5984_/X _5997_/X _6955_/Q _6169_/X VGND VGND VPWR VPWR _6170_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_124_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_3_csclk _6727_/CLK VGND VGND VPWR VPWR _6750_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_130_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2108 _6861_/Q VGND VGND VPWR VPWR hold782/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_124_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5121_ _5121_/A _5121_/B _5121_/C _5121_/D VGND VGND VPWR VPWR _5121_/X sky130_fd_sc_hd__and4_1
XFILLER_97_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2119 _7081_/Q VGND VGND VPWR VPWR hold740/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1407 hold327/X VGND VGND VPWR VPWR _4320_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_38_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1418 hold326/X VGND VGND VPWR VPWR _4290_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5052_ _5052_/A _5052_/B _5052_/C VGND VGND VPWR VPWR _5107_/B sky130_fd_sc_hd__and3_1
Xhold1429 _6587_/Q VGND VGND VPWR VPWR hold332/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4003_ hold579/X _5187_/A1 _4008_/S VGND VGND VPWR VPWR _6481_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5954_ _6583_/Q _5688_/X _5952_/X _5953_/X VGND VGND VPWR VPWR _5954_/X sky130_fd_sc_hd__a211o_1
XFILLER_179_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4905_ _4601_/A _4523_/Y _4491_/Y VGND VGND VPWR VPWR _4905_/X sky130_fd_sc_hd__a21o_1
XFILLER_178_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5885_ _3200_/Y _5872_/B _5677_/B VGND VGND VPWR VPWR _5885_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4836_ _4836_/A _4836_/B VGND VGND VPWR VPWR _4906_/B sky130_fd_sc_hd__nor2_1
XFILLER_138_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4767_ _4767_/A _4880_/B VGND VGND VPWR VPWR _4933_/C sky130_fd_sc_hd__and2_1
X_6506_ _7139_/CLK _6506_/D fanout478/X VGND VGND VPWR VPWR _6506_/Q sky130_fd_sc_hd__dfrtp_4
X_3718_ _6815_/Q _3391_/Y _3431_/Y input62/X _3717_/X VGND VGND VPWR VPWR _3725_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_147_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4698_ _4712_/A _4712_/B _4698_/C VGND VGND VPWR VPWR _4698_/Y sky130_fd_sc_hd__nand3_4
XFILLER_107_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6437_ _3958_/A1 _6437_/D _6392_/X VGND VGND VPWR VPWR _6437_/Q sky130_fd_sc_hd__dfrtp_4
X_3649_ _6734_/Q _4304_/A _3648_/Y _6818_/Q VGND VGND VPWR VPWR _3649_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6368_ _6684_/Q _6368_/A2 _6368_/B1 _4218_/Y _6367_/X VGND VGND VPWR VPWR _6368_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5319_ hold773/X _5571_/A1 _5325_/S VGND VGND VPWR VPWR _6902_/D sky130_fd_sc_hd__mux2_1
X_6299_ _6538_/Q _5983_/X _5993_/X _6622_/Q _6298_/X VGND VGND VPWR VPWR _6304_/B
+ sky130_fd_sc_hd__a221o_1
Xhold12 hold12/A VGND VGND VPWR VPWR hold12/X sky130_fd_sc_hd__buf_12
XFILLER_102_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold23 hold23/A VGND VGND VPWR VPWR hold23/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold34 hold34/A VGND VGND VPWR VPWR hold34/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold45 hold45/A VGND VGND VPWR VPWR hold45/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold56 hold56/A VGND VGND VPWR VPWR hold56/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold67 hold67/A VGND VGND VPWR VPWR hold67/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1930 _7015_/Q VGND VGND VPWR VPWR hold304/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1941 _7048_/Q VGND VGND VPWR VPWR hold537/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold78 hold78/A VGND VGND VPWR VPWR hold78/X sky130_fd_sc_hd__buf_12
XFILLER_28_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1952 _7135_/Q VGND VGND VPWR VPWR hold315/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1963 hold746/X VGND VGND VPWR VPWR _4264_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold89 hold89/A VGND VGND VPWR VPWR hold89/X sky130_fd_sc_hd__buf_2
Xhold1974 _4181_/X VGND VGND VPWR VPWR _6623_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1985 _6741_/Q VGND VGND VPWR VPWR hold97/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1996 _5501_/X VGND VGND VPWR VPWR _7064_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_9 _5389_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_2__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7186_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_121_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5670_ _5686_/A _5686_/B _5687_/C VGND VGND VPWR VPWR _5670_/X sky130_fd_sc_hd__and3b_4
XFILLER_176_836 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4621_ _4621_/A _5048_/A VGND VGND VPWR VPWR _5052_/A sky130_fd_sc_hd__nand2_1
XFILLER_30_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4552_ _5009_/A _4552_/B VGND VGND VPWR VPWR _5090_/C sky130_fd_sc_hd__nand2_1
XFILLER_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold504 hold504/A VGND VGND VPWR VPWR hold504/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold515 hold515/A VGND VGND VPWR VPWR hold515/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3503_ _6583_/Q _4128_/A _4334_/A _6761_/Q _3502_/X VGND VGND VPWR VPWR _3515_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold526 hold526/A VGND VGND VPWR VPWR hold526/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4483_ _4486_/A _4483_/B VGND VGND VPWR VPWR _4570_/D sky130_fd_sc_hd__nand2_8
Xhold537 hold537/A VGND VGND VPWR VPWR hold537/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold548 hold548/A VGND VGND VPWR VPWR _6536_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6222_ _6604_/Q _5982_/X _5987_/X _6727_/Q VGND VGND VPWR VPWR _6222_/X sky130_fd_sc_hd__a22o_1
Xhold559 hold559/A VGND VGND VPWR VPWR hold559/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3434_ input8/X _3315_/Y _3336_/Y input25/X VGND VGND VPWR VPWR _3434_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6153_ _6954_/Q _5997_/X _6004_/X _6882_/Q VGND VGND VPWR VPWR _6153_/X sky130_fd_sc_hd__a22o_1
X_3365_ _6980_/Q _5398_/A _3315_/Y input10/X _3362_/X VGND VGND VPWR VPWR _3368_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5104_ _4976_/B _4976_/A _5104_/C _5104_/D VGND VGND VPWR VPWR _5135_/D sky130_fd_sc_hd__and4bb_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ _7087_/Q _5638_/X _6015_/X _7015_/Q VGND VGND VPWR VPWR _6084_/X sky130_fd_sc_hd__a22o_1
Xhold1204 _6713_/Q VGND VGND VPWR VPWR hold220/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3296_ _3338_/A _3487_/A VGND VGND VPWR VPWR _5344_/A sky130_fd_sc_hd__nor2_8
Xhold1215 _6840_/Q VGND VGND VPWR VPWR hold182/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1226 _6824_/Q VGND VGND VPWR VPWR hold252/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1237 _6764_/Q VGND VGND VPWR VPWR hold37/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1248 hold117/X VGND VGND VPWR VPWR _4169_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5035_ _4683_/A _5029_/X _4961_/D _4529_/B VGND VGND VPWR VPWR _5151_/B sky130_fd_sc_hd__o211a_1
Xhold1259 _7193_/Q VGND VGND VPWR VPWR hold864/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6986_ _7125_/CLK _6986_/D fanout454/X VGND VGND VPWR VPWR _6986_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5937_ _6572_/Q _5674_/X _5680_/X _6710_/Q VGND VGND VPWR VPWR _5937_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5868_ _6752_/Q _5681_/X _5865_/X _5867_/X VGND VGND VPWR VPWR _5869_/C sky130_fd_sc_hd__a211o_1
XFILLER_178_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4819_ _4658_/A _4633_/B _4683_/A _4727_/Y _4818_/X VGND VGND VPWR VPWR _4820_/C
+ sky130_fd_sc_hd__o311a_1
XFILLER_166_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5799_ _6850_/Q _5842_/A2 _5662_/X _6898_/Q _5798_/X VGND VGND VPWR VPWR _5799_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_181_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput102 wb_adr_i[12] VGND VGND VPWR VPWR _4344_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput113 wb_adr_i[22] VGND VGND VPWR VPWR _4649_/D sky130_fd_sc_hd__buf_2
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput124 wb_adr_i[3] VGND VGND VPWR VPWR _4637_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput135 wb_dat_i[12] VGND VGND VPWR VPWR _6374_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput146 wb_dat_i[22] VGND VGND VPWR VPWR _6379_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2450 _7176_/Q VGND VGND VPWR VPWR _6141_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput157 wb_dat_i[3] VGND VGND VPWR VPWR _6371_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2461 _7178_/Q VGND VGND VPWR VPWR _6191_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput168 wb_sel_i[3] VGND VGND VPWR VPWR _6357_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2472 _7183_/Q VGND VGND VPWR VPWR _6316_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2483 _6435_/Q VGND VGND VPWR VPWR _3927_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2494 _6445_/Q VGND VGND VPWR VPWR _3870_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1760 _5355_/X VGND VGND VPWR VPWR _6934_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1771 _6746_/Q VGND VGND VPWR VPWR hold520/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_63_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1782 _6743_/Q VGND VGND VPWR VPWR hold585/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1793 hold470/X VGND VGND VPWR VPWR _3987_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_189_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6840_ _7121_/CLK _6840_/D _6399_/A VGND VGND VPWR VPWR _6840_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6771_ _6809_/CLK _6771_/D fanout444/X VGND VGND VPWR VPWR _6771_/Q sky130_fd_sc_hd__dfstp_2
X_3983_ hold202/X _4337_/A1 _3987_/S VGND VGND VPWR VPWR _6452_/D sky130_fd_sc_hd__mux2_1
X_5722_ _6902_/Q _5679_/X _5685_/X _7070_/Q _5721_/X VGND VGND VPWR VPWR _5727_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_149_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_21_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7135_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_148_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5653_ _5689_/A _5676_/B _5686_/B VGND VGND VPWR VPWR _5653_/X sky130_fd_sc_hd__and3b_4
X_4604_ _4580_/Y _4581_/X _4473_/A VGND VGND VPWR VPWR _4604_/X sky130_fd_sc_hd__o21ba_1
XFILLER_164_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5584_ hold42/X hold20/X _5586_/S VGND VGND VPWR VPWR _5584_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_36_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7140_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold301 hold301/A VGND VGND VPWR VPWR hold301/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4535_ _4463_/B _4570_/D _4533_/X _4534_/Y _4893_/A VGND VGND VPWR VPWR _4535_/X
+ sky130_fd_sc_hd__o2111a_1
Xhold312 hold312/A VGND VGND VPWR VPWR hold312/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold323 hold323/A VGND VGND VPWR VPWR hold323/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold334 hold334/A VGND VGND VPWR VPWR hold334/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold345 hold345/A VGND VGND VPWR VPWR hold345/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4466_ _4466_/A VGND VGND VPWR VPWR _4765_/B sky130_fd_sc_hd__inv_2
Xhold356 hold356/A VGND VGND VPWR VPWR hold356/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold367 hold367/A VGND VGND VPWR VPWR hold367/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold378 hold378/A VGND VGND VPWR VPWR hold378/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6205_ _7012_/Q _5993_/X _5994_/X _7068_/Q VGND VGND VPWR VPWR _6205_/X sky130_fd_sc_hd__a22o_1
XFILLER_89_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold389 hold389/A VGND VGND VPWR VPWR hold389/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3417_ input41/X _4056_/C _5308_/A _6899_/Q VGND VGND VPWR VPWR _3417_/X sky130_fd_sc_hd__a22o_1
XFILLER_132_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7185_ _7186_/CLK _7185_/D fanout465/X VGND VGND VPWR VPWR _7185_/Q sky130_fd_sc_hd__dfrtp_4
X_4397_ _4637_/A _4637_/B VGND VGND VPWR VPWR _4523_/A sky130_fd_sc_hd__and2_4
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6136_ _7049_/Q _5996_/X _6012_/X _7001_/Q _6135_/X VGND VGND VPWR VPWR _6136_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3348_ _6884_/Q _5290_/A _3347_/Y _7012_/Q VGND VGND VPWR VPWR _3348_/X sky130_fd_sc_hd__a22o_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1001 _5431_/X VGND VGND VPWR VPWR _7002_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1012 _4249_/X VGND VGND VPWR VPWR hold17/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_133_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1023 _5541_/X VGND VGND VPWR VPWR hold72/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1034 _6939_/Q VGND VGND VPWR VPWR hold348/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6067_ _6067_/A1 _6342_/S _6065_/X _6066_/X VGND VGND VPWR VPWR _6067_/X sky130_fd_sc_hd__o22a_1
XTAP_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3279_ _3277_/B hold53/A VGND VGND VPWR VPWR hold54/A sky130_fd_sc_hd__nand2b_2
Xhold1045 hold389/X VGND VGND VPWR VPWR _5459_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1056 _5558_/X VGND VGND VPWR VPWR _7115_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1067 hold429/X VGND VGND VPWR VPWR _5494_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5018_ _4664_/Y _5011_/X _4736_/Y VGND VGND VPWR VPWR _5018_/X sky130_fd_sc_hd__o21a_1
Xhold1078 hold433/X VGND VGND VPWR VPWR _5413_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1089 hold386/X VGND VGND VPWR VPWR _4248_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_54_720 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_207 _6432_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6969_ _7103_/CLK _6969_/D fanout472/X VGND VGND VPWR VPWR _6969_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_186_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_788 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold890 _3266_/X VGND VGND VPWR VPWR hold66/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_67_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2280 _5311_/X VGND VGND VPWR VPWR _6895_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2291 _7024_/Q VGND VGND VPWR VPWR hold697/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_92_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1590 _6916_/Q VGND VGND VPWR VPWR hold489/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_123_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4320_ _4320_/A0 _5303_/A1 _4321_/S VGND VGND VPWR VPWR _6745_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4251_ _4251_/A0 _5221_/A1 _4255_/S VGND VGND VPWR VPWR _4251_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3202_ _7136_/Q VGND VGND VPWR VPWR _3202_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4182_ _4182_/A _5229_/C VGND VGND VPWR VPWR _4187_/S sky130_fd_sc_hd__and2_4
XFILLER_94_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7157__486 VGND VGND VPWR VPWR _7157_/D _7157__486/LO sky130_fd_sc_hd__conb_1
XFILLER_36_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6823_ _6826_/CLK _6823_/D _6414_/A VGND VGND VPWR VPWR _6823_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_90_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6754_ _6760_/CLK _6754_/D _6433_/A VGND VGND VPWR VPWR _6754_/Q sky130_fd_sc_hd__dfstp_2
X_3966_ _6456_/Q _3966_/B VGND VGND VPWR VPWR _3966_/X sky130_fd_sc_hd__and2b_4
X_5705_ _6845_/Q _5653_/X _5702_/X _5704_/X VGND VGND VPWR VPWR _5705_/X sky130_fd_sc_hd__a211o_1
X_6685_ _7204_/CLK _6685_/D fanout484/X VGND VGND VPWR VPWR _6685_/Q sky130_fd_sc_hd__dfrtp_4
X_3897_ _4344_/C _4344_/D _4343_/A _4343_/B VGND VGND VPWR VPWR _3898_/C sky130_fd_sc_hd__nor4_1
XFILLER_31_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5636_ _5634_/B _5636_/A2 _5639_/B VGND VGND VPWR VPWR _7155_/D sky130_fd_sc_hd__a21oi_1
XFILLER_163_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5567_ _5567_/A0 _5585_/A1 _5568_/S VGND VGND VPWR VPWR _5567_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold120 hold120/A VGND VGND VPWR VPWR hold120/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold131 hold131/A VGND VGND VPWR VPWR hold131/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4518_ _4615_/B _4972_/A VGND VGND VPWR VPWR _5063_/A sky130_fd_sc_hd__nand2_1
Xhold142 hold142/A VGND VGND VPWR VPWR hold142/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5498_ hold806/X _5552_/A1 _5505_/S VGND VGND VPWR VPWR _5498_/X sky130_fd_sc_hd__mux2_1
Xhold153 hold153/A VGND VGND VPWR VPWR hold153/X sky130_fd_sc_hd__buf_12
XFILLER_132_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold164 hold164/A VGND VGND VPWR VPWR hold164/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold175 hold175/A VGND VGND VPWR VPWR hold175/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4449_ _4457_/A _4671_/A VGND VGND VPWR VPWR _4450_/B sky130_fd_sc_hd__nor2_1
Xhold186 hold186/A VGND VGND VPWR VPWR hold186/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold197 hold197/A VGND VGND VPWR VPWR wb_dat_o[26] sky130_fd_sc_hd__buf_12
XFILLER_144_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7168_ _7183_/CLK _7168_/D fanout466/X VGND VGND VPWR VPWR _7168_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6119_ _7089_/Q _5638_/X _5998_/X _6889_/Q _6118_/X VGND VGND VPWR VPWR _6119_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7099_ _7123_/CLK _7099_/D fanout477/X VGND VGND VPWR VPWR _7099_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3820_ _3846_/S VGND VGND VPWR VPWR _3835_/S sky130_fd_sc_hd__clkinv_2
XFILLER_33_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3751_ _6614_/Q _4170_/A _4176_/A _6619_/Q VGND VGND VPWR VPWR _3751_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6470_ _3958_/A1 _6470_/D _6420_/X VGND VGND VPWR VPWR _6470_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_9_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3682_ _6738_/Q _4310_/A _4274_/A _6708_/Q VGND VGND VPWR VPWR _3682_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5421_ _5421_/A0 _5556_/A1 _5424_/S VGND VGND VPWR VPWR _5421_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput203 _3935_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[35] sky130_fd_sc_hd__buf_12
XFILLER_161_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5352_ _5352_/A0 _5577_/A1 _5352_/S VGND VGND VPWR VPWR _5352_/X sky130_fd_sc_hd__mux2_1
Xoutput214 _3939_/X VGND VGND VPWR VPWR mgmt_gpio_out[10] sky130_fd_sc_hd__buf_12
Xoutput225 _7220_/X VGND VGND VPWR VPWR mgmt_gpio_out[22] sky130_fd_sc_hd__buf_12
Xoutput236 _3936_/X VGND VGND VPWR VPWR mgmt_gpio_out[32] sky130_fd_sc_hd__buf_12
XFILLER_99_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput247 _3941_/X VGND VGND VPWR VPWR mgmt_gpio_out[8] sky130_fd_sc_hd__buf_12
XFILLER_114_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput258 _6793_/Q VGND VGND VPWR VPWR pll90_sel[1] sky130_fd_sc_hd__buf_12
X_4303_ _4303_/A0 _5538_/A1 _4303_/S VGND VGND VPWR VPWR _4303_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput269 _6790_/Q VGND VGND VPWR VPWR pll_sel[1] sky130_fd_sc_hd__buf_12
X_5283_ hold754/X _5571_/A1 _5289_/S VGND VGND VPWR VPWR _5283_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7022_ _7126_/CLK _7022_/D fanout475/X VGND VGND VPWR VPWR _7022_/Q sky130_fd_sc_hd__dfstp_2
X_4234_ _4234_/A0 _4233_/X _4240_/S VGND VGND VPWR VPWR _6664_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4165_ _4165_/A0 _5221_/A1 _4169_/S VGND VGND VPWR VPWR _6609_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4096_ hold340/X _5303_/A1 _4097_/S VGND VGND VPWR VPWR _4096_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6806_ _6833_/CLK _6806_/D fanout454/X VGND VGND VPWR VPWR _6806_/Q sky130_fd_sc_hd__dfrtp_4
X_4998_ _4658_/A _4633_/B _4683_/A _4727_/Y _4885_/X VGND VGND VPWR VPWR _4999_/D
+ sky130_fd_sc_hd__o311a_1
X_6737_ _6822_/CLK _6737_/D fanout451/X VGND VGND VPWR VPWR _6737_/Q sky130_fd_sc_hd__dfrtp_4
X_3949_ _6508_/Q user_clock _6819_/Q VGND VGND VPWR VPWR _3949_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6668_ _7016_/CLK _6668_/D fanout481/X VGND VGND VPWR VPWR _7222_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_176_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5619_ _5686_/A _5639_/A VGND VGND VPWR VPWR _5619_/Y sky130_fd_sc_hd__nor2_1
XFILLER_192_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6599_ _6817_/CLK _6599_/D fanout451/X VGND VGND VPWR VPWR _6599_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_118_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout441 fanout450/X VGND VGND VPWR VPWR _3959_/B sky130_fd_sc_hd__clkbuf_16
Xfanout452 fanout453/X VGND VGND VPWR VPWR fanout452/X sky130_fd_sc_hd__buf_12
Xfanout463 fanout466/X VGND VGND VPWR VPWR _6414_/A sky130_fd_sc_hd__buf_8
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout474 fanout481/X VGND VGND VPWR VPWR fanout474/X sky130_fd_sc_hd__clkbuf_8
Xfanout485 _4637_/C VGND VGND VPWR VPWR _4575_/C sky130_fd_sc_hd__buf_12
XFILLER_74_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5970_ _5970_/A1 _6342_/S _5968_/X _5969_/X VGND VGND VPWR VPWR _7172_/D sky130_fd_sc_hd__o22a_1
XFILLER_18_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4921_ _4921_/A _4921_/B VGND VGND VPWR VPWR _4930_/C sky130_fd_sc_hd__nor2_1
XFILLER_178_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4852_ _4638_/Y _4688_/C _4625_/Y VGND VGND VPWR VPWR _5046_/A sky130_fd_sc_hd__o21a_1
XFILLER_21_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3803_ _3803_/A _3803_/B VGND VGND VPWR VPWR _3803_/Y sky130_fd_sc_hd__nand2_8
XFILLER_60_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4783_ _4384_/A _4658_/A _4417_/B _4986_/C VGND VGND VPWR VPWR _5044_/A sky130_fd_sc_hd__o31a_2
X_6522_ _6522_/CLK hold61/X fanout479/X VGND VGND VPWR VPWR _6522_/Q sky130_fd_sc_hd__dfrtp_1
X_3734_ input35/X _3315_/Y _3347_/Y _7006_/Q _3733_/X VGND VGND VPWR VPWR _3735_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6453_ _6691_/CLK _6453_/D fanout442/X VGND VGND VPWR VPWR _6453_/Q sky130_fd_sc_hd__dfrtp_4
X_3665_ _6895_/Q _5308_/A _4250_/A _6689_/Q VGND VGND VPWR VPWR _3665_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5404_ _5404_/A0 _5503_/A1 _5406_/S VGND VGND VPWR VPWR _6978_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6384_ _6383_/X hold967/X _6384_/S VGND VGND VPWR VPWR _7202_/D sky130_fd_sc_hd__mux2_1
X_3596_ _7032_/Q _5461_/A _4200_/A _6642_/Q VGND VGND VPWR VPWR _3596_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5335_ _5335_/A _5569_/B VGND VGND VPWR VPWR _5343_/S sky130_fd_sc_hd__and2_4
XFILLER_102_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5266_ hold144/X _5518_/A1 _5271_/S VGND VGND VPWR VPWR _5266_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7005_ _7077_/CLK _7005_/D fanout456/X VGND VGND VPWR VPWR _7005_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_87_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4217_ hold116/X _5538_/A1 _4217_/S VGND VGND VPWR VPWR _4217_/X sky130_fd_sc_hd__mux2_1
X_5197_ hold432/X _5503_/A1 _5199_/S VGND VGND VPWR VPWR _5197_/X sky130_fd_sc_hd__mux2_1
X_4148_ _4148_/A0 _5186_/A1 _4151_/S VGND VGND VPWR VPWR _6595_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4079_ _4079_/A0 _5186_/A1 _4082_/S VGND VGND VPWR VPWR _4079_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_1__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7194_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_79_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap416 _3738_/S VGND VGND VPWR VPWR _3857_/B sky130_fd_sc_hd__clkbuf_4
Xhold708 hold708/A VGND VGND VPWR VPWR hold708/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap427 _4672_/B VGND VGND VPWR VPWR _4698_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_7_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold719 hold719/A VGND VGND VPWR VPWR hold719/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3450_ _7058_/Q _5488_/A _3391_/Y _3428_/X VGND VGND VPWR VPWR _3450_/X sky130_fd_sc_hd__a22o_1
XFILLER_6_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3381_ _6868_/Q _5272_/A _5380_/A _6964_/Q VGND VGND VPWR VPWR _3381_/X sky130_fd_sc_hd__a22o_1
X_5120_ _4402_/Y _4523_/Y _4583_/B _4642_/Y _4839_/X VGND VGND VPWR VPWR _5121_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2109 _5273_/X VGND VGND VPWR VPWR _6861_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5051_ _4583_/B _4688_/B _4691_/Y _4638_/Y _4622_/C VGND VGND VPWR VPWR _5052_/C
+ sky130_fd_sc_hd__o221a_1
Xhold1408 _6523_/Q VGND VGND VPWR VPWR hold397/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1419 _4290_/X VGND VGND VPWR VPWR _6720_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4002_ hold737/X _5186_/A1 _4008_/S VGND VGND VPWR VPWR _6480_/D sky130_fd_sc_hd__mux2_1
XFILLER_38_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5953_ _6534_/Q _5653_/X _5662_/X _6588_/Q _5951_/X VGND VGND VPWR VPWR _5953_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_851 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4904_ _4879_/X _4892_/X _4903_/X _4561_/X VGND VGND VPWR VPWR _4906_/D sky130_fd_sc_hd__a31o_1
X_5884_ _6605_/Q _5684_/X _5686_/X _6620_/Q VGND VGND VPWR VPWR _5884_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4835_ _5114_/B _4834_/X _4716_/Y VGND VGND VPWR VPWR _4836_/B sky130_fd_sc_hd__a21oi_1
XFILLER_21_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4766_ _4735_/Y _4765_/Y _4407_/Y VGND VGND VPWR VPWR _4791_/C sky130_fd_sc_hd__a21o_1
XFILLER_147_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3717_ _6728_/Q _3509_/Y _4065_/A _6526_/Q VGND VGND VPWR VPWR _3717_/X sky130_fd_sc_hd__a22o_1
X_6505_ _6522_/CLK _6505_/D fanout478/X VGND VGND VPWR VPWR _7213_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_162_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4697_ _4712_/A _4712_/B _4751_/C VGND VGND VPWR VPWR _4702_/B sky130_fd_sc_hd__and3_1
XFILLER_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3648_ _3648_/A _3648_/B VGND VGND VPWR VPWR _3648_/Y sky130_fd_sc_hd__nor2_4
X_6436_ _6436_/CLK _6436_/D _3882_/X VGND VGND VPWR VPWR _6436_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_106_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6367_ _6686_/Q _6367_/A2 _6367_/B1 _6685_/Q VGND VGND VPWR VPWR _6367_/X sky130_fd_sc_hd__a22o_1
X_3579_ _6864_/Q _5272_/A _4122_/A _6577_/Q _3565_/X VGND VGND VPWR VPWR _3580_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_88_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5318_ hold785/X _5570_/A1 _5325_/S VGND VGND VPWR VPWR _6901_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6298_ _6572_/Q _5988_/X _6014_/X _6745_/Q VGND VGND VPWR VPWR _6298_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold13 hold13/A VGND VGND VPWR VPWR hold13/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold24 hold24/A VGND VGND VPWR VPWR hold24/X sky130_fd_sc_hd__buf_2
X_5249_ _5249_/A0 _5249_/A1 _5253_/S VGND VGND VPWR VPWR _6840_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold35 hold35/A VGND VGND VPWR VPWR hold35/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold46 hold46/A VGND VGND VPWR VPWR hold46/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1920 _6604_/Q VGND VGND VPWR VPWR hold656/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold57 hold57/A VGND VGND VPWR VPWR hold57/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1931 hold304/X VGND VGND VPWR VPWR _5446_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1942 hold537/X VGND VGND VPWR VPWR _5483_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold68 hold68/A VGND VGND VPWR VPWR hold68/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold79 hold79/A VGND VGND VPWR VPWR hold79/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1953 hold315/X VGND VGND VPWR VPWR _5581_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1964 _7077_/Q VGND VGND VPWR VPWR hold637/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1975 _6627_/Q VGND VGND VPWR VPWR hold658/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1986 _7211_/A VGND VGND VPWR VPWR hold660/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_16_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1997 _6943_/Q VGND VGND VPWR VPWR hold333/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4620_ _4625_/A _4621_/A VGND VGND VPWR VPWR _4622_/C sky130_fd_sc_hd__nand2_2
XFILLER_129_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4551_ _4601_/A _4491_/Y _4548_/X _5138_/A _4550_/Y VGND VGND VPWR VPWR _4553_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_190_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3502_ _7001_/Q _5425_/A _5461_/A _7033_/Q VGND VGND VPWR VPWR _3502_/X sky130_fd_sc_hd__a22o_1
XFILLER_156_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold505 hold505/A VGND VGND VPWR VPWR hold505/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold516 hold516/A VGND VGND VPWR VPWR hold516/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4482_ _4486_/A _4485_/B _4564_/B VGND VGND VPWR VPWR _4615_/B sky130_fd_sc_hd__and3_1
XFILLER_143_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold527 hold527/A VGND VGND VPWR VPWR hold527/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold538 hold538/A VGND VGND VPWR VPWR hold538/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6221_ _6548_/Q _5999_/X _6019_/X _6732_/Q _6220_/X VGND VGND VPWR VPWR _6238_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_104_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold549 hold549/A VGND VGND VPWR VPWR hold549/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3433_ _7042_/Q _5470_/A _5533_/A _7098_/Q VGND VGND VPWR VPWR _3433_/X sky130_fd_sc_hd__a22o_4
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ _6152_/A _6152_/B _6152_/C VGND VGND VPWR VPWR _6164_/C sky130_fd_sc_hd__nor3_1
XFILLER_131_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _6996_/Q _5416_/A _5470_/A _7044_/Q _3361_/X VGND VGND VPWR VPWR _3368_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_98_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _5103_/A _5103_/B _5103_/C VGND VGND VPWR VPWR _5104_/D sky130_fd_sc_hd__and3_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _6895_/Q _5989_/X _6013_/X _7079_/Q _6082_/X VGND VGND VPWR VPWR _6088_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ _3563_/A hold32/X VGND VGND VPWR VPWR hold33/A sky130_fd_sc_hd__nor2_8
Xhold1205 hold220/X VGND VGND VPWR VPWR _4282_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1216 hold182/X VGND VGND VPWR VPWR _5249_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1227 hold252/X VGND VGND VPWR VPWR _5231_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5034_ _5034_/A _5034_/B _5034_/C _5034_/D VGND VGND VPWR VPWR _5117_/C sky130_fd_sc_hd__and4_1
Xhold1238 hold37/X VGND VGND VPWR VPWR _3263_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1249 _4169_/X VGND VGND VPWR VPWR _6613_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_26_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6985_ _7121_/CLK _6985_/D _6399_/A VGND VGND VPWR VPWR _6985_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5936_ _6695_/Q _5658_/X _5664_/X _6760_/Q VGND VGND VPWR VPWR _5936_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5867_ _6697_/Q _5672_/X _5680_/X _6707_/Q _5866_/X VGND VGND VPWR VPWR _5867_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_139_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4818_ _4818_/A _4818_/B _5080_/A VGND VGND VPWR VPWR _4818_/X sky130_fd_sc_hd__and3_1
XFILLER_182_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5798_ _6882_/Q _5667_/X _5682_/X _7042_/Q VGND VGND VPWR VPWR _5798_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4749_ _4804_/A _4686_/X _4748_/X VGND VGND VPWR VPWR _4749_/X sky130_fd_sc_hd__a21o_1
XFILLER_181_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6419_ _6426_/A _6432_/B VGND VGND VPWR VPWR _6419_/X sky130_fd_sc_hd__and2_1
XFILLER_1_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput103 wb_adr_i[13] VGND VGND VPWR VPWR _4344_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput114 wb_adr_i[23] VGND VGND VPWR VPWR _4649_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput125 wb_adr_i[4] VGND VGND VPWR VPWR _4701_/A sky130_fd_sc_hd__buf_12
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput136 wb_dat_i[13] VGND VGND VPWR VPWR _6377_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2440 _6092_/X VGND VGND VPWR VPWR _7175_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2451 _7168_/Q VGND VGND VPWR VPWR _5903_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput147 wb_dat_i[23] VGND VGND VPWR VPWR _6383_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput158 wb_dat_i[4] VGND VGND VPWR VPWR _6373_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2462 _6167_/X VGND VGND VPWR VPWR _7178_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput169 wb_stb_i VGND VGND VPWR VPWR _3893_/D sky130_fd_sc_hd__buf_4
Xhold2473 _6458_/Q VGND VGND VPWR VPWR _3851_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2484 _3927_/Y VGND VGND VPWR VPWR _6657_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1750 _6696_/Q VGND VGND VPWR VPWR hold514/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2495 _3869_/Y VGND VGND VPWR VPWR _6446_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1761 _6638_/Q VGND VGND VPWR VPWR hold522/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1772 hold520/X VGND VGND VPWR VPWR _4321_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1783 hold585/X VGND VGND VPWR VPWR _4318_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1794 _6769_/Q VGND VGND VPWR VPWR hold605/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_2_csclk _6727_/CLK VGND VGND VPWR VPWR _6757_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6770_ _6794_/CLK _6770_/D fanout445/X VGND VGND VPWR VPWR _6770_/Q sky130_fd_sc_hd__dfrtp_4
X_3982_ _3982_/A0 hold73/X _3996_/S VGND VGND VPWR VPWR _3982_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5721_ _6910_/Q _5670_/X _5678_/B _6966_/Q _5707_/B VGND VGND VPWR VPWR _5721_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_176_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5652_ _7147_/Q _7146_/Q VGND VGND VPWR VPWR _5686_/B sky130_fd_sc_hd__and2b_4
XFILLER_148_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4603_ _4981_/A _4917_/D VGND VGND VPWR VPWR _4616_/B sky130_fd_sc_hd__nand2_1
XFILLER_191_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5583_ _5583_/A0 _5583_/A1 _5586_/S VGND VGND VPWR VPWR _7137_/D sky130_fd_sc_hd__mux2_1
XFILLER_190_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4534_ _4562_/A _4972_/A VGND VGND VPWR VPWR _4534_/Y sky130_fd_sc_hd__nand2_2
XFILLER_156_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold302 hold302/A VGND VGND VPWR VPWR hold302/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold313 hold313/A VGND VGND VPWR VPWR hold313/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold324 hold324/A VGND VGND VPWR VPWR hold324/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold335 hold335/A VGND VGND VPWR VPWR hold335/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4465_ _4363_/B _4465_/B VGND VGND VPWR VPWR _4466_/A sky130_fd_sc_hd__nand2b_4
Xhold346 hold346/A VGND VGND VPWR VPWR hold346/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold357 hold357/A VGND VGND VPWR VPWR _6859_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold368 hold368/A VGND VGND VPWR VPWR hold368/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6204_ _6204_/A _6204_/B _6204_/C _6204_/D VGND VGND VPWR VPWR _6204_/Y sky130_fd_sc_hd__nor4_1
X_3416_ _7027_/Q _5452_/A hold40/A _6851_/Q _3415_/X VGND VGND VPWR VPWR _3421_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold379 hold379/A VGND VGND VPWR VPWR hold379/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7184_ _7186_/CLK _7184_/D _6409_/A VGND VGND VPWR VPWR _7184_/Q sky130_fd_sc_hd__dfrtp_1
X_4396_ _4513_/A _5009_/A _4584_/A _4652_/A VGND VGND VPWR VPWR _4396_/X sky130_fd_sc_hd__and4_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6135_ _7065_/Q _5994_/X _6018_/X _6969_/Q VGND VGND VPWR VPWR _6135_/X sky130_fd_sc_hd__a22o_1
X_3347_ _3501_/A hold32/X VGND VGND VPWR VPWR _3347_/Y sky130_fd_sc_hd__nor2_8
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_824 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1002 _6844_/Q VGND VGND VPWR VPWR _5253_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1013 _7092_/Q VGND VGND VPWR VPWR hold35/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6066_ _6490_/Q _7173_/Q _5649_/Y VGND VGND VPWR VPWR _6066_/X sky130_fd_sc_hd__a21o_1
Xhold1024 _7003_/Q VGND VGND VPWR VPWR hold366/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_3278_ hold52/X _3302_/A VGND VGND VPWR VPWR hold53/A sky130_fd_sc_hd__nor2_4
Xhold1035 hold348/X VGND VGND VPWR VPWR _5360_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1046 _5459_/X VGND VGND VPWR VPWR _7027_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1057 _6467_/Q VGND VGND VPWR VPWR _3253_/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5017_ _4691_/Y _4995_/B _5016_/X _4818_/B VGND VGND VPWR VPWR _5080_/B sky130_fd_sc_hd__o211a_1
XFILLER_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1068 _5494_/X VGND VGND VPWR VPWR _7058_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1079 _6970_/Q VGND VGND VPWR VPWR hold435/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_732 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_208 hold153/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6968_ _7139_/CLK _6968_/D fanout478/X VGND VGND VPWR VPWR _6968_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5919_ _6532_/Q _5653_/X _5918_/X VGND VGND VPWR VPWR _5919_/X sky130_fd_sc_hd__a21o_1
X_6899_ _7139_/CLK _6899_/D fanout471/X VGND VGND VPWR VPWR _6899_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_10_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold880 _7204_/Q VGND VGND VPWR VPWR hold11/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold891 _3297_/Y VGND VGND VPWR VPWR hold39/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2270 _6598_/Q VGND VGND VPWR VPWR hold523/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2281 _6926_/Q VGND VGND VPWR VPWR hold751/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2292 hold697/X VGND VGND VPWR VPWR _5456_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1580 _5277_/X VGND VGND VPWR VPWR _6865_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1591 hold489/X VGND VGND VPWR VPWR _5334_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4250_ _4250_/A _5229_/C VGND VGND VPWR VPWR _4255_/S sky130_fd_sc_hd__and2_4
XFILLER_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3201_ _6719_/Q VGND VGND VPWR VPWR _3201_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4181_ _4181_/A0 _4339_/A1 _4181_/S VGND VGND VPWR VPWR _4181_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6822_ _6822_/CLK _6822_/D fanout451/X VGND VGND VPWR VPWR _6822_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6753_ _6761_/CLK _6753_/D _6426_/A VGND VGND VPWR VPWR _6753_/Q sky130_fd_sc_hd__dfrtp_4
X_3965_ _6457_/Q _3965_/B VGND VGND VPWR VPWR _3965_/X sky130_fd_sc_hd__and2b_4
XFILLER_10_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5704_ _6957_/Q _5680_/X _5686_/X _7005_/Q _5703_/X VGND VGND VPWR VPWR _5704_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3896_ _4343_/C _4343_/D _3896_/C VGND VGND VPWR VPWR _3898_/B sky130_fd_sc_hd__nor3_1
X_6684_ _7204_/CLK _6684_/D fanout484/X VGND VGND VPWR VPWR _6684_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_137_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5635_ _7155_/Q _5639_/A VGND VGND VPWR VPWR _5635_/Y sky130_fd_sc_hd__nor2_1
XFILLER_163_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5566_ hold930/X hold20/X _5568_/S VGND VGND VPWR VPWR _5566_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold110 hold110/A VGND VGND VPWR VPWR hold110/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold121 _4050_/X VGND VGND VPWR VPWR _6511_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_191_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4517_ _4812_/A _4948_/A VGND VGND VPWR VPWR _4959_/A sky130_fd_sc_hd__and2_1
Xhold132 hold132/A VGND VGND VPWR VPWR hold132/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5497_ _5497_/A _5551_/B VGND VGND VPWR VPWR _5505_/S sky130_fd_sc_hd__and2_4
Xhold143 hold143/A VGND VGND VPWR VPWR hold143/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold154 hold154/A VGND VGND VPWR VPWR hold154/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold165 hold165/A VGND VGND VPWR VPWR hold165/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold176 hold176/A VGND VGND VPWR VPWR hold176/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4448_ _4714_/B VGND VGND VPWR VPWR _4671_/A sky130_fd_sc_hd__inv_2
Xhold187 hold187/A VGND VGND VPWR VPWR hold187/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold198 hold198/A VGND VGND VPWR VPWR hold857/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4379_ _5001_/A _4717_/A _4717_/B VGND VGND VPWR VPWR _4811_/B sky130_fd_sc_hd__and3_4
X_7167_ _3950_/A1 _7167_/D _6409_/A VGND VGND VPWR VPWR _7167_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6118_ _6849_/Q _6007_/X _6019_/X _6985_/Q VGND VGND VPWR VPWR _6118_/X sky130_fd_sc_hd__a22o_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7098_ _7133_/CLK hold83/X fanout471/X VGND VGND VPWR VPWR _7098_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6049_ _6958_/Q _5992_/X _6019_/X _6982_/Q _6048_/X VGND VGND VPWR VPWR _6054_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_754 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_20_csclk _6850_/CLK VGND VGND VPWR VPWR _7008_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_49_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_35_csclk _6850_/CLK VGND VGND VPWR VPWR _7091_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3750_ _3750_/A _3750_/B _3750_/C _3750_/D VGND VGND VPWR VPWR _3770_/A sky130_fd_sc_hd__nor4_1
XFILLER_118_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3681_ _6926_/Q _5344_/A _5290_/A _6878_/Q _3680_/X VGND VGND VPWR VPWR _3684_/B
+ sky130_fd_sc_hd__a221o_1
X_5420_ _5420_/A0 _5582_/A1 _5424_/S VGND VGND VPWR VPWR _5420_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput204 _3934_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[36] sky130_fd_sc_hd__buf_12
X_5351_ _5351_/A0 _5576_/A1 _5352_/S VGND VGND VPWR VPWR _5351_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput215 _7212_/X VGND VGND VPWR VPWR mgmt_gpio_out[11] sky130_fd_sc_hd__buf_12
Xoutput226 _7221_/X VGND VGND VPWR VPWR mgmt_gpio_out[23] sky130_fd_sc_hd__buf_12
Xoutput237 _3937_/X VGND VGND VPWR VPWR mgmt_gpio_out[33] sky130_fd_sc_hd__buf_12
Xoutput248 _3959_/Y VGND VGND VPWR VPWR pad_flash_clk_oeb sky130_fd_sc_hd__buf_12
X_4302_ _4302_/A0 _5249_/A1 _4303_/S VGND VGND VPWR VPWR _4302_/X sky130_fd_sc_hd__mux2_1
Xoutput259 _6794_/Q VGND VGND VPWR VPWR pll90_sel[2] sky130_fd_sc_hd__buf_12
X_5282_ hold645/X _5561_/A1 _5289_/S VGND VGND VPWR VPWR _5282_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4233_ _5241_/A0 hold95/X _4239_/S VGND VGND VPWR VPWR _4233_/X sky130_fd_sc_hd__mux2_1
X_7021_ _7125_/CLK _7021_/D fanout454/X VGND VGND VPWR VPWR _7021_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_87_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4164_ _4164_/A hold13/A VGND VGND VPWR VPWR _4169_/S sky130_fd_sc_hd__and2_4
XFILLER_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4095_ _4095_/A0 _4337_/A1 _4097_/S VGND VGND VPWR VPWR _6550_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6805_ _6833_/CLK _6805_/D fanout454/X VGND VGND VPWR VPWR _6805_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_169_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4997_ _4997_/A _5104_/C VGND VGND VPWR VPWR _5139_/B sky130_fd_sc_hd__and2_1
XFILLER_168_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6736_ _6742_/CLK _6736_/D fanout439/X VGND VGND VPWR VPWR _6736_/Q sky130_fd_sc_hd__dfrtp_4
X_3948_ _3239_/Y input2/X input1/X VGND VGND VPWR VPWR _3948_/X sky130_fd_sc_hd__mux2_8
XFILLER_183_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6667_ _7084_/CLK _6667_/D fanout455/X VGND VGND VPWR VPWR _7211_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_136_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3879_ _3879_/A wire1/X VGND VGND VPWR VPWR _3879_/X sky130_fd_sc_hd__and2_1
XFILLER_192_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5618_ _5620_/S _5617_/X _5611_/Y VGND VGND VPWR VPWR _7149_/D sky130_fd_sc_hd__o21a_1
XFILLER_118_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6598_ _6788_/CLK _6598_/D _3959_/B VGND VGND VPWR VPWR _6598_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5549_ hold84/X hold78/X _5550_/S VGND VGND VPWR VPWR hold85/A sky130_fd_sc_hd__mux2_1
XFILLER_3_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_0__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _6568_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_160_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7219_ _7219_/A VGND VGND VPWR VPWR _7219_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_120_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout420 _7150_/Q VGND VGND VPWR VPWR _5872_/B sky130_fd_sc_hd__buf_12
Xfanout442 fanout445/X VGND VGND VPWR VPWR fanout442/X sky130_fd_sc_hd__buf_12
Xfanout453 fanout457/X VGND VGND VPWR VPWR fanout453/X sky130_fd_sc_hd__buf_8
Xfanout464 fanout466/X VGND VGND VPWR VPWR _6409_/A sky130_fd_sc_hd__buf_12
XFILLER_47_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout475 fanout476/X VGND VGND VPWR VPWR fanout475/X sky130_fd_sc_hd__buf_12
XFILLER_101_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4920_ _5114_/A _4920_/B _5114_/B VGND VGND VPWR VPWR _4929_/B sky130_fd_sc_hd__and3_1
XFILLER_61_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4851_ _4917_/D _5048_/B VGND VGND VPWR VPWR _4913_/A sky130_fd_sc_hd__nand2_1
X_3802_ _3774_/X _3802_/B _3802_/C _3802_/D VGND VGND VPWR VPWR _3803_/B sky130_fd_sc_hd__and4b_4
X_4782_ _4552_/B _4955_/D _4396_/X VGND VGND VPWR VPWR _4782_/X sky130_fd_sc_hd__a21o_1
XFILLER_20_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6521_ _6523_/CLK _6521_/D fanout479/X VGND VGND VPWR VPWR _6521_/Q sky130_fd_sc_hd__dfrtp_1
X_3733_ _6480_/Q _3357_/Y _4134_/A _6585_/Q VGND VGND VPWR VPWR _3733_/X sky130_fd_sc_hd__a22o_1
XFILLER_186_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6452_ _6809_/CLK _6452_/D fanout444/X VGND VGND VPWR VPWR _6452_/Q sky130_fd_sc_hd__dfstp_2
X_3664_ _3664_/A _3664_/B _3664_/C VGND VGND VPWR VPWR _3674_/C sky130_fd_sc_hd__nor3_1
XFILLER_109_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5403_ _5403_/A0 _5556_/A1 _5406_/S VGND VGND VPWR VPWR _6977_/D sky130_fd_sc_hd__mux2_1
X_6383_ _6684_/Q _6383_/A2 _6383_/B1 _4218_/Y _6382_/X VGND VGND VPWR VPWR _6383_/X
+ sky130_fd_sc_hd__a221o_1
X_3595_ _3595_/A _3595_/B _3595_/C _3595_/D VGND VGND VPWR VPWR _3615_/A sky130_fd_sc_hd__nor4_1
X_5334_ _5334_/A0 _5559_/A1 _5334_/S VGND VGND VPWR VPWR _5334_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5265_ hold499/X _5499_/A1 _5271_/S VGND VGND VPWR VPWR _5265_/X sky130_fd_sc_hd__mux2_1
X_7004_ _7084_/CLK _7004_/D fanout456/X VGND VGND VPWR VPWR _7004_/Q sky130_fd_sc_hd__dfrtp_4
X_4216_ hold146/X _5249_/A1 _4217_/S VGND VGND VPWR VPWR _4216_/X sky130_fd_sc_hd__mux2_1
X_5196_ hold443/X _5196_/A1 _5199_/S VGND VGND VPWR VPWR _6799_/D sky130_fd_sc_hd__mux2_1
X_4147_ _4147_/A0 _5208_/A1 _4151_/S VGND VGND VPWR VPWR _6594_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4078_ hold427/X _5208_/A1 _4082_/S VGND VGND VPWR VPWR _4078_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6719_ _6788_/CLK _6719_/D _3959_/B VGND VGND VPWR VPWR _6719_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_137_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold709 hold709/A VGND VGND VPWR VPWR hold709/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap428 _4684_/A VGND VGND VPWR VPWR _4726_/C sky130_fd_sc_hd__buf_2
XFILLER_109_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3380_ _6956_/Q _5371_/A _3330_/Y input51/X _3379_/X VGND VGND VPWR VPWR _3383_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_171_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5050_ _4510_/A _4523_/Y _4583_/B _4995_/A _4859_/X VGND VGND VPWR VPWR _5112_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_85_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1409 hold397/X VGND VGND VPWR VPWR _4063_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4001_ hold796/X _5208_/A1 _4008_/S VGND VGND VPWR VPWR _6479_/D sky130_fd_sc_hd__mux2_1
XFILLER_78_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5952_ _6578_/Q _5667_/X _5682_/X _6454_/Q VGND VGND VPWR VPWR _5952_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4903_ _5155_/A _4903_/B _4903_/C _4903_/D VGND VGND VPWR VPWR _4903_/X sky130_fd_sc_hd__and4_1
X_5883_ _6688_/Q _5659_/X _5687_/X _6600_/Q VGND VGND VPWR VPWR _5883_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4834_ _4834_/A _4834_/B _4834_/C VGND VGND VPWR VPWR _4834_/X sky130_fd_sc_hd__and3_1
XFILLER_166_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4765_ _4955_/C _4765_/B _4972_/A VGND VGND VPWR VPWR _4765_/Y sky130_fd_sc_hd__nand3_2
XFILLER_193_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6504_ _6522_/CLK _6504_/D fanout478/X VGND VGND VPWR VPWR _7212_/A sky130_fd_sc_hd__dfrtp_1
X_3716_ _3716_/A _3716_/B _3716_/C _3716_/D VGND VGND VPWR VPWR _3736_/B sky130_fd_sc_hd__nor4_1
XFILLER_146_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4696_ _4990_/B _4691_/Y _4692_/X _4694_/Y _4922_/B VGND VGND VPWR VPWR _4703_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_174_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6435_ _6658_/CLK _6435_/D _6391_/X VGND VGND VPWR VPWR _6435_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_134_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3647_ input5/X _3315_/Y _4310_/A _6739_/Q _3646_/X VGND VGND VPWR VPWR _3655_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_161_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6366_ _6365_/X _6366_/A1 _6384_/S VGND VGND VPWR VPWR _7196_/D sky130_fd_sc_hd__mux2_1
X_3578_ _6872_/Q _5281_/A _5389_/A _6968_/Q _3577_/X VGND VGND VPWR VPWR _3580_/C
+ sky130_fd_sc_hd__a221o_4
XFILLER_115_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5317_ _5317_/A _5569_/B VGND VGND VPWR VPWR _5325_/S sky130_fd_sc_hd__and2_4
XFILLER_142_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6297_ _6612_/Q _5976_/B _5995_/X _6602_/Q _6296_/X VGND VGND VPWR VPWR _6304_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold14 hold14/A VGND VGND VPWR VPWR hold14/X sky130_fd_sc_hd__buf_4
X_5248_ _5248_/A0 _5581_/A1 _5253_/S VGND VGND VPWR VPWR _6839_/D sky130_fd_sc_hd__mux2_1
Xhold25 hold25/A VGND VGND VPWR VPWR hold25/X sky130_fd_sc_hd__buf_4
Xhold36 hold36/A VGND VGND VPWR VPWR hold36/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1910 _6993_/Q VGND VGND VPWR VPWR hold422/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold47 hold47/A VGND VGND VPWR VPWR hold47/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1921 hold656/X VGND VGND VPWR VPWR _4159_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold58 hold58/A VGND VGND VPWR VPWR hold58/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold69 hold69/A VGND VGND VPWR VPWR hold69/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1932 _7008_/Q VGND VGND VPWR VPWR hold532/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5179_ _5179_/A0 _5208_/A1 _5183_/S VGND VGND VPWR VPWR _6784_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1943 _6571_/Q VGND VGND VPWR VPWR hold294/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1954 _6729_/Q VGND VGND VPWR VPWR hold313/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1965 _6889_/Q VGND VGND VPWR VPWR hold436/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1976 hold658/X VGND VGND VPWR VPWR _4186_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1987 hold660/X VGND VGND VPWR VPWR _4240_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1998 hold333/X VGND VGND VPWR VPWR _5365_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4550_ _4972_/A _4628_/A VGND VGND VPWR VPWR _4550_/Y sky130_fd_sc_hd__nand2_2
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3501_ _3501_/A _3523_/B VGND VGND VPWR VPWR _4334_/A sky130_fd_sc_hd__nor2_8
Xhold506 hold506/A VGND VGND VPWR VPWR hold506/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4481_ _4724_/C _4562_/A VGND VGND VPWR VPWR _4893_/A sky130_fd_sc_hd__nand2_2
Xhold517 hold517/A VGND VGND VPWR VPWR _6539_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold528 hold528/A VGND VGND VPWR VPWR hold528/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6220_ _6752_/Q _5638_/X _6015_/X _6757_/Q VGND VGND VPWR VPWR _6220_/X sky130_fd_sc_hd__a22o_1
Xhold539 hold539/A VGND VGND VPWR VPWR hold539/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3432_ _7138_/Q hold33/A _4241_/A input57/X VGND VGND VPWR VPWR _3432_/X sky130_fd_sc_hd__a22o_1
XFILLER_98_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3363_ _7052_/Q _5479_/A _5407_/A _6988_/Q _3359_/X VGND VGND VPWR VPWR _3368_/A
+ sky130_fd_sc_hd__a221o_1
X_6151_ _7034_/Q _5986_/X _5998_/X _6890_/Q _6150_/X VGND VGND VPWR VPWR _6152_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_124_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _5102_/A _5102_/B _5102_/C VGND VGND VPWR VPWR _5103_/C sky130_fd_sc_hd__and3_1
X_3294_ hold31/X _3430_/A VGND VGND VPWR VPWR hold32/A sky130_fd_sc_hd__nand2_2
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _6935_/Q _5980_/X _6017_/X _7071_/Q VGND VGND VPWR VPWR _6082_/X sky130_fd_sc_hd__a22o_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1206 _4282_/X VGND VGND VPWR VPWR _6713_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1217 _6572_/Q VGND VGND VPWR VPWR hold176/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1228 _5231_/X VGND VGND VPWR VPWR _6824_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5033_ _5033_/A _5033_/B VGND VGND VPWR VPWR _5089_/C sky130_fd_sc_hd__nand2_1
Xhold1239 _3263_/X VGND VGND VPWR VPWR hold38/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6984_ _7138_/CLK _6984_/D fanout480/X VGND VGND VPWR VPWR _6984_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_25_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5935_ _6637_/Q _5671_/X _5931_/X _5933_/X _5934_/X VGND VGND VPWR VPWR _5935_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_178_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5866_ _6609_/Q _5660_/X _5669_/X _6649_/Q VGND VGND VPWR VPWR _5866_/X sky130_fd_sc_hd__a22o_1
X_4817_ _4917_/A _4672_/Y _4812_/Y _4815_/X _5010_/A VGND VGND VPWR VPWR _4820_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_178_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5797_ _3242_/Y _5872_/B _5677_/B VGND VGND VPWR VPWR _5797_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4748_ _4637_/C _4719_/A _4686_/X _4747_/Y VGND VGND VPWR VPWR _4748_/X sky130_fd_sc_hd__a31o_1
XFILLER_107_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4679_ _5009_/B _4826_/A VGND VGND VPWR VPWR _4679_/Y sky130_fd_sc_hd__nor2_2
XFILLER_107_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6418_ _6426_/A _6432_/B VGND VGND VPWR VPWR _6418_/X sky130_fd_sc_hd__and2_1
XFILLER_162_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6349_ _3675_/Y hold852/A _6354_/S VGND VGND VPWR VPWR _7189_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput104 wb_adr_i[14] VGND VGND VPWR VPWR _4344_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput115 wb_adr_i[24] VGND VGND VPWR VPWR _3896_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput126 wb_adr_i[5] VGND VGND VPWR VPWR _4917_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_76_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2430 _7163_/Q VGND VGND VPWR VPWR _5794_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput137 wb_dat_i[14] VGND VGND VPWR VPWR _6379_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2441 _6655_/Q VGND VGND VPWR VPWR _3920_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput148 wb_dat_i[24] VGND VGND VPWR VPWR _6361_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2452 _5882_/X VGND VGND VPWR VPWR _7168_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput159 wb_dat_i[5] VGND VGND VPWR VPWR _6376_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2463 hold76/A VGND VGND VPWR VPWR _3873_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2474 _3851_/X VGND VGND VPWR VPWR _6458_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1740 _6806_/Q VGND VGND VPWR VPWR hold234/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2485 _6658_/Q VGND VGND VPWR VPWR _3926_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1751 hold514/X VGND VGND VPWR VPWR _4261_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2496 _7167_/Q VGND VGND VPWR VPWR _5860_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1762 hold522/X VGND VGND VPWR VPWR _4199_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1773 _6829_/Q VGND VGND VPWR VPWR hold651/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1784 _7207_/A VGND VGND VPWR VPWR hold426/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1795 hold605/X VGND VGND VPWR VPWR _5170_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_189_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3981_ _3981_/A0 _5193_/A1 _3987_/S VGND VGND VPWR VPWR _6451_/D sky130_fd_sc_hd__mux2_1
XFILLER_63_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5720_ _6974_/Q _5660_/X _5686_/X _7006_/Q _5719_/X VGND VGND VPWR VPWR _5727_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_94_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5651_ _5689_/A _5676_/B _5689_/B VGND VGND VPWR VPWR _5651_/X sky130_fd_sc_hd__and3b_4
XFILLER_149_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4602_ _4581_/X _4602_/B VGND VGND VPWR VPWR _4602_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_175_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5582_ _5582_/A0 _5582_/A1 _5586_/S VGND VGND VPWR VPWR _7136_/D sky130_fd_sc_hd__mux2_1
XFILLER_175_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4533_ _5034_/A _4533_/B _4533_/C _4533_/D VGND VGND VPWR VPWR _4533_/X sky130_fd_sc_hd__and4_1
XFILLER_117_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold303 _4066_/X VGND VGND VPWR VPWR _6525_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold314 hold314/A VGND VGND VPWR VPWR hold314/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold325 hold325/A VGND VGND VPWR VPWR hold325/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold336 _5246_/X VGND VGND VPWR VPWR _6837_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4464_ _4576_/A _4488_/B VGND VGND VPWR VPWR _4464_/Y sky130_fd_sc_hd__nand2_4
Xhold347 hold988/X VGND VGND VPWR VPWR hold989/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold358 hold358/A VGND VGND VPWR VPWR hold358/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6203_ _7036_/Q _5986_/X _5988_/X _6876_/Q _6202_/X VGND VGND VPWR VPWR _6204_/D
+ sky130_fd_sc_hd__a221o_1
Xhold369 hold369/A VGND VGND VPWR VPWR hold369/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3415_ _7043_/Q _5470_/A _5407_/A _6987_/Q VGND VGND VPWR VPWR _3415_/X sky130_fd_sc_hd__a22o_1
X_7183_ _7183_/CLK _7183_/D _6409_/A VGND VGND VPWR VPWR _7183_/Q sky130_fd_sc_hd__dfrtp_1
X_4395_ _4395_/A _4650_/B VGND VGND VPWR VPWR _4652_/A sky130_fd_sc_hd__nor2_4
XFILLER_98_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6134_ _7097_/Q _5984_/X _6013_/X _7081_/Q VGND VGND VPWR VPWR _6134_/X sky130_fd_sc_hd__a22o_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3346_ hold54/X hold32/X VGND VGND VPWR VPWR _5290_/A sky130_fd_sc_hd__nor2_8
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1003 _5253_/X VGND VGND VPWR VPWR hold28/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1014 _5532_/X VGND VGND VPWR VPWR hold36/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6065_ _6838_/Q _6339_/B _6064_/Y _6341_/S VGND VGND VPWR VPWR _6065_/X sky130_fd_sc_hd__o211a_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3277_ _3302_/A _3277_/B VGND VGND VPWR VPWR _3290_/B sky130_fd_sc_hd__nor2_2
Xhold1025 hold366/X VGND VGND VPWR VPWR _5432_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_100_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1036 _5360_/X VGND VGND VPWR VPWR _6939_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1047 _6907_/Q VGND VGND VPWR VPWR hold346/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1058 _3253_/Y VGND VGND VPWR VPWR hold1058/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5016_ _5011_/A _4590_/Y _4688_/B VGND VGND VPWR VPWR _5016_/X sky130_fd_sc_hd__a21o_1
Xhold1069 _7099_/Q VGND VGND VPWR VPWR hold404/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_39_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6967_ _7077_/CLK _6967_/D fanout456/X VGND VGND VPWR VPWR _6967_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5918_ _6576_/Q _5667_/X _5682_/X _6452_/Q VGND VGND VPWR VPWR _5918_/X sky130_fd_sc_hd__a22o_1
X_6898_ _7124_/CLK _6898_/D fanout459/X VGND VGND VPWR VPWR _6898_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5849_ _7028_/Q _5663_/X _5843_/X _5844_/X _5848_/X VGND VGND VPWR VPWR _5849_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_10_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold870 hold870/A VGND VGND VPWR VPWR hold870/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold881 hold11/X VGND VGND VPWR VPWR hold881/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold892 hold39/X VGND VGND VPWR VPWR _3425_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_1_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2260 _7096_/Q VGND VGND VPWR VPWR hold695/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2271 hold523/X VGND VGND VPWR VPWR _4151_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2282 hold751/X VGND VGND VPWR VPWR _5346_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2293 _5456_/X VGND VGND VPWR VPWR _7024_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1570 hold710/X VGND VGND VPWR VPWR _4172_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1581 _6556_/Q VGND VGND VPWR VPWR hold826/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1592 _5334_/X VGND VGND VPWR VPWR _6916_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_83_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3200_ _6718_/Q VGND VGND VPWR VPWR _3200_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4180_ _4180_/A0 _5195_/A1 _4181_/S VGND VGND VPWR VPWR _4180_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6821_ _6822_/CLK _6821_/D fanout451/X VGND VGND VPWR VPWR _6821_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_63_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6752_ _6759_/CLK _6752_/D _6426_/A VGND VGND VPWR VPWR _6752_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_16_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3964_ input85/X wire1/X _6457_/Q VGND VGND VPWR VPWR _3964_/X sky130_fd_sc_hd__mux2_4
XFILLER_149_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5703_ _6861_/Q _5673_/X _5687_/X _6917_/Q VGND VGND VPWR VPWR _5703_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6683_ _7203_/CLK _6683_/D _6346_/B VGND VGND VPWR VPWR _6683_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_149_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3895_ _4345_/C _4345_/D _4344_/A _4344_/B VGND VGND VPWR VPWR _3899_/C sky130_fd_sc_hd__nor4_1
XFILLER_149_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5634_ _5637_/A _5634_/B VGND VGND VPWR VPWR _5639_/B sky130_fd_sc_hd__nor2_1
XFILLER_191_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5565_ _5565_/A0 _5583_/A1 _5568_/S VGND VGND VPWR VPWR _7121_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold100 _5268_/X VGND VGND VPWR VPWR _6857_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold111 _3259_/B VGND VGND VPWR VPWR _3260_/C sky130_fd_sc_hd__dlygate4sd1_1
X_4516_ _4596_/A _4955_/D VGND VGND VPWR VPWR _4767_/A sky130_fd_sc_hd__nand2_1
Xhold122 hold122/A VGND VGND VPWR VPWR hold122/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5496_ _5496_/A0 _5559_/A1 _5496_/S VGND VGND VPWR VPWR _5496_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold133 hold133/A VGND VGND VPWR VPWR hold133/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold144 hold144/A VGND VGND VPWR VPWR hold144/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold155 hold155/A VGND VGND VPWR VPWR hold155/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4447_ _4663_/D _4447_/B VGND VGND VPWR VPWR _4714_/B sky130_fd_sc_hd__and2b_4
Xhold166 hold166/A VGND VGND VPWR VPWR _6710_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold177 hold177/A VGND VGND VPWR VPWR hold177/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold188 hold188/A VGND VGND VPWR VPWR hold845/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold199 hold199/A VGND VGND VPWR VPWR wb_dat_o[20] sky130_fd_sc_hd__buf_12
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7166_ _3950_/A1 _7166_/D fanout482/X VGND VGND VPWR VPWR _7166_/Q sky130_fd_sc_hd__dfrtp_1
X_4378_ _4917_/A _4701_/A VGND VGND VPWR VPWR _4717_/B sky130_fd_sc_hd__and2b_4
XFILLER_58_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_1_csclk _6727_/CLK VGND VGND VPWR VPWR _6588_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_86_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6117_ _6141_/A1 _6116_/X _6342_/S VGND VGND VPWR VPWR _7176_/D sky130_fd_sc_hd__mux2_1
X_3329_ _3430_/A _3390_/B VGND VGND VPWR VPWR _3648_/A sky130_fd_sc_hd__nand2_8
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7097_ _7097_/CLK _7097_/D fanout468/X VGND VGND VPWR VPWR _7097_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6048_ _6878_/Q _6004_/X _6005_/X _6942_/Q VGND VGND VPWR VPWR _6048_/X sky130_fd_sc_hd__a22o_1
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2090 _7029_/Q VGND VGND VPWR VPWR hold795/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_77_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3680_ _6580_/Q _4128_/A _4304_/A _6733_/Q VGND VGND VPWR VPWR _3680_/X sky130_fd_sc_hd__a22o_2
XFILLER_9_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5350_ hold984/X _5503_/A1 _5352_/S VGND VGND VPWR VPWR _5350_/X sky130_fd_sc_hd__mux2_1
Xoutput205 _3933_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[37] sky130_fd_sc_hd__buf_12
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput216 _7213_/X VGND VGND VPWR VPWR mgmt_gpio_out[12] sky130_fd_sc_hd__buf_12
Xoutput227 _7222_/X VGND VGND VPWR VPWR mgmt_gpio_out[24] sky130_fd_sc_hd__buf_12
XFILLER_114_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput238 _7230_/X VGND VGND VPWR VPWR mgmt_gpio_out[34] sky130_fd_sc_hd__buf_12
X_4301_ _4301_/A0 _5581_/A1 _4303_/S VGND VGND VPWR VPWR _6729_/D sky130_fd_sc_hd__mux2_1
Xoutput249 _3956_/X VGND VGND VPWR VPWR pad_flash_csb sky130_fd_sc_hd__buf_12
XFILLER_126_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5281_ _5281_/A _5569_/B VGND VGND VPWR VPWR _5289_/S sky130_fd_sc_hd__and2_4
X_7020_ _7020_/CLK _7020_/D fanout458/X VGND VGND VPWR VPWR _7020_/Q sky130_fd_sc_hd__dfrtp_4
X_4232_ _4232_/A0 _4231_/X _4240_/S VGND VGND VPWR VPWR _6663_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4163_ _4163_/A0 _5538_/A1 _4163_/S VGND VGND VPWR VPWR _4163_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4094_ _4094_/A0 _5193_/A1 _4097_/S VGND VGND VPWR VPWR _6549_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6804_ _7125_/CLK _6804_/D fanout454/X VGND VGND VPWR VPWR _6804_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_63_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4996_ _4691_/B _4990_/Y _5081_/B VGND VGND VPWR VPWR _4999_/B sky130_fd_sc_hd__a21oi_1
X_6735_ _6757_/CLK _6735_/D fanout447/X VGND VGND VPWR VPWR _6735_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3947_ _3238_/Y _6436_/Q _6432_/B VGND VGND VPWR VPWR _3947_/X sky130_fd_sc_hd__mux2_4
XFILLER_149_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6666_ _6809_/CLK _6666_/D fanout444/X VGND VGND VPWR VPWR _6666_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_137_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3878_ wire1/X hold133/A _3878_/S VGND VGND VPWR VPWR _6438_/D sky130_fd_sc_hd__mux2_1
X_5617_ _7148_/Q _5613_/B _7149_/Q VGND VGND VPWR VPWR _5617_/X sky130_fd_sc_hd__o21a_1
XFILLER_118_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6597_ _6747_/CLK _6597_/D fanout450/X VGND VGND VPWR VPWR _6597_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_191_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5548_ hold49/X hold20/X _5550_/S VGND VGND VPWR VPWR _5548_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5479_ _5479_/A _5551_/B VGND VGND VPWR VPWR _5487_/S sky130_fd_sc_hd__and2_4
XFILLER_105_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7218_ _7218_/A VGND VGND VPWR VPWR _7218_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout410 hold1304/X VGND VGND VPWR VPWR hold153/A sky130_fd_sc_hd__buf_6
XFILLER_160_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout421 _6659_/Q VGND VGND VPWR VPWR _3996_/S sky130_fd_sc_hd__buf_12
Xfanout443 fanout445/X VGND VGND VPWR VPWR fanout443/X sky130_fd_sc_hd__buf_6
Xfanout454 fanout457/X VGND VGND VPWR VPWR fanout454/X sky130_fd_sc_hd__buf_12
X_7149_ _7152_/CLK _7149_/D fanout468/X VGND VGND VPWR VPWR _7149_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_98_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout465 fanout466/X VGND VGND VPWR VPWR fanout465/X sky130_fd_sc_hd__buf_12
Xfanout476 fanout481/X VGND VGND VPWR VPWR fanout476/X sky130_fd_sc_hd__buf_12
XFILLER_19_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4850_ _4402_/Y _4570_/C _4638_/Y _4674_/Y VGND VGND VPWR VPWR _4870_/A sky130_fd_sc_hd__o22a_1
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3801_ _3801_/A _3801_/B _3801_/C _3801_/D VGND VGND VPWR VPWR _3802_/D sky130_fd_sc_hd__nor4_1
XFILLER_33_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4781_ _4368_/A _4477_/Y _4729_/A _4550_/Y VGND VGND VPWR VPWR _4802_/B sky130_fd_sc_hd__o31a_1
X_6520_ _6522_/CLK _6520_/D fanout479/X VGND VGND VPWR VPWR _6520_/Q sky130_fd_sc_hd__dfrtp_1
X_3732_ input21/X _3336_/Y _4200_/A _6640_/Q _3731_/X VGND VGND VPWR VPWR _3735_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_159_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6451_ _6794_/CLK _6451_/D fanout442/X VGND VGND VPWR VPWR _6451_/Q sky130_fd_sc_hd__dfrtp_4
X_3663_ _6919_/Q _5335_/A _3660_/X _3662_/X VGND VGND VPWR VPWR _3664_/C sky130_fd_sc_hd__a211o_1
XFILLER_174_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5402_ hold487/X _5555_/A1 _5406_/S VGND VGND VPWR VPWR _5402_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6382_ _6686_/Q _6382_/A2 _6382_/B1 _6685_/Q VGND VGND VPWR VPWR _6382_/X sky130_fd_sc_hd__a22o_1
X_3594_ _6787_/Q _5178_/A _4182_/A _6627_/Q _3593_/X VGND VGND VPWR VPWR _3595_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5333_ hold951/X hold78/X _5334_/S VGND VGND VPWR VPWR _5333_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5264_ hold646/X _5570_/A1 _5271_/S VGND VGND VPWR VPWR _5264_/X sky130_fd_sc_hd__mux2_1
X_7003_ _7138_/CLK _7003_/D fanout477/X VGND VGND VPWR VPWR _7003_/Q sky130_fd_sc_hd__dfrtp_4
X_4215_ hold257/X _5581_/A1 _4217_/S VGND VGND VPWR VPWR _4215_/X sky130_fd_sc_hd__mux2_1
X_5195_ hold599/X _5195_/A1 _5199_/S VGND VGND VPWR VPWR _6798_/D sky130_fd_sc_hd__mux2_1
X_4146_ _4146_/A _5220_/C VGND VGND VPWR VPWR _4151_/S sky130_fd_sc_hd__and2_4
XFILLER_28_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4077_ _4077_/A _5407_/B VGND VGND VPWR VPWR _4082_/S sky130_fd_sc_hd__and2_4
XFILLER_56_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4979_ _4510_/A _4570_/C _4564_/Y _4968_/Y VGND VGND VPWR VPWR _4983_/B sky130_fd_sc_hd__a31o_1
XFILLER_133_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6718_ _6749_/CLK _6718_/D fanout439/X VGND VGND VPWR VPWR _6718_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_7_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6649_ _6761_/CLK _6649_/D _6426_/A VGND VGND VPWR VPWR _6649_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_137_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_49_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7130_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_75_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4000_ _4000_/A _5220_/C VGND VGND VPWR VPWR _4008_/S sky130_fd_sc_hd__and2_4
XFILLER_38_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5951_ _6598_/Q _5670_/X _5685_/X _6773_/Q VGND VGND VPWR VPWR _5951_/X sky130_fd_sc_hd__a22o_1
XFILLER_92_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4902_ _4902_/A _5073_/C _5063_/C _5098_/B VGND VGND VPWR VPWR _4903_/D sky130_fd_sc_hd__and4_1
XFILLER_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5882_ _5903_/A1 _5881_/X _6342_/S VGND VGND VPWR VPWR _5882_/X sky130_fd_sc_hd__mux2_1
X_4833_ _4683_/A _4832_/X _5127_/B _5104_/C _5021_/A VGND VGND VPWR VPWR _4834_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_178_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4764_ _5150_/A _4764_/B VGND VGND VPWR VPWR _4791_/B sky130_fd_sc_hd__nand2_1
X_6503_ _7139_/CLK _6503_/D fanout478/X VGND VGND VPWR VPWR _6503_/Q sky130_fd_sc_hd__dfrtp_2
X_3715_ _6950_/Q _5371_/A _5488_/A _7054_/Q _3714_/X VGND VGND VPWR VPWR _3716_/D
+ sky130_fd_sc_hd__a221o_1
X_4695_ _4826_/A _4719_/B VGND VGND VPWR VPWR _4922_/B sky130_fd_sc_hd__nand2_2
XFILLER_119_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6434_ _6656_/CLK _6434_/D _6390_/X VGND VGND VPWR VPWR _6434_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_134_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3646_ _6983_/Q _5407_/A _3391_/Y _6812_/Q VGND VGND VPWR VPWR _3646_/X sky130_fd_sc_hd__a22o_1
X_6365_ _6686_/Q _6365_/A2 _6365_/B1 _6685_/Q _6364_/X VGND VGND VPWR VPWR _6365_/X
+ sky130_fd_sc_hd__a221o_1
X_3577_ _7136_/Q hold33/A _3311_/Y _7104_/Q VGND VGND VPWR VPWR _3577_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5316_ _5316_/A0 _5577_/A1 _5316_/S VGND VGND VPWR VPWR _5316_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6296_ _6715_/Q _5973_/X _5986_/X _6642_/Q VGND VGND VPWR VPWR _6296_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5247_ hold774/X _5580_/A1 _5253_/S VGND VGND VPWR VPWR _6838_/D sky130_fd_sc_hd__mux2_1
Xhold15 hold15/A VGND VGND VPWR VPWR hold15/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold26 hold26/A VGND VGND VPWR VPWR hold26/X sky130_fd_sc_hd__buf_12
XFILLER_69_761 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold37 hold37/A VGND VGND VPWR VPWR hold37/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1900 hold491/X VGND VGND VPWR VPWR _5393_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1911 hold422/X VGND VGND VPWR VPWR _5421_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1922 _6611_/Q VGND VGND VPWR VPWR hold334/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_152_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold48 hold48/A VGND VGND VPWR VPWR hold48/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5178_ _5178_/A _5220_/C VGND VGND VPWR VPWR _5183_/S sky130_fd_sc_hd__and2_2
Xhold1933 _6887_/Q VGND VGND VPWR VPWR hold283/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold59 hold59/A VGND VGND VPWR VPWR hold59/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1944 _4119_/X VGND VGND VPWR VPWR _6571_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1955 hold313/X VGND VGND VPWR VPWR _4301_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4129_ _4129_/A0 _5208_/A1 _4133_/S VGND VGND VPWR VPWR _6579_/D sky130_fd_sc_hd__mux2_1
Xhold1966 hold436/X VGND VGND VPWR VPWR _5304_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1977 _6869_/Q VGND VGND VPWR VPWR hold645/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1988 _7016_/Q VGND VGND VPWR VPWR hold690/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1999 _7113_/Q VGND VGND VPWR VPWR hold536/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3500_ _3540_/A _3523_/B VGND VGND VPWR VPWR _4128_/A sky130_fd_sc_hd__nor2_8
XFILLER_7_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4480_ _4486_/A _4491_/B VGND VGND VPWR VPWR _4570_/C sky130_fd_sc_hd__nand2_4
Xhold507 hold507/A VGND VGND VPWR VPWR hold507/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold518 hold518/A VGND VGND VPWR VPWR hold518/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold529 hold529/A VGND VGND VPWR VPWR hold529/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3431_ _3431_/A _3523_/B VGND VGND VPWR VPWR _3431_/Y sky130_fd_sc_hd__nor2_8
XFILLER_144_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6150_ _6978_/Q _5976_/B _5993_/X _7010_/Q VGND VGND VPWR VPWR _6150_/X sky130_fd_sc_hd__a22o_1
X_3362_ _7060_/Q _5488_/A _5497_/A _7068_/Q VGND VGND VPWR VPWR _3362_/X sky130_fd_sc_hd__a22o_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _5131_/A _5131_/B _5101_/C VGND VGND VPWR VPWR _5101_/X sky130_fd_sc_hd__and3_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _7119_/Q _5978_/X _5995_/X _6919_/Q _6080_/X VGND VGND VPWR VPWR _6088_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ _3343_/A _3563_/A VGND VGND VPWR VPWR _3293_/Y sky130_fd_sc_hd__nor2_4
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1207 _7010_/Q VGND VGND VPWR VPWR hold493/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5032_ _5032_/A _5032_/B _5032_/C VGND VGND VPWR VPWR _5086_/A sky130_fd_sc_hd__and3_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1218 hold176/X VGND VGND VPWR VPWR _4120_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1229 _7090_/Q VGND VGND VPWR VPWR hold503/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_66_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6983_ _6983_/CLK _6983_/D fanout459/X VGND VGND VPWR VPWR _6983_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5934_ _6750_/Q _5666_/X _5689_/X _6627_/Q VGND VGND VPWR VPWR _5934_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5865_ _6569_/Q _5674_/X _5687_/X _6599_/Q VGND VGND VPWR VPWR _5865_/X sky130_fd_sc_hd__a22o_1
X_4816_ _4729_/A _4688_/B _4688_/C _4583_/B VGND VGND VPWR VPWR _5080_/A sky130_fd_sc_hd__o22a_1
XFILLER_167_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5796_ _6994_/Q _5929_/B VGND VGND VPWR VPWR _5796_/X sky130_fd_sc_hd__and2_1
XFILLER_193_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4747_ _4415_/B _4714_/Y _4746_/Y VGND VGND VPWR VPWR _4747_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_31_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4678_ _4638_/Y _4674_/Y _4676_/Y _4633_/B _5049_/A VGND VGND VPWR VPWR _4678_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_162_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6417_ _6432_/A _6433_/B VGND VGND VPWR VPWR _6417_/X sky130_fd_sc_hd__and2_1
XFILLER_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3629_ _6601_/Q _4152_/A _4164_/A _6611_/Q _3628_/X VGND VGND VPWR VPWR _3636_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6348_ _3737_/Y hold844/A _6354_/S VGND VGND VPWR VPWR _7188_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput105 wb_adr_i[15] VGND VGND VPWR VPWR _4344_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_6279_ _6279_/A _6279_/B _6279_/C _6279_/D VGND VGND VPWR VPWR _6289_/B sky130_fd_sc_hd__nor4_1
Xinput116 wb_adr_i[25] VGND VGND VPWR VPWR _3898_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2420 _6779_/Q VGND VGND VPWR VPWR _3464_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput127 wb_adr_i[6] VGND VGND VPWR VPWR _4447_/B sky130_fd_sc_hd__buf_12
XFILLER_88_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2431 _5773_/X VGND VGND VPWR VPWR _7163_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput138 wb_dat_i[15] VGND VGND VPWR VPWR _6382_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2442 _3920_/X VGND VGND VPWR VPWR _6655_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput149 wb_dat_i[25] VGND VGND VPWR VPWR _6365_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2453 _7161_/Q VGND VGND VPWR VPWR _5750_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2464 _7170_/Q VGND VGND VPWR VPWR _5947_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1730 _7047_/Q VGND VGND VPWR VPWR _5482_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2475 _6489_/Q VGND VGND VPWR VPWR _5611_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1741 hold234/X VGND VGND VPWR VPWR _5205_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2486 _3926_/X VGND VGND VPWR VPWR _6658_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1752 _4261_/X VGND VGND VPWR VPWR _6696_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2497 _6463_/Q VGND VGND VPWR VPWR _3838_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1763 _4199_/X VGND VGND VPWR VPWR _6638_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1774 hold651/X VGND VGND VPWR VPWR _5237_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1785 hold426/X VGND VGND VPWR VPWR _4230_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1796 _5170_/X VGND VGND VPWR VPWR _6769_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_112_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_720 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3980_ _3980_/A0 hold148/X _3996_/S VGND VGND VPWR VPWR _3980_/X sky130_fd_sc_hd__mux2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5650_ _7146_/Q _7147_/Q VGND VGND VPWR VPWR _5689_/B sky130_fd_sc_hd__and2b_4
XFILLER_30_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4601_ _4601_/A _4601_/B VGND VGND VPWR VPWR _4602_/B sky130_fd_sc_hd__nor2_1
XFILLER_175_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5581_ _5581_/A0 _5581_/A1 _5586_/S VGND VGND VPWR VPWR _7135_/D sky130_fd_sc_hd__mux2_1
XFILLER_191_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4532_ _4607_/B _4934_/B _4981_/A VGND VGND VPWR VPWR _4533_/D sky130_fd_sc_hd__o21ai_1
XFILLER_190_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold304 hold304/A VGND VGND VPWR VPWR hold304/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold315 hold315/A VGND VGND VPWR VPWR hold315/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold326 hold326/A VGND VGND VPWR VPWR hold326/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4463_ _4718_/A _4463_/B VGND VGND VPWR VPWR _4607_/B sky130_fd_sc_hd__nor2_8
Xhold337 hold337/A VGND VGND VPWR VPWR hold337/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold348 hold348/A VGND VGND VPWR VPWR hold348/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6202_ _6860_/Q _5983_/X _6007_/X _6852_/Q VGND VGND VPWR VPWR _6202_/X sky130_fd_sc_hd__a22o_1
XFILLER_104_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold359 hold359/A VGND VGND VPWR VPWR hold359/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3414_ _6875_/Q _5281_/A _5389_/A _6971_/Q _3413_/X VGND VGND VPWR VPWR _3421_/A
+ sky130_fd_sc_hd__a221o_2
X_7182_ _7183_/CLK _7182_/D _6409_/A VGND VGND VPWR VPWR _7182_/Q sky130_fd_sc_hd__dfrtp_1
X_4394_ _4394_/A _4650_/B VGND VGND VPWR VPWR _4394_/Y sky130_fd_sc_hd__nor2_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6133_ _7025_/Q _5971_/X _5990_/X _7057_/Q _6132_/X VGND VGND VPWR VPWR _6133_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3345_ _3487_/A _3470_/A VGND VGND VPWR VPWR _5335_/A sky130_fd_sc_hd__nor2_8
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1004 _6948_/Q VGND VGND VPWR VPWR hold62/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6064_ _6045_/X _6064_/B _6064_/C VGND VGND VPWR VPWR _6064_/Y sky130_fd_sc_hd__nand3b_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3276_ hold88/X _3302_/C VGND VGND VPWR VPWR _3277_/B sky130_fd_sc_hd__nand2_1
Xhold1015 _6956_/Q VGND VGND VPWR VPWR hold45/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_86_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1026 _5432_/X VGND VGND VPWR VPWR _7003_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1037 _6465_/Q VGND VGND VPWR VPWR _3832_/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5015_ _4702_/B _4990_/Y _5014_/X _4822_/Y VGND VGND VPWR VPWR _5015_/X sky130_fd_sc_hd__a211o_1
XFILLER_100_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1048 hold346/X VGND VGND VPWR VPWR _5324_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1059 _3254_/X VGND VGND VPWR VPWR hold87/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_54_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6966_ _7135_/CLK _6966_/D fanout474/X VGND VGND VPWR VPWR _6966_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_53_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5917_ _6734_/Q _5656_/X _5672_/X _6699_/Q _5916_/X VGND VGND VPWR VPWR _5917_/X
+ sky130_fd_sc_hd__a221o_1
X_6897_ _7008_/CLK _6897_/D fanout474/X VGND VGND VPWR VPWR _6897_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5848_ _6876_/Q _5674_/X _5845_/X _5847_/X VGND VGND VPWR VPWR _5848_/X sky130_fd_sc_hd__a211o_1
XFILLER_10_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5779_ _6945_/Q _5658_/X _5666_/X _7001_/Q VGND VGND VPWR VPWR _5779_/X sky130_fd_sc_hd__a22o_1
XFILLER_5_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold860 hold860/A VGND VGND VPWR VPWR hold860/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold871 hold871/A VGND VGND VPWR VPWR hold871/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold882 _3976_/X VGND VGND VPWR VPWR hold12/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold893 _3298_/Y VGND VGND VPWR VPWR _3726_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_150_558 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2250 _7120_/Q VGND VGND VPWR VPWR hold688/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2261 hold695/X VGND VGND VPWR VPWR _5537_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2272 _7072_/Q VGND VGND VPWR VPWR hold696/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2283 _5346_/X VGND VGND VPWR VPWR _6926_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_123_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2294 _7023_/Q VGND VGND VPWR VPWR hold555/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1560 _4273_/X VGND VGND VPWR VPWR _6706_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1571 _6854_/Q VGND VGND VPWR VPWR hold499/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1582 hold826/X VGND VGND VPWR VPWR hold239/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1593 _6553_/Q VGND VGND VPWR VPWR hold840/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6820_ _7103_/CLK _6820_/D fanout472/X VGND VGND VPWR VPWR _6820_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3963_ _3963_/A VGND VGND VPWR VPWR _3963_/Y sky130_fd_sc_hd__inv_2
X_6751_ _6757_/CLK _6751_/D fanout446/X VGND VGND VPWR VPWR _6751_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_189_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5702_ _6893_/Q _5662_/X _5672_/X _6949_/Q VGND VGND VPWR VPWR _5702_/X sky130_fd_sc_hd__a22o_1
X_6682_ _7204_/CLK _6682_/D fanout484/X VGND VGND VPWR VPWR _6682_/Q sky130_fd_sc_hd__dfrtp_4
X_3894_ input118/X input119/X _3894_/C _3894_/D VGND VGND VPWR VPWR _3900_/C sky130_fd_sc_hd__and4bb_1
XFILLER_31_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5633_ _5633_/A1 _5611_/Y _5634_/B _5632_/X VGND VGND VPWR VPWR _7154_/D sky130_fd_sc_hd__a31o_1
XFILLER_176_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5564_ _5564_/A0 _5582_/A1 _5568_/S VGND VGND VPWR VPWR _7120_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold101 hold908/X VGND VGND VPWR VPWR hold909/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4515_ _4462_/Y _4464_/Y _4466_/A _4570_/A _4947_/B VGND VGND VPWR VPWR _5151_/D
+ sky130_fd_sc_hd__o32a_1
Xhold112 _3261_/B VGND VGND VPWR VPWR _3313_/B sky130_fd_sc_hd__buf_2
X_5495_ _5495_/A0 _5585_/A1 _5496_/S VGND VGND VPWR VPWR _5495_/X sky130_fd_sc_hd__mux2_1
Xhold123 hold123/A VGND VGND VPWR VPWR hold123/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold134 hold134/A VGND VGND VPWR VPWR hold134/X sky130_fd_sc_hd__buf_4
XFILLER_144_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold145 hold145/A VGND VGND VPWR VPWR _6855_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4446_ _4498_/B _4663_/D VGND VGND VPWR VPWR _4450_/A sky130_fd_sc_hd__and2b_1
Xhold156 hold156/A VGND VGND VPWR VPWR hold156/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold167 hold167/A VGND VGND VPWR VPWR hold167/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold178 _5238_/X VGND VGND VPWR VPWR _6830_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold189 hold189/A VGND VGND VPWR VPWR wb_dat_o[25] sky130_fd_sc_hd__buf_12
X_7165_ _3950_/A1 _7165_/D fanout473/X VGND VGND VPWR VPWR _7165_/Q sky130_fd_sc_hd__dfrtp_1
X_4377_ _4447_/B _4663_/D VGND VGND VPWR VPWR _4717_/A sky130_fd_sc_hd__nor2_8
XFILLER_86_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116_ _6116_/A0 _6115_/X _6166_/S VGND VGND VPWR VPWR _6116_/X sky130_fd_sc_hd__mux2_1
X_3328_ _3429_/A hold66/X _3390_/B VGND VGND VPWR VPWR _3328_/X sky130_fd_sc_hd__and3_2
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7096_ _7126_/CLK _7096_/D fanout475/X VGND VGND VPWR VPWR _7096_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6047_ _6926_/Q _5982_/X _6016_/X _7038_/Q _6046_/X VGND VGND VPWR VPWR _6054_/A
+ sky130_fd_sc_hd__a221o_1
X_3259_ hold88/X _3259_/B VGND VGND VPWR VPWR hold89/A sky130_fd_sc_hd__and2_1
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6949_ _7132_/CLK _6949_/D fanout459/X VGND VGND VPWR VPWR _6949_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_53_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold690 hold690/A VGND VGND VPWR VPWR hold690/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2080 _6909_/Q VGND VGND VPWR VPWR hold813/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_92_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2091 _6789_/Q VGND VGND VPWR VPWR hold776/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1390 _6517_/Q VGND VGND VPWR VPWR hold215/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput206 _3185_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[3] sky130_fd_sc_hd__buf_12
Xoutput217 _3951_/X VGND VGND VPWR VPWR mgmt_gpio_out[13] sky130_fd_sc_hd__buf_12
X_4300_ _4300_/A0 _5544_/A1 _4303_/S VGND VGND VPWR VPWR _4300_/X sky130_fd_sc_hd__mux2_1
Xoutput228 _7223_/X VGND VGND VPWR VPWR mgmt_gpio_out[25] sky130_fd_sc_hd__buf_12
XFILLER_153_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput239 _3938_/X VGND VGND VPWR VPWR mgmt_gpio_out[35] sky130_fd_sc_hd__buf_12
X_5280_ _5280_/A0 _5559_/A1 _5280_/S VGND VGND VPWR VPWR _5280_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4231_ _5240_/A0 _5303_/A1 _4239_/S VGND VGND VPWR VPWR _4231_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4162_ _4162_/A0 _5249_/A1 _4163_/S VGND VGND VPWR VPWR _4162_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4093_ _4093_/A0 _5208_/A1 _4097_/S VGND VGND VPWR VPWR _6548_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6803_ _6822_/CLK _6803_/D fanout451/X VGND VGND VPWR VPWR _6803_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4995_ _4995_/A _4995_/B VGND VGND VPWR VPWR _5081_/B sky130_fd_sc_hd__nor2_1
X_6734_ _6742_/CLK _6734_/D fanout440/X VGND VGND VPWR VPWR _6734_/Q sky130_fd_sc_hd__dfstp_4
X_3946_ _6660_/Q input3/X input1/X VGND VGND VPWR VPWR _3946_/X sky130_fd_sc_hd__mux2_8
XFILLER_51_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6665_ _7084_/CLK _6665_/D fanout455/X VGND VGND VPWR VPWR _7210_/A sky130_fd_sc_hd__dfrtp_1
X_3877_ hold133/A hold1/A _3878_/S VGND VGND VPWR VPWR _6439_/D sky130_fd_sc_hd__mux2_1
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5616_ _6491_/Q _5679_/B _5676_/B VGND VGND VPWR VPWR _5620_/S sky130_fd_sc_hd__and3_1
XFILLER_191_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6596_ _6792_/CLK _6596_/D fanout442/X VGND VGND VPWR VPWR _6596_/Q sky130_fd_sc_hd__dfstp_2
X_5547_ _5547_/A0 _5556_/A1 _5550_/S VGND VGND VPWR VPWR _7105_/D sky130_fd_sc_hd__mux2_1
XFILLER_155_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5478_ hold992/X hold6/X _5478_/S VGND VGND VPWR VPWR _5478_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7217_ _7217_/A VGND VGND VPWR VPWR _7217_/X sky130_fd_sc_hd__clkbuf_2
X_4429_ _4637_/A _4575_/C _4637_/D VGND VGND VPWR VPWR _4808_/B sky130_fd_sc_hd__and3_4
Xfanout400 hold134/X VGND VGND VPWR VPWR hold135/A sky130_fd_sc_hd__buf_6
Xfanout411 _5229_/C VGND VGND VPWR VPWR _5220_/C sky130_fd_sc_hd__buf_8
XFILLER_132_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout444 fanout445/X VGND VGND VPWR VPWR fanout444/X sky130_fd_sc_hd__buf_12
X_7148_ _7204_/CLK _7148_/D fanout468/X VGND VGND VPWR VPWR _7148_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout455 fanout456/X VGND VGND VPWR VPWR fanout455/X sky130_fd_sc_hd__buf_12
Xfanout466 fanout482/X VGND VGND VPWR VPWR fanout466/X sky130_fd_sc_hd__clkbuf_16
Xfanout477 fanout479/X VGND VGND VPWR VPWR fanout477/X sky130_fd_sc_hd__buf_12
XFILLER_47_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7079_ _7079_/CLK _7079_/D fanout470/X VGND VGND VPWR VPWR _7079_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3800_ _6925_/Q _5344_/A _3311_/Y _7101_/Q _3799_/X VGND VGND VPWR VPWR _3801_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4780_ _4947_/A _4688_/A _4544_/Y VGND VGND VPWR VPWR _4800_/C sky130_fd_sc_hd__o21a_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3731_ _6693_/Q _4256_/A _4262_/A _6698_/Q VGND VGND VPWR VPWR _3731_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_0_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6742_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_174_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6450_ _6794_/CLK _6450_/D fanout444/X VGND VGND VPWR VPWR _6450_/Q sky130_fd_sc_hd__dfrtp_4
X_3662_ _6879_/Q _5290_/A _4128_/A _6581_/Q _3661_/X VGND VGND VPWR VPWR _3662_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5401_ _5401_/A0 _5518_/A1 _5406_/S VGND VGND VPWR VPWR _6975_/D sky130_fd_sc_hd__mux2_1
X_6381_ _6380_/X hold897/X _6384_/S VGND VGND VPWR VPWR _7201_/D sky130_fd_sc_hd__mux2_1
X_3593_ _7040_/Q _5470_/A _5497_/A _7064_/Q VGND VGND VPWR VPWR _3593_/X sky130_fd_sc_hd__a22o_2
X_5332_ _5332_/A0 _5503_/A1 _5334_/S VGND VGND VPWR VPWR _5332_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5263_ _5263_/A _5407_/B VGND VGND VPWR VPWR _5271_/S sky130_fd_sc_hd__and2_4
XFILLER_87_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7002_ _7100_/CLK _7002_/D fanout458/X VGND VGND VPWR VPWR _7002_/Q sky130_fd_sc_hd__dfrtp_4
X_4214_ _4214_/A0 _5544_/A1 _4217_/S VGND VGND VPWR VPWR _4214_/X sky130_fd_sc_hd__mux2_1
X_5194_ hold173/X _5518_/A1 _5199_/S VGND VGND VPWR VPWR _6797_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4145_ _4145_/A0 _5196_/A1 _4145_/S VGND VGND VPWR VPWR _6593_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4076_ _4076_/A0 _5196_/A1 _4076_/S VGND VGND VPWR VPWR _4076_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4978_ _4491_/Y _4655_/A _4581_/X _4969_/B _4905_/X VGND VGND VPWR VPWR _5103_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_51_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6717_ _6788_/CLK _6717_/D _3959_/B VGND VGND VPWR VPWR _6717_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_177_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3929_ _6655_/Q _6658_/Q VGND VGND VPWR VPWR _3929_/Y sky130_fd_sc_hd__nor2_1
XFILLER_177_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6648_ _6648_/CLK _6648_/D fanout449/X VGND VGND VPWR VPWR _6648_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_166_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6579_ _6808_/CLK _6579_/D fanout439/X VGND VGND VPWR VPWR _6579_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_105_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5950_ _3241_/Y _5872_/B _5677_/B VGND VGND VPWR VPWR _5950_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_65_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4901_ _5149_/A _4901_/B VGND VGND VPWR VPWR _5098_/B sky130_fd_sc_hd__and2_1
X_5881_ _7167_/Q _5880_/X _6341_/S VGND VGND VPWR VPWR _5881_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4832_ _4831_/X _4832_/B _4832_/C _4832_/D VGND VGND VPWR VPWR _4832_/X sky130_fd_sc_hd__and4b_1
XANTENNA_190 _5303_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4763_ _4477_/C _4765_/B _4972_/A _4955_/D _5150_/C VGND VGND VPWR VPWR _4764_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_147_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6502_ _6522_/CLK _6502_/D fanout478/X VGND VGND VPWR VPWR _6502_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_159_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3714_ _6966_/Q _5389_/A _4158_/A _6605_/Q VGND VGND VPWR VPWR _3714_/X sky130_fd_sc_hd__a22o_1
X_4694_ _4811_/B _4988_/A _4693_/B VGND VGND VPWR VPWR _4694_/Y sky130_fd_sc_hd__o21ai_1
X_6433_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6433_/X sky130_fd_sc_hd__and2_1
X_3645_ _3645_/A _3645_/B _3645_/C _3645_/D VGND VGND VPWR VPWR _3674_/A sky130_fd_sc_hd__nor4_1
XFILLER_174_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6364_ _6684_/Q _6364_/A2 _6364_/B1 _4218_/Y VGND VGND VPWR VPWR _6364_/X sky130_fd_sc_hd__a22o_1
X_3576_ _6944_/Q _5362_/A _5202_/A _6807_/Q _3568_/X VGND VGND VPWR VPWR _3580_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_136_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5315_ _5315_/A0 _5576_/A1 _5316_/S VGND VGND VPWR VPWR _5315_/X sky130_fd_sc_hd__mux2_1
X_6295_ _6725_/Q _5978_/X _6008_/X _6740_/Q _6294_/X VGND VGND VPWR VPWR _6295_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_114_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5246_ hold335/X hold153/X _5253_/S VGND VGND VPWR VPWR _5246_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold16 hold16/A VGND VGND VPWR VPWR hold16/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1901 _6700_/Q VGND VGND VPWR VPWR hold644/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold27 hold27/A VGND VGND VPWR VPWR hold27/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold38 hold38/A VGND VGND VPWR VPWR hold38/X sky130_fd_sc_hd__buf_2
X_5177_ hold757/X _5186_/A1 _5177_/S VGND VGND VPWR VPWR _5177_/X sky130_fd_sc_hd__mux2_1
Xhold49 hold49/A VGND VGND VPWR VPWR hold49/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1912 _5421_/X VGND VGND VPWR VPWR _6993_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1923 _6649_/Q VGND VGND VPWR VPWR hold659/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1934 hold283/X VGND VGND VPWR VPWR _5302_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1945 _6530_/Q VGND VGND VPWR VPWR hold619/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4128_ _4128_/A _5229_/C VGND VGND VPWR VPWR _4133_/S sky130_fd_sc_hd__and2_4
Xhold1956 _6761_/Q VGND VGND VPWR VPWR hold554/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1967 _7087_/Q VGND VGND VPWR VPWR hold324/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1978 _5282_/X VGND VGND VPWR VPWR _6869_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1989 hold690/X VGND VGND VPWR VPWR _5447_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4059_ hold540/X _5572_/A1 hold14/X VGND VGND VPWR VPWR _4059_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold508 hold508/A VGND VGND VPWR VPWR hold508/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3430_ _3430_/A _3430_/B VGND VGND VPWR VPWR _3523_/B sky130_fd_sc_hd__nand2_8
Xhold519 hold519/A VGND VGND VPWR VPWR hold519/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3361_ _6852_/Q hold40/A _4241_/A input60/X VGND VGND VPWR VPWR _3361_/X sky130_fd_sc_hd__a22o_1
XFILLER_98_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5100_ _5099_/X _5100_/B _5100_/C _5100_/D VGND VGND VPWR VPWR _5101_/C sky130_fd_sc_hd__and4b_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6080_ _7103_/Q _6008_/X _6016_/X _7039_/Q VGND VGND VPWR VPWR _6080_/X sky130_fd_sc_hd__a22o_1
XFILLER_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3292_ _3349_/A _3354_/A VGND VGND VPWR VPWR _5425_/A sky130_fd_sc_hd__nor2_8
XFILLER_112_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _4596_/A _4812_/A _4392_/X VGND VGND VPWR VPWR _5032_/C sky130_fd_sc_hd__a21oi_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1208 hold493/X VGND VGND VPWR VPWR _5440_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1219 _4120_/X VGND VGND VPWR VPWR _6572_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_66_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6982_ _7126_/CLK _6982_/D fanout474/X VGND VGND VPWR VPWR _6982_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_81_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5933_ _6622_/Q _5686_/X _5929_/X _5932_/X VGND VGND VPWR VPWR _5933_/X sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_33_csclk _6850_/CLK VGND VGND VPWR VPWR _7123_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_40_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5864_ _6644_/Q _5668_/X _5686_/X _6619_/Q _5863_/X VGND VGND VPWR VPWR _5869_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4815_ _4583_/B _4676_/Y _4688_/A _4729_/A VGND VGND VPWR VPWR _4815_/X sky130_fd_sc_hd__o22a_1
X_5795_ _5816_/A1 _5794_/X _6342_/S VGND VGND VPWR VPWR _7164_/D sky130_fd_sc_hd__mux2_1
XFILLER_119_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4746_ _4746_/A _4746_/B VGND VGND VPWR VPWR _4746_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_48_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7020_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_119_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4677_ _4726_/C _4677_/B VGND VGND VPWR VPWR _5049_/A sky130_fd_sc_hd__nand2_1
XFILLER_162_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6416_ _6432_/A _6433_/B VGND VGND VPWR VPWR _6416_/X sky130_fd_sc_hd__and2_1
XFILLER_174_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3628_ _6694_/Q _4256_/A _4182_/A _6626_/Q VGND VGND VPWR VPWR _3628_/X sky130_fd_sc_hd__a22o_1
X_6347_ _3803_/Y hold848/A _6354_/S VGND VGND VPWR VPWR _7187_/D sky130_fd_sc_hd__mux2_1
XFILLER_162_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3559_ _3618_/A1 _4112_/A0 _3857_/B VGND VGND VPWR VPWR _3559_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6278_ _6754_/Q _5638_/X _6007_/X _6532_/Q _6277_/X VGND VGND VPWR VPWR _6279_/D
+ sky130_fd_sc_hd__a221o_1
Xhold2410 hold750/X VGND VGND VPWR VPWR _5376_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput106 wb_adr_i[16] VGND VGND VPWR VPWR _4343_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput117 wb_adr_i[26] VGND VGND VPWR VPWR _3894_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2421 _3464_/X VGND VGND VPWR VPWR _6779_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput128 wb_adr_i[7] VGND VGND VPWR VPWR _4663_/D sky130_fd_sc_hd__buf_12
XFILLER_102_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2432 _7182_/Q VGND VGND VPWR VPWR _6291_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput139 wb_dat_i[16] VGND VGND VPWR VPWR _6362_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2443 _7198_/Q VGND VGND VPWR VPWR _6372_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5229_ hold90/A _5229_/B _5229_/C VGND VGND VPWR VPWR hold91/A sky130_fd_sc_hd__and3_2
XFILLER_88_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2454 _6680_/Q VGND VGND VPWR VPWR _3188_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1720 _5528_/X VGND VGND VPWR VPWR _7088_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2465 _5926_/X VGND VGND VPWR VPWR _7170_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1731 _5482_/X VGND VGND VPWR VPWR hold75/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2476 _3923_/Y VGND VGND VPWR VPWR _6489_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1742 _6880_/Q VGND VGND VPWR VPWR hold452/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2487 _6685_/Q VGND VGND VPWR VPWR _3918_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2498 _6459_/Q VGND VGND VPWR VPWR _3850_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1753 _7112_/Q VGND VGND VPWR VPWR hold453/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1764 _6452_/Q VGND VGND VPWR VPWR hold202/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1775 _6634_/Q VGND VGND VPWR VPWR hold711/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1786 _4230_/X VGND VGND VPWR VPWR _6662_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1797 _6645_/Q VGND VGND VPWR VPWR hold566/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_90 _3881_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4600_ _4402_/Y _4570_/A _4658_/B _4564_/Y VGND VGND VPWR VPWR _4609_/B sky130_fd_sc_hd__o22a_1
XFILLER_176_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5580_ hold775/X _5580_/A1 _5586_/S VGND VGND VPWR VPWR _7134_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4531_ _5117_/A _4531_/B _5095_/A VGND VGND VPWR VPWR _4533_/C sky130_fd_sc_hd__and3_1
XFILLER_184_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold305 hold305/A VGND VGND VPWR VPWR hold305/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold316 hold316/A VGND VGND VPWR VPWR hold316/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4462_ _4477_/A _4477_/B _4955_/C VGND VGND VPWR VPWR _4462_/Y sky130_fd_sc_hd__nand3_4
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold327 hold327/A VGND VGND VPWR VPWR hold327/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold338 _6508_/Q VGND VGND VPWR VPWR hold338/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6201_ _6980_/Q _5976_/B _5978_/X _7124_/Q _6200_/X VGND VGND VPWR VPWR _6204_/C
+ sky130_fd_sc_hd__a221o_1
Xhold349 hold981/X VGND VGND VPWR VPWR hold982/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3413_ _7123_/Q hold67/A _5362_/A _6947_/Q VGND VGND VPWR VPWR _3413_/X sky130_fd_sc_hd__a22o_1
X_4393_ _4720_/C _4649_/B VGND VGND VPWR VPWR _4650_/B sky130_fd_sc_hd__nor2_8
X_7181_ _7203_/CLK _7181_/D _6409_/A VGND VGND VPWR VPWR _7181_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3344_ _3563_/A _3764_/A VGND VGND VPWR VPWR _4241_/A sky130_fd_sc_hd__nor2_8
X_6132_ _6905_/Q _5985_/X _5989_/X _6897_/Q VGND VGND VPWR VPWR _6132_/X sky130_fd_sc_hd__a22o_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ _3501_/A _3343_/A VGND VGND VPWR VPWR _5452_/A sky130_fd_sc_hd__nor2_8
XFILLER_98_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6063_ _6056_/X _6058_/X _6063_/C _6339_/B VGND VGND VPWR VPWR _6064_/C sky130_fd_sc_hd__and4bb_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1005 hold62/X VGND VGND VPWR VPWR _5370_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1016 hold45/X VGND VGND VPWR VPWR _5379_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_112_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1027 _6440_/Q VGND VGND VPWR VPWR hold8/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1038 _3250_/X VGND VGND VPWR VPWR _3252_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5014_ _5009_/A _5009_/B _4719_/B VGND VGND VPWR VPWR _5014_/X sky130_fd_sc_hd__o21a_1
Xhold1049 _5324_/X VGND VGND VPWR VPWR _6907_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6965_ _7053_/CLK _6965_/D fanout454/X VGND VGND VPWR VPWR _6965_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_54_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5916_ _6641_/Q _5655_/X _5663_/X _6631_/Q _5905_/Y VGND VGND VPWR VPWR _5916_/X
+ sky130_fd_sc_hd__a221o_1
X_6896_ _7091_/CLK _6896_/D fanout471/X VGND VGND VPWR VPWR _6896_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5847_ _6956_/Q _5672_/X _5679_/X _6908_/Q _5846_/X VGND VGND VPWR VPWR _5847_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5778_ _7033_/Q _5655_/X _5668_/X _7057_/Q VGND VGND VPWR VPWR _5778_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4729_ _4729_/A _4995_/A VGND VGND VPWR VPWR _5081_/A sky130_fd_sc_hd__nor2_1
XFILLER_147_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold850 hold850/A VGND VGND VPWR VPWR hold850/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold861 hold861/A VGND VGND VPWR VPWR hold861/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold872 hold872/A VGND VGND VPWR VPWR hold872/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold883 hold12/X VGND VGND VPWR VPWR _5407_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold894 _3311_/Y VGND VGND VPWR VPWR _5542_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2240 _7040_/Q VGND VGND VPWR VPWR hold681/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2251 hold688/X VGND VGND VPWR VPWR _5564_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2262 _6870_/Q VGND VGND VPWR VPWR hold754/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2273 hold696/X VGND VGND VPWR VPWR _5510_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_184_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2284 _7119_/Q VGND VGND VPWR VPWR hold559/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1550 hold709/X VGND VGND VPWR VPWR _4269_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2295 hold555/X VGND VGND VPWR VPWR _5455_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1561 _7004_/Q VGND VGND VPWR VPWR hold528/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1572 _5265_/X VGND VGND VPWR VPWR hold500/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1583 _6557_/Q VGND VGND VPWR VPWR hold858/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1594 hold840/X VGND VGND VPWR VPWR hold265/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6750_ _6750_/CLK _6750_/D fanout446/X VGND VGND VPWR VPWR _6750_/Q sky130_fd_sc_hd__dfrtp_4
X_3962_ _6456_/Q _3962_/B VGND VGND VPWR VPWR _3963_/A sky130_fd_sc_hd__nor2_4
XFILLER_51_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5701_ _6981_/Q _5656_/X _5663_/X _7021_/Q _5700_/X VGND VGND VPWR VPWR _5701_/X
+ sky130_fd_sc_hd__a221o_1
X_6681_ _7152_/CLK _6681_/D fanout484/X VGND VGND VPWR VPWR _6681_/Q sky130_fd_sc_hd__dfrtp_4
X_3893_ input123/X input122/X _3893_/C _3893_/D VGND VGND VPWR VPWR _3900_/B sky130_fd_sc_hd__and4bb_1
XFILLER_188_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5632_ _6491_/Q _6015_/B _6014_/A VGND VGND VPWR VPWR _5632_/X sky130_fd_sc_hd__and3_1
XFILLER_148_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5563_ _5563_/A0 _5572_/A1 _5568_/S VGND VGND VPWR VPWR _7119_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4514_ _4729_/A _4514_/B VGND VGND VPWR VPWR _4514_/Y sky130_fd_sc_hd__nor2_1
Xhold102 _3272_/A VGND VGND VPWR VPWR _3285_/B sky130_fd_sc_hd__clkbuf_2
X_5494_ _5494_/A0 _5503_/A1 _5496_/S VGND VGND VPWR VPWR _5494_/X sky130_fd_sc_hd__mux2_1
Xhold113 hold113/A VGND VGND VPWR VPWR _6756_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold124 hold935/X VGND VGND VPWR VPWR hold936/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold135 hold135/A VGND VGND VPWR VPWR hold135/X sky130_fd_sc_hd__buf_8
XFILLER_160_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7233_ _7233_/A VGND VGND VPWR VPWR _7233_/X sky130_fd_sc_hd__buf_2
XFILLER_105_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold146 hold146/A VGND VGND VPWR VPWR hold146/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4445_ _4598_/A _4564_/B VGND VGND VPWR VPWR _4483_/B sky130_fd_sc_hd__and2_4
Xhold157 hold157/A VGND VGND VPWR VPWR hold157/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold168 hold168/A VGND VGND VPWR VPWR hold168/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold179 hold179/A VGND VGND VPWR VPWR hold179/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7164_ _7204_/CLK _7164_/D fanout468/X VGND VGND VPWR VPWR _7164_/Q sky130_fd_sc_hd__dfrtp_1
X_4376_ _4649_/B _4560_/A VGND VGND VPWR VPWR _4384_/A sky130_fd_sc_hd__nand2_8
XFILLER_113_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6115_ _6840_/Q _6011_/Y _6114_/X VGND VGND VPWR VPWR _6115_/X sky130_fd_sc_hd__o21ba_1
X_3327_ _3338_/A _3535_/A VGND VGND VPWR VPWR _5488_/A sky130_fd_sc_hd__nor2_8
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7095_ _7111_/CLK _7095_/D fanout472/X VGND VGND VPWR VPWR _7095_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ _7078_/Q _6013_/X _6017_/X _7070_/Q VGND VGND VPWR VPWR _6046_/X sky130_fd_sc_hd__a22o_1
XFILLER_37_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3258_ _3260_/C VGND VGND VPWR VPWR _3302_/C sky130_fd_sc_hd__inv_2
XFILLER_100_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3189_ _6680_/D VGND VGND VPWR VPWR _3189_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6948_ _7020_/CLK hold63/X fanout458/X VGND VGND VPWR VPWR _6948_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6879_ _7135_/CLK _6879_/D fanout473/X VGND VGND VPWR VPWR _6879_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold680 hold680/A VGND VGND VPWR VPWR hold680/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold691 hold691/A VGND VGND VPWR VPWR hold691/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2070 hold354/X VGND VGND VPWR VPWR _4052_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2081 _7103_/Q VGND VGND VPWR VPWR hold563/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2092 hold776/X VGND VGND VPWR VPWR _5185_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_94_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1380 _6507_/Q VGND VGND VPWR VPWR hold581/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1391 hold215/X VGND VGND VPWR VPWR _4057_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput207 _3236_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[4] sky130_fd_sc_hd__buf_12
XFILLER_142_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput218 _7214_/X VGND VGND VPWR VPWR mgmt_gpio_out[16] sky130_fd_sc_hd__buf_12
Xoutput229 _7224_/X VGND VGND VPWR VPWR mgmt_gpio_out[26] sky130_fd_sc_hd__buf_12
XFILLER_154_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4230_ _4230_/A0 _4229_/X _4240_/S VGND VGND VPWR VPWR _4230_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4161_ hold203/X _4337_/A1 _4163_/S VGND VGND VPWR VPWR _4161_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4092_ _4092_/A _5229_/C VGND VGND VPWR VPWR _4097_/S sky130_fd_sc_hd__and2_4
XFILLER_76_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6802_ _7013_/CLK _6802_/D fanout452/X VGND VGND VPWR VPWR _6802_/Q sky130_fd_sc_hd__dfstp_2
X_4994_ _4676_/Y _4812_/Y _4993_/Y _5138_/B VGND VGND VPWR VPWR _5010_/B sky130_fd_sc_hd__o211a_1
X_6733_ _6742_/CLK _6733_/D fanout440/X VGND VGND VPWR VPWR _6733_/Q sky130_fd_sc_hd__dfrtp_4
X_3945_ _3944_/X _3966_/B _6456_/Q VGND VGND VPWR VPWR _3945_/X sky130_fd_sc_hd__mux2_4
XFILLER_189_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6664_ _7116_/CLK _6664_/D fanout455/X VGND VGND VPWR VPWR _7209_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_176_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3876_ hold1/A hold8/A _3878_/S VGND VGND VPWR VPWR _6440_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5615_ _7149_/Q _7148_/Q VGND VGND VPWR VPWR _5676_/B sky130_fd_sc_hd__nor2_8
X_6595_ _6691_/CLK _6595_/D fanout443/X VGND VGND VPWR VPWR _6595_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5546_ _5546_/A0 _5582_/A1 _5550_/S VGND VGND VPWR VPWR _7104_/D sky130_fd_sc_hd__mux2_1
XFILLER_191_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5477_ _5477_/A0 _5585_/A1 _5478_/S VGND VGND VPWR VPWR _5477_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7216_ _7216_/A VGND VGND VPWR VPWR _7216_/X sky130_fd_sc_hd__clkbuf_2
X_4428_ _4637_/B _4637_/A VGND VGND VPWR VPWR _4463_/B sky130_fd_sc_hd__nand2b_4
Xfanout401 _5499_/A1 VGND VGND VPWR VPWR _5580_/A1 sky130_fd_sc_hd__buf_8
Xfanout412 _5407_/B VGND VGND VPWR VPWR _5229_/C sky130_fd_sc_hd__buf_12
Xclkbuf_2_3__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _3940_/A1
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_160_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7147_ _7203_/CLK _7147_/D _6399_/A VGND VGND VPWR VPWR _7147_/Q sky130_fd_sc_hd__dfstp_4
X_4359_ _4682_/A _4365_/B _4447_/B VGND VGND VPWR VPWR _4360_/B sky130_fd_sc_hd__a21o_1
Xfanout445 fanout450/X VGND VGND VPWR VPWR fanout445/X sky130_fd_sc_hd__buf_8
XFILLER_86_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout456 fanout457/X VGND VGND VPWR VPWR fanout456/X sky130_fd_sc_hd__buf_12
XFILLER_58_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout467 fanout468/X VGND VGND VPWR VPWR _6399_/A sky130_fd_sc_hd__clkbuf_16
Xfanout478 fanout479/X VGND VGND VPWR VPWR fanout478/X sky130_fd_sc_hd__buf_12
X_7078_ _7138_/CLK _7078_/D fanout477/X VGND VGND VPWR VPWR _7078_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6029_ _7093_/Q _5984_/X _6020_/X _6024_/X _6028_/X VGND VGND VPWR VPWR _6029_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_104_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3730_ _7094_/Q _5533_/A _5178_/A _6785_/Q _3729_/X VGND VGND VPWR VPWR _3735_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_159_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3661_ _6550_/Q _4092_/A _4134_/A _6586_/Q VGND VGND VPWR VPWR _3661_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5400_ hold545/X _5499_/A1 _5406_/S VGND VGND VPWR VPWR _6974_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6380_ _6686_/Q _6380_/A2 _6380_/B1 _4218_/Y _6379_/X VGND VGND VPWR VPWR _6380_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3592_ _7000_/Q _5425_/A _4304_/A _6735_/Q _3591_/X VGND VGND VPWR VPWR _3595_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_802 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5331_ _5331_/A0 _5583_/A1 _5334_/S VGND VGND VPWR VPWR _6913_/D sky130_fd_sc_hd__mux2_1
XFILLER_126_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5262_ hold997/X hold6/X _5262_/S VGND VGND VPWR VPWR _5262_/X sky130_fd_sc_hd__mux2_1
X_7001_ _7134_/CLK _7001_/D fanout476/X VGND VGND VPWR VPWR _7001_/Q sky130_fd_sc_hd__dfrtp_4
X_4213_ _4213_/A0 _5221_/A1 _4217_/S VGND VGND VPWR VPWR _4213_/X sky130_fd_sc_hd__mux2_1
X_5193_ hold529/X _5193_/A1 _5199_/S VGND VGND VPWR VPWR _6796_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4144_ _4144_/A0 _5195_/A1 _4145_/S VGND VGND VPWR VPWR _6592_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4075_ _4075_/A0 _5195_/A1 _4076_/S VGND VGND VPWR VPWR _4075_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_4_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_4_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4977_ _4569_/C _4968_/Y _4971_/Y _4972_/Y VGND VGND VPWR VPWR _4984_/B sky130_fd_sc_hd__o211a_1
X_6716_ _6729_/CLK _6716_/D fanout465/X VGND VGND VPWR VPWR _6716_/Q sky130_fd_sc_hd__dfstp_2
X_3928_ _6657_/Q _3904_/A _3904_/Y _6656_/Q VGND VGND VPWR VPWR _6656_/D sky130_fd_sc_hd__a22o_1
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6647_ _6761_/CLK _6647_/D _6426_/A VGND VGND VPWR VPWR _6647_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_149_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3859_ _6470_/Q _3879_/A _6468_/Q _6654_/Q VGND VGND VPWR VPWR _3860_/S sky130_fd_sc_hd__and4b_1
X_6578_ _6808_/CLK _6578_/D fanout439/X VGND VGND VPWR VPWR _6578_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_166_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5529_ _5529_/A0 _5583_/A1 _5532_/S VGND VGND VPWR VPWR _5529_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4900_ _4947_/B _4570_/D _4616_/A VGND VGND VPWR VPWR _5063_/C sky130_fd_sc_hd__o21a_1
XFILLER_18_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5880_ _5869_/Y wire350/X _6525_/Q _5678_/Y VGND VGND VPWR VPWR _5880_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_61_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4831_ _4955_/D _4718_/C _5026_/C _4812_/A VGND VGND VPWR VPWR _4831_/X sky130_fd_sc_hd__a22o_1
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_180 _6502_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_191 _5303_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4762_ _4402_/Y _4583_/B _4426_/Y VGND VGND VPWR VPWR _4791_/A sky130_fd_sc_hd__a21o_1
X_6501_ _7140_/CLK _6501_/D fanout471/X VGND VGND VPWR VPWR _6501_/Q sky130_fd_sc_hd__dfrtp_2
X_3713_ _6894_/Q _5308_/A _3539_/Y _6531_/Q _3712_/X VGND VGND VPWR VPWR _3716_/C
+ sky130_fd_sc_hd__a221o_1
X_4693_ _4811_/B _4693_/B VGND VGND VPWR VPWR _5108_/A sky130_fd_sc_hd__nand2_1
XFILLER_147_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6432_ _6432_/A _6432_/B VGND VGND VPWR VPWR _6432_/X sky130_fd_sc_hd__and2_1
XFILLER_119_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3644_ _7023_/Q _5452_/A _5236_/C wire1/A _3643_/X VGND VGND VPWR VPWR _3645_/D sky130_fd_sc_hd__a221o_2
XFILLER_174_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6363_ _6362_/X hold151/A _6384_/S VGND VGND VPWR VPWR _7195_/D sky130_fd_sc_hd__mux2_1
X_3575_ _6725_/Q _4292_/A _4164_/A _6612_/Q _3574_/X VGND VGND VPWR VPWR _3580_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_127_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5314_ _5314_/A0 _5575_/A1 _5316_/S VGND VGND VPWR VPWR _5314_/X sky130_fd_sc_hd__mux2_1
X_6294_ _6705_/Q _5977_/X _6007_/X _6533_/Q _6293_/X VGND VGND VPWR VPWR _6294_/X
+ sky130_fd_sc_hd__a221o_1
X_5245_ hold27/X hold13/A VGND VGND VPWR VPWR _5245_/X sky130_fd_sc_hd__and2_4
XFILLER_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold17 hold17/A VGND VGND VPWR VPWR hold17/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold28 hold28/A VGND VGND VPWR VPWR hold28/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1902 hold644/X VGND VGND VPWR VPWR _4266_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1913 _7031_/Q VGND VGND VPWR VPWR hold276/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5176_ _5176_/A0 _5208_/A1 _5177_/S VGND VGND VPWR VPWR _5176_/X sky130_fd_sc_hd__mux2_1
Xhold39 hold39/A VGND VGND VPWR VPWR hold39/X sky130_fd_sc_hd__buf_8
XFILLER_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1924 hold659/X VGND VGND VPWR VPWR _4213_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1935 _6693_/Q VGND VGND VPWR VPWR hold613/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4127_ _4127_/A0 _5196_/A1 _4127_/S VGND VGND VPWR VPWR _4127_/X sky130_fd_sc_hd__mux2_1
Xhold1946 hold619/X VGND VGND VPWR VPWR _4072_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1957 hold554/X VGND VGND VPWR VPWR _4339_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1968 hold324/X VGND VGND VPWR VPWR _5527_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1979 _6588_/Q VGND VGND VPWR VPWR hold590/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_83_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4058_ _4058_/A0 _5571_/A1 hold14/X VGND VGND VPWR VPWR _4058_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold509 hold509/A VGND VGND VPWR VPWR hold509/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3360_ _6802_/Q _3319_/Y _3336_/Y input28/X VGND VGND VPWR VPWR _3360_/X sky130_fd_sc_hd__a22o_1
XFILLER_124_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3291_ _3764_/A _3487_/A VGND VGND VPWR VPWR _5371_/A sky130_fd_sc_hd__nor2_8
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _4417_/B _4688_/B _4774_/X _4963_/A _4894_/A VGND VGND VPWR VPWR _5149_/B
+ sky130_fd_sc_hd__o2111a_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1209 _6526_/Q VGND VGND VPWR VPWR hold254/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6981_ _7053_/CLK _6981_/D fanout452/X VGND VGND VPWR VPWR _6981_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_53_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5932_ _6647_/Q _5668_/X _5684_/X _6607_/Q VGND VGND VPWR VPWR _5932_/X sky130_fd_sc_hd__a22o_1
XFILLER_18_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5863_ _6535_/Q _5651_/X _5658_/X _6692_/Q VGND VGND VPWR VPWR _5863_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4814_ _4583_/B _4688_/B _4691_/Y _4729_/A VGND VGND VPWR VPWR _4818_/B sky130_fd_sc_hd__o22a_1
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5794_ _5794_/A0 _5793_/X _6166_/S VGND VGND VPWR VPWR _5794_/X sky130_fd_sc_hd__mux2_1
X_4745_ _5011_/A _4947_/A _4714_/Y VGND VGND VPWR VPWR _4746_/B sky130_fd_sc_hd__a21oi_1
XFILLER_175_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4676_ _4751_/B _4726_/C VGND VGND VPWR VPWR _4676_/Y sky130_fd_sc_hd__nand2_4
XFILLER_119_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6415_ _6432_/A _6433_/B VGND VGND VPWR VPWR _6415_/X sky130_fd_sc_hd__and2_1
XFILLER_134_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3627_ _3627_/A _3627_/B _3627_/C _3627_/D VGND VGND VPWR VPWR _3675_/A sky130_fd_sc_hd__nor4_2
X_6346_ _6677_/Q _6346_/B VGND VGND VPWR VPWR _6354_/S sky130_fd_sc_hd__nand2_8
X_3558_ _3558_/A _3558_/B _3558_/C VGND VGND VPWR VPWR _3558_/Y sky130_fd_sc_hd__nand3_2
XFILLER_103_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6277_ _6626_/Q _6013_/X _6015_/X _6759_/Q VGND VGND VPWR VPWR _6277_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3489_ _6711_/Q _4274_/A _4256_/A _6696_/Q VGND VGND VPWR VPWR _3489_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2400 hold716/X VGND VGND VPWR VPWR _5511_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput107 wb_adr_i[17] VGND VGND VPWR VPWR _4343_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2411 _6929_/Q VGND VGND VPWR VPWR hold752/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput118 wb_adr_i[27] VGND VGND VPWR VPWR input118/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2422 _6683_/Q VGND VGND VPWR VPWR _6680_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5228_ _5228_/A0 hold135/X _5228_/S VGND VGND VPWR VPWR _5228_/X sky130_fd_sc_hd__mux2_1
Xinput129 wb_adr_i[8] VGND VGND VPWR VPWR _4345_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2433 _6267_/X VGND VGND VPWR VPWR _7182_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2444 _6447_/Q VGND VGND VPWR VPWR _3867_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1710 _6904_/Q VGND VGND VPWR VPWR hold446/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2455 _3922_/Y VGND VGND VPWR VPWR _6676_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1721 _7049_/Q VGND VGND VPWR VPWR hold130/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2466 _7174_/Q VGND VGND VPWR VPWR _6067_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1732 _7046_/Q VGND VGND VPWR VPWR hold502/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2477 _7166_/Q VGND VGND VPWR VPWR _5838_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1743 hold452/X VGND VGND VPWR VPWR _5294_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5159_ _5157_/X _5158_/X _5127_/X VGND VGND VPWR VPWR _5159_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_29_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2488 _7179_/Q VGND VGND VPWR VPWR _6192_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2499 _6464_/Q VGND VGND VPWR VPWR _3831_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1754 hold453/X VGND VGND VPWR VPWR _5555_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1765 _6450_/Q VGND VGND VPWR VPWR hold614/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1776 hold711/X VGND VGND VPWR VPWR _4195_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1787 _6661_/Q VGND VGND VPWR VPWR hold430/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1798 hold566/X VGND VGND VPWR VPWR _4208_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_71_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_80 input37/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_91 _3973_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4530_ _4575_/C _4463_/B _4510_/A _4509_/Y _4529_/X VGND VGND VPWR VPWR _4533_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4461_ _4506_/A _4461_/B VGND VGND VPWR VPWR _4955_/C sky130_fd_sc_hd__nor2_4
Xhold306 hold306/A VGND VGND VPWR VPWR hold306/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold317 hold317/A VGND VGND VPWR VPWR _6569_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold328 hold328/A VGND VGND VPWR VPWR hold328/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6200_ _6932_/Q _5982_/X _5999_/X _6868_/Q VGND VGND VPWR VPWR _6200_/X sky130_fd_sc_hd__a22o_1
Xhold339 hold339/A VGND VGND VPWR VPWR _6508_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3412_ _6963_/Q _5380_/A _3407_/X _3409_/X _3411_/X VGND VGND VPWR VPWR _3422_/B
+ sky130_fd_sc_hd__a2111oi_4
X_7180_ _3950_/A1 _7180_/D fanout468/X VGND VGND VPWR VPWR _7180_/Q sky130_fd_sc_hd__dfrtp_1
X_4392_ _4955_/A _5009_/A _4584_/A VGND VGND VPWR VPWR _4392_/X sky130_fd_sc_hd__and3_1
XFILLER_125_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6131_ _7113_/Q _5987_/X _6004_/X _6881_/Q _6130_/X VGND VGND VPWR VPWR _6131_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_125_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _3343_/A _3487_/A VGND VGND VPWR VPWR _5380_/A sky130_fd_sc_hd__nor2_8
XFILLER_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _6902_/Q _5985_/X _6059_/X _6061_/X VGND VGND VPWR VPWR _6063_/C sky130_fd_sc_hd__a211oi_1
X_3274_ _3355_/A hold31/X VGND VGND VPWR VPWR _3343_/A sky130_fd_sc_hd__nand2_8
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1006 _5370_/X VGND VGND VPWR VPWR hold63/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1017 _5379_/X VGND VGND VPWR VPWR hold46/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _4688_/C _4995_/B _5012_/X _4820_/A VGND VGND VPWR VPWR _5023_/C sky130_fd_sc_hd__o211a_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1028 hold8/X VGND VGND VPWR VPWR _3984_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_66_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1039 _3252_/Y VGND VGND VPWR VPWR hold24/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_94_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6964_ _7131_/CLK hold44/X fanout469/X VGND VGND VPWR VPWR _6964_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5915_ _6689_/Q _5659_/X _5687_/X _6601_/Q VGND VGND VPWR VPWR _5915_/X sky130_fd_sc_hd__a22o_1
X_6895_ _7079_/CLK _6895_/D fanout469/X VGND VGND VPWR VPWR _6895_/Q sky130_fd_sc_hd__dfrtp_4
X_5846_ _6940_/Q _5659_/X _5687_/X _6924_/Q VGND VGND VPWR VPWR _5846_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5777_ _6881_/Q _5667_/X _5673_/X _6865_/Q _5776_/X VGND VGND VPWR VPWR _5782_/B
+ sky130_fd_sc_hd__a221o_1
X_4728_ _5150_/B _4730_/B VGND VGND VPWR VPWR _4728_/Y sky130_fd_sc_hd__nand2_1
XFILLER_163_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4659_ _4652_/Y _4677_/B VGND VGND VPWR VPWR _4704_/C sky130_fd_sc_hd__nand2b_1
XFILLER_174_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold840 hold840/A VGND VGND VPWR VPWR hold840/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold851 hold851/A VGND VGND VPWR VPWR hold851/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold862 hold862/A VGND VGND VPWR VPWR hold862/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold873 hold973/X VGND VGND VPWR VPWR hold974/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6329_ _6711_/Q _5992_/X _6012_/X _6751_/Q _6328_/X VGND VGND VPWR VPWR _6329_/X
+ sky130_fd_sc_hd__a221o_1
Xhold884 _5245_/X VGND VGND VPWR VPWR _5253_/S sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_115_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold895 _5548_/X VGND VGND VPWR VPWR hold50/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_107_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2230 _5454_/X VGND VGND VPWR VPWR _7022_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2241 hold681/X VGND VGND VPWR VPWR _5474_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2252 _6629_/Q VGND VGND VPWR VPWR hold804/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_67_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2263 _5283_/X VGND VGND VPWR VPWR _6870_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2274 _5510_/X VGND VGND VPWR VPWR _7072_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2285 hold559/X VGND VGND VPWR VPWR _5563_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1540 hold830/X VGND VGND VPWR VPWR hold242/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1551 _4269_/X VGND VGND VPWR VPWR _6702_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2296 _5455_/X VGND VGND VPWR VPWR _7023_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1562 hold528/X VGND VGND VPWR VPWR _5433_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1573 _6545_/Q VGND VGND VPWR VPWR hold824/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1584 hold858/X VGND VGND VPWR VPWR hold281/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1595 _6546_/Q VGND VGND VPWR VPWR hold822/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_32_csclk _6850_/CLK VGND VGND VPWR VPWR _7139_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_106_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_47_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7100_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_180_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3961_ _3961_/A VGND VGND VPWR VPWR _3961_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5700_ _7013_/Q _5664_/X _5666_/X _6997_/Q VGND VGND VPWR VPWR _5700_/X sky130_fd_sc_hd__a22o_1
XFILLER_149_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6680_ _7152_/CLK _6680_/D _6346_/B VGND VGND VPWR VPWR _6680_/Q sky130_fd_sc_hd__dfrtp_1
X_3892_ _4720_/C _4649_/B _4649_/C _4649_/D VGND VGND VPWR VPWR _4395_/A sky130_fd_sc_hd__a211o_4
XFILLER_189_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5631_ _5631_/A _6017_/B VGND VGND VPWR VPWR _5634_/B sky130_fd_sc_hd__nand2_1
XFILLER_31_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5562_ hold714/X _5571_/A1 _5568_/S VGND VGND VPWR VPWR _7118_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4513_ _4513_/A _4513_/B _4652_/A VGND VGND VPWR VPWR _4514_/B sky130_fd_sc_hd__nand3_4
Xhold103 hold960/X VGND VGND VPWR VPWR _6477_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5493_ _5493_/A0 _5583_/A1 _5496_/S VGND VGND VPWR VPWR _5493_/X sky130_fd_sc_hd__mux2_1
Xhold114 hold927/X VGND VGND VPWR VPWR hold928/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold125 hold125/A VGND VGND VPWR VPWR hold125/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7232_ _7232_/A VGND VGND VPWR VPWR _7232_/X sky130_fd_sc_hd__buf_2
Xhold136 hold136/A VGND VGND VPWR VPWR _6822_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4444_ _4506_/A _4469_/B VGND VGND VPWR VPWR _4564_/B sky130_fd_sc_hd__nor2_4
XFILLER_171_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold147 _4216_/X VGND VGND VPWR VPWR _6652_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold158 hold158/A VGND VGND VPWR VPWR _6612_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold169 _4338_/X VGND VGND VPWR VPWR _6760_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7163_ _3950_/A1 _7163_/D fanout468/X VGND VGND VPWR VPWR _7163_/Q sky130_fd_sc_hd__dfrtp_1
X_4375_ _4649_/B _4560_/A VGND VGND VPWR VPWR _5001_/A sky130_fd_sc_hd__and2_4
XFILLER_59_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6114_ _6105_/X _6339_/B _6114_/C _6114_/D VGND VGND VPWR VPWR _6114_/X sky130_fd_sc_hd__and4b_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3326_ _3535_/A _3470_/A VGND VGND VPWR VPWR _5479_/A sky130_fd_sc_hd__nor2_8
XFILLER_100_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7094_ _7102_/CLK _7094_/D fanout465/X VGND VGND VPWR VPWR _7094_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_113_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _7054_/Q _5990_/X _5997_/X _6950_/Q _6044_/X VGND VGND VPWR VPWR _6045_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ _3256_/X _3257_/A1 _3996_/S VGND VGND VPWR VPWR _3257_/X sky130_fd_sc_hd__mux2_2
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3188_ _3188_/A VGND VGND VPWR VPWR _4222_/B sky130_fd_sc_hd__inv_2
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6947_ _7123_/CLK _6947_/D fanout478/X VGND VGND VPWR VPWR _6947_/Q sky130_fd_sc_hd__dfrtp_4
X_6878_ _7137_/CLK _6878_/D fanout476/X VGND VGND VPWR VPWR _6878_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_22_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5829_ _7067_/Q _5671_/X _5678_/B _6971_/Q _5707_/B VGND VGND VPWR VPWR _5829_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_139_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold670 hold670/A VGND VGND VPWR VPWR hold670/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold681 hold681/A VGND VGND VPWR VPWR hold681/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold692 hold692/A VGND VGND VPWR VPWR hold692/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2060 hold615/X VGND VGND VPWR VPWR _4192_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2071 _7225_/A VGND VGND VPWR VPWR hold674/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2082 hold563/X VGND VGND VPWR VPWR _5545_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2093 _5185_/X VGND VGND VPWR VPWR _6789_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_64_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1370 _5225_/X VGND VGND VPWR VPWR hold249/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1381 hold581/X VGND VGND VPWR VPWR _4044_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1392 _6802_/Q VGND VGND VPWR VPWR hold376/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput208 _3235_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[5] sky130_fd_sc_hd__buf_12
Xoutput219 _7215_/X VGND VGND VPWR VPWR mgmt_gpio_out[17] sky130_fd_sc_hd__buf_12
XFILLER_126_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4160_ hold167/X _5544_/A1 _4163_/S VGND VGND VPWR VPWR _4160_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4091_ _3385_/Y hold830/A _4091_/S VGND VGND VPWR VPWR _6547_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6801_ _7013_/CLK _6801_/D fanout452/X VGND VGND VPWR VPWR _6801_/Q sky130_fd_sc_hd__dfstp_4
X_4993_ _4993_/A _4993_/B VGND VGND VPWR VPWR _4993_/Y sky130_fd_sc_hd__nand2_1
X_6732_ _6747_/CLK _6732_/D _3959_/B VGND VGND VPWR VPWR _6732_/Q sky130_fd_sc_hd__dfrtp_4
X_3944_ _3943_/X input38/X _6458_/Q VGND VGND VPWR VPWR _3944_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6663_ _7116_/CLK _6663_/D fanout455/X VGND VGND VPWR VPWR _7208_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_149_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3875_ hold8/A hold93/A _3878_/S VGND VGND VPWR VPWR _6441_/D sky130_fd_sc_hd__mux2_1
XFILLER_177_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5614_ _5614_/A1 _5613_/B _5611_/Y _5613_/Y VGND VGND VPWR VPWR _7148_/D sky130_fd_sc_hd__a31o_1
XFILLER_176_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6594_ _6792_/CLK _6594_/D fanout442/X VGND VGND VPWR VPWR _6594_/Q sky130_fd_sc_hd__dfrtp_4
X_5545_ _5545_/A0 _5572_/A1 _5550_/S VGND VGND VPWR VPWR _7103_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_0_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_0_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5476_ hold69/X hold20/X _5478_/S VGND VGND VPWR VPWR _5476_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4427_ _4637_/B _4637_/A VGND VGND VPWR VPWR _4488_/B sky130_fd_sc_hd__and2b_4
X_7215_ _7215_/A VGND VGND VPWR VPWR _7215_/X sky130_fd_sc_hd__clkbuf_2
Xfanout402 _5499_/A1 VGND VGND VPWR VPWR _5571_/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout413 _5407_/B VGND VGND VPWR VPWR _5551_/B sky130_fd_sc_hd__buf_12
X_7146_ _7152_/CLK _7146_/D _6399_/A VGND VGND VPWR VPWR _7146_/Q sky130_fd_sc_hd__dfrtp_4
X_4358_ _4513_/A _4560_/A VGND VGND VPWR VPWR _4955_/A sky130_fd_sc_hd__and2b_4
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout435 _6423_/B VGND VGND VPWR VPWR _6433_/B sky130_fd_sc_hd__buf_6
Xfanout446 fanout449/X VGND VGND VPWR VPWR fanout446/X sky130_fd_sc_hd__buf_12
Xfanout457 fanout482/X VGND VGND VPWR VPWR fanout457/X sky130_fd_sc_hd__buf_12
XFILLER_86_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3309_ _3309_/A _3430_/B VGND VGND VPWR VPWR _3531_/B sky130_fd_sc_hd__nand2_8
Xfanout468 fanout482/X VGND VGND VPWR VPWR fanout468/X sky130_fd_sc_hd__buf_12
X_7077_ _7077_/CLK _7077_/D fanout456/X VGND VGND VPWR VPWR _7077_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_59_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4289_ hold606/X _5187_/A1 _4291_/S VGND VGND VPWR VPWR _6719_/D sky130_fd_sc_hd__mux2_1
XFILLER_100_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout479 fanout481/X VGND VGND VPWR VPWR fanout479/X sky130_fd_sc_hd__buf_6
XFILLER_58_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6028_ _7101_/Q _6008_/X _6026_/X _6027_/X _5976_/X VGND VGND VPWR VPWR _6028_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_46_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3660_ _6935_/Q _5353_/A _5202_/A _6806_/Q VGND VGND VPWR VPWR _3660_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3591_ _6647_/Q _4206_/A _4194_/A _6637_/Q VGND VGND VPWR VPWR _3591_/X sky130_fd_sc_hd__a22o_1
XFILLER_127_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5330_ _5330_/A0 _5555_/A1 _5334_/S VGND VGND VPWR VPWR _6912_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5261_ _5261_/A0 _5585_/A1 _5262_/S VGND VGND VPWR VPWR _5261_/X sky130_fd_sc_hd__mux2_1
X_7000_ _7136_/CLK _7000_/D fanout476/X VGND VGND VPWR VPWR _7000_/Q sky130_fd_sc_hd__dfrtp_4
X_4212_ _4212_/A hold13/A VGND VGND VPWR VPWR _4217_/S sky130_fd_sc_hd__and2_4
XFILLER_87_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5192_ hold779/X _5552_/A1 _5199_/S VGND VGND VPWR VPWR _6795_/D sky130_fd_sc_hd__mux2_1
X_4143_ hold557/X _5187_/A1 _4145_/S VGND VGND VPWR VPWR _6591_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4074_ _4074_/A0 _5187_/A1 _4076_/S VGND VGND VPWR VPWR _4074_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4976_ _4976_/A _4976_/B VGND VGND VPWR VPWR _4985_/C sky130_fd_sc_hd__nor2_1
X_6715_ _6731_/CLK _6715_/D fanout465/X VGND VGND VPWR VPWR _6715_/Q sky130_fd_sc_hd__dfstp_2
X_3927_ _3927_/A1 _6437_/Q _3850_/S _3904_/A _3862_/A VGND VGND VPWR VPWR _3927_/Y
+ sky130_fd_sc_hd__o32ai_2
XFILLER_177_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6646_ _6750_/CLK _6646_/D fanout446/X VGND VGND VPWR VPWR _6646_/Q sky130_fd_sc_hd__dfstp_2
X_3858_ wire1/X _3858_/A1 _3858_/S VGND VGND VPWR VPWR _6449_/D sky130_fd_sc_hd__mux2_1
XFILLER_164_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6577_ _6588_/CLK _6577_/D fanout446/X VGND VGND VPWR VPWR _6577_/Q sky130_fd_sc_hd__dfrtp_4
X_3789_ _6917_/Q _5335_/A _4274_/A _6707_/Q _3788_/X VGND VGND VPWR VPWR _3792_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_3_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5528_ _5528_/A0 _5555_/A1 _5532_/S VGND VGND VPWR VPWR _5528_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5459_ _5459_/A0 _5585_/A1 _5460_/S VGND VGND VPWR VPWR _5459_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7129_ _7135_/CLK _7129_/D fanout473/X VGND VGND VPWR VPWR _7129_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_115_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_170 _6958_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4830_ _4417_/B _4633_/B _4384_/A _4658_/A VGND VGND VPWR VPWR _5127_/B sky130_fd_sc_hd__a211o_2
XFILLER_178_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_181 _7172_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_192 _5221_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4761_ _4625_/A _5033_/A _4976_/A VGND VGND VPWR VPWR _5108_/B sky130_fd_sc_hd__a21oi_2
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6500_ _7016_/CLK _6500_/D fanout475/X VGND VGND VPWR VPWR _7221_/A sky130_fd_sc_hd__dfrtp_1
X_3712_ _6723_/Q _4292_/A _4146_/A _6595_/Q VGND VGND VPWR VPWR _3712_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4692_ _4676_/Y _4688_/X _4691_/Y _5011_/B VGND VGND VPWR VPWR _4692_/X sky130_fd_sc_hd__a31o_1
XFILLER_174_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6431_ _6432_/A _6432_/B VGND VGND VPWR VPWR _6431_/X sky130_fd_sc_hd__and2_1
X_3643_ _6991_/Q _5416_/A _3330_/Y input45/X VGND VGND VPWR VPWR _3643_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6362_ _6684_/Q _6362_/A2 _6362_/B1 _4218_/Y _6361_/X VGND VGND VPWR VPWR _6362_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3574_ input46/X _4047_/C hold67/A _7120_/Q VGND VGND VPWR VPWR _3574_/X sky130_fd_sc_hd__a22o_2
XFILLER_115_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5313_ _5313_/A0 _5583_/A1 _5316_/S VGND VGND VPWR VPWR _5313_/X sky130_fd_sc_hd__mux2_1
X_6293_ _6617_/Q _5984_/X _5998_/X _6582_/Q VGND VGND VPWR VPWR _6293_/X sky130_fd_sc_hd__a22o_1
XFILLER_114_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5244_ _5244_/A0 _5559_/A1 _5244_/S VGND VGND VPWR VPWR _5244_/X sky130_fd_sc_hd__mux2_1
Xhold18 hold18/A VGND VGND VPWR VPWR hold18/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5175_ _5175_/A _5220_/C VGND VGND VPWR VPWR _5177_/S sky130_fd_sc_hd__and2_2
Xhold29 hold29/A VGND VGND VPWR VPWR hold29/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1903 _6583_/Q VGND VGND VPWR VPWR hold538/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1914 hold276/X VGND VGND VPWR VPWR _5464_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1925 _4213_/X VGND VGND VPWR VPWR _6649_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_4126_ _4126_/A0 _5195_/A1 _4127_/S VGND VGND VPWR VPWR _4126_/X sky130_fd_sc_hd__mux2_1
Xhold1936 hold613/X VGND VGND VPWR VPWR _4258_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1947 _4072_/X VGND VGND VPWR VPWR _6530_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1958 _6509_/Q VGND VGND VPWR VPWR _4014_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1969 _5527_/X VGND VGND VPWR VPWR _7087_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4057_ _4057_/A0 hold153/X hold14/X VGND VGND VPWR VPWR _4057_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4959_ _4959_/A _4959_/B VGND VGND VPWR VPWR _5042_/A sky130_fd_sc_hd__nor2_1
XFILLER_177_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6629_ _6788_/CLK _6629_/D _3959_/B VGND VGND VPWR VPWR _6629_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_137_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3290_ hold52/X _3290_/B VGND VGND VPWR VPWR _3550_/A sky130_fd_sc_hd__nand2_8
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6980_ _7084_/CLK _6980_/D fanout455/X VGND VGND VPWR VPWR _6980_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5931_ _6533_/Q _5653_/X _5662_/X _6587_/Q _5930_/X VGND VGND VPWR VPWR _5931_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5862_ _6574_/Q _5667_/X _5688_/X _6579_/Q _5861_/X VGND VGND VPWR VPWR _5869_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4813_ _5009_/A _4607_/B _4811_/B VGND VGND VPWR VPWR _5104_/C sky130_fd_sc_hd__o21ai_4
XFILLER_167_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5793_ _5782_/Y _5792_/Y _6841_/Q _5678_/Y VGND VGND VPWR VPWR _5793_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_166_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4744_ _4415_/B _4713_/Y _4743_/Y VGND VGND VPWR VPWR _4746_/A sky130_fd_sc_hd__o21ai_1
XFILLER_193_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4675_ _4675_/A _4683_/A VGND VGND VPWR VPWR _4725_/B sky130_fd_sc_hd__nor2_1
XFILLER_174_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3626_ _3971_/A _3431_/Y _4158_/A _6606_/Q _3625_/X VGND VGND VPWR VPWR _3627_/D
+ sky130_fd_sc_hd__a221o_1
X_6414_ _6414_/A _6433_/B VGND VGND VPWR VPWR _6414_/X sky130_fd_sc_hd__and2_1
XFILLER_147_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3557_ _3557_/A _3557_/B _3557_/C _3557_/D VGND VGND VPWR VPWR _3558_/C sky130_fd_sc_hd__and4_2
X_6345_ _6683_/D _3922_/B _6344_/Y _6345_/B2 VGND VGND VPWR VPWR _7186_/D sky130_fd_sc_hd__a22o_1
XFILLER_143_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6276_ _6729_/Q _5987_/X _6014_/X _6744_/Q _6275_/X VGND VGND VPWR VPWR _6279_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3488_ _3550_/A _3553_/B VGND VGND VPWR VPWR _4256_/A sky130_fd_sc_hd__nor2_8
Xhold2401 _6961_/Q VGND VGND VPWR VPWR hold748/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput108 wb_adr_i[18] VGND VGND VPWR VPWR _4343_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5227_ _5227_/A0 _5552_/A1 _5228_/S VGND VGND VPWR VPWR _5227_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2412 hold752/X VGND VGND VPWR VPWR _5349_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput119 wb_adr_i[28] VGND VGND VPWR VPWR input119/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2423 _6780_/Q VGND VGND VPWR VPWR _3424_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2434 hold86/A VGND VGND VPWR VPWR _3829_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1700 hold699/X VGND VGND VPWR VPWR _5203_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2445 _3867_/X VGND VGND VPWR VPWR _6447_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1711 hold446/X VGND VGND VPWR VPWR _5321_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2456 _6684_/Q VGND VGND VPWR VPWR _3917_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1722 hold130/X VGND VGND VPWR VPWR _5484_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5158_ _4583_/B _4691_/Y _5058_/C _5121_/X VGND VGND VPWR VPWR _5158_/X sky130_fd_sc_hd__o211a_1
Xhold2467 _6067_/X VGND VGND VPWR VPWR _7174_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1733 _6810_/Q VGND VGND VPWR VPWR hold139/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2478 _5838_/X VGND VGND VPWR VPWR _7166_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1744 _5294_/X VGND VGND VPWR VPWR _6880_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2489 _7165_/Q VGND VGND VPWR VPWR _5817_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1755 _7210_/A VGND VGND VPWR VPWR hold667/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1766 hold614/X VGND VGND VPWR VPWR _3979_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4109_ _3737_/Y hold870/A _4115_/S VGND VGND VPWR VPWR _6562_/D sky130_fd_sc_hd__mux2_1
Xhold1777 _4195_/X VGND VGND VPWR VPWR _6634_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5089_ _5089_/A _5089_/B _5089_/C VGND VGND VPWR VPWR _5136_/C sky130_fd_sc_hd__and3_1
Xhold1788 hold430/X VGND VGND VPWR VPWR _4228_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1799 _4208_/X VGND VGND VPWR VPWR _6645_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_112_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_70 _7097_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_81 input38/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_92 input72/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4460_ _4473_/A _4564_/C _4881_/A VGND VGND VPWR VPWR _4570_/A sky130_fd_sc_hd__nand3_4
Xhold307 hold307/A VGND VGND VPWR VPWR hold307/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold318 hold318/A VGND VGND VPWR VPWR hold318/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold329 hold329/A VGND VGND VPWR VPWR _6538_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3411_ _6801_/Q _3319_/Y _5479_/A _7051_/Q _3410_/X VGND VGND VPWR VPWR _3411_/X
+ sky130_fd_sc_hd__a221o_4
X_4391_ _5009_/A _4584_/A VGND VGND VPWR VPWR _4391_/Y sky130_fd_sc_hd__nand2_2
X_6130_ _6913_/Q _5991_/X _6005_/X _6945_/Q VGND VGND VPWR VPWR _6130_/X sky130_fd_sc_hd__a22o_1
X_3342_ _3343_/A hold54/X VGND VGND VPWR VPWR _5308_/A sky130_fd_sc_hd__nor2_8
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _7134_/Q _5977_/X _5995_/X _6918_/Q _6060_/X VGND VGND VPWR VPWR _6061_/X
+ sky130_fd_sc_hd__a221o_1
X_3273_ _3355_/A hold31/X VGND VGND VPWR VPWR _5226_/A sky130_fd_sc_hd__and2_2
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1007 _6922_/Q VGND VGND VPWR VPWR hold388/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_100_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5012_ _5011_/A _4590_/Y _4688_/A VGND VGND VPWR VPWR _5012_/X sky130_fd_sc_hd__a21o_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1018 _7043_/Q VGND VGND VPWR VPWR hold368/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1029 _3984_/X VGND VGND VPWR VPWR hold171/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_38_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6963_ _7123_/CLK _6963_/D fanout477/X VGND VGND VPWR VPWR _6963_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5914_ _6550_/Q _5673_/X _5909_/X _5911_/X _5913_/X VGND VGND VPWR VPWR _5914_/X
+ sky130_fd_sc_hd__a2111o_1
X_6894_ _7138_/CLK _6894_/D fanout477/X VGND VGND VPWR VPWR _6894_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_22_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5845_ _6980_/Q _5660_/X _5669_/X _7052_/Q VGND VGND VPWR VPWR _5845_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5776_ _7049_/Q _5669_/X _5687_/X _6921_/Q VGND VGND VPWR VPWR _5776_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4727_ _4727_/A _4993_/B VGND VGND VPWR VPWR _4727_/Y sky130_fd_sc_hd__nand2_2
XFILLER_135_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4658_ _4658_/A _4658_/B VGND VGND VPWR VPWR _4677_/B sky130_fd_sc_hd__nor2_2
XFILLER_163_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput90 spimemio_flash_io2_oeb VGND VGND VPWR VPWR input90/X sky130_fd_sc_hd__clkbuf_2
X_3609_ _7008_/Q _3347_/Y _4188_/A _6632_/Q VGND VGND VPWR VPWR _3609_/X sky130_fd_sc_hd__a22o_1
Xhold830 hold830/A VGND VGND VPWR VPWR hold830/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold841 hold841/A VGND VGND VPWR VPWR hold841/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4589_ _4637_/D _5011_/B VGND VGND VPWR VPWR _5009_/B sky130_fd_sc_hd__nor2_8
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold852 hold852/A VGND VGND VPWR VPWR hold852/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold863 hold863/A VGND VGND VPWR VPWR hold863/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6328_ _6701_/Q _5997_/X _6004_/X _6578_/Q VGND VGND VPWR VPWR _6328_/X sky130_fd_sc_hd__a22o_1
Xhold874 _6509_/Q VGND VGND VPWR VPWR hold874/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold885 _5251_/X VGND VGND VPWR VPWR _6842_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold896 hold50/X VGND VGND VPWR VPWR _7106_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_67_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6259_ _6738_/Q _6008_/X _6016_/X _6451_/Q VGND VGND VPWR VPWR _6259_/X sky130_fd_sc_hd__a22o_1
Xhold2220 hold465/X VGND VGND VPWR VPWR _4193_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_190_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2231 _7126_/Q VGND VGND VPWR VPWR hold722/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2242 _6960_/Q VGND VGND VPWR VPWR hold689/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2253 hold804/X VGND VGND VPWR VPWR _4189_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2264 _7071_/Q VGND VGND VPWR VPWR hold556/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1530 hold219/X VGND VGND VPWR VPWR _5204_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2275 _6990_/Q VGND VGND VPWR VPWR hold741/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2286 _6719_/Q VGND VGND VPWR VPWR hold606/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1541 _6559_/Q VGND VGND VPWR VPWR hold828/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1552 _6975_/Q VGND VGND VPWR VPWR hold345/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2297 _6992_/Q VGND VGND VPWR VPWR hold702/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1563 _6940_/Q VGND VGND VPWR VPWR hold483/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_123_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1574 hold824/X VGND VGND VPWR VPWR hold223/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1585 _6540_/Q VGND VGND VPWR VPWR hold846/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1596 hold822/X VGND VGND VPWR VPWR hold217/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3960_ _6457_/Q _3960_/B VGND VGND VPWR VPWR _3961_/A sky130_fd_sc_hd__nand2b_4
XFILLER_51_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3891_ _4649_/C _4649_/D VGND VGND VPWR VPWR _4720_/B sky130_fd_sc_hd__nor2_2
XFILLER_31_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5630_ _7154_/Q _7153_/Q VGND VGND VPWR VPWR _6017_/B sky130_fd_sc_hd__and2_4
XFILLER_188_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5561_ hold672/X _5561_/A1 _5568_/S VGND VGND VPWR VPWR _7117_/D sky130_fd_sc_hd__mux2_1
XFILLER_191_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4512_ _4719_/A _4638_/B VGND VGND VPWR VPWR _4729_/A sky130_fd_sc_hd__nand2_8
XFILLER_145_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5492_ _5492_/A0 _5582_/A1 _5496_/S VGND VGND VPWR VPWR _5492_/X sky130_fd_sc_hd__mux2_1
Xhold104 _6485_/Q VGND VGND VPWR VPWR hold104/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold115 hold115/A VGND VGND VPWR VPWR hold115/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7231_ _7231_/A VGND VGND VPWR VPWR _7231_/X sky130_fd_sc_hd__clkbuf_2
Xhold126 _5241_/X VGND VGND VPWR VPWR _6833_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4443_ _4486_/A _4598_/A _4598_/B VGND VGND VPWR VPWR _4569_/A sky130_fd_sc_hd__nand3_4
Xhold137 hold137/A VGND VGND VPWR VPWR hold137/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold148 _7196_/Q VGND VGND VPWR VPWR hold148/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold159 hold159/A VGND VGND VPWR VPWR hold159/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7162_ _3950_/A1 _7162_/D fanout468/X VGND VGND VPWR VPWR _7162_/Q sky130_fd_sc_hd__dfrtp_1
X_4374_ _4370_/Y _5011_/A _6686_/Q VGND VGND VPWR VPWR _4374_/Y sky130_fd_sc_hd__o21ai_2
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3325_ _3726_/A _3535_/A VGND VGND VPWR VPWR _5470_/A sky130_fd_sc_hd__nor2_8
X_6113_ _6113_/A _6113_/B _6113_/C _6113_/D VGND VGND VPWR VPWR _6114_/D sky130_fd_sc_hd__nor4_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7093_ _7093_/CLK _7093_/D fanout460/X VGND VGND VPWR VPWR _7093_/Q sky130_fd_sc_hd__dfstp_2
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ _3832_/A _6657_/Q hold86/X VGND VGND VPWR VPWR _3256_/X sky130_fd_sc_hd__a21o_1
X_6044_ _6910_/Q _5991_/X _5993_/X _7006_/Q _6043_/X VGND VGND VPWR VPWR _6044_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3187_ _6766_/Q VGND VGND VPWR VPWR _3187_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6946_ _7020_/CLK hold81/X fanout470/X VGND VGND VPWR VPWR _6946_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6877_ _6903_/CLK _6877_/D fanout460/X VGND VGND VPWR VPWR _6877_/Q sky130_fd_sc_hd__dfstp_2
X_5828_ _6995_/Q _5929_/B _5681_/X _7091_/Q _5827_/X VGND VGND VPWR VPWR _5835_/A
+ sky130_fd_sc_hd__a221o_1
X_5759_ _6888_/Q _5688_/X _5756_/X _5758_/X VGND VGND VPWR VPWR _5760_/C sky130_fd_sc_hd__a211o_1
XFILLER_154_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold660 hold660/A VGND VGND VPWR VPWR hold660/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold671 _4243_/X VGND VGND VPWR VPWR _6669_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold682 hold682/A VGND VGND VPWR VPWR hold682/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold693 hold693/A VGND VGND VPWR VPWR hold693/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2050 _7136_/Q VGND VGND VPWR VPWR hold758/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2061 _6736_/Q VGND VGND VPWR VPWR hold458/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2072 hold674/X VGND VGND VPWR VPWR _4245_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_58_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2083 _7085_/Q VGND VGND VPWR VPWR hold665/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2094 _7109_/Q VGND VGND VPWR VPWR hold809/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1360 _6439_/Q VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_18_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1371 _6974_/Q VGND VGND VPWR VPWR hold545/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1382 _4044_/X VGND VGND VPWR VPWR _6507_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1393 _6725_/Q VGND VGND VPWR VPWR hold321/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput209 _3234_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[6] sky130_fd_sc_hd__buf_12
XFILLER_181_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4090_ _3422_/Y hold822/A _4091_/S VGND VGND VPWR VPWR _6546_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6800_ _6822_/CLK _6800_/D fanout451/X VGND VGND VPWR VPWR _6800_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_91_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4992_ _4701_/B _4995_/B _4991_/X _5083_/B _5021_/B VGND VGND VPWR VPWR _5000_/A
+ sky130_fd_sc_hd__o2111a_1
XFILLER_90_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6731_ _6731_/CLK _6731_/D fanout465/X VGND VGND VPWR VPWR _6731_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_189_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3943_ _6661_/Q _6781_/Q _6432_/B VGND VGND VPWR VPWR _3943_/X sky130_fd_sc_hd__mux2_1
X_6662_ _7116_/CLK _6662_/D fanout454/X VGND VGND VPWR VPWR _7207_/A sky130_fd_sc_hd__dfrtp_1
X_3874_ hold93/A _3874_/A1 _3878_/S VGND VGND VPWR VPWR _6442_/D sky130_fd_sc_hd__mux2_1
XFILLER_149_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5613_ _7148_/Q _5613_/B VGND VGND VPWR VPWR _5613_/Y sky130_fd_sc_hd__nor2_1
X_6593_ _6747_/CLK _6593_/D _3959_/B VGND VGND VPWR VPWR _6593_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_191_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5544_ hold284/X _5544_/A1 _5550_/S VGND VGND VPWR VPWR _7102_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5475_ _5475_/A0 _5583_/A1 _5478_/S VGND VGND VPWR VPWR _7041_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7214_ _7214_/A VGND VGND VPWR VPWR _7214_/X sky130_fd_sc_hd__clkbuf_2
X_4426_ _4513_/B _5150_/A VGND VGND VPWR VPWR _4426_/Y sky130_fd_sc_hd__nand2_1
XFILLER_160_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout403 _5544_/A1 VGND VGND VPWR VPWR _5499_/A1 sky130_fd_sc_hd__buf_6
XFILLER_98_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout414 hold13/A VGND VGND VPWR VPWR _5569_/B sky130_fd_sc_hd__buf_12
X_7145_ _7203_/CLK _7145_/D _6414_/A VGND VGND VPWR VPWR _7145_/Q sky130_fd_sc_hd__dfrtp_2
X_4357_ _4649_/B _4357_/B VGND VGND VPWR VPWR _4513_/A sky130_fd_sc_hd__xor2_4
XFILLER_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout436 wire438/X VGND VGND VPWR VPWR _6423_/B sky130_fd_sc_hd__buf_8
Xfanout447 fanout449/X VGND VGND VPWR VPWR fanout447/X sky130_fd_sc_hd__buf_6
X_3308_ _3305_/A hold30/X VGND VGND VPWR VPWR _3308_/X sky130_fd_sc_hd__and2b_4
Xfanout458 fanout460/X VGND VGND VPWR VPWR fanout458/X sky130_fd_sc_hd__buf_12
X_4288_ _4288_/A0 _5186_/A1 _4291_/S VGND VGND VPWR VPWR _6718_/D sky130_fd_sc_hd__mux2_1
X_7076_ _7124_/CLK _7076_/D fanout459/X VGND VGND VPWR VPWR _7076_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout469 fanout470/X VGND VGND VPWR VPWR fanout469/X sky130_fd_sc_hd__buf_12
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6027_ _6901_/Q _5985_/X _6016_/X _7037_/Q VGND VGND VPWR VPWR _6027_/X sky130_fd_sc_hd__a22o_1
X_3239_ _6840_/Q VGND VGND VPWR VPWR _3239_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_27_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6929_ _7135_/CLK _6929_/D fanout473/X VGND VGND VPWR VPWR _6929_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_31_csclk _6850_/CLK VGND VGND VPWR VPWR _6522_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_168_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_46_csclk _7093_/CLK VGND VGND VPWR VPWR _7047_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_109_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold490 hold490/A VGND VGND VPWR VPWR hold490/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1190 _7026_/Q VGND VGND VPWR VPWR hold497/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3590_ _7096_/Q _5533_/A _3391_/Y _6811_/Q _3589_/X VGND VGND VPWR VPWR _3595_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5260_ hold982/X hold20/X _5262_/S VGND VGND VPWR VPWR _6850_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4211_ _4211_/A0 _4339_/A1 _4211_/S VGND VGND VPWR VPWR _4211_/X sky130_fd_sc_hd__mux2_1
X_5191_ _5207_/A _5220_/B _5220_/C VGND VGND VPWR VPWR _5198_/S sky130_fd_sc_hd__and3_4
X_4142_ _4142_/A0 _5186_/A1 _4145_/S VGND VGND VPWR VPWR _6590_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4073_ _4073_/A0 _5186_/A1 _4076_/S VGND VGND VPWR VPWR _4073_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_810 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4975_ _4564_/B _4934_/B _4881_/B _4572_/Y _4886_/A VGND VGND VPWR VPWR _4976_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_189_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6714_ _6731_/CLK _6714_/D fanout465/X VGND VGND VPWR VPWR _6714_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3926_ _6437_/Q _6654_/Q _3904_/A _3926_/B1 VGND VGND VPWR VPWR _3926_/X sky130_fd_sc_hd__a31o_1
XFILLER_149_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6645_ _6759_/CLK _6645_/D _6426_/A VGND VGND VPWR VPWR _6645_/Q sky130_fd_sc_hd__dfrtp_4
X_3857_ _6654_/Q _3857_/B VGND VGND VPWR VPWR _3858_/S sky130_fd_sc_hd__nand2_1
XFILLER_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6576_ _6747_/CLK _6576_/D fanout443/X VGND VGND VPWR VPWR _6576_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_166_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3788_ _7037_/Q _5470_/A _4065_/A _6525_/Q VGND VGND VPWR VPWR _3788_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5527_ _5527_/A0 _5581_/A1 _5532_/S VGND VGND VPWR VPWR _5527_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5458_ _5458_/A0 _5503_/A1 _5460_/S VGND VGND VPWR VPWR _5458_/X sky130_fd_sc_hd__mux2_1
X_4409_ _4575_/C _4637_/D VGND VGND VPWR VPWR _4638_/B sky130_fd_sc_hd__nor2_8
X_5389_ _5389_/A _5551_/B VGND VGND VPWR VPWR _5397_/S sky130_fd_sc_hd__and2_4
XFILLER_120_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7128_ _7137_/CLK _7128_/D fanout475/X VGND VGND VPWR VPWR _7128_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7059_ _7139_/CLK _7059_/D fanout478/X VGND VGND VPWR VPWR _7059_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_86_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_160 _5684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_171 _6984_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_182 _7159_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_193 fanout472/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4760_ _4759_/X _4558_/X _5139_/A hold29/A VGND VGND VPWR VPWR _6762_/D sky130_fd_sc_hd__o2bb2a_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3711_ _6846_/Q hold40/A _5461_/A _7030_/Q _3710_/X VGND VGND VPWR VPWR _3716_/B
+ sky130_fd_sc_hd__a221o_1
X_4691_ _4713_/A _4691_/B VGND VGND VPWR VPWR _4691_/Y sky130_fd_sc_hd__nand2_8
XFILLER_174_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6430_ _6432_/A _6433_/B VGND VGND VPWR VPWR _6430_/X sky130_fd_sc_hd__and2_1
X_3642_ _6724_/Q _4292_/A _3539_/Y _6532_/Q _3641_/X VGND VGND VPWR VPWR _3645_/C
+ sky130_fd_sc_hd__a221o_1
X_6361_ _6686_/Q _6361_/A2 _6361_/B1 _6685_/Q VGND VGND VPWR VPWR _6361_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3573_ _6920_/Q _5335_/A _4274_/A _6710_/Q _3572_/X VGND VGND VPWR VPWR _3573_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_114_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5312_ _5312_/A0 _5555_/A1 _5316_/S VGND VGND VPWR VPWR _5312_/X sky130_fd_sc_hd__mux2_1
X_6292_ _6316_/A1 _6342_/S _6290_/X _6291_/X VGND VGND VPWR VPWR _7183_/D sky130_fd_sc_hd__o22a_1
X_5243_ hold928/X hold78/X _5244_/S VGND VGND VPWR VPWR _5243_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold19 hold19/A VGND VGND VPWR VPWR hold19/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5174_ _5174_/A0 _5196_/A1 _5174_/S VGND VGND VPWR VPWR _5174_/X sky130_fd_sc_hd__mux2_1
Xhold1904 hold538/X VGND VGND VPWR VPWR _4133_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1915 _6622_/Q VGND VGND VPWR VPWR hold654/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4125_ _4125_/A0 _5187_/A1 _4127_/S VGND VGND VPWR VPWR _4125_/X sky130_fd_sc_hd__mux2_1
Xhold1926 _6753_/Q VGND VGND VPWR VPWR hold600/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_110_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1937 _4258_/X VGND VGND VPWR VPWR _6693_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1948 _6839_/Q VGND VGND VPWR VPWR hold311/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1959 _4014_/X VGND VGND VPWR VPWR _4015_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4056_ _6432_/B hold13/A _4056_/C VGND VGND VPWR VPWR hold14/A sky130_fd_sc_hd__and3b_1
XFILLER_37_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_840 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4958_ _5044_/A _5044_/B _5032_/B _4958_/D VGND VGND VPWR VPWR _4961_/B sky130_fd_sc_hd__and4_1
XFILLER_61_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3909_ _6019_/A _6015_/B _6008_/A VGND VGND VPWR VPWR _3909_/X sky130_fd_sc_hd__and3_1
X_4889_ _5138_/A _4889_/B VGND VGND VPWR VPWR _5130_/A sky130_fd_sc_hd__and2_1
XFILLER_177_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6628_ _6759_/CLK _6628_/D fanout449/X VGND VGND VPWR VPWR _6628_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6559_ _6568_/CLK _6559_/D VGND VGND VPWR VPWR _6559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire431 _4637_/Y VGND VGND VPWR VPWR _4732_/B sky130_fd_sc_hd__buf_2
XFILLER_11_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5930_ _6577_/Q _5667_/X _5682_/X _6453_/Q VGND VGND VPWR VPWR _5930_/X sky130_fd_sc_hd__a22o_1
XFILLER_19_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5861_ _6687_/Q _5659_/X _5684_/X _6604_/Q VGND VGND VPWR VPWR _5861_/X sky130_fd_sc_hd__a22o_1
XFILLER_33_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4812_ _4812_/A _4826_/A VGND VGND VPWR VPWR _4812_/Y sky130_fd_sc_hd__nor2_2
XFILLER_22_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5792_ _5792_/A _5792_/B _5792_/C _5792_/D VGND VGND VPWR VPWR _5792_/Y sky130_fd_sc_hd__nor4_1
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4743_ _4719_/A _4719_/B _4741_/Y _4742_/Y VGND VGND VPWR VPWR _4743_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_147_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4674_ _4682_/A _4691_/B VGND VGND VPWR VPWR _4674_/Y sky130_fd_sc_hd__nand2_4
XFILLER_190_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6413_ _6414_/A _6423_/B VGND VGND VPWR VPWR _6413_/X sky130_fd_sc_hd__and2_1
X_3625_ input26/X _3307_/Y _4286_/A _6719_/Q VGND VGND VPWR VPWR _3625_/X sky130_fd_sc_hd__a22o_2
XFILLER_134_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6344_ _6344_/A VGND VGND VPWR VPWR _6344_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3556_ _3556_/A _3556_/B _3556_/C _3556_/D VGND VGND VPWR VPWR _3557_/D sky130_fd_sc_hd__nor4_2
XFILLER_143_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6275_ _6714_/Q _5973_/X _5988_/X _6571_/Q VGND VGND VPWR VPWR _6275_/X sky130_fd_sc_hd__a22o_1
X_3487_ _3487_/A _3648_/A VGND VGND VPWR VPWR _4274_/A sky130_fd_sc_hd__nor2_8
XFILLER_102_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2402 hold748/X VGND VGND VPWR VPWR _5385_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput109 wb_adr_i[19] VGND VGND VPWR VPWR _4343_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_5226_ _5226_/A _5226_/B _5551_/B VGND VGND VPWR VPWR _5228_/S sky130_fd_sc_hd__and3_1
Xhold2413 _5349_/X VGND VGND VPWR VPWR _6929_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2424 _6777_/Q VGND VGND VPWR VPWR _3618_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2435 _7181_/Q VGND VGND VPWR VPWR _6242_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1701 _7007_/Q VGND VGND VPWR VPWR hold181/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2446 _6449_/Q VGND VGND VPWR VPWR _3858_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2457 hold73/A VGND VGND VPWR VPWR _6369_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1712 _6983_/Q VGND VGND VPWR VPWR hold344/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1723 _6737_/Q VGND VGND VPWR VPWR hold698/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5157_ _4570_/C _4523_/Y _4870_/A _4925_/A _5113_/B VGND VGND VPWR VPWR _5157_/X
+ sky130_fd_sc_hd__o2111a_1
Xhold2468 _7173_/Q VGND VGND VPWR VPWR _6042_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1734 hold139/X VGND VGND VPWR VPWR _5212_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2479 _7184_/Q VGND VGND VPWR VPWR _6341_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_186_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1745 _6694_/Q VGND VGND VPWR VPWR hold291/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1756 hold667/X VGND VGND VPWR VPWR _4236_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4108_ _3803_/Y hold868/A _4115_/S VGND VGND VPWR VPWR _6561_/D sky130_fd_sc_hd__mux2_1
Xhold1767 _6833_/Q VGND VGND VPWR VPWR hold125/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1778 _6646_/Q VGND VGND VPWR VPWR hold310/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5088_ _4477_/Y _4938_/X _5027_/X _5087_/X _4791_/B VGND VGND VPWR VPWR _5088_/X
+ sky130_fd_sc_hd__o2111a_1
Xhold1789 _6636_/Q VGND VGND VPWR VPWR hold298/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4039_ _4061_/A0 _5556_/A1 _4056_/C VGND VGND VPWR VPWR _4039_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_60 _6744_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_71 _7128_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_82 input38/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_93 _3966_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold308 hold308/A VGND VGND VPWR VPWR hold308/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold319 hold319/A VGND VGND VPWR VPWR hold319/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3410_ input32/X _3307_/Y _5461_/A _7035_/Q VGND VGND VPWR VPWR _3410_/X sky130_fd_sc_hd__a22o_1
XFILLER_171_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4390_ _4717_/A _4712_/A VGND VGND VPWR VPWR _4658_/A sky130_fd_sc_hd__nand2_8
XFILLER_131_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3341_ _3487_/A hold32/X VGND VGND VPWR VPWR _5362_/A sky130_fd_sc_hd__nor2_8
XFILLER_124_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6060_ _7094_/Q _5984_/X _5986_/X _7030_/Q VGND VGND VPWR VPWR _6060_/X sky130_fd_sc_hd__a22o_1
XFILLER_140_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ _3272_/A _3305_/B VGND VGND VPWR VPWR hold31/A sky130_fd_sc_hd__nor2_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _5011_/A _5011_/B VGND VGND VPWR VPWR _5011_/X sky130_fd_sc_hd__and2_1
Xhold1008 hold388/X VGND VGND VPWR VPWR _5341_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1019 hold368/X VGND VGND VPWR VPWR _5477_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_26_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6962_ _7020_/CLK _6962_/D fanout458/X VGND VGND VPWR VPWR _6962_/Q sky130_fd_sc_hd__dfrtp_4
X_5913_ _6611_/Q _5660_/X _5669_/X _6651_/Q _5912_/X VGND VGND VPWR VPWR _5913_/X
+ sky130_fd_sc_hd__a221o_1
X_6893_ _7077_/CLK _6893_/D fanout456/X VGND VGND VPWR VPWR _6893_/Q sky130_fd_sc_hd__dfstp_2
X_5844_ _7036_/Q _5655_/X _5656_/X _6988_/Q _5839_/Y VGND VGND VPWR VPWR _5844_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5775_ _6913_/Q _5670_/X _5671_/X _7065_/Q _5774_/X VGND VGND VPWR VPWR _5782_/A
+ sky130_fd_sc_hd__a221o_1
X_4726_ _4808_/A _4732_/B _4726_/C VGND VGND VPWR VPWR _5083_/A sky130_fd_sc_hd__nand3_2
XFILLER_108_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4657_ _4500_/Y _4640_/Y _5047_/A VGND VGND VPWR VPWR _5124_/B sky130_fd_sc_hd__o21a_1
Xinput80 spi_sck VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__clkbuf_4
X_3608_ _6992_/Q _5416_/A _3310_/Y input14/X _3607_/X VGND VGND VPWR VPWR _3614_/B
+ sky130_fd_sc_hd__a221o_2
Xhold820 hold820/A VGND VGND VPWR VPWR hold820/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput91 spimemio_flash_io3_do VGND VGND VPWR VPWR input91/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold831 hold831/A VGND VGND VPWR VPWR hold831/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4588_ _4596_/A _4972_/A VGND VGND VPWR VPWR _4986_/C sky130_fd_sc_hd__nand2_4
Xhold842 hold842/A VGND VGND VPWR VPWR hold842/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold853 hold853/A VGND VGND VPWR VPWR hold853/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6327_ _6327_/A _6327_/B _6327_/C VGND VGND VPWR VPWR _6339_/C sky130_fd_sc_hd__nor3_1
Xhold864 hold864/A VGND VGND VPWR VPWR hold864/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3539_ _3549_/B _3648_/B VGND VGND VPWR VPWR _3539_/Y sky130_fd_sc_hd__nor2_4
Xmgmt_gpio_15_buff_inst _3949_/X VGND VGND VPWR VPWR mgmt_gpio_out[15] sky130_fd_sc_hd__clkbuf_8
Xhold875 _7200_/Q VGND VGND VPWR VPWR hold875/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold886 _7227_/A VGND VGND VPWR VPWR hold886/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_103_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold897 _7201_/Q VGND VGND VPWR VPWR hold897/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_67_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6258_ _6713_/Q _5973_/X _5988_/X _6570_/Q _6257_/X VGND VGND VPWR VPWR _6258_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2210 _7118_/Q VGND VGND VPWR VPWR hold714/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2221 _7215_/A VGND VGND VPWR VPWR hold814/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2232 hold722/X VGND VGND VPWR VPWR _5571_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5209_ hold649/X _5221_/A1 _5209_/S VGND VGND VPWR VPWR _5210_/B sky130_fd_sc_hd__mux2_1
XFILLER_76_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2243 hold689/X VGND VGND VPWR VPWR _5384_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2254 _6723_/Q VGND VGND VPWR VPWR hold747/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6189_ _6170_/X _6189_/B _6189_/C VGND VGND VPWR VPWR _6189_/Y sky130_fd_sc_hd__nand3b_2
Xhold1520 _5307_/X VGND VGND VPWR VPWR _6892_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2265 hold556/X VGND VGND VPWR VPWR _5509_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1531 _5204_/X VGND VGND VPWR VPWR _6805_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2276 hold741/X VGND VGND VPWR VPWR _5418_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1542 hold828/X VGND VGND VPWR VPWR hold235/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2287 _6952_/Q VGND VGND VPWR VPWR hold703/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1553 hold345/X VGND VGND VPWR VPWR _5401_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2298 hold702/X VGND VGND VPWR VPWR _5420_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1564 hold483/X VGND VGND VPWR VPWR _5361_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1575 _6863_/Q VGND VGND VPWR VPWR hold138/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1586 hold846/X VGND VGND VPWR VPWR hold274/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1597 _6651_/Q VGND VGND VPWR VPWR hold257/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3890_ _4720_/C _4649_/B VGND VGND VPWR VPWR _3890_/Y sky130_fd_sc_hd__nand2_2
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5560_ hold67/X _5569_/B VGND VGND VPWR VPWR _5568_/S sky130_fd_sc_hd__and2_4
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4511_ _4719_/A _4638_/B VGND VGND VPWR VPWR _4955_/D sky130_fd_sc_hd__and2_4
XFILLER_156_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5491_ _5491_/A0 _5518_/A1 _5496_/S VGND VGND VPWR VPWR _5491_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7230_ _7230_/A VGND VGND VPWR VPWR _7230_/X sky130_fd_sc_hd__clkbuf_2
Xhold105 _6801_/Q VGND VGND VPWR VPWR hold105/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold116 hold116/A VGND VGND VPWR VPWR hold116/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4442_ _4486_/A _4485_/B _4598_/B VGND VGND VPWR VPWR _4971_/A sky130_fd_sc_hd__and3_4
Xhold127 hold127/A VGND VGND VPWR VPWR hold127/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold138 hold138/A VGND VGND VPWR VPWR hold138/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold149 hold149/A VGND VGND VPWR VPWR hold149/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7161_ _3950_/A1 _7161_/D fanout468/X VGND VGND VPWR VPWR _7161_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_172_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4373_ _4576_/A _4719_/A VGND VGND VPWR VPWR _5011_/A sky130_fd_sc_hd__nand2_8
XFILLER_171_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6112_ _7136_/Q _5977_/X _5984_/X _7096_/Q _6111_/X VGND VGND VPWR VPWR _6113_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3324_ _3764_/A _3535_/A VGND VGND VPWR VPWR _5515_/A sky130_fd_sc_hd__nor2_8
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7092_ _7131_/CLK hold36/X fanout470/X VGND VGND VPWR VPWR _7092_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_113_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6043_ _7086_/Q _5638_/X _6012_/X _6998_/Q VGND VGND VPWR VPWR _6043_/X sky130_fd_sc_hd__a22o_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _3996_/S _3255_/B VGND VGND VPWR VPWR _3255_/Y sky130_fd_sc_hd__nand2b_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ _6657_/Q VGND VGND VPWR VPWR _3862_/A sky130_fd_sc_hd__inv_2
XFILLER_66_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6945_ _6945_/CLK _6945_/D _6399_/A VGND VGND VPWR VPWR _6945_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6876_ _7130_/CLK _6876_/D fanout458/X VGND VGND VPWR VPWR _6876_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5827_ _6859_/Q _5651_/X _5688_/X _6891_/Q VGND VGND VPWR VPWR _5827_/X sky130_fd_sc_hd__a22o_1
X_5758_ _7032_/Q _5655_/X _5667_/X _6880_/Q _5757_/X VGND VGND VPWR VPWR _5758_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_136_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4709_ _4495_/B _4638_/B _4507_/Y _4704_/X _4708_/X VGND VGND VPWR VPWR _4709_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_185_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5689_ _5689_/A _5689_/B _5689_/C VGND VGND VPWR VPWR _5689_/X sky130_fd_sc_hd__and3_4
XFILLER_147_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold650 hold650/A VGND VGND VPWR VPWR hold650/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold661 hold661/A VGND VGND VPWR VPWR hold661/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold672 hold672/A VGND VGND VPWR VPWR hold672/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold683 hold683/A VGND VGND VPWR VPWR hold683/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold694 hold694/A VGND VGND VPWR VPWR hold694/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2040 _6531_/Q VGND VGND VPWR VPWR hold727/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2051 hold758/X VGND VGND VPWR VPWR _5582_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2062 hold458/X VGND VGND VPWR VPWR _4309_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2073 _6941_/Q VGND VGND VPWR VPWR hold593/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_182_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2084 _5525_/X VGND VGND VPWR VPWR _7085_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2095 _6474_/Q VGND VGND VPWR VPWR hold631/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1350 _6996_/Q VGND VGND VPWR VPWR hold350/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_18_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1361 hold1/X VGND VGND VPWR VPWR _3982_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1372 _6750_/Q VGND VGND VPWR VPWR hold312/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1383 _6903_/Q VGND VGND VPWR VPWR _5320_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1394 hold321/X VGND VGND VPWR VPWR _4296_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4991_ _4668_/Y _4688_/A _4995_/B VGND VGND VPWR VPWR _4991_/X sky130_fd_sc_hd__a21o_1
X_6730_ _6731_/CLK _6730_/D fanout465/X VGND VGND VPWR VPWR _6730_/Q sky130_fd_sc_hd__dfrtp_4
X_3942_ _6666_/Q input77/X _3970_/B VGND VGND VPWR VPWR _3942_/X sky130_fd_sc_hd__mux2_8
XFILLER_90_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6661_ _7013_/CLK _6661_/D fanout452/X VGND VGND VPWR VPWR _6661_/Q sky130_fd_sc_hd__dfrtp_4
X_3873_ _3874_/A1 _3873_/A1 _3878_/S VGND VGND VPWR VPWR _6443_/D sky130_fd_sc_hd__mux2_1
X_5612_ _5647_/B _5679_/B _5684_/B _5612_/B1 _5605_/Y VGND VGND VPWR VPWR _7147_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_177_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6592_ _6742_/CLK _6592_/D fanout440/X VGND VGND VPWR VPWR _6592_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_118_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5543_ hold817/X _5552_/A1 _5550_/S VGND VGND VPWR VPWR _7101_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5474_ _5474_/A0 _5582_/A1 _5478_/S VGND VGND VPWR VPWR _7040_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7213_ _7213_/A VGND VGND VPWR VPWR _7213_/X sky130_fd_sc_hd__clkbuf_2
X_4425_ _4513_/B _5150_/A VGND VGND VPWR VPWR _4552_/B sky130_fd_sc_hd__and2_1
XFILLER_144_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7144_ _7183_/CLK _7144_/D _6414_/A VGND VGND VPWR VPWR _7144_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout404 hold1127/X VGND VGND VPWR VPWR _5544_/A1 sky130_fd_sc_hd__buf_6
X_4356_ _4492_/B _4356_/B VGND VGND VPWR VPWR _4357_/B sky130_fd_sc_hd__nand2_2
XFILLER_98_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout415 _5407_/B VGND VGND VPWR VPWR hold13/A sky130_fd_sc_hd__buf_12
XFILLER_86_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout437 _3881_/Y VGND VGND VPWR VPWR _6432_/B sky130_fd_sc_hd__buf_12
XFILLER_59_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3307_ _3764_/B _3553_/B VGND VGND VPWR VPWR _3307_/Y sky130_fd_sc_hd__nor2_8
Xfanout448 fanout449/X VGND VGND VPWR VPWR _6426_/A sky130_fd_sc_hd__buf_8
XFILLER_101_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout459 fanout460/X VGND VGND VPWR VPWR fanout459/X sky130_fd_sc_hd__buf_12
X_7075_ _7123_/CLK _7075_/D fanout477/X VGND VGND VPWR VPWR _7075_/Q sky130_fd_sc_hd__dfrtp_4
X_4287_ _4287_/A0 _5208_/A1 _4291_/S VGND VGND VPWR VPWR _6717_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6026_ _6997_/Q _6012_/X _6019_/X _6981_/Q _6025_/X VGND VGND VPWR VPWR _6026_/X
+ sky130_fd_sc_hd__a221o_1
X_3238_ _6848_/Q VGND VGND VPWR VPWR _3238_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6928_ _7139_/CLK _6928_/D fanout478/X VGND VGND VPWR VPWR _6928_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_154_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6859_ _7140_/CLK _6859_/D fanout469/X VGND VGND VPWR VPWR _6859_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_168_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold480 hold480/A VGND VGND VPWR VPWR hold480/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold491 hold491/A VGND VGND VPWR VPWR hold491/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1180 hold94/X VGND VGND VPWR VPWR hold1180/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1191 hold497/X VGND VGND VPWR VPWR _5458_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_61_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4210_ _4210_/A0 _5303_/A1 _4211_/S VGND VGND VPWR VPWR _4210_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5190_ _5190_/A0 _5503_/A1 _5190_/S VGND VGND VPWR VPWR _5190_/X sky130_fd_sc_hd__mux2_1
X_4141_ _4141_/A0 _5208_/A1 _4145_/S VGND VGND VPWR VPWR _6589_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4072_ _4072_/A0 _5221_/A1 _4076_/S VGND VGND VPWR VPWR _4072_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4974_ _5114_/A _4986_/C _5114_/B VGND VGND VPWR VPWR _5061_/B sky130_fd_sc_hd__and3_1
X_6713_ _6731_/CLK _6713_/D _6409_/A VGND VGND VPWR VPWR _6713_/Q sky130_fd_sc_hd__dfrtp_4
X_3925_ _6341_/S _3912_/B _5647_/B VGND VGND VPWR VPWR _6490_/D sky130_fd_sc_hd__o21ai_1
XFILLER_32_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6644_ _6750_/CLK _6644_/D fanout446/X VGND VGND VPWR VPWR _6644_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3856_ _3807_/B _3904_/A _3855_/X _3856_/B2 _3903_/A VGND VGND VPWR VPWR _6455_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_149_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6575_ _6742_/CLK _6575_/D fanout439/X VGND VGND VPWR VPWR _6575_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_166_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3787_ _6965_/Q _5389_/A _5308_/A _6893_/Q _3786_/X VGND VGND VPWR VPWR _3792_/B
+ sky130_fd_sc_hd__a221o_1
X_5526_ hold769/X _5580_/A1 _5532_/S VGND VGND VPWR VPWR _5526_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5457_ _5457_/A0 _5583_/A1 _5460_/S VGND VGND VPWR VPWR _5457_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4408_ _4391_/Y _4969_/A _4407_/Y VGND VGND VPWR VPWR _4529_/B sky130_fd_sc_hd__a21o_1
XFILLER_182_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5388_ hold43/X hold6/X _5388_/S VGND VGND VPWR VPWR _5388_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7127_ _7127_/CLK _7127_/D fanout477/X VGND VGND VPWR VPWR _7127_/Q sky130_fd_sc_hd__dfrtp_4
X_4339_ _4339_/A0 _4339_/A1 _4339_/S VGND VGND VPWR VPWR _6761_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7058_ _7116_/CLK _7058_/D fanout455/X VGND VGND VPWR VPWR _7058_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_86_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6009_ _5637_/A _6017_/A _6019_/C _5980_/X _5995_/X VGND VGND VPWR VPWR _6010_/C
+ sky130_fd_sc_hd__a311o_1
XFILLER_55_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_150 _3703_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_161 _5685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_172 _7000_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_183 input1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_194 hold2/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3710_ _6472_/Q _3339_/Y _3977_/A _6451_/Q VGND VGND VPWR VPWR _3710_/X sky130_fd_sc_hd__a22o_2
XFILLER_81_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4690_ _4638_/Y _4668_/Y _4688_/X _4990_/B _4689_/Y VGND VGND VPWR VPWR _4703_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_147_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3641_ input54/X _4241_/A _3509_/Y _6729_/Q VGND VGND VPWR VPWR _3641_/X sky130_fd_sc_hd__a22o_2
XFILLER_146_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6360_ _6684_/Q _6358_/Y _6359_/X _6355_/Y VGND VGND VPWR VPWR _6384_/S sky130_fd_sc_hd__a211o_4
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3572_ _6912_/Q _5326_/A _3569_/X _3571_/X VGND VGND VPWR VPWR _3572_/X sky130_fd_sc_hd__a211o_1
XFILLER_155_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5311_ _5311_/A0 _5572_/A1 _5316_/S VGND VGND VPWR VPWR _5311_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6291_ _6490_/Q _6291_/A2 _5649_/Y VGND VGND VPWR VPWR _6291_/X sky130_fd_sc_hd__a21o_1
XFILLER_142_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5242_ _5242_/A0 _5503_/A1 _5244_/S VGND VGND VPWR VPWR _5242_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_30_csclk _6850_/CLK VGND VGND VPWR VPWR _6523_/CLK sky130_fd_sc_hd__clkbuf_16
X_5173_ _5173_/A0 _5195_/A1 _5174_/S VGND VGND VPWR VPWR _5173_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1905 _6862_/Q VGND VGND VPWR VPWR hold539/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4124_ _4124_/A0 _5186_/A1 _4127_/S VGND VGND VPWR VPWR _4124_/X sky130_fd_sc_hd__mux2_1
Xhold1916 hold654/X VGND VGND VPWR VPWR _4180_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1927 hold600/X VGND VGND VPWR VPWR _4330_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1938 _6935_/Q VGND VGND VPWR VPWR hold308/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1949 hold311/X VGND VGND VPWR VPWR _5248_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput1 debug_mode VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__clkbuf_4
XFILLER_68_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4055_ hold974/X hold6/X _4055_/S VGND VGND VPWR VPWR _4055_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_45_csclk _7093_/CLK VGND VGND VPWR VPWR _7018_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_37_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4957_ _5067_/A _5023_/A _4957_/C _5034_/C VGND VGND VPWR VPWR _4958_/D sky130_fd_sc_hd__and4_1
XFILLER_178_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3908_ _5637_/A _7156_/Q VGND VGND VPWR VPWR _6008_/A sky130_fd_sc_hd__and2_2
XFILLER_193_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4888_ _4575_/C _4463_/B _4568_/Y _4878_/Y _4491_/Y VGND VGND VPWR VPWR _4892_/C
+ sky130_fd_sc_hd__o32a_1
X_6627_ _6761_/CLK _6627_/D _6426_/A VGND VGND VPWR VPWR _6627_/Q sky130_fd_sc_hd__dfrtp_4
X_3839_ _6460_/Q _6657_/Q _3835_/S _6461_/Q VGND VGND VPWR VPWR _3841_/A sky130_fd_sc_hd__o211a_1
XFILLER_192_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6558_ _6568_/CLK _6558_/D VGND VGND VPWR VPWR _6558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5509_ _5509_/A0 _5572_/A1 _5514_/S VGND VGND VPWR VPWR _5509_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6489_ _7203_/CLK _6489_/D _6409_/A VGND VGND VPWR VPWR _6489_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_126_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5860_ _5860_/A1 _6342_/S _5858_/X _5859_/X VGND VGND VPWR VPWR _7167_/D sky130_fd_sc_hd__o22a_1
XFILLER_61_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4811_ _4679_/Y _4811_/B VGND VGND VPWR VPWR _5021_/A sky130_fd_sc_hd__nand2b_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5791_ _6849_/Q _5842_/A2 _5674_/X _6873_/Q _5790_/X VGND VGND VPWR VPWR _5792_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4742_ _5011_/A _4947_/A _4713_/Y VGND VGND VPWR VPWR _4742_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_193_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4673_ _4682_/A _4714_/B _4698_/C VGND VGND VPWR VPWR _4719_/B sky130_fd_sc_hd__and3_4
XFILLER_147_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6412_ _6414_/A _6433_/B VGND VGND VPWR VPWR _6412_/X sky130_fd_sc_hd__and2_1
X_3624_ _7135_/Q hold33/A _3347_/Y _7007_/Q _3623_/X VGND VGND VPWR VPWR _3627_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6343_ _6676_/Q _6677_/Q _6680_/Q _6683_/Q _3922_/B VGND VGND VPWR VPWR _6344_/A
+ sky130_fd_sc_hd__o41a_1
X_3555_ _7113_/Q _5551_/A _3336_/Y input24/X _3554_/X VGND VGND VPWR VPWR _3556_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6274_ _6704_/Q _5977_/X _5990_/X _6646_/Q _6273_/X VGND VGND VPWR VPWR _6279_/B
+ sky130_fd_sc_hd__a221o_1
X_3486_ _3686_/B _3516_/B VGND VGND VPWR VPWR _3486_/Y sky130_fd_sc_hd__nor2_2
XFILLER_130_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5225_ hold248/X hold153/X _5225_/S VGND VGND VPWR VPWR _5225_/X sky130_fd_sc_hd__mux2_1
Xhold2403 _5385_/X VGND VGND VPWR VPWR _6961_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2414 _6921_/Q VGND VGND VPWR VPWR hold756/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2425 _6774_/Q VGND VGND VPWR VPWR _3805_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2436 _6242_/X VGND VGND VPWR VPWR _7181_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1702 hold181/X VGND VGND VPWR VPWR _5437_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2447 _7199_/Q VGND VGND VPWR VPWR _6375_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5156_ _5156_/A _5156_/B _5156_/C VGND VGND VPWR VPWR _5156_/Y sky130_fd_sc_hd__nand3_1
Xhold1713 hold344/X VGND VGND VPWR VPWR _5410_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2458 hold18/A VGND VGND VPWR VPWR _3874_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1724 hold698/X VGND VGND VPWR VPWR _4311_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2469 _6781_/Q VGND VGND VPWR VPWR _3388_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1735 _6836_/Q VGND VGND VPWR VPWR hold372/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1746 hold291/X VGND VGND VPWR VPWR _4259_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4107_ _6679_/Q _6346_/B VGND VGND VPWR VPWR _4115_/S sky130_fd_sc_hd__nand2_8
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1757 _6610_/Q VGND VGND VPWR VPWR hold576/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_110_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5087_ _4417_/B _4668_/Y _4777_/X _5117_/B _5117_/A VGND VGND VPWR VPWR _5087_/X
+ sky130_fd_sc_hd__o2111a_1
Xhold1768 hold125/X VGND VGND VPWR VPWR _5241_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1779 _4209_/X VGND VGND VPWR VPWR _6646_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_4038_ _4038_/A0 _4037_/X _4046_/S VGND VGND VPWR VPWR _4038_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5989_ _6015_/B _6014_/A _6007_/C VGND VGND VPWR VPWR _5989_/X sky130_fd_sc_hd__and3_4
XFILLER_169_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_50 _5997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_61 _6744_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 _6436_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_83 input51/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_94 input90/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput190 _3216_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[23] sky130_fd_sc_hd__buf_12
XFILLER_121_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold309 hold309/A VGND VGND VPWR VPWR hold309/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3340_ _3487_/A _3563_/B VGND VGND VPWR VPWR _5389_/A sky130_fd_sc_hd__nor2_8
XFILLER_98_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _3270_/X hold955/X _3996_/S VGND VGND VPWR VPWR _3271_/X sky130_fd_sc_hd__mux2_2
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5010_ _5010_/A _5010_/B VGND VGND VPWR VPWR _5083_/C sky130_fd_sc_hd__and2_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1009 _5341_/X VGND VGND VPWR VPWR _6922_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_66_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6961_ _7105_/CLK _6961_/D fanout473/X VGND VGND VPWR VPWR _6961_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5912_ _6571_/Q _5674_/X _5680_/X _6709_/Q VGND VGND VPWR VPWR _5912_/X sky130_fd_sc_hd__a22o_1
X_6892_ _7084_/CLK _6892_/D fanout459/X VGND VGND VPWR VPWR _6892_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_34_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5843_ _6916_/Q _5670_/X _5685_/X _7076_/Q _5842_/X VGND VGND VPWR VPWR _5843_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5774_ _6953_/Q _5672_/X _5682_/X _7041_/Q VGND VGND VPWR VPWR _5774_/X sky130_fd_sc_hd__a22o_1
X_4725_ _5026_/B _4725_/B VGND VGND VPWR VPWR _5138_/B sky130_fd_sc_hd__nand2_2
XFILLER_30_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4656_ _4652_/Y _4656_/B VGND VGND VPWR VPWR _5047_/A sky130_fd_sc_hd__nand2b_1
XFILLER_190_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3607_ _6740_/Q _4310_/A _3539_/Y _6533_/Q VGND VGND VPWR VPWR _3607_/X sky130_fd_sc_hd__a22o_1
Xinput70 mgmt_gpio_in[7] VGND VGND VPWR VPWR _3973_/B sky130_fd_sc_hd__clkbuf_4
Xinput81 spi_sdo VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__clkbuf_4
Xhold810 hold810/A VGND VGND VPWR VPWR hold810/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold821 hold821/A VGND VGND VPWR VPWR hold821/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4587_ _4621_/A _4693_/B VGND VGND VPWR VPWR _4901_/B sky130_fd_sc_hd__nand2_2
Xinput92 spimemio_flash_io3_oeb VGND VGND VPWR VPWR input92/X sky130_fd_sc_hd__clkbuf_2
Xhold832 hold832/A VGND VGND VPWR VPWR hold832/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold843 hold843/A VGND VGND VPWR VPWR hold843/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6326_ _6643_/Q _5986_/X _5998_/X _6583_/Q _6325_/X VGND VGND VPWR VPWR _6327_/C
+ sky130_fd_sc_hd__a221o_1
X_3538_ _6937_/Q _5353_/A _4170_/A _6618_/Q _3537_/X VGND VGND VPWR VPWR _3543_/B
+ sky130_fd_sc_hd__a221o_1
Xhold854 hold854/A VGND VGND VPWR VPWR hold854/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold865 hold865/A VGND VGND VPWR VPWR hold865/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold876 _3994_/X VGND VGND VPWR VPWR hold19/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold887 _4247_/X VGND VGND VPWR VPWR hold21/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold898 _3996_/X VGND VGND VPWR VPWR hold77/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6257_ _6708_/Q _5992_/X _6012_/X _6748_/Q _6256_/X VGND VGND VPWR VPWR _6257_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3469_ _3563_/A _3516_/B VGND VGND VPWR VPWR _4292_/A sky130_fd_sc_hd__nor2_4
XFILLER_77_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2200 _5428_/X VGND VGND VPWR VPWR _6999_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2211 _6590_/Q VGND VGND VPWR VPWR hold720/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2222 hold814/X VGND VGND VPWR VPWR _4017_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5208_ _5208_/A0 _5208_/A1 _5208_/S VGND VGND VPWR VPWR _5208_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2233 _5571_/X VGND VGND VPWR VPWR _7126_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_6188_ _6181_/X _6183_/X _6188_/C _6339_/B VGND VGND VPWR VPWR _6189_/C sky130_fd_sc_hd__and4bb_1
Xhold2244 _5384_/X VGND VGND VPWR VPWR _6960_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2255 hold747/X VGND VGND VPWR VPWR _4294_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1510 _6652_/Q VGND VGND VPWR VPWR hold146/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1521 _6823_/Q VGND VGND VPWR VPWR hold330/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2266 _5509_/X VGND VGND VPWR VPWR _7071_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1532 _6760_/Q VGND VGND VPWR VPWR hold168/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2277 _5418_/X VGND VGND VPWR VPWR _6990_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5139_ _5139_/A _5139_/B _5139_/C VGND VGND VPWR VPWR _5140_/C sky130_fd_sc_hd__and3_1
Xhold1543 _6558_/Q VGND VGND VPWR VPWR hold836/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2288 hold703/X VGND VGND VPWR VPWR _5375_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1554 _6560_/Q VGND VGND VPWR VPWR hold842/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2299 _5420_/X VGND VGND VPWR VPWR _6992_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1565 _5361_/X VGND VGND VPWR VPWR _6940_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1576 hold138/X VGND VGND VPWR VPWR _5275_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1587 _6616_/Q VGND VGND VPWR VPWR hold193/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1598 _4215_/X VGND VGND VPWR VPWR _6651_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_53_750 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_811 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4510_ _4510_/A _4510_/B VGND VGND VPWR VPWR _4776_/A sky130_fd_sc_hd__nor2_1
XFILLER_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5490_ hold683/X _5580_/A1 _5496_/S VGND VGND VPWR VPWR _5490_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4441_ _4457_/A _4457_/C _4469_/B VGND VGND VPWR VPWR _4598_/B sky130_fd_sc_hd__a21boi_4
XFILLER_171_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold106 _7199_/Q VGND VGND VPWR VPWR hold106/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold117 hold117/A VGND VGND VPWR VPWR hold117/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold128 hold128/A VGND VGND VPWR VPWR hold128/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold139 hold139/A VGND VGND VPWR VPWR hold139/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7160_ _3950_/A1 _7160_/D fanout466/X VGND VGND VPWR VPWR _7160_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_160_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4372_ _4576_/A _4719_/A VGND VGND VPWR VPWR _5009_/A sky130_fd_sc_hd__and2_4
XFILLER_98_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6111_ _6928_/Q _5982_/X _5987_/X _7112_/Q VGND VGND VPWR VPWR _6111_/X sky130_fd_sc_hd__a22o_1
X_3323_ _3333_/A _3563_/B VGND VGND VPWR VPWR _5317_/A sky130_fd_sc_hd__nor2_8
XFILLER_98_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7091_ _7091_/CLK _7091_/D fanout481/X VGND VGND VPWR VPWR _7091_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6042_ _6042_/A1 _5649_/Y _6041_/X VGND VGND VPWR VPWR _7173_/D sky130_fd_sc_hd__a21o_1
X_3254_ hold86/X _6657_/Q hold1058/X VGND VGND VPWR VPWR _3254_/X sky130_fd_sc_hd__a21bo_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3185_ _6864_/Q VGND VGND VPWR VPWR _3185_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6944_ _7091_/CLK _6944_/D fanout471/X VGND VGND VPWR VPWR _6944_/Q sky130_fd_sc_hd__dfrtp_4
X_6875_ _7091_/CLK _6875_/D fanout471/X VGND VGND VPWR VPWR _6875_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_169_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5826_ _5826_/A _5826_/B _5826_/C VGND VGND VPWR VPWR _5826_/Y sky130_fd_sc_hd__nor3_1
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5757_ _6856_/Q _5651_/X _5679_/X _6904_/Q VGND VGND VPWR VPWR _5757_/X sky130_fd_sc_hd__a22o_1
XFILLER_182_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4708_ _4370_/Y _4947_/A _5067_/A _4707_/X VGND VGND VPWR VPWR _4708_/X sky130_fd_sc_hd__o211a_1
XFILLER_163_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5688_ _5689_/A _5689_/B _5688_/C VGND VGND VPWR VPWR _5688_/X sky130_fd_sc_hd__and3b_4
XFILLER_135_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4639_ _4650_/B _4394_/A _4639_/S VGND VGND VPWR VPWR _4640_/B sky130_fd_sc_hd__mux2_1
XFILLER_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold640 hold640/A VGND VGND VPWR VPWR hold640/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold651 hold651/A VGND VGND VPWR VPWR hold651/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold662 hold662/A VGND VGND VPWR VPWR hold662/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap370 _3868_/B VGND VGND VPWR VPWR _3866_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_150_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold673 hold673/A VGND VGND VPWR VPWR hold673/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6309_ _6627_/Q _6013_/X _6015_/X _6760_/Q VGND VGND VPWR VPWR _6309_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold684 hold684/A VGND VGND VPWR VPWR hold684/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold695 hold695/A VGND VGND VPWR VPWR hold695/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2030 _6533_/Q VGND VGND VPWR VPWR hold628/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_131_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2041 hold727/X VGND VGND VPWR VPWR _4073_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2052 _7104_/Q VGND VGND VPWR VPWR hold700/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2063 _6482_/Q VGND VGND VPWR VPWR hold618/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2074 _7005_/Q VGND VGND VPWR VPWR hold805/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2085 _7053_/Q VGND VGND VPWR VPWR hold807/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1340 _7097_/Q VGND VGND VPWR VPWR hold185/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1351 hold350/X VGND VGND VPWR VPWR _5424_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2096 _6816_/Q VGND VGND VPWR VPWR hold420/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1362 _3982_/X VGND VGND VPWR VPWR hold74/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1373 hold312/X VGND VGND VPWR VPWR _4326_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1384 _5320_/X VGND VGND VPWR VPWR hold3/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_150_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1395 _4296_/X VGND VGND VPWR VPWR _6725_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4990_ _5150_/B _4990_/B VGND VGND VPWR VPWR _4990_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_51_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3941_ _6501_/Q _3881_/C _6459_/Q VGND VGND VPWR VPWR _3941_/X sky130_fd_sc_hd__mux2_2
XFILLER_32_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6660_ _6822_/CLK _6660_/D fanout451/X VGND VGND VPWR VPWR _6660_/Q sky130_fd_sc_hd__dfrtp_4
X_3872_ hold76/A _3872_/A1 _3878_/S VGND VGND VPWR VPWR _3872_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5611_ _5611_/A _5647_/B VGND VGND VPWR VPWR _5611_/Y sky130_fd_sc_hd__nand2_2
XFILLER_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6591_ _6747_/CLK _6591_/D fanout439/X VGND VGND VPWR VPWR _6591_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_129_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5542_ _5542_/A hold13/A VGND VGND VPWR VPWR _5550_/S sky130_fd_sc_hd__and2_4
XFILLER_145_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5473_ _5473_/A0 _5572_/A1 _5478_/S VGND VGND VPWR VPWR _7039_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7212_ _7212_/A VGND VGND VPWR VPWR _7212_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_144_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4424_ _4384_/A _4658_/A _4417_/B _4522_/B _4370_/Y VGND VGND VPWR VPWR _4704_/A
+ sky130_fd_sc_hd__o32a_1
X_4355_ _4447_/B _4663_/D _4682_/A _4365_/B VGND VGND VPWR VPWR _4362_/A sky130_fd_sc_hd__nand4_4
X_7143_ _7203_/CLK _7143_/D _6414_/A VGND VGND VPWR VPWR _7143_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout405 _5221_/A1 VGND VGND VPWR VPWR _5208_/A1 sky130_fd_sc_hd__buf_8
XFILLER_141_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3306_ _3309_/A _3390_/B VGND VGND VPWR VPWR _3553_/B sky130_fd_sc_hd__nand2_8
X_7074_ _7084_/CLK _7074_/D fanout456/X VGND VGND VPWR VPWR _7074_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_86_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4286_ _4286_/A _5220_/C VGND VGND VPWR VPWR _4291_/S sky130_fd_sc_hd__and2_4
Xfanout449 fanout450/X VGND VGND VPWR VPWR fanout449/X sky130_fd_sc_hd__buf_8
XFILLER_59_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6025_ _7085_/Q _5638_/X _6018_/X _6965_/Q VGND VGND VPWR VPWR _6025_/X sky130_fd_sc_hd__a22o_1
X_3237_ _6856_/Q VGND VGND VPWR VPWR _3237_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6927_ _7119_/CLK _6927_/D fanout470/X VGND VGND VPWR VPWR _6927_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_120_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6858_ _7132_/CLK _6858_/D fanout459/X VGND VGND VPWR VPWR _6858_/Q sky130_fd_sc_hd__dfrtp_4
X_5809_ _7034_/Q _5655_/X _5656_/X _6986_/Q _5797_/Y VGND VGND VPWR VPWR _5809_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6789_ _6793_/CLK _6789_/D fanout442/X VGND VGND VPWR VPWR _6789_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold470 hold470/A VGND VGND VPWR VPWR hold470/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold481 hold481/A VGND VGND VPWR VPWR hold481/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold492 hold492/A VGND VGND VPWR VPWR hold492/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1170 _6890_/Q VGND VGND VPWR VPWR hold474/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_46_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1181 _4217_/X VGND VGND VPWR VPWR _6653_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1192 _5458_/X VGND VGND VPWR VPWR _7026_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_783 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4140_ _4140_/A _5220_/C VGND VGND VPWR VPWR _4145_/S sky130_fd_sc_hd__and2_4
XFILLER_141_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4071_ _5220_/B _5226_/B _5220_/C VGND VGND VPWR VPWR _4076_/S sky130_fd_sc_hd__and3_4
XFILLER_83_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4973_ _5136_/A _4997_/A _4973_/C VGND VGND VPWR VPWR _5135_/A sky130_fd_sc_hd__and3_1
X_6712_ _6729_/CLK _6712_/D fanout465/X VGND VGND VPWR VPWR _6712_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3924_ _6490_/Q _5643_/A VGND VGND VPWR VPWR _3924_/Y sky130_fd_sc_hd__nand2_8
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6643_ _6747_/CLK _6643_/D fanout443/X VGND VGND VPWR VPWR _6643_/Q sky130_fd_sc_hd__dfrtp_4
X_3855_ _6657_/Q _6656_/Q _6448_/Q VGND VGND VPWR VPWR _3855_/X sky130_fd_sc_hd__o21a_1
XFILLER_149_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6574_ _6747_/CLK _6574_/D fanout439/X VGND VGND VPWR VPWR _6574_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3786_ _6687_/Q _4250_/A _4158_/A _6604_/Q VGND VGND VPWR VPWR _3786_/X sky130_fd_sc_hd__a22o_1
XFILLER_164_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5525_ hold665/X _5561_/A1 _5532_/S VGND VGND VPWR VPWR _5525_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5456_ _5456_/A0 _5582_/A1 _5460_/S VGND VGND VPWR VPWR _5456_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4407_ _4477_/A _4477_/B VGND VGND VPWR VPWR _4407_/Y sky130_fd_sc_hd__nand2_4
XFILLER_121_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5387_ _5387_/A0 _5585_/A1 _5388_/S VGND VGND VPWR VPWR _5387_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7126_ _7126_/CLK _7126_/D fanout475/X VGND VGND VPWR VPWR _7126_/Q sky130_fd_sc_hd__dfstp_2
X_4338_ hold168/X _5249_/A1 _4339_/S VGND VGND VPWR VPWR _4338_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4269_ _4269_/A0 _5552_/A1 _4273_/S VGND VGND VPWR VPWR _4269_/X sky130_fd_sc_hd__mux2_1
X_7057_ _7121_/CLK _7057_/D fanout473/X VGND VGND VPWR VPWR _7057_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_87_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6008_ _6008_/A _6017_/A _6019_/C VGND VGND VPWR VPWR _6008_/X sky130_fd_sc_hd__and3_4
XFILLER_28_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_140 _5320_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_151 _5451_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_162 _5686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_173 _6632_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_184 input24/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_195 hold9/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3640_ _7055_/Q _5488_/A _3977_/A _6452_/Q _3639_/X VGND VGND VPWR VPWR _3645_/B
+ sky130_fd_sc_hd__a221o_1
X_3571_ input38/X _3293_/Y _3509_/Y _6730_/Q _3570_/X VGND VGND VPWR VPWR _3571_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5310_ hold701/X _5580_/A1 _5316_/S VGND VGND VPWR VPWR _5310_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6290_ _6527_/Q _6339_/B _6289_/Y _6341_/S VGND VGND VPWR VPWR _6290_/X sky130_fd_sc_hd__o211a_1
XFILLER_114_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5241_ _5241_/A0 hold95/X _5244_/S VGND VGND VPWR VPWR _5241_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5172_ _5172_/A0 _5187_/A1 _5174_/S VGND VGND VPWR VPWR _5172_/X sky130_fd_sc_hd__mux2_1
X_4123_ _4123_/A0 _5208_/A1 _4127_/S VGND VGND VPWR VPWR _4123_/X sky130_fd_sc_hd__mux2_1
Xhold1906 hold539/X VGND VGND VPWR VPWR _5274_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1917 _4180_/X VGND VGND VPWR VPWR _6622_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1928 _4330_/X VGND VGND VPWR VPWR _6753_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1939 hold308/X VGND VGND VPWR VPWR _5356_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4054_ _4054_/A0 _5585_/A1 _4055_/S VGND VGND VPWR VPWR _4054_/X sky130_fd_sc_hd__mux2_1
Xinput2 debug_oeb VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4956_ _4466_/A _4477_/Y _4934_/Y _4784_/X VGND VGND VPWR VPWR _5034_/C sky130_fd_sc_hd__o31a_1
X_3907_ _7154_/Q _7153_/Q VGND VGND VPWR VPWR _6015_/B sky130_fd_sc_hd__and2b_4
X_4887_ _4947_/B _4570_/A _4986_/C _4885_/X _5023_/A VGND VGND VPWR VPWR _4892_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_165_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6626_ _6750_/CLK _6626_/D fanout446/X VGND VGND VPWR VPWR _6626_/Q sky130_fd_sc_hd__dfstp_2
X_3838_ _3838_/A1 _3835_/S _3837_/X VGND VGND VPWR VPWR _6463_/D sky130_fd_sc_hd__o21a_1
X_6557_ _6568_/CLK _6557_/D VGND VGND VPWR VPWR _6557_/Q sky130_fd_sc_hd__dfxtp_1
X_3769_ _3769_/A _3769_/B _3769_/C _3769_/D VGND VGND VPWR VPWR _3770_/C sky130_fd_sc_hd__nor4_1
XFILLER_118_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5508_ hold706/X _5580_/A1 _5514_/S VGND VGND VPWR VPWR _5508_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6488_ _7013_/CLK _6488_/D fanout452/X VGND VGND VPWR VPWR _6488_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5439_ _5439_/A0 _5556_/A1 _5442_/S VGND VGND VPWR VPWR _7009_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7109_ _7109_/CLK _7109_/D fanout453/X VGND VGND VPWR VPWR _7109_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_74_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4810_ _4583_/B _4688_/A _4688_/C _4729_/A VGND VGND VPWR VPWR _4820_/A sky130_fd_sc_hd__o22a_1
XFILLER_178_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5790_ _6977_/Q _5660_/X _5662_/X _6897_/Q VGND VGND VPWR VPWR _5790_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4741_ _4415_/B _4712_/Y _4740_/X VGND VGND VPWR VPWR _4741_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4672_ _4714_/B _4672_/B VGND VGND VPWR VPWR _4672_/Y sky130_fd_sc_hd__nand2_1
XFILLER_175_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6411_ _6414_/A _6423_/B VGND VGND VPWR VPWR _6411_/X sky130_fd_sc_hd__and2_1
X_3623_ _7071_/Q _5506_/A _4328_/A _6754_/Q VGND VGND VPWR VPWR _3623_/X sky130_fd_sc_hd__a22o_1
XFILLER_190_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6342_ _6342_/A0 _6341_/X _6342_/S VGND VGND VPWR VPWR _7185_/D sky130_fd_sc_hd__mux2_1
X_3554_ _7057_/Q _5488_/A _4176_/A _6623_/Q VGND VGND VPWR VPWR _3554_/X sky130_fd_sc_hd__a22o_1
X_6273_ _6596_/Q _5991_/X _5997_/X _6699_/Q VGND VGND VPWR VPWR _6273_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3485_ _6929_/Q _5344_/A _4047_/C input48/X _3484_/X VGND VGND VPWR VPWR _3499_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_143_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5224_ hold273/X _5544_/A1 _5224_/S VGND VGND VPWR VPWR _5224_/X sky130_fd_sc_hd__mux2_1
Xhold2404 _6905_/Q VGND VGND VPWR VPWR hold749/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2415 hold756/X VGND VGND VPWR VPWR _5340_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2426 _6681_/Q VGND VGND VPWR VPWR _3919_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2437 _6682_/Q VGND VGND VPWR VPWR _3968_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1703 _6886_/Q VGND VGND VPWR VPWR hold481/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5155_ _5155_/A _5155_/B _5155_/C _5155_/D VGND VGND VPWR VPWR _5156_/C sky130_fd_sc_hd__and4_1
Xhold2448 hold4/A VGND VGND VPWR VPWR _3872_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1714 _6689_/Q VGND VGND VPWR VPWR hold280/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2459 _6676_/Q VGND VGND VPWR VPWR _3921_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1725 _6832_/Q VGND VGND VPWR VPWR hold299/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1736 hold372/X VGND VGND VPWR VPWR _5244_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4106_ _3385_/Y hold842/A _4106_/S VGND VGND VPWR VPWR _6560_/D sky130_fd_sc_hd__mux2_1
Xhold1747 _4259_/X VGND VGND VPWR VPWR _6694_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5086_ _5086_/A _5086_/B VGND VGND VPWR VPWR _5086_/Y sky130_fd_sc_hd__nand2_1
Xhold1758 hold576/X VGND VGND VPWR VPWR _4166_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1769 _6451_/Q VGND VGND VPWR VPWR hold524/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4037_ hold704/X _5582_/A1 _4056_/C VGND VGND VPWR VPWR _4037_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5988_ _6015_/B _6018_/B _6007_/C VGND VGND VPWR VPWR _5988_/X sky130_fd_sc_hd__and3_4
XFILLER_40_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4939_ _4936_/Y _4938_/X _4776_/Y VGND VGND VPWR VPWR _5117_/B sky130_fd_sc_hd__o21a_1
XFILLER_138_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_40 _5688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_51 _5998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 _6531_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 _7212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_84 input59/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6609_ _6648_/CLK _6609_/D _6426_/A VGND VGND VPWR VPWR _6609_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_95 input93/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput180 _3226_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[14] sky130_fd_sc_hd__buf_12
Xoutput191 _3215_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[24] sky130_fd_sc_hd__buf_12
XFILLER_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_44_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _6903_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_140_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3270_ _6460_/Q wire1/X _6657_/Q VGND VGND VPWR VPWR _3270_/X sky130_fd_sc_hd__mux2_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_59_csclk _7093_/CLK VGND VGND VPWR VPWR _7117_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6960_ _7138_/CLK _6960_/D fanout477/X VGND VGND VPWR VPWR _6960_/Q sky130_fd_sc_hd__dfrtp_4
X_5911_ _6754_/Q _5681_/X _5910_/X VGND VGND VPWR VPWR _5911_/X sky130_fd_sc_hd__a21o_1
XFILLER_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6891_ _7131_/CLK _6891_/D fanout469/X VGND VGND VPWR VPWR _6891_/Q sky130_fd_sc_hd__dfrtp_4
X_5842_ _6852_/Q _5842_/A2 _5840_/X _5841_/X VGND VGND VPWR VPWR _5842_/X sky130_fd_sc_hd__a211o_1
XFILLER_179_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5773_ _5794_/A0 _5772_/X _6342_/S VGND VGND VPWR VPWR _5773_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4724_ _5001_/A _4724_/B _4724_/C VGND VGND VPWR VPWR _4920_/B sky130_fd_sc_hd__nand3_2
XFILLER_159_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4655_ _4655_/A _4655_/B VGND VGND VPWR VPWR _4656_/B sky130_fd_sc_hd__nor2_1
XFILLER_107_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput60 mgmt_gpio_in[31] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__buf_2
Xhold800 hold800/A VGND VGND VPWR VPWR hold800/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3606_ _6840_/Q hold27/A _4212_/A _6652_/Q _3605_/X VGND VGND VPWR VPWR _3614_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_190_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput71 mgmt_gpio_in[8] VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__clkbuf_2
Xhold811 hold811/A VGND VGND VPWR VPWR hold811/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput82 spi_sdoenb VGND VGND VPWR VPWR input82/X sky130_fd_sc_hd__buf_4
X_4586_ _4625_/A _4628_/A VGND VGND VPWR VPWR _4586_/Y sky130_fd_sc_hd__nand2_2
Xinput93 trap VGND VGND VPWR VPWR input93/X sky130_fd_sc_hd__buf_6
Xhold822 hold822/A VGND VGND VPWR VPWR hold822/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold833 hold833/A VGND VGND VPWR VPWR hold833/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6325_ _6613_/Q _5976_/B _5993_/X _6623_/Q VGND VGND VPWR VPWR _6325_/X sky130_fd_sc_hd__a22o_1
XFILLER_89_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold844 hold844/A VGND VGND VPWR VPWR hold844/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3537_ _7049_/Q _5479_/A _4268_/A _6706_/Q VGND VGND VPWR VPWR _3537_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold855 hold855/A VGND VGND VPWR VPWR hold855/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold866 hold866/A VGND VGND VPWR VPWR hold866/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold877 hold19/X VGND VGND VPWR VPWR hold877/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold888 _6765_/Q VGND VGND VPWR VPWR hold65/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6256_ _6698_/Q _5997_/X _6004_/X _6575_/Q VGND VGND VPWR VPWR _6256_/X sky130_fd_sc_hd__a22o_1
Xhold899 hold77/X VGND VGND VPWR VPWR hold899/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_3468_ _7073_/Q _5506_/A _4250_/A _6691_/Q _3466_/X VGND VGND VPWR VPWR _3481_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2201 _6591_/Q VGND VGND VPWR VPWR hold557/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2212 hold720/X VGND VGND VPWR VPWR _4142_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2223 _4017_/X VGND VGND VPWR VPWR _6494_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5207_ _5207_/A _5222_/A _5220_/C VGND VGND VPWR VPWR _5208_/S sky130_fd_sc_hd__and3_1
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2234 _6991_/Q VGND VGND VPWR VPWR hold549/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6187_ _6923_/Q _5995_/X _6184_/X _6186_/X VGND VGND VPWR VPWR _6188_/C sky130_fd_sc_hd__a211oi_1
XFILLER_97_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3399_ _6955_/Q _5371_/A _5326_/A _6915_/Q VGND VGND VPWR VPWR _3399_/X sky130_fd_sc_hd__a22o_1
Xhold2245 _7070_/Q VGND VGND VPWR VPWR hold706/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1500 _6985_/Q VGND VGND VPWR VPWR hold682/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2256 _6721_/Q VGND VGND VPWR VPWR hold475/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1511 _7052_/Q VGND VGND VPWR VPWR hold501/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1522 hold330/X VGND VGND VPWR VPWR _5230_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2267 _7212_/A VGND VGND VPWR VPWR hold808/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1533 _7108_/Q VGND VGND VPWR VPWR hold518/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2278 _6895_/Q VGND VGND VPWR VPWR hold580/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5138_ _5138_/A _5138_/B _5138_/C VGND VGND VPWR VPWR _5148_/C sky130_fd_sc_hd__and3_1
Xhold1544 hold836/X VGND VGND VPWR VPWR hold260/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2289 _6717_/Q VGND VGND VPWR VPWR hold803/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1555 hold842/X VGND VGND VPWR VPWR hold267/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1566 _7068_/Q VGND VGND VPWR VPWR hold505/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1577 _5275_/X VGND VGND VPWR VPWR _6863_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_123_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1588 _6544_/Q VGND VGND VPWR VPWR hold856/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5069_ _5069_/A _5069_/B VGND VGND VPWR VPWR _5072_/C sky130_fd_sc_hd__and2_1
Xhold1599 _6855_/Q VGND VGND VPWR VPWR hold144/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_53_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4440_ _4701_/A _4808_/B _4917_/A VGND VGND VPWR VPWR _4457_/C sky130_fd_sc_hd__a21o_2
XFILLER_7_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold107 hold107/A VGND VGND VPWR VPWR hold107/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold118 hold118/A VGND VGND VPWR VPWR hold118/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold129 hold129/A VGND VGND VPWR VPWR hold129/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4371_ _4637_/A _4637_/B VGND VGND VPWR VPWR _4719_/A sky130_fd_sc_hd__and2b_4
XFILLER_125_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6110_ _6864_/Q _5999_/X _6019_/X _6984_/Q _6109_/X VGND VGND VPWR VPWR _6113_/C
+ sky130_fd_sc_hd__a221o_1
X_3322_ _3355_/A _3322_/B VGND VGND VPWR VPWR _3353_/A sky130_fd_sc_hd__nand2_8
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7090_ _7124_/CLK _7090_/D fanout459/X VGND VGND VPWR VPWR _7090_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6041_ _6837_/Q _6339_/B _6029_/X _6040_/Y _5647_/Y VGND VGND VPWR VPWR _6041_/X
+ sky130_fd_sc_hd__o221a_2
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _3253_/A _3862_/A VGND VGND VPWR VPWR _3253_/Y sky130_fd_sc_hd__nand2_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3184_ _3921_/A VGND VGND VPWR VPWR _3184_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6943_ _6945_/CLK _6943_/D _6409_/A VGND VGND VPWR VPWR _6943_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6874_ _7020_/CLK _6874_/D fanout458/X VGND VGND VPWR VPWR _6874_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5825_ _6955_/Q _5672_/X _5822_/X _5824_/X VGND VGND VPWR VPWR _5826_/C sky130_fd_sc_hd__a211o_1
XFILLER_50_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5756_ _6936_/Q _5659_/X _5669_/X _7048_/Q VGND VGND VPWR VPWR _5756_/X sky130_fd_sc_hd__a22o_1
X_4707_ _4391_/Y _4969_/A _4705_/Y _4832_/D _4640_/Y VGND VGND VPWR VPWR _4707_/X
+ sky130_fd_sc_hd__a41o_1
X_5687_ _5686_/A _5689_/B _5687_/C VGND VGND VPWR VPWR _5687_/X sky130_fd_sc_hd__and3b_4
XFILLER_108_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4638_ _4638_/A _4638_/B VGND VGND VPWR VPWR _4638_/Y sky130_fd_sc_hd__nand2_8
Xhold630 hold630/A VGND VGND VPWR VPWR hold630/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold641 hold641/A VGND VGND VPWR VPWR hold641/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4569_ _4569_/A _4569_/B _4569_/C VGND VGND VPWR VPWR _4569_/X sky130_fd_sc_hd__and3_1
XFILLER_162_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold652 _5237_/X VGND VGND VPWR VPWR _6829_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap360 hold54/X VGND VGND VPWR VPWR _3333_/A sky130_fd_sc_hd__buf_12
Xhold663 hold663/A VGND VGND VPWR VPWR hold663/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold674 hold674/A VGND VGND VPWR VPWR hold674/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6308_ _6632_/Q _5971_/X _5990_/X _6647_/Q _6307_/X VGND VGND VPWR VPWR _6308_/X
+ sky130_fd_sc_hd__a221o_1
Xhold685 hold685/A VGND VGND VPWR VPWR hold685/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold696 hold696/A VGND VGND VPWR VPWR hold696/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6239_ _6233_/X _6339_/B _6239_/C _6239_/D VGND VGND VPWR VPWR _6239_/X sky130_fd_sc_hd__and4b_1
XFILLER_77_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2020 hold601/X VGND VGND VPWR VPWR _4144_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_58_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2031 hold628/X VGND VGND VPWR VPWR _4075_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_103_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2042 _4073_/X VGND VGND VPWR VPWR _6531_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_131_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2053 hold700/X VGND VGND VPWR VPWR _5546_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2064 _6798_/Q VGND VGND VPWR VPWR hold599/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1330 _6876_/Q VGND VGND VPWR VPWR hold343/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2075 _7137_/Q VGND VGND VPWR VPWR hold712/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2086 _5489_/X VGND VGND VPWR VPWR _7053_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1341 hold185/X VGND VGND VPWR VPWR _5538_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2097 _7061_/Q VGND VGND VPWR VPWR hold806/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1352 _5424_/X VGND VGND VPWR VPWR _6996_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1363 hold74/X VGND VGND VPWR VPWR hold2/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1374 _4326_/X VGND VGND VPWR VPWR _6750_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_150_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1385 _6637_/Q VGND VGND VPWR VPWR hold323/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1396 _7221_/A VGND VGND VPWR VPWR hold160/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3940_ _6502_/Q _3940_/A1 _6458_/Q VGND VGND VPWR VPWR _3940_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3871_ wire1/X _3866_/A _3869_/A _3903_/A _3870_/X VGND VGND VPWR VPWR _6445_/D sky130_fd_sc_hd__a221o_1
XFILLER_32_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5610_ _5610_/A _5610_/B VGND VGND VPWR VPWR _5639_/A sky130_fd_sc_hd__nor2_2
X_6590_ _6742_/CLK _6590_/D fanout440/X VGND VGND VPWR VPWR _6590_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5541_ _5541_/A0 hold6/X _5541_/S VGND VGND VPWR VPWR _5541_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5472_ hold759/X _5580_/A1 _5478_/S VGND VGND VPWR VPWR _7038_/D sky130_fd_sc_hd__mux2_1
X_7211_ _7211_/A VGND VGND VPWR VPWR _7211_/X sky130_fd_sc_hd__clkbuf_2
X_4423_ _4575_/C _4523_/A VGND VGND VPWR VPWR _4522_/B sky130_fd_sc_hd__nand2b_4
XFILLER_172_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7142_ _7183_/CLK _7142_/D _6414_/A VGND VGND VPWR VPWR _7142_/Q sky130_fd_sc_hd__dfrtp_4
X_4354_ _4447_/B _4663_/D _4682_/A _4365_/B VGND VGND VPWR VPWR _4356_/B sky130_fd_sc_hd__and4_2
XFILLER_125_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout406 hold153/X VGND VGND VPWR VPWR _5221_/A1 sky130_fd_sc_hd__buf_12
XFILLER_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout417 _6166_/S VGND VGND VPWR VPWR _6341_/S sky130_fd_sc_hd__buf_12
X_3305_ _3305_/A _3305_/B VGND VGND VPWR VPWR _3390_/B sky130_fd_sc_hd__and2_4
Xfanout439 fanout440/X VGND VGND VPWR VPWR fanout439/X sky130_fd_sc_hd__buf_12
X_7073_ _7137_/CLK _7073_/D fanout476/X VGND VGND VPWR VPWR _7073_/Q sky130_fd_sc_hd__dfrtp_4
X_4285_ _4285_/A0 _5538_/A1 _4285_/S VGND VGND VPWR VPWR _4285_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6024_ _7077_/Q _6013_/X _6017_/X _7069_/Q _6023_/X VGND VGND VPWR VPWR _6024_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_140_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3236_ _6872_/Q VGND VGND VPWR VPWR _3236_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_67_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6926_ _7127_/CLK _6926_/D fanout477/X VGND VGND VPWR VPWR _6926_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_23_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6857_ _6941_/CLK _6857_/D fanout460/X VGND VGND VPWR VPWR _6857_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5808_ _7090_/Q _5681_/X _5803_/X _5804_/X _5807_/X VGND VGND VPWR VPWR _5808_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_167_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6788_ _6788_/CLK _6788_/D _3959_/B VGND VGND VPWR VPWR _6788_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_183_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5739_ _6871_/Q _5674_/X _5736_/X _5738_/X VGND VGND VPWR VPWR _5739_/X sky130_fd_sc_hd__a211o_1
XFILLER_182_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold460 hold460/A VGND VGND VPWR VPWR hold460/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold471 hold471/A VGND VGND VPWR VPWR hold471/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold482 hold482/A VGND VGND VPWR VPWR hold482/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold493 hold493/A VGND VGND VPWR VPWR hold493/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1160 _5342_/X VGND VGND VPWR VPWR _6923_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1171 hold474/X VGND VGND VPWR VPWR _5305_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1182 _7034_/Q VGND VGND VPWR VPWR hold472/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_18_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1193 _7050_/Q VGND VGND VPWR VPWR hold494/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_2__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _6656_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4070_ hold122/X _5538_/A1 _4070_/S VGND VGND VPWR VPWR _6529_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4972_ _4972_/A _4972_/B VGND VGND VPWR VPWR _4972_/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6711_ _6711_/CLK _6711_/D _6432_/A VGND VGND VPWR VPWR _6711_/Q sky130_fd_sc_hd__dfrtp_4
X_3923_ _6816_/Q _5610_/A _3197_/Y _3915_/Y VGND VGND VPWR VPWR _3923_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_149_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6642_ _6747_/CLK _6642_/D fanout450/X VGND VGND VPWR VPWR _6642_/Q sky130_fd_sc_hd__dfrtp_4
X_3854_ _3903_/A _3926_/B1 _3807_/B _3854_/B1 VGND VGND VPWR VPWR _6456_/D sky130_fd_sc_hd__a31o_1
XFILLER_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6573_ _6816_/CLK _6573_/D _6409_/A VGND VGND VPWR VPWR _6573_/Q sky130_fd_sc_hd__dfrtp_4
X_3785_ _6479_/Q _3357_/Y _4304_/A _6732_/Q _3784_/X VGND VGND VPWR VPWR _3792_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5524_ _5524_/A _5569_/B VGND VGND VPWR VPWR _5532_/S sky130_fd_sc_hd__and2_4
XFILLER_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5455_ _5455_/A0 _5572_/A1 _5460_/S VGND VGND VPWR VPWR _5455_/X sky130_fd_sc_hd__mux2_1
X_4406_ _4477_/A _4477_/B VGND VGND VPWR VPWR _5150_/A sky130_fd_sc_hd__and2_2
XFILLER_160_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5386_ hold979/X _5575_/A1 _5388_/S VGND VGND VPWR VPWR _5386_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7125_ _7125_/CLK _7125_/D fanout454/X VGND VGND VPWR VPWR _7125_/Q sky130_fd_sc_hd__dfstp_2
X_4337_ hold307/X _4337_/A1 _4339_/S VGND VGND VPWR VPWR _6759_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7056_ _7136_/CLK _7056_/D fanout475/X VGND VGND VPWR VPWR _7056_/Q sky130_fd_sc_hd__dfrtp_4
X_4268_ _4268_/A _5551_/B VGND VGND VPWR VPWR _4273_/S sky130_fd_sc_hd__and2_4
XFILLER_115_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6007_ _6017_/A _6019_/C _6007_/C VGND VGND VPWR VPWR _6007_/X sky130_fd_sc_hd__and3_4
X_3219_ _7000_/Q VGND VGND VPWR VPWR _3219_/Y sky130_fd_sc_hd__inv_2
X_4199_ _4199_/A0 _4339_/A1 _4199_/S VGND VGND VPWR VPWR _4199_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6909_ _7013_/CLK _6909_/D fanout452/X VGND VGND VPWR VPWR _6909_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_168_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold290 hold290/A VGND VGND VPWR VPWR hold290/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_130 _3940_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_141 _4309_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_152 _5451_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_163 _5687_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 _7048_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_185 _3974_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_196 hold135/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3570_ _6597_/Q _4146_/A _4134_/A _6587_/Q VGND VGND VPWR VPWR _3570_/X sky130_fd_sc_hd__a22o_2
XFILLER_127_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5240_ _5240_/A0 _5303_/A1 _5244_/S VGND VGND VPWR VPWR _5240_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_702 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5171_ _5171_/A0 _5193_/A1 _5174_/S VGND VGND VPWR VPWR _5171_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4122_ _4122_/A _5220_/C VGND VGND VPWR VPWR _4127_/S sky130_fd_sc_hd__and2_4
Xhold1907 _5274_/X VGND VGND VPWR VPWR _6862_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1918 _6579_/Q VGND VGND VPWR VPWR hold735/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1929 _7037_/Q VGND VGND VPWR VPWR hold639/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4053_ hold925/X hold20/X _4055_/S VGND VGND VPWR VPWR _4053_/X sky130_fd_sc_hd__mux2_1
Xinput3 debug_out VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4955_ _4955_/A _4955_/B _4955_/C _4955_/D VGND VGND VPWR VPWR _4957_/C sky130_fd_sc_hd__nand4_1
XFILLER_178_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3906_ _7151_/Q _7152_/Q VGND VGND VPWR VPWR _6019_/A sky130_fd_sc_hd__and2b_4
X_4886_ _4886_/A _4976_/A VGND VGND VPWR VPWR _5023_/A sky130_fd_sc_hd__nor2_4
XFILLER_193_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6625_ _6759_/CLK _6625_/D fanout449/X VGND VGND VPWR VPWR _6625_/Q sky130_fd_sc_hd__dfrtp_4
X_3837_ _6462_/Q _6657_/Q _3830_/Y _3836_/X _3846_/S VGND VGND VPWR VPWR _3837_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6556_ _6568_/CLK _6556_/D VGND VGND VPWR VPWR _6556_/Q sky130_fd_sc_hd__dfxtp_1
X_3768_ _6869_/Q _5281_/A _4334_/A _6757_/Q _3767_/X VGND VGND VPWR VPWR _3769_/D
+ sky130_fd_sc_hd__a221o_1
X_5507_ hold816/X _5552_/A1 _5514_/S VGND VGND VPWR VPWR _7069_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6487_ _7013_/CLK _6487_/D fanout452/X VGND VGND VPWR VPWR _6487_/Q sky130_fd_sc_hd__dfstp_2
X_3699_ _6822_/Q _5226_/A _5226_/B _5202_/A _6805_/Q VGND VGND VPWR VPWR _3699_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_106_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5438_ hold532/X _5555_/A1 _5442_/S VGND VGND VPWR VPWR _7008_/D sky130_fd_sc_hd__mux2_1
Xoutput340 hold1347/X VGND VGND VPWR VPWR hold272/A sky130_fd_sc_hd__buf_6
XFILLER_161_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5369_ _5369_/A0 _5585_/A1 _5370_/S VGND VGND VPWR VPWR _5369_/X sky130_fd_sc_hd__mux2_1
X_7108_ _7124_/CLK _7108_/D fanout459/X VGND VGND VPWR VPWR _7108_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_75_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7039_ _7137_/CLK _7039_/D fanout476/X VGND VGND VPWR VPWR _7039_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_142_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire434 _4808_/A VGND VGND VPWR VPWR _4584_/A sky130_fd_sc_hd__buf_2
XFILLER_7_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ _4411_/Y _4712_/Y _4728_/Y _4737_/Y _4739_/X VGND VGND VPWR VPWR _4740_/X
+ sky130_fd_sc_hd__o2111a_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4671_ _4671_/A _4683_/A VGND VGND VPWR VPWR _4691_/B sky130_fd_sc_hd__nor2_8
XFILLER_175_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6410_ _6414_/A _6433_/B VGND VGND VPWR VPWR _6410_/X sky130_fd_sc_hd__and2_1
X_3622_ _7015_/Q _5443_/A _5362_/A _6943_/Q _3621_/X VGND VGND VPWR VPWR _3627_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6341_ _6341_/A0 _6340_/X _6341_/S VGND VGND VPWR VPWR _6341_/X sky130_fd_sc_hd__mux2_1
X_3553_ _3553_/A _3553_/B VGND VGND VPWR VPWR _4176_/A sky130_fd_sc_hd__nor2_8
X_6272_ _6601_/Q _5995_/X _6019_/X _6734_/Q _6271_/X VGND VGND VPWR VPWR _6279_/A
+ sky130_fd_sc_hd__a221o_1
X_3484_ _6633_/Q _4188_/A _4316_/A _6746_/Q VGND VGND VPWR VPWR _3484_/X sky130_fd_sc_hd__a22o_2
XFILLER_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5223_ _5223_/A0 _5572_/A1 _5224_/S VGND VGND VPWR VPWR _6818_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2405 hold749/X VGND VGND VPWR VPWR _5322_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2416 _7069_/Q VGND VGND VPWR VPWR hold816/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2427 _6678_/Q VGND VGND VPWR VPWR _3917_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5154_ _4402_/Y _4570_/C _4570_/D _4968_/Y _4534_/Y VGND VGND VPWR VPWR _5155_/D
+ sky130_fd_sc_hd__o221a_1
Xhold2438 _7196_/Q VGND VGND VPWR VPWR _6366_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1704 _6830_/Q VGND VGND VPWR VPWR hold177/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2449 _3872_/X VGND VGND VPWR VPWR _6444_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1715 hold280/X VGND VGND VPWR VPWR _4253_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1726 hold299/X VGND VGND VPWR VPWR _5240_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4105_ _3422_/Y hold828/A _4106_/S VGND VGND VPWR VPWR _6559_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1737 _7065_/Q VGND VGND VPWR VPWR hold131/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1748 _7189_/Q VGND VGND VPWR VPWR hold852/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5085_ _5143_/A _5139_/C _5165_/B _5006_/Y VGND VGND VPWR VPWR _5085_/X sky130_fd_sc_hd__a31o_1
Xhold1759 _6934_/Q VGND VGND VPWR VPWR hold508/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_110_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4036_ hold405/X _4036_/A1 _4046_/S VGND VGND VPWR VPWR _4036_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5987_ _6019_/A _6008_/A _6019_/C VGND VGND VPWR VPWR _5987_/X sky130_fd_sc_hd__and3_4
XFILLER_24_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4938_ _5011_/A _4601_/A _4466_/A VGND VGND VPWR VPWR _4938_/X sky130_fd_sc_hd__a21o_2
XFILLER_21_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_30 _5660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_41 _5688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4869_ _4570_/C _4655_/A _4590_/Y _4713_/Y VGND VGND VPWR VPWR _4870_/D sky130_fd_sc_hd__o22a_1
XANTENNA_52 _6012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_63 _6750_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6608_ _6711_/CLK _6608_/D fanout465/X VGND VGND VPWR VPWR _6608_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_74 _6508_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_85 input59/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_96 input95/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6539_ _6757_/CLK _6539_/D fanout446/X VGND VGND VPWR VPWR _6539_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_146_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput181 _3225_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[15] sky130_fd_sc_hd__buf_12
Xoutput192 _3214_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[25] sky130_fd_sc_hd__buf_12
XFILLER_88_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5910_ _6694_/Q _5658_/X _5664_/X _6759_/Q VGND VGND VPWR VPWR _5910_/X sky130_fd_sc_hd__a22o_1
X_6890_ _7035_/CLK _6890_/D fanout455/X VGND VGND VPWR VPWR _6890_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5841_ _6860_/Q _5651_/X _5662_/X _6900_/Q VGND VGND VPWR VPWR _5841_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5772_ _6490_/Q _7162_/Q _5771_/X VGND VGND VPWR VPWR _5772_/X sky130_fd_sc_hd__a21bo_1
XFILLER_148_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4723_ _4812_/A _4725_/B VGND VGND VPWR VPWR _4770_/B sky130_fd_sc_hd__nand2_1
XFILLER_147_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4654_ _4917_/C _4838_/B _4917_/B VGND VGND VPWR VPWR _4655_/B sky130_fd_sc_hd__nand3b_2
XFILLER_174_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput50 mgmt_gpio_in[22] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__clkbuf_2
X_3605_ _7056_/Q _5488_/A _4328_/A _6755_/Q VGND VGND VPWR VPWR _3605_/X sky130_fd_sc_hd__a22o_1
Xinput61 mgmt_gpio_in[32] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__buf_2
Xhold801 hold801/A VGND VGND VPWR VPWR hold801/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput72 mgmt_gpio_in[9] VGND VGND VPWR VPWR input72/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4585_ _4948_/A _4724_/C VGND VGND VPWR VPWR _4973_/C sky130_fd_sc_hd__nand2_1
Xhold812 hold812/A VGND VGND VPWR VPWR hold812/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold823 hold823/A VGND VGND VPWR VPWR hold823/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput83 spimemio_flash_clk VGND VGND VPWR VPWR input83/X sky130_fd_sc_hd__clkbuf_4
Xinput94 uart_enabled VGND VGND VPWR VPWR _3970_/B sky130_fd_sc_hd__clkbuf_2
X_6324_ _6633_/Q _5971_/X _6007_/X _6534_/Q _6323_/X VGND VGND VPWR VPWR _6327_/B
+ sky130_fd_sc_hd__a221o_1
Xhold834 hold834/A VGND VGND VPWR VPWR hold834/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3536_ _3563_/A _3553_/B VGND VGND VPWR VPWR _4268_/A sky130_fd_sc_hd__nor2_4
XFILLER_116_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold845 hold845/A VGND VGND VPWR VPWR hold845/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold856 hold856/A VGND VGND VPWR VPWR hold856/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold867 hold867/A VGND VGND VPWR VPWR hold867/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold878 hold878/A VGND VGND VPWR VPWR hold20/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6255_ _6255_/A _6255_/B _6255_/C VGND VGND VPWR VPWR _6264_/C sky130_fd_sc_hd__nor3_2
Xhold889 hold65/X VGND VGND VPWR VPWR hold889/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_3467_ _3550_/A _3531_/B VGND VGND VPWR VPWR _4250_/A sky130_fd_sc_hd__nor2_8
XFILLER_103_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2202 _6643_/Q VGND VGND VPWR VPWR hold442/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5206_ _5206_/A0 _5303_/A1 _5206_/S VGND VGND VPWR VPWR _5206_/X sky130_fd_sc_hd__mux2_1
Xhold2213 _6808_/Q VGND VGND VPWR VPWR hold728/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2224 _6783_/Q VGND VGND VPWR VPWR hold757/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6186_ _6851_/Q _6007_/X _6019_/X _6987_/Q _6185_/X VGND VGND VPWR VPWR _6186_/X
+ sky130_fd_sc_hd__a221o_1
X_3398_ _6891_/Q _5299_/A _3389_/Y _3395_/X _3397_/X VGND VGND VPWR VPWR _3406_/A
+ sky130_fd_sc_hd__a2111o_1
Xhold2235 hold549/X VGND VGND VPWR VPWR _5419_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2246 _5508_/X VGND VGND VPWR VPWR _7070_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1501 hold682/X VGND VGND VPWR VPWR _5412_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1512 hold501/X VGND VGND VPWR VPWR _5487_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2257 hold475/X VGND VGND VPWR VPWR _4291_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5137_ _5086_/Y _5137_/B _5137_/C VGND VGND VPWR VPWR _5137_/X sky130_fd_sc_hd__and3b_1
Xhold1523 _5230_/X VGND VGND VPWR VPWR hold331/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2268 hold808/X VGND VGND VPWR VPWR _4038_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1534 hold518/X VGND VGND VPWR VPWR _5550_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2279 hold580/X VGND VGND VPWR VPWR _5311_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1545 _6568_/Q VGND VGND VPWR VPWR hold850/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1556 _6555_/Q VGND VGND VPWR VPWR hold832/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1567 hold505/X VGND VGND VPWR VPWR _5505_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5068_ _4391_/Y _4580_/Y _4584_/Y _4765_/Y _4438_/Y VGND VGND VPWR VPWR _5069_/B
+ sky130_fd_sc_hd__a41o_1
Xhold1578 _6865_/Q VGND VGND VPWR VPWR hold109/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1589 hold856/X VGND VGND VPWR VPWR hold198/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4019_ _4019_/A0 _4018_/X _4029_/S VGND VGND VPWR VPWR _4019_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold108 hold108/A VGND VGND VPWR VPWR _6711_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold119 hold119/A VGND VGND VPWR VPWR hold119/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4370_ _4955_/A _4513_/B VGND VGND VPWR VPWR _4370_/Y sky130_fd_sc_hd__nand2_2
XFILLER_98_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3321_ _3563_/A _3470_/A VGND VGND VPWR VPWR _5551_/A sky130_fd_sc_hd__nor2_8
XFILLER_113_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6032_/X _6040_/B _6339_/B VGND VGND VPWR VPWR _6040_/Y sky130_fd_sc_hd__nand3b_2
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _3996_/S _3252_/A2 hold23/X VGND VGND VPWR VPWR _3252_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_140_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3183_ _6437_/Q VGND VGND VPWR VPWR _3183_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6942_ _7134_/CLK _6942_/D fanout476/X VGND VGND VPWR VPWR _6942_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6873_ _7111_/CLK _6873_/D fanout472/X VGND VGND VPWR VPWR _6873_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5824_ _6987_/Q _5656_/X _5668_/X _7059_/Q _5823_/X VGND VGND VPWR VPWR _5824_/X
+ sky130_fd_sc_hd__a221o_1
X_5755_ _6992_/Q _5929_/B _5682_/X _7040_/Q _5754_/X VGND VGND VPWR VPWR _5760_/B
+ sky130_fd_sc_hd__a221o_1
X_4706_ _4826_/A _4735_/B VGND VGND VPWR VPWR _4832_/D sky130_fd_sc_hd__nand2_1
X_5686_ _5686_/A _5686_/B _5688_/C VGND VGND VPWR VPWR _5686_/X sky130_fd_sc_hd__and3_4
X_4637_ _4637_/A _4637_/B _4637_/C _4637_/D VGND VGND VPWR VPWR _4637_/Y sky130_fd_sc_hd__nor4_1
XFILLER_190_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold620 hold620/A VGND VGND VPWR VPWR hold620/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold631 hold631/A VGND VGND VPWR VPWR hold631/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4568_ _4568_/A _4881_/B VGND VGND VPWR VPWR _4568_/Y sky130_fd_sc_hd__nand2_1
Xhold642 hold642/A VGND VGND VPWR VPWR hold642/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold653 hold653/A VGND VGND VPWR VPWR hold653/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap361 hold54/X VGND VGND VPWR VPWR _3540_/A sky130_fd_sc_hd__buf_12
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold664 hold664/A VGND VGND VPWR VPWR hold664/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3519_ _6552_/Q _4092_/A _5169_/A _6773_/Q _3518_/X VGND VGND VPWR VPWR _3529_/A
+ sky130_fd_sc_hd__a221o_2
X_6307_ _6592_/Q _5985_/X _5999_/X _6551_/Q VGND VGND VPWR VPWR _6307_/X sky130_fd_sc_hd__a22o_1
Xhold675 _4245_/X VGND VGND VPWR VPWR _6671_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4499_ _4682_/A _4693_/B _4447_/B VGND VGND VPWR VPWR _4499_/Y sky130_fd_sc_hd__a21oi_2
Xhold686 hold686/A VGND VGND VPWR VPWR hold686/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold697 hold697/A VGND VGND VPWR VPWR hold697/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6238_ _6238_/A _6238_/B _6238_/C _6238_/D VGND VGND VPWR VPWR _6239_/D sky130_fd_sc_hd__nor4_2
Xhold2010 hold120/X VGND VGND VPWR VPWR _4050_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2021 _6642_/Q VGND VGND VPWR VPWR hold597/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2032 _4075_/X VGND VGND VPWR VPWR _6533_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2043 _6838_/Q VGND VGND VPWR VPWR hold774/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2054 _7223_/A VGND VGND VPWR VPWR hold670/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6169_ _6899_/Q _5989_/X _5994_/X _7067_/Q _6168_/X VGND VGND VPWR VPWR _6169_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2065 _6732_/Q VGND VGND VPWR VPWR hold781/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1320 _6868_/Q VGND VGND VPWR VPWR hold342/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1331 hold343/X VGND VGND VPWR VPWR _5289_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2076 hold712/X VGND VGND VPWR VPWR _5583_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_27_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2087 _6933_/Q VGND VGND VPWR VPWR hold784/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1342 _6858_/Q VGND VGND VPWR VPWR hold551/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2098 _5498_/X VGND VGND VPWR VPWR _7061_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1353 _6841_/Q VGND VGND VPWR VPWR hold156/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1364 hold2/X VGND VGND VPWR VPWR _5320_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1375 _6807_/Q VGND VGND VPWR VPWR hold309/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1386 hold323/X VGND VGND VPWR VPWR _4198_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1397 hold160/X VGND VGND VPWR VPWR _4029_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_43_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _6941_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_58_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7077_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3870_ _3870_/A _3870_/B VGND VGND VPWR VPWR _3870_/X sky130_fd_sc_hd__and2_1
XFILLER_71_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5540_ _5540_/A0 _5585_/A1 _5541_/S VGND VGND VPWR VPWR _7099_/D sky130_fd_sc_hd__mux2_1
XFILLER_192_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5471_ hold639/X _5561_/A1 _5478_/S VGND VGND VPWR VPWR _7037_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7210_ _7210_/A VGND VGND VPWR VPWR _7210_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_145_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4422_ _4575_/C _4495_/B VGND VGND VPWR VPWR _4610_/A sky130_fd_sc_hd__nor2_2
XFILLER_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7141_ _7203_/CLK _7141_/D _6409_/A VGND VGND VPWR VPWR _7141_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_132_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4353_ _4447_/B _4682_/A _4365_/B VGND VGND VPWR VPWR _4360_/A sky130_fd_sc_hd__nand3_2
XFILLER_125_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout407 _5570_/A1 VGND VGND VPWR VPWR _5552_/A1 sky130_fd_sc_hd__buf_8
X_3304_ hold52/X hold25/X VGND VGND VPWR VPWR _3686_/B sky130_fd_sc_hd__nand2b_4
XFILLER_59_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout418 _5686_/A VGND VGND VPWR VPWR _5689_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_140_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7072_ _7126_/CLK _7072_/D fanout475/X VGND VGND VPWR VPWR _7072_/Q sky130_fd_sc_hd__dfrtp_4
X_4284_ _4284_/A0 _5249_/A1 _4285_/S VGND VGND VPWR VPWR _4284_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6023_ _6877_/Q _6004_/X _6007_/X _6845_/Q VGND VGND VPWR VPWR _6023_/X sky130_fd_sc_hd__a22o_1
X_3235_ _6880_/Q VGND VGND VPWR VPWR _3235_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6925_ _6983_/CLK _6925_/D fanout459/X VGND VGND VPWR VPWR _6925_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_120_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6856_ _7124_/CLK _6856_/D fanout458/X VGND VGND VPWR VPWR _6856_/Q sky130_fd_sc_hd__dfrtp_4
X_5807_ _6866_/Q _5673_/X _5805_/X _5806_/X VGND VGND VPWR VPWR _5807_/X sky130_fd_sc_hd__a211o_1
XFILLER_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6787_ _6788_/CLK _6787_/D _3959_/B VGND VGND VPWR VPWR _6787_/Q sky130_fd_sc_hd__dfrtp_4
X_3999_ hold394/X _5559_/A1 _3999_/S VGND VGND VPWR VPWR _6478_/D sky130_fd_sc_hd__mux2_1
XFILLER_109_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5738_ _6951_/Q _5672_/X _5679_/X _6903_/Q _5737_/X VGND VGND VPWR VPWR _5738_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5669_ _5686_/A _5689_/B _5687_/C VGND VGND VPWR VPWR _5669_/X sky130_fd_sc_hd__and3_4
XFILLER_129_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold450 hold450/A VGND VGND VPWR VPWR hold450/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold461 hold461/A VGND VGND VPWR VPWR hold461/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold472 hold472/A VGND VGND VPWR VPWR hold472/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold483 hold483/A VGND VGND VPWR VPWR hold483/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold494 hold494/A VGND VGND VPWR VPWR hold494/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1150 hold385/X VGND VGND VPWR VPWR _5504_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1161 _6898_/Q VGND VGND VPWR VPWR hold482/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_100_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1172 _5305_/X VGND VGND VPWR VPWR _6890_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1183 hold472/X VGND VGND VPWR VPWR _5467_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1194 hold494/X VGND VGND VPWR VPWR _5485_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4971_ _4971_/A _4981_/B VGND VGND VPWR VPWR _4971_/Y sky130_fd_sc_hd__nand2_1
X_6710_ _6711_/CLK _6710_/D fanout465/X VGND VGND VPWR VPWR _6710_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3922_ _4222_/B _3922_/B VGND VGND VPWR VPWR _3922_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6641_ _6793_/CLK _6641_/D fanout442/X VGND VGND VPWR VPWR _6641_/Q sky130_fd_sc_hd__dfstp_2
X_3853_ _3853_/A0 _3880_/A0 _3853_/S VGND VGND VPWR VPWR _6457_/D sky130_fd_sc_hd__mux2_1
X_3784_ _7029_/Q _5461_/A _4009_/A _6487_/Q VGND VGND VPWR VPWR _3784_/X sky130_fd_sc_hd__a22o_1
X_6572_ _6711_/CLK _6572_/D fanout465/X VGND VGND VPWR VPWR _6572_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_118_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5523_ _5523_/A0 _5577_/A1 _5523_/S VGND VGND VPWR VPWR _7084_/D sky130_fd_sc_hd__mux2_1
XFILLER_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5454_ _5454_/A0 _5571_/A1 _5460_/S VGND VGND VPWR VPWR _5454_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4405_ _3890_/Y _4492_/B _4356_/B _4341_/X VGND VGND VPWR VPWR _4477_/B sky130_fd_sc_hd__a31oi_4
XFILLER_132_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5385_ _5385_/A0 _5583_/A1 _5388_/S VGND VGND VPWR VPWR _5385_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7124_ _7124_/CLK _7124_/D fanout459/X VGND VGND VPWR VPWR _7124_/Q sky130_fd_sc_hd__dfrtp_4
X_4336_ _4336_/A0 _5193_/A1 _4339_/S VGND VGND VPWR VPWR _6758_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7055_ _7117_/CLK _7055_/D fanout457/X VGND VGND VPWR VPWR _7055_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4267_ _4267_/A0 _4339_/A1 _4267_/S VGND VGND VPWR VPWR _6701_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6006_ _5637_/A _6015_/B _6017_/A _5985_/X _6005_/X VGND VGND VPWR VPWR _6010_/B
+ sky130_fd_sc_hd__a311o_1
X_3218_ _7008_/Q VGND VGND VPWR VPWR _3218_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4198_ _4198_/A0 _5303_/A1 _4199_/S VGND VGND VPWR VPWR _4198_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6908_ _7124_/CLK _6908_/D fanout459/X VGND VGND VPWR VPWR _6908_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6839_ _7121_/CLK _6839_/D fanout473/X VGND VGND VPWR VPWR _6839_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold280 hold280/A VGND VGND VPWR VPWR hold280/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold291 hold291/A VGND VGND VPWR VPWR hold291/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_120 _5581_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 hold2/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_142 _6660_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_153 _5469_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_164 _5689_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_175 _6625_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_186 _7233_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_197 _5308_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5170_ _5170_/A0 _5221_/A1 _5174_/S VGND VGND VPWR VPWR _5170_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4121_ _4121_/A0 _5538_/A1 _4121_/S VGND VGND VPWR VPWR _4121_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1908 _6527_/Q VGND VGND VPWR VPWR hold287/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1919 hold735/X VGND VGND VPWR VPWR _4129_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4052_ _4052_/A0 _5556_/A1 _4055_/S VGND VGND VPWR VPWR _4052_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput4 mask_rev_in[0] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4954_ _4954_/A _5117_/B _5038_/B _4954_/D VGND VGND VPWR VPWR _4962_/B sky130_fd_sc_hd__and4_1
XFILLER_189_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3905_ _6656_/Q _3904_/A _3904_/B _3903_/Y VGND VGND VPWR VPWR _6654_/D sky130_fd_sc_hd__a31o_1
X_4885_ _4391_/Y _4584_/Y _4683_/A VGND VGND VPWR VPWR _4885_/X sky130_fd_sc_hd__a21o_1
XFILLER_193_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6624_ _6742_/CLK _6624_/D fanout440/X VGND VGND VPWR VPWR _6624_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3836_ _6462_/Q _6461_/Q _6460_/Q _6463_/Q VGND VGND VPWR VPWR _3836_/X sky130_fd_sc_hd__a31o_1
XFILLER_137_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3767_ _6803_/Q _3303_/X _5229_/B _5452_/A _7021_/Q VGND VGND VPWR VPWR _3767_/X
+ sky130_fd_sc_hd__a32o_1
X_6555_ _6568_/CLK _6555_/D VGND VGND VPWR VPWR _6555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5506_ _5506_/A _5569_/B VGND VGND VPWR VPWR _5514_/S sky130_fd_sc_hd__and2_4
X_6486_ _6809_/CLK _6486_/D fanout451/X VGND VGND VPWR VPWR _6486_/Q sky130_fd_sc_hd__dfstp_4
X_3698_ _6743_/Q _4316_/A _4122_/A _6575_/Q _3697_/X VGND VGND VPWR VPWR _3703_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5437_ _5437_/A0 _5518_/A1 _5442_/S VGND VGND VPWR VPWR _7007_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput330 hold849/X VGND VGND VPWR VPWR hold192/A sky130_fd_sc_hd__buf_6
XFILLER_160_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput341 hold861/X VGND VGND VPWR VPWR hold286/A sky130_fd_sc_hd__buf_6
XFILLER_133_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5368_ hold922/X hold20/X _5370_/S VGND VGND VPWR VPWR _5368_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7107_ _7130_/CLK hold85/X fanout460/X VGND VGND VPWR VPWR _7107_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4319_ hold314/X _4337_/A1 _4321_/S VGND VGND VPWR VPWR _6744_/D sky130_fd_sc_hd__mux2_1
X_5299_ _5299_/A _5551_/B VGND VGND VPWR VPWR _5307_/S sky130_fd_sc_hd__and2_4
XFILLER_87_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7038_ _7136_/CLK _7038_/D fanout476/X VGND VGND VPWR VPWR _7038_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_101_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4670_ _4637_/A _4637_/B _4667_/X _4669_/X _4387_/Y VGND VGND VPWR VPWR _4703_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_187_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3621_ _6786_/Q _5178_/A _4206_/A _6646_/Q VGND VGND VPWR VPWR _3621_/X sky130_fd_sc_hd__a22o_2
XFILLER_186_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3552_ _6953_/Q _5371_/A _3427_/Y _6793_/Q _3551_/X VGND VGND VPWR VPWR _3556_/C
+ sky130_fd_sc_hd__a221o_2
X_6340_ _6529_/Q _6339_/B _6339_/X VGND VGND VPWR VPWR _6340_/X sky130_fd_sc_hd__o21ba_1
XFILLER_6_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6271_ _6586_/Q _5989_/X _5999_/X _6550_/Q VGND VGND VPWR VPWR _6271_/X sky130_fd_sc_hd__a22o_1
X_3483_ _3553_/A _3516_/B VGND VGND VPWR VPWR _4316_/A sky130_fd_sc_hd__nor2_8
XFILLER_115_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5222_ _5222_/A _5226_/B _5229_/C VGND VGND VPWR VPWR _5225_/S sky130_fd_sc_hd__and3_4
XFILLER_170_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2406 _7089_/Q VGND VGND VPWR VPWR hold739/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2417 _6775_/Q VGND VGND VPWR VPWR _3739_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5153_ _5137_/X _5152_/Y _5147_/X _5146_/X VGND VGND VPWR VPWR _6767_/D sky130_fd_sc_hd__a211o_1
XFILLER_97_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2428 _6679_/Q VGND VGND VPWR VPWR _3918_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2439 _7175_/Q VGND VGND VPWR VPWR _6116_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1705 hold177/X VGND VGND VPWR VPWR _5238_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1716 _4253_/X VGND VGND VPWR VPWR _6689_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_4104_ _3462_/Y hold836/A _4106_/S VGND VGND VPWR VPWR _6558_/D sky130_fd_sc_hd__mux2_1
Xhold1727 _6644_/Q VGND VGND VPWR VPWR hold642/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5084_ _4698_/Y _5011_/X _5022_/C _5081_/Y VGND VGND VPWR VPWR _5165_/B sky130_fd_sc_hd__o211a_1
Xhold1738 hold131/X VGND VGND VPWR VPWR _5502_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1749 hold852/X VGND VGND VPWR VPWR hold196/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_2_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4035_ hold540/A _5581_/A1 _4056_/C VGND VGND VPWR VPWR _4035_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5986_ _6019_/B _6018_/B _6016_/C VGND VGND VPWR VPWR _5986_/X sky130_fd_sc_hd__and3_4
XFILLER_52_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4937_ _4729_/A _4688_/B _4935_/X _4936_/Y _4539_/Y VGND VGND VPWR VPWR _4954_/A
+ sky130_fd_sc_hd__o221a_1
XANTENNA_20 _3658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_31 _5664_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4868_ _4638_/Y _4712_/Y _4922_/C _4867_/X _5063_/B VGND VGND VPWR VPWR _4870_/C
+ sky130_fd_sc_hd__o2111a_1
XANTENNA_42 _5971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 _6013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6607_ _6711_/CLK _6607_/D _6433_/A VGND VGND VPWR VPWR _6607_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_64 _7000_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_75 _7141_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3819_ _6654_/Q _3816_/Y _3904_/B _3840_/B VGND VGND VPWR VPWR _3846_/S sky130_fd_sc_hd__o31a_4
XFILLER_165_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_86 _3971_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4799_ _4729_/A _4714_/Y _4779_/X _4798_/X _4539_/Y VGND VGND VPWR VPWR _4800_/D
+ sky130_fd_sc_hd__o2111a_1
XANTENNA_97 input95/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6538_ _6757_/CLK _6538_/D fanout446/X VGND VGND VPWR VPWR _6538_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6469_ _3958_/A1 _6469_/D _6419_/X VGND VGND VPWR VPWR _6469_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_121_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput171 _3972_/X VGND VGND VPWR VPWR debug_in sky130_fd_sc_hd__buf_12
Xoutput182 _5763_/A VGND VGND VPWR VPWR mgmt_gpio_oeb[16] sky130_fd_sc_hd__buf_12
Xoutput193 _3213_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[26] sky130_fd_sc_hd__buf_12
XFILLER_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5840_ _6884_/Q _5667_/X _5682_/X _7044_/Q VGND VGND VPWR VPWR _5840_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5771_ _3239_/Y _5707_/B _5760_/Y _5770_/Y _6490_/Q VGND VGND VPWR VPWR _5771_/X
+ sky130_fd_sc_hd__a221o_1
X_4722_ _5001_/A _4732_/B _4722_/C VGND VGND VPWR VPWR _4722_/X sky130_fd_sc_hd__and3_1
XFILLER_148_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4653_ _4682_/A _4693_/B _4504_/X VGND VGND VPWR VPWR _4838_/B sky130_fd_sc_hd__a21o_1
Xinput40 mgmt_gpio_in[13] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__clkbuf_2
X_3604_ _3604_/A _3604_/B _3604_/C _3604_/D VGND VGND VPWR VPWR _3615_/B sky130_fd_sc_hd__nor4_1
Xinput51 mgmt_gpio_in[23] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__clkbuf_4
Xinput62 mgmt_gpio_in[33] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__buf_2
Xhold802 hold802/A VGND VGND VPWR VPWR hold802/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4584_ _4584_/A _4710_/A VGND VGND VPWR VPWR _4584_/Y sky130_fd_sc_hd__nand2_2
Xinput73 pad_flash_io0_di VGND VGND VPWR VPWR _3965_/B sky130_fd_sc_hd__clkbuf_2
Xhold813 hold813/A VGND VGND VPWR VPWR hold813/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput84 spimemio_flash_csb VGND VGND VPWR VPWR input84/X sky130_fd_sc_hd__clkbuf_4
Xinput95 usr1_vcc_pwrgood VGND VGND VPWR VPWR input95/X sky130_fd_sc_hd__clkbuf_4
X_6323_ _6539_/Q _5983_/X _6005_/X _6696_/Q VGND VGND VPWR VPWR _6323_/X sky130_fd_sc_hd__a22o_1
Xhold824 hold824/A VGND VGND VPWR VPWR hold824/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3535_ _3535_/A _3550_/B VGND VGND VPWR VPWR _4170_/A sky130_fd_sc_hd__nor2_8
Xhold835 hold835/A VGND VGND VPWR VPWR hold835/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold846 hold846/A VGND VGND VPWR VPWR hold846/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold857 hold857/A VGND VGND VPWR VPWR hold857/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold868 hold868/A VGND VGND VPWR VPWR hold868/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3466_ input7/X _3315_/Y _4152_/A _6603_/Q VGND VGND VPWR VPWR _3466_/X sky130_fd_sc_hd__a22o_1
X_6254_ _6610_/Q _5976_/B _5993_/X _6620_/Q _6253_/X VGND VGND VPWR VPWR _6255_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_107_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold879 _5584_/X VGND VGND VPWR VPWR _7138_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_170_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2203 hold442/X VGND VGND VPWR VPWR _4205_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5205_ _5205_/A0 _5518_/A1 _5206_/S VGND VGND VPWR VPWR _6806_/D sky130_fd_sc_hd__mux2_1
XFILLER_103_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2214 hold728/X VGND VGND VPWR VPWR _5208_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_3397_ _6995_/Q _5416_/A _3357_/Y _6485_/Q _3396_/X VGND VGND VPWR VPWR _3397_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6185_ _6963_/Q _5992_/X _6012_/X _7003_/Q VGND VGND VPWR VPWR _6185_/X sky130_fd_sc_hd__a22o_1
Xhold2225 _5177_/X VGND VGND VPWR VPWR _6783_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2236 _5419_/X VGND VGND VPWR VPWR _6991_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2247 _6595_/Q VGND VGND VPWR VPWR hold733/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1502 _6864_/Q VGND VGND VPWR VPWR _5276_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2258 _6724_/Q VGND VGND VPWR VPWR hold591/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1513 _7076_/Q VGND VGND VPWR VPWR hold513/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5136_ _5136_/A _5136_/B _5136_/C VGND VGND VPWR VPWR _5137_/C sky130_fd_sc_hd__and3_1
Xhold1524 _6541_/Q VGND VGND VPWR VPWR hold838/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_123_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2269 _4038_/X VGND VGND VPWR VPWR _6504_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1535 _6542_/Q VGND VGND VPWR VPWR hold818/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1546 hold850/X VGND VGND VPWR VPWR hold277/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1557 hold832/X VGND VGND VPWR VPWR hold250/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5067_ _5067_/A _5067_/B VGND VGND VPWR VPWR _5102_/C sky130_fd_sc_hd__and2_1
Xhold1568 _5505_/X VGND VGND VPWR VPWR _7068_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1579 hold109/X VGND VGND VPWR VPWR _5277_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4018_ _4050_/A0 _5581_/A1 _4047_/C VGND VGND VPWR VPWR _4018_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5969_ _5969_/A1 _3924_/Y _5647_/Y VGND VGND VPWR VPWR _5969_/X sky130_fd_sc_hd__o21ba_1
XFILLER_166_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold109 hold109/A VGND VGND VPWR VPWR hold109/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3320_ _3322_/B _3425_/A VGND VGND VPWR VPWR _3470_/A sky130_fd_sc_hd__nand2_8
XFILLER_125_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3251_ hold22/X _3996_/S VGND VGND VPWR VPWR hold23/A sky130_fd_sc_hd__nand2b_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3182_ _6460_/Q VGND VGND VPWR VPWR _3182_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6941_ _6941_/CLK _6941_/D fanout460/X VGND VGND VPWR VPWR _6941_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_81_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6872_ _7140_/CLK _6872_/D fanout471/X VGND VGND VPWR VPWR _6872_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5823_ _6979_/Q _5660_/X _5669_/X _7051_/Q VGND VGND VPWR VPWR _5823_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5754_ _7016_/Q _5664_/X _5686_/X _7008_/Q VGND VGND VPWR VPWR _5754_/X sky130_fd_sc_hd__a22o_1
X_4705_ _5009_/B _5150_/C VGND VGND VPWR VPWR _4705_/Y sky130_fd_sc_hd__nand2_1
XFILLER_148_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5685_ _5686_/A _5686_/B _5689_/C VGND VGND VPWR VPWR _5685_/X sky130_fd_sc_hd__and3_4
XFILLER_190_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4636_ _4663_/D _4840_/A _4498_/X _3969_/A VGND VGND VPWR VPWR _4636_/X sky130_fd_sc_hd__a31o_2
XFILLER_118_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold610 hold610/A VGND VGND VPWR VPWR hold610/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold621 hold621/A VGND VGND VPWR VPWR hold621/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4567_ _4980_/A _4693_/B VGND VGND VPWR VPWR _5100_/C sky130_fd_sc_hd__nand2_2
Xhold632 hold632/A VGND VGND VPWR VPWR hold632/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap351 _4239_/S VGND VGND VPWR VPWR _5236_/C sky130_fd_sc_hd__buf_8
Xhold643 hold643/A VGND VGND VPWR VPWR hold643/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap362 _3501_/A VGND VGND VPWR VPWR _3349_/A sky130_fd_sc_hd__buf_12
Xhold654 hold654/A VGND VGND VPWR VPWR hold654/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6306_ _6730_/Q _5987_/X _6004_/X _6577_/Q _6305_/X VGND VGND VPWR VPWR _6306_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3518_ _6865_/Q _5272_/A _3357_/Y _6483_/Q VGND VGND VPWR VPWR _3518_/X sky130_fd_sc_hd__a22o_1
Xhold665 hold665/A VGND VGND VPWR VPWR hold665/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold676 hold676/A VGND VGND VPWR VPWR hold676/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4498_ _4637_/B _4498_/B VGND VGND VPWR VPWR _4498_/X sky130_fd_sc_hd__and2_1
Xhold687 hold687/A VGND VGND VPWR VPWR _6803_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold698 hold698/A VGND VGND VPWR VPWR hold698/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6237_ _6584_/Q _5989_/X _6013_/X _6624_/Q _6236_/X VGND VGND VPWR VPWR _6238_/D
+ sky130_fd_sc_hd__a221o_1
X_3449_ _3449_/A _3449_/B _3449_/C VGND VGND VPWR VPWR _3461_/A sky130_fd_sc_hd__nor3_1
Xhold2000 hold536/X VGND VGND VPWR VPWR _5556_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2011 _7105_/Q VGND VGND VPWR VPWR hold535/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2022 hold597/X VGND VGND VPWR VPWR _4204_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2033 _7045_/Q VGND VGND VPWR VPWR hold788/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2044 _6734_/Q VGND VGND VPWR VPWR hold558/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _7123_/Q _5978_/X _6016_/X _7043_/Q VGND VGND VPWR VPWR _6168_/X sky130_fd_sc_hd__a22o_1
Xhold2055 hold670/X VGND VGND VPWR VPWR _4243_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1310 _6528_/Q VGND VGND VPWR VPWR hold262/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2066 hold781/X VGND VGND VPWR VPWR _4305_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1321 hold342/X VGND VGND VPWR VPWR _5280_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2077 _6925_/Q VGND VGND VPWR VPWR hold669/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1332 _5289_/X VGND VGND VPWR VPWR _6876_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2088 _5354_/X VGND VGND VPWR VPWR _6933_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1343 hold551/X VGND VGND VPWR VPWR _5269_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5119_ _5119_/A _5119_/B _5119_/C VGND VGND VPWR VPWR _6766_/D sky130_fd_sc_hd__nand3_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1354 hold156/X VGND VGND VPWR VPWR _5250_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2099 _7117_/Q VGND VGND VPWR VPWR hold672/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_27_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6099_ _7024_/Q _5971_/X _6007_/X _6848_/Q _6098_/X VGND VGND VPWR VPWR _6102_/B
+ sky130_fd_sc_hd__a221o_1
Xhold1365 _4080_/X VGND VGND VPWR VPWR hold445/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1376 hold309/X VGND VGND VPWR VPWR _5206_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1387 _4198_/X VGND VGND VPWR VPWR _6637_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1398 _4029_/X VGND VGND VPWR VPWR hold161/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5470_ _5470_/A _5569_/B VGND VGND VPWR VPWR _5478_/S sky130_fd_sc_hd__and2_4
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4421_ _4955_/A _4955_/B _4477_/C VGND VGND VPWR VPWR _5033_/A sky130_fd_sc_hd__and3_4
XFILLER_172_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7140_ _7140_/CLK hold34/X fanout469/X VGND VGND VPWR VPWR _7140_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_113_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4352_ _4682_/A _4365_/B VGND VGND VPWR VPWR _4420_/A sky130_fd_sc_hd__nand2_1
XFILLER_125_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout408 _5561_/A1 VGND VGND VPWR VPWR _5570_/A1 sky130_fd_sc_hd__buf_6
X_3303_ hold52/X hold25/X VGND VGND VPWR VPWR _3303_/X sky130_fd_sc_hd__and2b_4
XFILLER_141_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7071_ _7103_/CLK _7071_/D fanout472/X VGND VGND VPWR VPWR _7071_/Q sky130_fd_sc_hd__dfrtp_4
X_4283_ _4283_/A0 _5581_/A1 _4285_/S VGND VGND VPWR VPWR _4283_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout419 _5872_/B VGND VGND VPWR VPWR _5686_/A sky130_fd_sc_hd__buf_6
XFILLER_98_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6022_ _6853_/Q _5983_/X _5995_/X _6917_/Q _6021_/X VGND VGND VPWR VPWR _6039_/A
+ sky130_fd_sc_hd__a221o_1
X_3234_ _6888_/Q VGND VGND VPWR VPWR _3234_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6924_ _7124_/CLK _6924_/D fanout459/X VGND VGND VPWR VPWR _6924_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6855_ _6941_/CLK _6855_/D fanout460/X VGND VGND VPWR VPWR _6855_/Q sky130_fd_sc_hd__dfrtp_4
X_5806_ _6978_/Q _5660_/X _5669_/X _7050_/Q VGND VGND VPWR VPWR _5806_/X sky130_fd_sc_hd__a22o_1
XFILLER_167_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6786_ _6788_/CLK _6786_/D _3959_/B VGND VGND VPWR VPWR _6786_/Q sky130_fd_sc_hd__dfstp_4
X_3998_ hold4/X hold967/X _6659_/Q VGND VGND VPWR VPWR _3998_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5737_ _6935_/Q _5659_/X _5687_/X _6919_/Q VGND VGND VPWR VPWR _5737_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5668_ _5689_/A _5684_/B _5687_/C VGND VGND VPWR VPWR _5668_/X sky130_fd_sc_hd__and3_4
XFILLER_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4619_ _4570_/C _4655_/A _4922_/A _4617_/X _4618_/Y VGND VGND VPWR VPWR _4622_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_191_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5599_ _7142_/Q _7143_/Q _7144_/Q _5599_/D VGND VGND VPWR VPWR _5601_/B sky130_fd_sc_hd__nand4_2
XFILLER_151_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold440 hold440/A VGND VGND VPWR VPWR hold440/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold451 hold451/A VGND VGND VPWR VPWR hold451/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold462 hold462/A VGND VGND VPWR VPWR hold462/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold473 hold473/A VGND VGND VPWR VPWR hold473/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold484 hold484/A VGND VGND VPWR VPWR hold484/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold495 hold495/A VGND VGND VPWR VPWR hold495/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1140 _4276_/X VGND VGND VPWR VPWR _6708_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_100_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1151 _5504_/X VGND VGND VPWR VPWR _7067_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1162 hold482/X VGND VGND VPWR VPWR _5314_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1173 _6971_/Q VGND VGND VPWR VPWR hold391/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1184 _6666_/Q VGND VGND VPWR VPWR hold418/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1195 _7082_/Q VGND VGND VPWR VPWR hold480/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4970_ _4598_/A _5001_/B _4883_/X VGND VGND VPWR VPWR _5069_/A sky130_fd_sc_hd__a21boi_1
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3921_ _3921_/A _3921_/B VGND VGND VPWR VPWR _3922_/B sky130_fd_sc_hd__nand2_2
XFILLER_177_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6640_ _6793_/CLK _6640_/D fanout443/X VGND VGND VPWR VPWR _6640_/Q sky130_fd_sc_hd__dfrtp_4
X_3852_ _6468_/Q _3852_/B VGND VGND VPWR VPWR _3853_/S sky130_fd_sc_hd__nor2_2
XFILLER_20_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6571_ _6731_/CLK _6571_/D _6409_/A VGND VGND VPWR VPWR _6571_/Q sky130_fd_sc_hd__dfstp_2
X_3783_ _3783_/A _3783_/B _3783_/C _3783_/D VGND VGND VPWR VPWR _3802_/B sky130_fd_sc_hd__nor4_1
X_5522_ _5522_/A0 _5576_/A1 _5523_/S VGND VGND VPWR VPWR _5522_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5453_ _5453_/A0 _5552_/A1 _5460_/S VGND VGND VPWR VPWR _5453_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4404_ _4492_/B _4356_/B _4650_/B VGND VGND VPWR VPWR _4477_/A sky130_fd_sc_hd__a21o_4
Xclkbuf_leaf_42_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7065_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_145_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5384_ _5384_/A0 _5582_/A1 _5388_/S VGND VGND VPWR VPWR _5384_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7123_ _7123_/CLK _7123_/D fanout479/X VGND VGND VPWR VPWR _7123_/Q sky130_fd_sc_hd__dfrtp_4
X_4335_ _4335_/A0 _5221_/A1 _4339_/S VGND VGND VPWR VPWR _6757_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7054_ _7126_/CLK _7054_/D fanout474/X VGND VGND VPWR VPWR _7054_/Q sky130_fd_sc_hd__dfstp_2
X_4266_ _4266_/A0 _5195_/A1 _4267_/S VGND VGND VPWR VPWR _6700_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_57_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7125_/CLK sky130_fd_sc_hd__clkbuf_16
X_6005_ _6017_/A _6017_/B _6007_/C VGND VGND VPWR VPWR _6005_/X sky130_fd_sc_hd__and3_4
X_3217_ _7016_/Q VGND VGND VPWR VPWR _3217_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4197_ _4197_/A0 _4337_/A1 _4199_/S VGND VGND VPWR VPWR _4197_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6907_ _7140_/CLK _6907_/D fanout471/X VGND VGND VPWR VPWR _6907_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_168_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6838_ _7134_/CLK _6838_/D fanout476/X VGND VGND VPWR VPWR _6838_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_50_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6769_ _6809_/CLK _6769_/D fanout444/X VGND VGND VPWR VPWR _6769_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_183_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold270 hold270/A VGND VGND VPWR VPWR hold270/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold281 hold281/A VGND VGND VPWR VPWR hold859/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold292 hold292/A VGND VGND VPWR VPWR hold292/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_110 _5842_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_121 _5221_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_132 hold20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_143 _5569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_154 _5577_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 _5971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_176 _7102_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_187 _3974_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_198 _5673_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4120_ _4120_/A0 _5249_/A1 _4121_/S VGND VGND VPWR VPWR _4120_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1909 hold287/X VGND VGND VPWR VPWR _4068_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4051_ _4051_/A0 _5555_/A1 _4055_/S VGND VGND VPWR VPWR _4051_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput5 mask_rev_in[10] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4953_ _4368_/B _4407_/Y _4938_/X _4786_/X VGND VGND VPWR VPWR _4954_/D sky130_fd_sc_hd__o31a_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3904_ _3904_/A _3904_/B VGND VGND VPWR VPWR _3904_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4884_ _4658_/B _4564_/Y _4965_/C _5102_/B _4883_/X VGND VGND VPWR VPWR _4892_/A
+ sky130_fd_sc_hd__o2111a_1
XFILLER_178_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6623_ _6648_/CLK _6623_/D fanout449/X VGND VGND VPWR VPWR _6623_/Q sky130_fd_sc_hd__dfrtp_4
X_3835_ _3831_/B _3834_/X _3835_/S VGND VGND VPWR VPWR _6464_/D sky130_fd_sc_hd__mux2_1
XFILLER_165_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6554_ _6568_/CLK _6554_/D VGND VGND VPWR VPWR _6554_/Q sky130_fd_sc_hd__dfxtp_1
X_3766_ _7117_/Q hold67/A _4322_/A _6747_/Q _3765_/X VGND VGND VPWR VPWR _3769_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5505_ _5505_/A0 _5559_/A1 _5505_/S VGND VGND VPWR VPWR _5505_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6485_ _6809_/CLK _6485_/D fanout451/X VGND VGND VPWR VPWR _6485_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_173_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3697_ _7086_/Q _5524_/A _5470_/A _7038_/Q VGND VGND VPWR VPWR _3697_/X sky130_fd_sc_hd__a22o_2
XFILLER_118_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5436_ hold141/X hold135/X _5442_/S VGND VGND VPWR VPWR _5436_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput320 hold843/X VGND VGND VPWR VPWR hold268/A sky130_fd_sc_hd__buf_6
Xoutput331 hold845/X VGND VGND VPWR VPWR hold189/A sky130_fd_sc_hd__buf_6
Xoutput342 hold863/X VGND VGND VPWR VPWR hold289/A sky130_fd_sc_hd__buf_6
XFILLER_133_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5367_ _5367_/A0 _5538_/A1 _5370_/S VGND VGND VPWR VPWR _5367_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7106_ _7140_/CLK _7106_/D fanout470/X VGND VGND VPWR VPWR hold49/A sky130_fd_sc_hd__dfrtp_2
X_4318_ _4318_/A0 _5193_/A1 _4321_/S VGND VGND VPWR VPWR _6743_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5298_ _5298_/A0 _5559_/A1 _5298_/S VGND VGND VPWR VPWR _5298_/X sky130_fd_sc_hd__mux2_1
X_7037_ _7065_/CLK _7037_/D fanout460/X VGND VGND VPWR VPWR _7037_/Q sky130_fd_sc_hd__dfstp_2
X_4249_ _4249_/A0 hold6/X _4249_/S VGND VGND VPWR VPWR _4249_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3620_ _6911_/Q _5326_/A _4194_/A _6636_/Q _3619_/X VGND VGND VPWR VPWR _3627_/A
+ sky130_fd_sc_hd__a221o_1
X_3551_ _6454_/Q _3977_/A _4286_/A _6721_/Q VGND VGND VPWR VPWR _3551_/X sky130_fd_sc_hd__a22o_1
XFILLER_155_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6270_ _6636_/Q _5994_/X _5996_/X _6651_/Q _6269_/X VGND VGND VPWR VPWR _6270_/X
+ sky130_fd_sc_hd__a221o_1
X_3482_ _3553_/A _3648_/A VGND VGND VPWR VPWR _4188_/A sky130_fd_sc_hd__nor2_8
XFILLER_170_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5221_ _5221_/A0 _5221_/A1 _5221_/S VGND VGND VPWR VPWR _5221_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2407 hold739/X VGND VGND VPWR VPWR _5529_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2418 _3739_/X VGND VGND VPWR VPWR _6775_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5152_ _5152_/A _5152_/B VGND VGND VPWR VPWR _5152_/Y sky130_fd_sc_hd__nand2_1
Xhold2429 _6677_/Q VGND VGND VPWR VPWR _6683_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_4103_ _4112_/A0 hold858/A _4106_/S VGND VGND VPWR VPWR _6557_/D sky130_fd_sc_hd__mux2_1
Xhold1706 _6872_/Q VGND VGND VPWR VPWR hold451/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1717 _6739_/Q VGND VGND VPWR VPWR hold183/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1728 hold642/X VGND VGND VPWR VPWR _4207_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5083_ _5083_/A _5083_/B _5083_/C _5083_/D VGND VGND VPWR VPWR _5139_/C sky130_fd_sc_hd__and4_1
Xhold1739 _5502_/X VGND VGND VPWR VPWR _7065_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_4034_ _4034_/A0 _4033_/X _4046_/S VGND VGND VPWR VPWR _4034_/X sky130_fd_sc_hd__mux2_1
XFILLER_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5985_ _6018_/B _6007_/C _6016_/C VGND VGND VPWR VPWR _5985_/X sky130_fd_sc_hd__and3_4
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4936_ _5150_/A _4936_/B VGND VGND VPWR VPWR _4936_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_10 _5335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_21 _3697_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4867_ _4590_/Y _4712_/Y _4866_/X _4616_/B VGND VGND VPWR VPWR _4867_/X sky130_fd_sc_hd__o211a_1
XANTENNA_32 _5669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 _5985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6606_ _6760_/CLK _6606_/D _6433_/A VGND VGND VPWR VPWR _6606_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA_54 _6014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3818_ _6445_/Q _3863_/A VGND VGND VPWR VPWR _3904_/B sky130_fd_sc_hd__and2_1
XFILLER_193_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_65 _7008_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4798_ _4947_/A _4714_/Y _4797_/X _4536_/Y VGND VGND VPWR VPWR _4798_/X sky130_fd_sc_hd__o211a_1
XFILLER_21_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_87 _3971_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_98 input97/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6537_ _6691_/CLK _6537_/D fanout443/X VGND VGND VPWR VPWR _6537_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_192_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3749_ _6609_/Q _4164_/A _3562_/Y input98/X _3748_/X VGND VGND VPWR VPWR _3750_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_134_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6468_ _3958_/A1 _6468_/D _6418_/X VGND VGND VPWR VPWR _6468_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_133_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5419_ _5419_/A0 _5572_/A1 _5424_/S VGND VGND VPWR VPWR _5419_/X sky130_fd_sc_hd__mux2_1
X_6399_ _6399_/A _6432_/B VGND VGND VPWR VPWR _6399_/X sky130_fd_sc_hd__and2_1
Xoutput172 _7206_/X VGND VGND VPWR VPWR irq[0] sky130_fd_sc_hd__buf_12
Xoutput183 _3222_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[17] sky130_fd_sc_hd__buf_12
Xoutput194 _3212_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[27] sky130_fd_sc_hd__buf_12
XFILLER_153_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5770_ _5770_/A _5770_/B _5770_/C _5770_/D VGND VGND VPWR VPWR _5770_/Y sky130_fd_sc_hd__nor4_2
XFILLER_15_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4721_ _4808_/A _4989_/B _4993_/B VGND VGND VPWR VPWR _5010_/A sky130_fd_sc_hd__nand3_1
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4652_ _4652_/A _4652_/B VGND VGND VPWR VPWR _4652_/Y sky130_fd_sc_hd__nand2_2
XFILLER_175_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3603_ _6745_/Q _4316_/A _3977_/A _6453_/Q _3602_/X VGND VGND VPWR VPWR _3604_/D
+ sky130_fd_sc_hd__a221o_1
Xinput30 mask_rev_in[4] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput41 mgmt_gpio_in[14] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput52 mgmt_gpio_in[24] VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4583_ _4658_/A _4583_/B VGND VGND VPWR VPWR _4993_/A sky130_fd_sc_hd__nor2_1
Xinput63 mgmt_gpio_in[34] VGND VGND VPWR VPWR _3971_/A sky130_fd_sc_hd__buf_6
Xhold803 hold803/A VGND VGND VPWR VPWR hold803/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput74 pad_flash_io1_di VGND VGND VPWR VPWR _3966_/B sky130_fd_sc_hd__buf_4
X_6322_ _6746_/Q _6014_/X _6320_/X _6321_/X VGND VGND VPWR VPWR _6327_/A sky130_fd_sc_hd__a211o_1
Xhold814 hold814/A VGND VGND VPWR VPWR hold814/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3534_ _6475_/Q _3339_/Y _4304_/A _6736_/Q _3532_/X VGND VGND VPWR VPWR _3543_/A
+ sky130_fd_sc_hd__a221o_2
Xhold825 hold825/A VGND VGND VPWR VPWR hold825/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput85 spimemio_flash_io0_do VGND VGND VPWR VPWR input85/X sky130_fd_sc_hd__clkbuf_4
Xinput96 usr1_vdd_pwrgood VGND VGND VPWR VPWR input96/X sky130_fd_sc_hd__buf_2
XFILLER_115_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold836 hold836/A VGND VGND VPWR VPWR hold836/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold847 hold847/A VGND VGND VPWR VPWR hold847/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold858 hold858/A VGND VGND VPWR VPWR hold858/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6253_ _6640_/Q _5986_/X _5998_/X _6580_/Q VGND VGND VPWR VPWR _6253_/X sky130_fd_sc_hd__a22o_1
Xhold869 hold869/A VGND VGND VPWR VPWR hold869/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3465_ _3550_/A _3533_/B VGND VGND VPWR VPWR _4152_/A sky130_fd_sc_hd__nor2_8
XFILLER_88_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5204_ _5204_/A0 hold135/X _5206_/S VGND VGND VPWR VPWR _5204_/X sky130_fd_sc_hd__mux2_1
Xhold2204 _6782_/Q VGND VGND VPWR VPWR hold794/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6184_ _6939_/Q _5980_/X _6008_/X _7107_/Q VGND VGND VPWR VPWR _6184_/X sky130_fd_sc_hd__a22o_1
Xhold2215 _6726_/Q VGND VGND VPWR VPWR hold466/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_3396_ _7139_/Q hold33/A _5533_/A _7099_/Q VGND VGND VPWR VPWR _3396_/X sky130_fd_sc_hd__a22o_2
Xhold2226 _6594_/Q VGND VGND VPWR VPWR hold798/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2237 _6475_/Q VGND VGND VPWR VPWR hold486/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1503 _5276_/X VGND VGND VPWR VPWR hold172/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5135_ _5135_/A _5135_/B _5135_/C _5135_/D VGND VGND VPWR VPWR _5135_/X sky130_fd_sc_hd__and4_1
Xhold2248 hold733/X VGND VGND VPWR VPWR _4148_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2259 _6483_/Q VGND VGND VPWR VPWR hold473/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1514 hold513/X VGND VGND VPWR VPWR _5514_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1525 hold838/X VGND VGND VPWR VPWR hold263/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1536 hold818/X VGND VGND VPWR VPWR hold204/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1547 _6566_/Q VGND VGND VPWR VPWR hold860/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1558 _6706_/Q VGND VGND VPWR VPWR hold118/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5066_ _5155_/B _5130_/B _5131_/A VGND VGND VPWR VPWR _5066_/X sky130_fd_sc_hd__and3_1
Xhold1569 _6615_/Q VGND VGND VPWR VPWR hold710/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4017_ _4017_/A0 _4016_/X _4029_/S VGND VGND VPWR VPWR _4017_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5968_ _6529_/Q _5678_/Y _5959_/X _5967_/X _6341_/S VGND VGND VPWR VPWR _5968_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4919_ _5115_/B _5047_/C _4919_/C VGND VGND VPWR VPWR _5126_/B sky130_fd_sc_hd__and3_1
X_5899_ _6536_/Q _5651_/X _5653_/X _6531_/Q VGND VGND VPWR VPWR _5899_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _3832_/A _6464_/Q _6657_/Q VGND VGND VPWR VPWR _3250_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3181_ _6468_/Q VGND VGND VPWR VPWR _3181_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6940_ _7084_/CLK _6940_/D fanout455/X VGND VGND VPWR VPWR _6940_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_66_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6871_ _7079_/CLK _6871_/D fanout470/X VGND VGND VPWR VPWR _6871_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5822_ _6963_/Q _5680_/X _5685_/X _7075_/Q VGND VGND VPWR VPWR _5822_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5753_ _6960_/Q _5680_/X _5685_/X _7072_/Q _5752_/X VGND VGND VPWR VPWR _5760_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_188_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4704_ _4704_/A _5124_/B _4704_/C _4704_/D VGND VGND VPWR VPWR _4704_/X sky130_fd_sc_hd__and4_1
XFILLER_148_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5684_ _5689_/A _5684_/B _5687_/C VGND VGND VPWR VPWR _5684_/X sky130_fd_sc_hd__and3b_4
XFILLER_147_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4635_ _4986_/C _4880_/B _4632_/X _4965_/B _4561_/X VGND VGND VPWR VPWR _4759_/B
+ sky130_fd_sc_hd__a41o_1
XFILLER_147_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold600 hold600/A VGND VGND VPWR VPWR hold600/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold611 hold611/A VGND VGND VPWR VPWR hold611/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4566_ _4981_/A _4693_/B VGND VGND VPWR VPWR _4616_/A sky130_fd_sc_hd__nand2_1
Xhold622 hold622/A VGND VGND VPWR VPWR hold622/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_851 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold633 hold633/A VGND VGND VPWR VPWR hold633/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold644 hold644/A VGND VGND VPWR VPWR hold644/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6305_ _6597_/Q _5991_/X _6005_/X _6695_/Q VGND VGND VPWR VPWR _6305_/X sky130_fd_sc_hd__a22o_1
Xmax_cap352 _3330_/Y VGND VGND VPWR VPWR _4047_/C sky130_fd_sc_hd__buf_12
XFILLER_150_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3517_ _3553_/B _3535_/A VGND VGND VPWR VPWR _5169_/A sky130_fd_sc_hd__nor2_8
Xmax_cap363 _3501_/A VGND VGND VPWR VPWR _3553_/A sky130_fd_sc_hd__buf_12
Xhold655 hold655/A VGND VGND VPWR VPWR hold655/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold666 hold666/A VGND VGND VPWR VPWR hold666/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4497_ _4701_/A _4693_/B VGND VGND VPWR VPWR _4643_/D sky130_fd_sc_hd__nand2_1
Xhold677 hold677/A VGND VGND VPWR VPWR hold677/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold688 hold688/A VGND VGND VPWR VPWR hold688/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6236_ _6687_/Q _5980_/X _6017_/X _6769_/Q VGND VGND VPWR VPWR _6236_/X sky130_fd_sc_hd__a22o_1
Xhold699 hold699/A VGND VGND VPWR VPWR hold699/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3448_ _6994_/Q _5416_/A _5308_/A _6898_/Q _3434_/X VGND VGND VPWR VPWR _3449_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2001 _6534_/Q VGND VGND VPWR VPWR hold455/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2012 hold535/X VGND VGND VPWR VPWR _5547_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_58_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2023 _6873_/Q VGND VGND VPWR VPWR hold546/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2034 _7013_/Q VGND VGND VPWR VPWR hold778/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6167_ _6191_/A2 _6166_/X _6342_/S VGND VGND VPWR VPWR _6167_/X sky130_fd_sc_hd__mux2_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2045 _6597_/Q VGND VGND VPWR VPWR hold598/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_58_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3379_ _6876_/Q _5281_/A _5362_/A _6948_/Q VGND VGND VPWR VPWR _3379_/X sky130_fd_sc_hd__a22o_1
Xhold1300 _5233_/X VGND VGND VPWR VPWR _6826_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_134_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1311 _6811_/Q VGND VGND VPWR VPWR hold231/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2056 _6792_/Q VGND VGND VPWR VPWR hold611/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1322 _5280_/X VGND VGND VPWR VPWR _6868_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2067 _6787_/Q VGND VGND VPWR VPWR hold620/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5118_ _4417_/B _4688_/C _4779_/X _4954_/A VGND VGND VPWR VPWR _5149_/C sky130_fd_sc_hd__o211a_1
Xhold1333 _6705_/Q VGND VGND VPWR VPWR hold279/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2078 _5345_/X VGND VGND VPWR VPWR _6925_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1344 _5269_/X VGND VGND VPWR VPWR _6858_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2089 _6845_/Q VGND VGND VPWR VPWR hold666/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6098_ _6856_/Q _5983_/X _6005_/X _6944_/Q VGND VGND VPWR VPWR _6098_/X sky130_fd_sc_hd__a22o_1
XFILLER_85_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1355 _6977_/Q VGND VGND VPWR VPWR hold434/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1366 _6973_/Q VGND VGND VPWR VPWR hold657/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1377 _5206_/X VGND VGND VPWR VPWR _6807_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5049_ _5049_/A _5049_/B _5049_/C _5049_/D VGND VGND VPWR VPWR _5121_/C sky130_fd_sc_hd__and4_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1388 _6617_/Q VGND VGND VPWR VPWR hold318/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1399 _6988_/Q VGND VGND VPWR VPWR hold413/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_702 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4420_ _4420_/A _4461_/B _4420_/C VGND VGND VPWR VPWR _4477_/C sky130_fd_sc_hd__and3_2
XFILLER_172_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4351_ _4637_/A _4637_/B _4575_/C _4637_/D VGND VGND VPWR VPWR _4365_/B sky130_fd_sc_hd__o211a_4
XFILLER_125_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3302_ _3302_/A hold88/A _3302_/C VGND VGND VPWR VPWR _3302_/X sky130_fd_sc_hd__and3_1
XFILLER_99_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout409 hold153/X VGND VGND VPWR VPWR _5561_/A1 sky130_fd_sc_hd__buf_6
X_7070_ _7127_/CLK _7070_/D fanout477/X VGND VGND VPWR VPWR _7070_/Q sky130_fd_sc_hd__dfstp_2
X_4282_ _4282_/A0 _5544_/A1 _4285_/S VGND VGND VPWR VPWR _4282_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6021_ _6893_/Q _5989_/X _6015_/X _7013_/Q VGND VGND VPWR VPWR _6021_/X sky130_fd_sc_hd__a22o_1
XFILLER_101_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3233_ _6896_/Q VGND VGND VPWR VPWR _3233_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6923_ _7091_/CLK _6923_/D fanout471/X VGND VGND VPWR VPWR _6923_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6854_ _7140_/CLK _6854_/D fanout469/X VGND VGND VPWR VPWR _6854_/Q sky130_fd_sc_hd__dfstp_2
X_5805_ _6874_/Q _5674_/X _5680_/X _6962_/Q VGND VGND VPWR VPWR _5805_/X sky130_fd_sc_hd__a22o_1
X_6785_ _6793_/CLK _6785_/D _3959_/B VGND VGND VPWR VPWR _6785_/Q sky130_fd_sc_hd__dfrtp_4
X_3997_ _6477_/Q hold78/X _3999_/S VGND VGND VPWR VPWR _3997_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5736_ _6975_/Q _5660_/X _5669_/X _7047_/Q VGND VGND VPWR VPWR _5736_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5667_ _5689_/A _5686_/B _5688_/C VGND VGND VPWR VPWR _5667_/X sky130_fd_sc_hd__and3b_4
XFILLER_136_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4618_ _4625_/A _5048_/A _4562_/A VGND VGND VPWR VPWR _4618_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_190_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5598_ _5598_/A1 _5591_/Y _5641_/B _5597_/X VGND VGND VPWR VPWR _7143_/D sky130_fd_sc_hd__a22o_1
XFILLER_190_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold430 hold430/A VGND VGND VPWR VPWR hold430/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4549_ _4724_/C _4628_/A VGND VGND VPWR VPWR _5138_/A sky130_fd_sc_hd__nand2_1
Xhold441 hold441/A VGND VGND VPWR VPWR hold441/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold452 hold452/A VGND VGND VPWR VPWR hold452/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold463 hold463/A VGND VGND VPWR VPWR _6501_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold474 hold474/A VGND VGND VPWR VPWR hold474/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold485 hold485/A VGND VGND VPWR VPWR hold485/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold496 hold496/A VGND VGND VPWR VPWR hold496/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6219_ _6644_/Q _5990_/X _5996_/X _6649_/Q VGND VGND VPWR VPWR _6219_/X sky130_fd_sc_hd__a22o_1
XFILLER_104_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7199_ _7204_/CLK _7199_/D fanout484/X VGND VGND VPWR VPWR _7199_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1130 hold437/X VGND VGND VPWR VPWR _5190_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_161_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1141 _7083_/Q VGND VGND VPWR VPWR hold367/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1152 _6899_/Q VGND VGND VPWR VPWR hold379/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_161_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1163 _5314_/X VGND VGND VPWR VPWR _6898_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1174 hold391/X VGND VGND VPWR VPWR _5396_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1185 hold418/X VGND VGND VPWR VPWR _4238_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1196 hold480/X VGND VGND VPWR VPWR _5521_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3920_ _6435_/Q _3183_/Y _6654_/Q _3904_/A _3920_/B1 VGND VGND VPWR VPWR _3920_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_32_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3851_ _3920_/B1 _3199_/Y _3814_/B _3851_/B1 VGND VGND VPWR VPWR _3851_/X sky130_fd_sc_hd__a31o_1
XFILLER_20_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6570_ _6731_/CLK _6570_/D _6409_/A VGND VGND VPWR VPWR _6570_/Q sky130_fd_sc_hd__dfrtp_4
X_3782_ _6949_/Q _5371_/A _4056_/C input71/X _3781_/X VGND VGND VPWR VPWR _3783_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_164_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5521_ _5521_/A0 _5575_/A1 _5523_/S VGND VGND VPWR VPWR _5521_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5452_ _5452_/A _5569_/B VGND VGND VPWR VPWR _5460_/S sky130_fd_sc_hd__and2_4
XFILLER_173_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4403_ _4724_/B _4625_/A VGND VGND VPWR VPWR _4969_/A sky130_fd_sc_hd__nand2_4
XFILLER_114_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5383_ _5383_/A0 _5572_/A1 _5388_/S VGND VGND VPWR VPWR _5383_/X sky130_fd_sc_hd__mux2_1
X_7122_ _7127_/CLK hold68/X fanout477/X VGND VGND VPWR VPWR _7122_/Q sky130_fd_sc_hd__dfrtp_4
X_4334_ _4334_/A _5229_/C VGND VGND VPWR VPWR _4339_/S sky130_fd_sc_hd__and2_4
XFILLER_99_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7053_ _7053_/CLK _7053_/D fanout452/X VGND VGND VPWR VPWR _7053_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_115_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4265_ hold584/X _5187_/A1 _4267_/S VGND VGND VPWR VPWR _6699_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6004_ _6015_/B _6017_/A _6007_/C VGND VGND VPWR VPWR _6004_/X sky130_fd_sc_hd__and3_4
X_3216_ _7024_/Q VGND VGND VPWR VPWR _3216_/Y sky130_fd_sc_hd__inv_2
X_4196_ _4196_/A0 _5193_/A1 _4199_/S VGND VGND VPWR VPWR _4196_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6906_ _7130_/CLK _6906_/D fanout458/X VGND VGND VPWR VPWR _6906_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6837_ _7102_/CLK _6837_/D _6409_/A VGND VGND VPWR VPWR _6837_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_23_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6768_ _7183_/CLK _6768_/D _6346_/B VGND VGND VPWR VPWR _6768_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5719_ _6942_/Q _5658_/X _5681_/X _7086_/Q VGND VGND VPWR VPWR _5719_/X sky130_fd_sc_hd__a22o_1
X_6699_ _6742_/CLK _6699_/D fanout439/X VGND VGND VPWR VPWR _6699_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_136_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold260 hold260/A VGND VGND VPWR VPWR hold837/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold271 hold271/A VGND VGND VPWR VPWR hold271/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold282 hold282/A VGND VGND VPWR VPWR wb_dat_o[12] sky130_fd_sc_hd__buf_12
XFILLER_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold293 hold293/A VGND VGND VPWR VPWR _7133_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_100 _3893_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 _5559_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 _5221_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_133 hold20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_144 _5488_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_155 _5662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_166 _6015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_177 _7128_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_188 _5559_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_199 _5673_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_749 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4050_ _4050_/A0 _5581_/A1 _4055_/S VGND VGND VPWR VPWR _4050_/X sky130_fd_sc_hd__mux2_1
Xinput6 mask_rev_in[11] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4952_ _4601_/A _4491_/Y _4514_/B _4947_/A _4802_/B VGND VGND VPWR VPWR _5038_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3903_ _3903_/A _3904_/A VGND VGND VPWR VPWR _3903_/Y sky130_fd_sc_hd__nor2_1
X_4883_ _4438_/Y _4601_/A _4601_/B _4580_/Y _4581_/X VGND VGND VPWR VPWR _4883_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_177_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6622_ _6761_/CLK _6622_/D fanout449/X VGND VGND VPWR VPWR _6622_/Q sky130_fd_sc_hd__dfrtp_4
X_3834_ _3248_/X _3247_/Y _3834_/S VGND VGND VPWR VPWR _3834_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6553_ _6568_/CLK _6553_/D VGND VGND VPWR VPWR _6553_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3765_ input11/X _3310_/Y _5209_/S _7206_/A VGND VGND VPWR VPWR _3765_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5504_ _5504_/A0 _5576_/A1 _5505_/S VGND VGND VPWR VPWR _5504_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6484_ _6809_/CLK _6484_/D fanout444/X VGND VGND VPWR VPWR _6484_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_118_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3696_ _6796_/Q _3319_/Y _4164_/A _6610_/Q _3695_/X VGND VGND VPWR VPWR _3703_/A
+ sky130_fd_sc_hd__a221o_2
Xpad_flashh_clk_buff_inst _3958_/X VGND VGND VPWR VPWR pad_flash_clk sky130_fd_sc_hd__clkbuf_8
X_5435_ hold805/X _5552_/A1 _5442_/S VGND VGND VPWR VPWR _7005_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput310 _3966_/X VGND VGND VPWR VPWR spimemio_flash_io1_di sky130_fd_sc_hd__buf_12
Xoutput321 hold847/X VGND VGND VPWR VPWR hold275/A sky130_fd_sc_hd__buf_6
Xoutput332 hold853/X VGND VGND VPWR VPWR hold197/A sky130_fd_sc_hd__buf_6
XFILLER_105_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput343 hold851/X VGND VGND VPWR VPWR hold278/A sky130_fd_sc_hd__buf_6
X_5366_ _5366_/A0 _5555_/A1 _5370_/S VGND VGND VPWR VPWR _5366_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4317_ _4317_/A0 _5208_/A1 _4321_/S VGND VGND VPWR VPWR _6742_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_824 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7105_ _7105_/CLK _7105_/D fanout473/X VGND VGND VPWR VPWR _7105_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_113_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5297_ _5297_/A0 _5585_/A1 _5298_/S VGND VGND VPWR VPWR _5297_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7036_ _7116_/CLK _7036_/D fanout455/X VGND VGND VPWR VPWR _7036_/Q sky130_fd_sc_hd__dfrtp_4
X_4248_ _4248_/A0 _5585_/A1 _4249_/S VGND VGND VPWR VPWR _4248_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4179_ _4179_/A0 _4337_/A1 _4181_/S VGND VGND VPWR VPWR _4179_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_41_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7103_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_56_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _6833_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_186_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3550_ _3550_/A _3550_/B VGND VGND VPWR VPWR _4286_/A sky130_fd_sc_hd__nor2_8
XFILLER_128_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3481_ _3481_/A _3481_/B _3481_/C _3481_/D VGND VGND VPWR VPWR _3558_/A sky130_fd_sc_hd__nor4_2
XFILLER_127_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5220_ hold90/X _5220_/B _5220_/C VGND VGND VPWR VPWR _5221_/S sky130_fd_sc_hd__and3_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5151_ _5150_/X _5151_/B _5151_/C _5151_/D VGND VGND VPWR VPWR _5152_/B sky130_fd_sc_hd__and4b_1
Xhold2408 _5529_/X VGND VGND VPWR VPWR _7089_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2419 _6776_/Q VGND VGND VPWR VPWR _3677_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4102_ _3616_/Y hold826/A _4106_/S VGND VGND VPWR VPWR _6556_/D sky130_fd_sc_hd__mux2_1
Xhold1707 hold451/X VGND VGND VPWR VPWR _5285_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5082_ _4578_/A _4990_/B _5108_/A _5023_/A VGND VGND VPWR VPWR _5083_/D sky130_fd_sc_hd__o211a_1
XFILLER_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1718 _7088_/Q VGND VGND VPWR VPWR hold441/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1729 _4207_/X VGND VGND VPWR VPWR _6644_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4033_ hold742/X _5571_/A1 _4056_/C VGND VGND VPWR VPWR _4033_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5984_ _6008_/A _6018_/B _6019_/C VGND VGND VPWR VPWR _5984_/X sky130_fd_sc_hd__and3_4
X_4935_ _5011_/A _4601_/A _4663_/D _4465_/B VGND VGND VPWR VPWR _4935_/X sky130_fd_sc_hd__a211o_2
XFILLER_21_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_7_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR _6850_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_11 _3347_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 _3699_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4866_ _4638_/Y _4995_/A _4924_/C _4865_/X _5095_/B VGND VGND VPWR VPWR _4866_/X
+ sky130_fd_sc_hd__o2111a_1
XANTENNA_33 _5670_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_44 _5989_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6605_ _6711_/CLK _6605_/D _6433_/A VGND VGND VPWR VPWR _6605_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_193_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3817_ _6447_/Q _6446_/Q VGND VGND VPWR VPWR _3863_/A sky130_fd_sc_hd__nor2_1
XANTENNA_55 _6015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_66 _7072_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4797_ _4729_/A _4713_/Y _4796_/X _4534_/Y VGND VGND VPWR VPWR _4797_/X sky130_fd_sc_hd__o211a_1
XFILLER_165_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_808 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_77 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_88 _7232_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_99 input97/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6536_ _6808_/CLK _6536_/D fanout439/X VGND VGND VPWR VPWR _6536_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3748_ _7133_/Q hold33/A _3431_/Y input61/X VGND VGND VPWR VPWR _3748_/X sky130_fd_sc_hd__a22o_2
XFILLER_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6467_ _6658_/CLK _6467_/D _6417_/X VGND VGND VPWR VPWR _6467_/Q sky130_fd_sc_hd__dfrtp_1
X_3679_ _6918_/Q _5335_/A _4280_/A _6713_/Q _3678_/X VGND VGND VPWR VPWR _3684_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5418_ _5418_/A0 _5571_/A1 _5424_/S VGND VGND VPWR VPWR _5418_/X sky130_fd_sc_hd__mux2_1
X_6398_ _6399_/A _6423_/B VGND VGND VPWR VPWR _6398_/X sky130_fd_sc_hd__and2_1
XFILLER_133_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput173 _3973_/X VGND VGND VPWR VPWR irq[1] sky130_fd_sc_hd__buf_12
XFILLER_121_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput184 _3221_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[18] sky130_fd_sc_hd__buf_12
X_5349_ _5349_/A0 _5583_/A1 _5352_/S VGND VGND VPWR VPWR _5349_/X sky130_fd_sc_hd__mux2_1
Xoutput195 _3211_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[28] sky130_fd_sc_hd__buf_12
XFILLER_75_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7019_ _7140_/CLK _7019_/D fanout471/X VGND VGND VPWR VPWR _7019_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _4649_/B _4720_/B _4720_/C VGND VGND VPWR VPWR _4993_/B sky130_fd_sc_hd__and3b_2
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4651_ _4590_/Y _4648_/Y _4683_/A _5121_/A VGND VGND VPWR VPWR _4651_/X sky130_fd_sc_hd__o31a_1
XFILLER_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput20 mask_rev_in[24] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__clkbuf_2
X_3602_ input29/X _3307_/Y _3315_/Y input6/X VGND VGND VPWR VPWR _3602_/X sky130_fd_sc_hd__a22o_2
Xinput31 mask_rev_in[5] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4582_ _4582_/A _4724_/C VGND VGND VPWR VPWR _4969_/B sky130_fd_sc_hd__nand2_2
XFILLER_190_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput42 mgmt_gpio_in[15] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput53 mgmt_gpio_in[25] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput64 mgmt_gpio_in[35] VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__buf_2
XFILLER_190_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6321_ _6598_/Q _5991_/X _6018_/X _6721_/Q _6318_/X VGND VGND VPWR VPWR _6321_/X
+ sky130_fd_sc_hd__a221o_1
X_3533_ _3553_/A _3533_/B VGND VGND VPWR VPWR _4304_/A sky130_fd_sc_hd__nor2_8
Xhold804 hold804/A VGND VGND VPWR VPWR hold804/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput75 porb VGND VGND VPWR VPWR input75/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold815 hold815/A VGND VGND VPWR VPWR hold815/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput86 spimemio_flash_io0_oeb VGND VGND VPWR VPWR _3960_/B sky130_fd_sc_hd__buf_4
Xhold826 hold826/A VGND VGND VPWR VPWR hold826/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput97 usr2_vcc_pwrgood VGND VGND VPWR VPWR input97/X sky130_fd_sc_hd__clkbuf_4
Xhold837 hold837/A VGND VGND VPWR VPWR hold837/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold848 hold848/A VGND VGND VPWR VPWR hold848/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6252_ _6630_/Q _5971_/X _6007_/X _6531_/Q _6251_/X VGND VGND VPWR VPWR _6255_/B
+ sky130_fd_sc_hd__a221o_1
Xhold859 hold859/A VGND VGND VPWR VPWR hold859/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3464_ _3463_/X _3464_/A1 _3739_/S VGND VGND VPWR VPWR _3464_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5203_ _5203_/A0 _5570_/A1 _5206_/S VGND VGND VPWR VPWR _6804_/D sky130_fd_sc_hd__mux2_1
X_6183_ _7131_/Q _5973_/X _5986_/X _7035_/Q _6182_/X VGND VGND VPWR VPWR _6183_/X
+ sky130_fd_sc_hd__a221o_1
Xhold2205 hold794/X VGND VGND VPWR VPWR _5176_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_3395_ _7115_/Q _5551_/A _5263_/A _6859_/Q VGND VGND VPWR VPWR _3395_/X sky130_fd_sc_hd__a22o_1
XFILLER_97_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2216 hold466/X VGND VGND VPWR VPWR _4297_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2227 hold798/X VGND VGND VPWR VPWR _4147_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5134_ _5134_/A _5155_/C VGND VGND VPWR VPWR _5134_/Y sky130_fd_sc_hd__nand2_1
Xhold2238 hold486/X VGND VGND VPWR VPWR _3993_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2249 _6631_/Q VGND VGND VPWR VPWR hold587/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1504 _6837_/Q VGND VGND VPWR VPWR hold335/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1515 _6543_/Q VGND VGND VPWR VPWR hold820/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1526 _7124_/Q VGND VGND VPWR VPWR hold519/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1537 _6487_/Q VGND VGND VPWR VPWR hold668/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5065_ _4570_/C _4968_/Y _4903_/B _4622_/C _4539_/Y VGND VGND VPWR VPWR _5131_/A
+ sky130_fd_sc_hd__o2111a_1
Xhold1548 hold860/X VGND VGND VPWR VPWR hold285/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1559 hold118/X VGND VGND VPWR VPWR _4273_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4016_ _4049_/A0 _5571_/A1 _4047_/C VGND VGND VPWR VPWR _4016_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5967_ _6539_/Q _5651_/X _5962_/X _5966_/X VGND VGND VPWR VPWR _5967_/X sky130_fd_sc_hd__a211o_1
X_4918_ _4365_/B _4988_/A _4840_/A _4917_/X VGND VGND VPWR VPWR _4919_/C sky130_fd_sc_hd__a22oi_4
X_5898_ _6575_/Q _5667_/X _5682_/X _6451_/Q VGND VGND VPWR VPWR _5898_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4849_ _5009_/A _4710_/A _4811_/B VGND VGND VPWR VPWR _5089_/B sky130_fd_sc_hd__o21ai_2
XFILLER_21_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6519_ _6522_/CLK _6519_/D fanout478/X VGND VGND VPWR VPWR _6519_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3180_ _6469_/Q VGND VGND VPWR VPWR _3879_/A sky130_fd_sc_hd__clkinv_2
XFILLER_93_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6870_ _7127_/CLK _6870_/D fanout477/X VGND VGND VPWR VPWR _6870_/Q sky130_fd_sc_hd__dfstp_2
X_5821_ _6883_/Q _5667_/X _5687_/X _6923_/Q _5820_/X VGND VGND VPWR VPWR _5826_/B
+ sky130_fd_sc_hd__a221o_1
X_5752_ _7056_/Q _5668_/X _5681_/X _7088_/Q VGND VGND VPWR VPWR _5752_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4703_ _4703_/A _4703_/B _4703_/C _4703_/D VGND VGND VPWR VPWR _4704_/D sky130_fd_sc_hd__and4_1
XFILLER_187_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5683_ _7085_/Q _5681_/X _5682_/X _7037_/Q VGND VGND VPWR VPWR _5683_/X sky130_fd_sc_hd__a22o_1
XFILLER_175_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4634_ _5001_/A _4731_/A VGND VGND VPWR VPWR _4965_/B sky130_fd_sc_hd__nand2_2
XFILLER_175_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold601 hold601/A VGND VGND VPWR VPWR hold601/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4565_ _4971_/A _4693_/B VGND VGND VPWR VPWR _4898_/B sky130_fd_sc_hd__nand2_1
Xhold612 hold612/A VGND VGND VPWR VPWR hold612/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold623 hold623/A VGND VGND VPWR VPWR hold623/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold634 hold634/A VGND VGND VPWR VPWR hold634/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6304_ _6304_/A _6304_/B _6304_/C _6304_/D VGND VGND VPWR VPWR _6314_/B sky130_fd_sc_hd__nor4_1
XFILLER_144_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold645 hold645/A VGND VGND VPWR VPWR hold645/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3516_ _3540_/A _3516_/B VGND VGND VPWR VPWR _4092_/A sky130_fd_sc_hd__nor2_4
Xmax_cap353 _3293_/Y VGND VGND VPWR VPWR _4056_/C sky130_fd_sc_hd__buf_12
XFILLER_143_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold656 hold656/A VGND VGND VPWR VPWR hold656/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4496_ _4576_/A _4523_/A VGND VGND VPWR VPWR _4658_/B sky130_fd_sc_hd__nand2_4
Xhold667 hold667/A VGND VGND VPWR VPWR hold667/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold678 hold678/A VGND VGND VPWR VPWR hold678/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3447_ _6890_/Q _5299_/A _5497_/A _7066_/Q _3435_/X VGND VGND VPWR VPWR _3449_/B
+ sky130_fd_sc_hd__a221o_1
X_6235_ _6722_/Q _5978_/X _5995_/X _6599_/Q _6234_/X VGND VGND VPWR VPWR _6238_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold689 hold689/A VGND VGND VPWR VPWR hold689/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2002 hold455/X VGND VGND VPWR VPWR _4076_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2013 _6818_/Q VGND VGND VPWR VPWR hold641/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2024 hold546/X VGND VGND VPWR VPWR _5286_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_3378_ _7028_/Q _5452_/A _3307_/Y input33/X _3348_/X VGND VGND VPWR VPWR _3383_/B
+ sky130_fd_sc_hd__a221o_1
Xhold2035 _6532_/Q VGND VGND VPWR VPWR hold589/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6166_ _7177_/Q _6165_/X _6166_/S VGND VGND VPWR VPWR _6166_/X sky130_fd_sc_hd__mux2_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2046 hold598/X VGND VGND VPWR VPWR _4150_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1301 _7195_/Q VGND VGND VPWR VPWR hold151/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1312 hold231/X VGND VGND VPWR VPWR _5213_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2057 hold611/X VGND VGND VPWR VPWR _5188_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1323 _6740_/Q VGND VGND VPWR VPWR hold269/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2068 hold620/X VGND VGND VPWR VPWR _5182_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5117_ _5117_/A _5117_/B _5117_/C VGND VGND VPWR VPWR _5117_/X sky130_fd_sc_hd__and3_1
Xhold1334 hold279/X VGND VGND VPWR VPWR _4272_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2079 _6965_/Q VGND VGND VPWR VPWR hold810/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6097_ _6992_/Q _6014_/X _6095_/X _6096_/X VGND VGND VPWR VPWR _6102_/A sky130_fd_sc_hd__a211o_1
Xhold1345 _6565_/Q VGND VGND VPWR VPWR hold872/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1356 hold434/X VGND VGND VPWR VPWR _5403_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1367 _7020_/Q VGND VGND VPWR VPWR hold358/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5048_ _5048_/A _5048_/B VGND VGND VPWR VPWR _5049_/D sky130_fd_sc_hd__nand2_1
Xhold1378 _6853_/Q VGND VGND VPWR VPWR hold646/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1389 hold318/X VGND VGND VPWR VPWR _4174_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6999_ _7126_/CLK _6999_/D fanout475/X VGND VGND VPWR VPWR _6999_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_43_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1890 _6757_/Q VGND VGND VPWR VPWR hold653/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_90_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4350_ _4637_/A _4637_/B VGND VGND VPWR VPWR _4638_/A sky130_fd_sc_hd__nor2_8
XFILLER_125_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3301_ _3349_/A _3726_/A VGND VGND VPWR VPWR _5398_/A sky130_fd_sc_hd__nor2_8
X_4281_ _4281_/A0 hold153/X _4285_/S VGND VGND VPWR VPWR _4281_/X sky130_fd_sc_hd__mux2_1
X_6020_ _6861_/Q _5999_/X _6005_/X _6941_/Q VGND VGND VPWR VPWR _6020_/X sky130_fd_sc_hd__a22o_1
X_3232_ _6904_/Q VGND VGND VPWR VPWR _3232_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6922_ _7020_/CLK _6922_/D fanout458/X VGND VGND VPWR VPWR _6922_/Q sky130_fd_sc_hd__dfrtp_4
X_6853_ _7125_/CLK _6853_/D fanout454/X VGND VGND VPWR VPWR _6853_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_120_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5804_ _6946_/Q _5658_/X _5664_/X _7018_/Q VGND VGND VPWR VPWR _5804_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6784_ _6793_/CLK _6784_/D _3959_/B VGND VGND VPWR VPWR _6784_/Q sky130_fd_sc_hd__dfrtp_4
X_3996_ hold76/X hold897/X _3996_/S VGND VGND VPWR VPWR _3996_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5735_ _6983_/Q _5656_/X _5663_/X _7023_/Q _5734_/X VGND VGND VPWR VPWR _5735_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5666_ _5689_/A _5679_/B _5688_/C VGND VGND VPWR VPWR _5666_/X sky130_fd_sc_hd__and3_4
X_4617_ _4522_/B _4570_/D _4614_/X _4616_/X VGND VGND VPWR VPWR _4617_/X sky130_fd_sc_hd__o211a_1
XFILLER_117_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5597_ _7142_/Q _7143_/Q _6490_/Q _6492_/Q _3924_/Y VGND VGND VPWR VPWR _5597_/X
+ sky130_fd_sc_hd__o221a_1
Xhold420 hold420/A VGND VGND VPWR VPWR hold420/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold431 hold431/A VGND VGND VPWR VPWR hold431/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4548_ _4575_/C _4463_/B _4569_/B _4546_/X _4770_/A VGND VGND VPWR VPWR _4548_/X
+ sky130_fd_sc_hd__o311a_1
Xhold442 hold442/A VGND VGND VPWR VPWR hold442/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold453 hold453/A VGND VGND VPWR VPWR hold453/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold464 hold464/A VGND VGND VPWR VPWR hold464/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold475 hold475/A VGND VGND VPWR VPWR hold475/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold486 hold486/A VGND VGND VPWR VPWR hold486/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4479_ _4486_/A _4485_/B _4881_/A VGND VGND VPWR VPWR _4562_/A sky130_fd_sc_hd__and3_2
Xhold497 hold497/A VGND VGND VPWR VPWR hold497/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6218_ _6594_/Q _5991_/X _6018_/X _6717_/Q VGND VGND VPWR VPWR _6218_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7198_ _7204_/CLK _7198_/D fanout484/X VGND VGND VPWR VPWR _7198_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6149_ _7026_/Q _5971_/X _6007_/X _6850_/Q _6148_/X VGND VGND VPWR VPWR _6152_/B
+ sky130_fd_sc_hd__a221o_1
Xhold1120 _6947_/Q VGND VGND VPWR VPWR hold407/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1131 _5190_/X VGND VGND VPWR VPWR _6794_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1142 hold367/X VGND VGND VPWR VPWR _5522_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1153 hold379/X VGND VGND VPWR VPWR _5315_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1164 _6570_/Q VGND VGND VPWR VPWR hold194/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_161_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1175 _5396_/X VGND VGND VPWR VPWR _6971_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1186 _4238_/X VGND VGND VPWR VPWR _6666_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1197 _5521_/X VGND VGND VPWR VPWR _7082_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3850_ _3927_/A1 _3850_/A1 _3850_/S VGND VGND VPWR VPWR _6459_/D sky130_fd_sc_hd__mux2_1
X_3781_ _6957_/Q _5380_/A _4152_/A _6599_/Q VGND VGND VPWR VPWR _3781_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5520_ _5520_/A0 _5583_/A1 _5523_/S VGND VGND VPWR VPWR _7081_/D sky130_fd_sc_hd__mux2_1
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5451_ _5451_/A0 _5559_/A1 _5451_/S VGND VGND VPWR VPWR _7020_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4402_ _4523_/A _4590_/B VGND VGND VPWR VPWR _4402_/Y sky130_fd_sc_hd__nand2_4
X_5382_ hold764/X _5580_/A1 _5388_/S VGND VGND VPWR VPWR _5382_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7121_ _7121_/CLK _7121_/D fanout473/X VGND VGND VPWR VPWR _7121_/Q sky130_fd_sc_hd__dfrtp_4
X_4333_ _4333_/A0 _5538_/A1 _4333_/S VGND VGND VPWR VPWR _4333_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4264_ _4264_/A0 _5186_/A1 _4267_/S VGND VGND VPWR VPWR _6698_/D sky130_fd_sc_hd__mux2_1
X_7052_ _7084_/CLK _7052_/D fanout456/X VGND VGND VPWR VPWR _7052_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6003_ _7151_/Q _6007_/C _6016_/C _5989_/X _5997_/X VGND VGND VPWR VPWR _6010_/A
+ sky130_fd_sc_hd__a311o_1
X_3215_ _7032_/Q VGND VGND VPWR VPWR _3215_/Y sky130_fd_sc_hd__clkinv_2
X_4195_ _4195_/A0 _5208_/A1 _4199_/S VGND VGND VPWR VPWR _4195_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6905_ _7135_/CLK _6905_/D fanout473/X VGND VGND VPWR VPWR _6905_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6836_ _7116_/CLK _6836_/D fanout457/X VGND VGND VPWR VPWR _6836_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_51_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6767_ _7183_/CLK _6767_/D _6346_/B VGND VGND VPWR VPWR hold22/A sky130_fd_sc_hd__dfrtp_1
XFILLER_149_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3979_ _3979_/A0 _5221_/A1 _3987_/S VGND VGND VPWR VPWR _6450_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5718_ _5718_/A _5718_/B _5718_/C VGND VGND VPWR VPWR _5718_/Y sky130_fd_sc_hd__nor3_1
XFILLER_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6698_ _6808_/CLK _6698_/D fanout440/X VGND VGND VPWR VPWR _6698_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5649_ _5730_/S VGND VGND VPWR VPWR _5649_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_136_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold250 hold250/A VGND VGND VPWR VPWR hold833/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold261 hold261/A VGND VGND VPWR VPWR wb_dat_o[13] sky130_fd_sc_hd__buf_12
XFILLER_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold272 hold272/A VGND VGND VPWR VPWR wb_dat_o[4] sky130_fd_sc_hd__buf_12
Xhold283 hold283/A VGND VGND VPWR VPWR hold283/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold294 hold294/A VGND VGND VPWR VPWR hold294/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 _3893_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_112 _5559_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_123 _5561_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 hold135/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 _5362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 _5663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_167 _6018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_178 _6574_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_189 _5503_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput7 mask_rev_in[12] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4951_ _4368_/A _4462_/Y _4934_/Y _5041_/A _4800_/B VGND VGND VPWR VPWR _5148_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3902_ _3968_/A _3969_/B _3901_/Y _3921_/A VGND VGND VPWR VPWR _6682_/D sky130_fd_sc_hd__a22o_1
X_4882_ _4934_/B _4972_/B VGND VGND VPWR VPWR _5102_/B sky130_fd_sc_hd__nand2_1
XFILLER_177_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6621_ _6759_/CLK _6621_/D _6426_/A VGND VGND VPWR VPWR _6621_/Q sky130_fd_sc_hd__dfstp_2
X_3833_ _3833_/A _3833_/B VGND VGND VPWR VPWR _6465_/D sky130_fd_sc_hd__xnor2_1
XFILLER_193_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6552_ _6757_/CLK _6552_/D fanout446/X VGND VGND VPWR VPWR _6552_/Q sky130_fd_sc_hd__dfrtp_4
X_3764_ _3764_/A _3764_/B VGND VGND VPWR VPWR _5209_/S sky130_fd_sc_hd__nor2_2
X_5503_ _5503_/A0 _5503_/A1 _5505_/S VGND VGND VPWR VPWR _5503_/X sky130_fd_sc_hd__mux2_1
X_6483_ _6792_/CLK _6483_/D fanout442/X VGND VGND VPWR VPWR _6483_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_145_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3695_ _6630_/Q _4188_/A _4322_/A _6748_/Q VGND VGND VPWR VPWR _3695_/X sky130_fd_sc_hd__a22o_1
Xoutput300 _6807_/Q VGND VGND VPWR VPWR pwr_ctrl_out[3] sky130_fd_sc_hd__buf_12
X_5434_ _5434_/A _5551_/B VGND VGND VPWR VPWR _5442_/S sky130_fd_sc_hd__and2_4
XFILLER_161_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput311 _7232_/X VGND VGND VPWR VPWR spimemio_flash_io2_di sky130_fd_sc_hd__buf_12
Xoutput322 hold839/X VGND VGND VPWR VPWR hold264/A sky130_fd_sc_hd__buf_6
XFILLER_133_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput333 hold855/X VGND VGND VPWR VPWR hold201/A sky130_fd_sc_hd__buf_6
Xoutput344 hold841/X VGND VGND VPWR VPWR hold266/A sky130_fd_sc_hd__buf_6
XFILLER_160_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5365_ _5365_/A0 _5581_/A1 _5370_/S VGND VGND VPWR VPWR _6943_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_3_3_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR _7093_/CLK sky130_fd_sc_hd__clkbuf_8
X_7104_ _7138_/CLK _7104_/D fanout480/X VGND VGND VPWR VPWR _7104_/Q sky130_fd_sc_hd__dfrtp_4
X_4316_ _4316_/A _5229_/C VGND VGND VPWR VPWR _4321_/S sky130_fd_sc_hd__and2_4
XFILLER_141_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5296_ hold919/X hold20/X _5298_/S VGND VGND VPWR VPWR _5296_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7035_ _7035_/CLK _7035_/D fanout456/X VGND VGND VPWR VPWR _7035_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4247_ hold886/X hold20/X _4249_/S VGND VGND VPWR VPWR _4247_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4178_ _4178_/A0 _5193_/A1 _4181_/S VGND VGND VPWR VPWR _4178_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6819_ _7102_/CLK _6819_/D fanout465/X VGND VGND VPWR VPWR _6819_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_168_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire438 _3881_/Y VGND VGND VPWR VPWR wire438/X sky130_fd_sc_hd__buf_4
XFILLER_183_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3480_ input56/X _4241_/A _4158_/A _6608_/Q _3478_/X VGND VGND VPWR VPWR _3481_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_155_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5150_ _5150_/A _5150_/B _5150_/C VGND VGND VPWR VPWR _5150_/X sky130_fd_sc_hd__and3_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2409 _6953_/Q VGND VGND VPWR VPWR hold750/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4101_ _3675_/Y hold832/A _4106_/S VGND VGND VPWR VPWR _6555_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5081_ _5081_/A _5081_/B VGND VGND VPWR VPWR _5081_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1708 _5285_/X VGND VGND VPWR VPWR _6872_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1719 hold441/X VGND VGND VPWR VPWR _5528_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4032_ _4032_/A0 _4031_/X _4046_/S VGND VGND VPWR VPWR _4032_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5983_ _6019_/A _6019_/C _6007_/C VGND VGND VPWR VPWR _5983_/X sky130_fd_sc_hd__and3_4
X_4934_ _5009_/A _4934_/B VGND VGND VPWR VPWR _4934_/Y sky130_fd_sc_hd__nor2_1
XFILLER_178_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4865_ _4402_/Y _4570_/A _4651_/X _4856_/X _4864_/X VGND VGND VPWR VPWR _4865_/X
+ sky130_fd_sc_hd__o2111a_1
XANTENNA_12 hold27/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 _3783_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 _5673_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6604_ _6759_/CLK _6604_/D fanout447/X VGND VGND VPWR VPWR _6604_/Q sky130_fd_sc_hd__dfrtp_4
X_3816_ _6656_/Q _3904_/A VGND VGND VPWR VPWR _3816_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_45 _5989_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 _6016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4796_ _4796_/A _4796_/B _4796_/C VGND VGND VPWR VPWR _4796_/X sky130_fd_sc_hd__and3_1
XFILLER_20_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_67 _6856_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_78 wb_clk_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_89 _7233_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6535_ _6747_/CLK _6535_/D fanout439/X VGND VGND VPWR VPWR _6535_/Q sky130_fd_sc_hd__dfrtp_4
X_3747_ _3303_/X _3328_/X _3745_/Y _3746_/X VGND VGND VPWR VPWR _3750_/C sky130_fd_sc_hd__a31o_1
XFILLER_21_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6466_ _6658_/CLK _6466_/D _6416_/X VGND VGND VPWR VPWR hold86/A sky130_fd_sc_hd__dfrtp_1
X_3678_ _6650_/Q _4212_/A _3562_/Y input96/X VGND VGND VPWR VPWR _3678_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5417_ hold792/X _5570_/A1 _5424_/S VGND VGND VPWR VPWR _5417_/X sky130_fd_sc_hd__mux2_1
X_6397_ _6399_/A _6423_/B VGND VGND VPWR VPWR _6397_/X sky130_fd_sc_hd__and2_1
Xoutput174 _3974_/X VGND VGND VPWR VPWR irq[2] sky130_fd_sc_hd__buf_12
XFILLER_0_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5348_ _5348_/A0 _5555_/A1 _5352_/S VGND VGND VPWR VPWR _5348_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput185 _3220_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[19] sky130_fd_sc_hd__buf_12
Xoutput196 _3210_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[29] sky130_fd_sc_hd__buf_12
XFILLER_0_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5279_ _5279_/A0 _5576_/A1 _5280_/S VGND VGND VPWR VPWR _5279_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7018_ _7018_/CLK _7018_/D fanout459/X VGND VGND VPWR VPWR _7018_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout390 _5555_/A1 VGND VGND VPWR VPWR _5582_/A1 sky130_fd_sc_hd__buf_8
XFILLER_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4650_ _4720_/B _4650_/B VGND VGND VPWR VPWR _4683_/A sky130_fd_sc_hd__nand2_8
XFILLER_187_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput10 mask_rev_in[15] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3601_ _6984_/Q _5407_/A _4176_/A _6622_/Q _3600_/X VGND VGND VPWR VPWR _3604_/C
+ sky130_fd_sc_hd__a221o_1
Xinput21 mask_rev_in[25] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__buf_2
Xinput32 mask_rev_in[6] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4581_ _4560_/B _4560_/C _4652_/A VGND VGND VPWR VPWR _4581_/X sky130_fd_sc_hd__a21bo_4
Xinput43 mgmt_gpio_in[16] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__clkbuf_2
Xinput54 mgmt_gpio_in[26] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__clkbuf_4
X_6320_ _6648_/Q _5990_/X _5996_/X _6653_/Q VGND VGND VPWR VPWR _6320_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput65 mgmt_gpio_in[36] VGND VGND VPWR VPWR _7232_/A sky130_fd_sc_hd__buf_4
Xhold805 hold805/A VGND VGND VPWR VPWR hold805/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3532_ _6638_/Q _4194_/A _4322_/A _6751_/Q VGND VGND VPWR VPWR _3532_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput76 qspi_enabled VGND VGND VPWR VPWR _3934_/S sky130_fd_sc_hd__buf_8
Xhold816 hold816/A VGND VGND VPWR VPWR hold816/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput87 spimemio_flash_io1_do VGND VGND VPWR VPWR _7231_/A sky130_fd_sc_hd__buf_4
Xinput98 usr2_vdd_pwrgood VGND VGND VPWR VPWR input98/X sky130_fd_sc_hd__buf_2
Xhold827 hold827/A VGND VGND VPWR VPWR hold827/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold838 hold838/A VGND VGND VPWR VPWR hold838/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6251_ _6536_/Q _5983_/X _6005_/X _6693_/Q VGND VGND VPWR VPWR _6251_/X sky130_fd_sc_hd__a22o_1
Xhold849 hold849/A VGND VGND VPWR VPWR hold849/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3463_ _6778_/Q _3462_/Y _3857_/B VGND VGND VPWR VPWR _3463_/X sky130_fd_sc_hd__mux2_1
X_5202_ _5202_/A _5551_/B VGND VGND VPWR VPWR _5206_/S sky130_fd_sc_hd__and2_2
X_6182_ _7091_/Q _5638_/X _5999_/X _6867_/Q VGND VGND VPWR VPWR _6182_/X sky130_fd_sc_hd__a22o_1
X_3394_ _7107_/Q _3311_/Y _3336_/Y input27/X VGND VGND VPWR VPWR _3394_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2206 _5176_/X VGND VGND VPWR VPWR _6782_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2217 _6894_/Q VGND VGND VPWR VPWR hold701/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5133_ _4564_/Y _4968_/Y _5072_/C _5132_/X _4609_/B VGND VGND VPWR VPWR _5155_/C
+ sky130_fd_sc_hd__o2111a_1
Xhold2228 _7022_/Q VGND VGND VPWR VPWR hold723/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2239 _6596_/Q VGND VGND VPWR VPWR hold572/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1505 _7084_/Q VGND VGND VPWR VPWR hold510/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1516 hold820/X VGND VGND VPWR VPWR hold209/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1527 hold519/X VGND VGND VPWR VPWR _5568_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1538 _6976_/Q VGND VGND VPWR VPWR hold487/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5064_ _4569_/B _4510_/B _4625_/Y _4902_/A _4971_/Y VGND VGND VPWR VPWR _5130_/B
+ sky130_fd_sc_hd__o2111a_1
Xhold1549 _6702_/Q VGND VGND VPWR VPWR hold709/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4015_ hold439/X _4015_/A1 _4029_/S VGND VGND VPWR VPWR _4015_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5966_ _6701_/Q _5672_/X _5963_/X _5965_/X VGND VGND VPWR VPWR _5966_/X sky130_fd_sc_hd__a211o_1
X_4917_ _4917_/A _4917_/B _4917_/C _4917_/D VGND VGND VPWR VPWR _4917_/X sky130_fd_sc_hd__and4_1
X_5897_ _6743_/Q _5929_/B _5668_/X _6645_/Q _5884_/X VGND VGND VPWR VPWR _5897_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_32_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4848_ _4391_/Y _4580_/Y _4640_/Y VGND VGND VPWR VPWR _5049_/B sky130_fd_sc_hd__a21o_1
XFILLER_138_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4779_ _4464_/Y _4569_/C _4688_/C _4947_/A VGND VGND VPWR VPWR _4779_/X sky130_fd_sc_hd__o22a_1
XFILLER_165_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6518_ _6522_/CLK _6518_/D fanout478/X VGND VGND VPWR VPWR _6518_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6449_ _6656_/CLK _6449_/D _6404_/X VGND VGND VPWR VPWR _6449_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_40_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7119_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_115_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_55_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7116_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_91_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5820_ _7035_/Q _5655_/X _5679_/X _6907_/Q VGND VGND VPWR VPWR _5820_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5751_ _5751_/A1 _5730_/S _5749_/X _5750_/X VGND VGND VPWR VPWR _7162_/D sky130_fd_sc_hd__o22a_1
XFILLER_15_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4702_ _5009_/B _4702_/B VGND VGND VPWR VPWR _4702_/Y sky130_fd_sc_hd__nand2_1
XFILLER_148_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5682_ _5686_/A _5686_/B _5687_/C VGND VGND VPWR VPWR _5682_/X sky130_fd_sc_hd__and3_4
XFILLER_148_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4633_ _4658_/A _4633_/B VGND VGND VPWR VPWR _4731_/A sky130_fd_sc_hd__nor2_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4564_ _4579_/B _4564_/B _4564_/C VGND VGND VPWR VPWR _4564_/Y sky130_fd_sc_hd__nand3_4
Xhold602 hold602/A VGND VGND VPWR VPWR hold602/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold613 hold613/A VGND VGND VPWR VPWR hold613/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6303_ _6690_/Q _5980_/X _6016_/X _6453_/Q _6302_/X VGND VGND VPWR VPWR _6304_/D
+ sky130_fd_sc_hd__a221o_1
Xhold624 hold624/A VGND VGND VPWR VPWR hold624/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3515_ _3515_/A _3515_/B _3515_/C _3515_/D VGND VGND VPWR VPWR _3557_/A sky130_fd_sc_hd__nor4_1
Xhold635 hold635/A VGND VGND VPWR VPWR hold635/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap354 _3550_/A VGND VGND VPWR VPWR _3487_/A sky130_fd_sc_hd__buf_12
Xhold646 hold646/A VGND VGND VPWR VPWR hold646/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4495_ _4718_/A _4495_/B VGND VGND VPWR VPWR _4693_/B sky130_fd_sc_hd__nor2_8
Xhold657 hold657/A VGND VGND VPWR VPWR hold657/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap365 _4473_/A VGND VGND VPWR VPWR _4485_/B sky130_fd_sc_hd__clkbuf_4
Xhold668 hold668/A VGND VGND VPWR VPWR hold668/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6234_ _6737_/Q _6008_/X _6016_/X _6450_/Q VGND VGND VPWR VPWR _6234_/X sky130_fd_sc_hd__a22o_1
Xhold679 hold679/A VGND VGND VPWR VPWR hold679/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3446_ _6954_/Q _5371_/A _5236_/C _3970_/A _3445_/X VGND VGND VPWR VPWR _3449_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2003 _4076_/X VGND VGND VPWR VPWR _6534_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2014 hold641/X VGND VGND VPWR VPWR _5223_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6165_ _6842_/Q _6011_/Y _6164_/X VGND VGND VPWR VPWR _6165_/X sky130_fd_sc_hd__o21ba_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3377_ _7124_/Q hold67/A _5353_/A _6940_/Q _3376_/X VGND VGND VPWR VPWR _3383_/A
+ sky130_fd_sc_hd__a221o_1
Xhold2025 _5286_/X VGND VGND VPWR VPWR _6873_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2036 hold589/X VGND VGND VPWR VPWR _4074_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2047 _6957_/Q VGND VGND VPWR VPWR hold663/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1302 hold151/X VGND VGND VPWR VPWR _3978_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1313 _6562_/Q VGND VGND VPWR VPWR hold870/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5116_ _5110_/Y _5113_/Y _5115_/X VGND VGND VPWR VPWR _5119_/C sky130_fd_sc_hd__o21ai_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2058 _5188_/X VGND VGND VPWR VPWR _6792_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2069 _6513_/Q VGND VGND VPWR VPWR hold354/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1324 hold269/X VGND VGND VPWR VPWR _4314_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6096_ _6904_/Q _5985_/X _5994_/X _7064_/Q _6094_/X VGND VGND VPWR VPWR _6096_/X
+ sky130_fd_sc_hd__a221o_1
Xhold1335 _4272_/X VGND VGND VPWR VPWR _6705_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1346 hold872/X VGND VGND VPWR VPWR hold271/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1357 _6945_/Q VGND VGND VPWR VPWR hold190/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1368 hold358/X VGND VGND VPWR VPWR _5451_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5047_ _5047_/A _5126_/A _5047_/C VGND VGND VPWR VPWR _5110_/A sky130_fd_sc_hd__and3_1
XFILLER_26_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1379 _5264_/X VGND VGND VPWR VPWR _6853_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6998_ _7137_/CLK _6998_/D fanout473/X VGND VGND VPWR VPWR _6998_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_41_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5949_ _6608_/Q _5684_/X _5686_/X _6623_/Q VGND VGND VPWR VPWR _5949_/X sky130_fd_sc_hd__a22o_1
XFILLER_40_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1880 hold425/X VGND VGND VPWR VPWR _5394_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1891 hold653/X VGND VGND VPWR VPWR _4335_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3300_ _3349_/A _3338_/A VGND VGND VPWR VPWR _5416_/A sky130_fd_sc_hd__nor2_8
X_4280_ _4280_/A hold13/A VGND VGND VPWR VPWR _4285_/S sky130_fd_sc_hd__and2_2
X_3231_ _6912_/Q VGND VGND VPWR VPWR _3231_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6921_ _7105_/CLK _6921_/D fanout473/X VGND VGND VPWR VPWR _6921_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6852_ _7131_/CLK hold41/X fanout469/X VGND VGND VPWR VPWR _6852_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5803_ _7066_/Q _5671_/X _5799_/X _5801_/X _5802_/X VGND VGND VPWR VPWR _5803_/X
+ sky130_fd_sc_hd__a2111o_1
X_6783_ _6788_/CLK _6783_/D _3959_/B VGND VGND VPWR VPWR _6783_/Q sky130_fd_sc_hd__dfstp_4
X_3995_ hold411/X _5503_/A1 _3999_/S VGND VGND VPWR VPWR _6476_/D sky130_fd_sc_hd__mux2_1
XFILLER_167_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5734_ _7031_/Q _5655_/X _5678_/B _6967_/Q _5707_/B VGND VGND VPWR VPWR _5734_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5665_ _5689_/A _5684_/B _5676_/B VGND VGND VPWR VPWR _5929_/B sky130_fd_sc_hd__and3_4
XFILLER_148_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4616_ _4616_/A _4616_/B _5063_/B VGND VGND VPWR VPWR _4616_/X sky130_fd_sc_hd__and3_1
XFILLER_190_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5596_ _7142_/Q _7143_/Q VGND VGND VPWR VPWR _5641_/B sky130_fd_sc_hd__nand2_1
XFILLER_191_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold410 hold410/A VGND VGND VPWR VPWR hold410/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold421 _5218_/X VGND VGND VPWR VPWR _5219_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4547_ _4625_/B _4607_/B VGND VGND VPWR VPWR _4770_/A sky130_fd_sc_hd__nand2_1
Xhold432 _6800_/Q VGND VGND VPWR VPWR hold432/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold443 hold443/A VGND VGND VPWR VPWR hold443/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold454 hold454/A VGND VGND VPWR VPWR hold454/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold465 hold465/A VGND VGND VPWR VPWR hold465/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold476 hold476/A VGND VGND VPWR VPWR hold476/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4478_ _4724_/C _4611_/A VGND VGND VPWR VPWR _5034_/A sky130_fd_sc_hd__nand2_2
Xhold487 hold487/A VGND VGND VPWR VPWR hold487/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold498 hold498/A VGND VGND VPWR VPWR hold498/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6217_ _6217_/A1 _5730_/S _6215_/X _6216_/X VGND VGND VPWR VPWR _6217_/X sky130_fd_sc_hd__o22a_1
X_3429_ _3429_/A hold66/X _3430_/B VGND VGND VPWR VPWR _5229_/B sky130_fd_sc_hd__and3_2
X_7197_ _7204_/CLK _7197_/D fanout484/X VGND VGND VPWR VPWR hold73/A sky130_fd_sc_hd__dfrtp_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6148_ _6858_/Q _5983_/X _6005_/X _6946_/Q VGND VGND VPWR VPWR _6148_/X sky130_fd_sc_hd__a22o_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1110 hold410/X VGND VGND VPWR VPWR _5297_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_161_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1121 hold407/X VGND VGND VPWR VPWR _5369_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_161_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1132 _6891_/Q VGND VGND VPWR VPWR hold392/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1143 _5522_/X VGND VGND VPWR VPWR _7083_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_161_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6079_ _7127_/Q _5973_/X _5988_/X _6871_/Q _6078_/X VGND VGND VPWR VPWR _6079_/X
+ sky130_fd_sc_hd__a221o_1
Xhold1154 _5315_/X VGND VGND VPWR VPWR _6899_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1165 hold194/X VGND VGND VPWR VPWR _4118_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1176 _6441_/Q VGND VGND VPWR VPWR hold93/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1187 _6875_/Q VGND VGND VPWR VPWR hold382/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1198 _6938_/Q VGND VGND VPWR VPWR hold459/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3780_ _6837_/Q hold27/A _5202_/A _6804_/Q _3779_/X VGND VGND VPWR VPWR _3783_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5450_ _5450_/A0 _5576_/A1 _5451_/S VGND VGND VPWR VPWR _5450_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4401_ _4495_/B _4454_/A VGND VGND VPWR VPWR _4625_/A sky130_fd_sc_hd__nor2_8
X_5381_ _5381_/A0 _5561_/A1 _5388_/S VGND VGND VPWR VPWR _5381_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7120_ _7126_/CLK _7120_/D fanout475/X VGND VGND VPWR VPWR _7120_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4332_ _4332_/A0 _5249_/A1 _4333_/S VGND VGND VPWR VPWR _4332_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7051_ _7131_/CLK _7051_/D fanout469/X VGND VGND VPWR VPWR _7051_/Q sky130_fd_sc_hd__dfrtp_4
X_4263_ _4263_/A0 _5221_/A1 _4267_/S VGND VGND VPWR VPWR _6697_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6002_ _5637_/A _6001_/X _6000_/X _5992_/X _6019_/B VGND VGND VPWR VPWR _6002_/X
+ sky130_fd_sc_hd__a2111o_1
X_3214_ _7040_/Q VGND VGND VPWR VPWR _3214_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4194_ _4194_/A _5229_/C VGND VGND VPWR VPWR _4199_/S sky130_fd_sc_hd__and2_4
XFILLER_67_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6904_ _7140_/CLK _6904_/D fanout469/X VGND VGND VPWR VPWR _6904_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6835_ _7053_/CLK _6835_/D fanout452/X VGND VGND VPWR VPWR _6835_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6766_ _7183_/CLK _6766_/D _6346_/B VGND VGND VPWR VPWR _6766_/Q sky130_fd_sc_hd__dfrtp_1
X_3978_ wire1/X _3978_/A1 _3996_/S VGND VGND VPWR VPWR _3978_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5717_ _6878_/Q _5667_/X _5714_/X _5716_/X VGND VGND VPWR VPWR _5718_/C sky130_fd_sc_hd__a211o_1
XFILLER_164_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6697_ _6808_/CLK _6697_/D fanout440/X VGND VGND VPWR VPWR _6697_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_1__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _6658_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_136_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5648_ _6490_/Q _5643_/A _5647_/Y VGND VGND VPWR VPWR _5730_/S sky130_fd_sc_hd__a21o_4
XFILLER_108_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5579_ hold292/X hold153/X _5586_/S VGND VGND VPWR VPWR _5579_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold240 hold240/A VGND VGND VPWR VPWR wb_dat_o[11] sky130_fd_sc_hd__buf_12
Xhold251 hold251/A VGND VGND VPWR VPWR wb_dat_o[10] sky130_fd_sc_hd__buf_12
Xhold262 hold262/A VGND VGND VPWR VPWR hold262/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold273 hold273/A VGND VGND VPWR VPWR hold273/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold284 hold284/A VGND VGND VPWR VPWR hold284/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold295 hold295/A VGND VGND VPWR VPWR hold295/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 _6792_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 _5585_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_124 hold13/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_135 hold153/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_146 _5308_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 _5929_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_179 _6582_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput8 mask_rev_in[13] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4950_ _4955_/A _4955_/B _4955_/C _4955_/D _4949_/Y VGND VGND VPWR VPWR _4950_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_64_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3901_ _3921_/B VGND VGND VPWR VPWR _3901_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4881_ _4881_/A _4881_/B VGND VGND VPWR VPWR _4972_/B sky130_fd_sc_hd__and2_1
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6620_ _6750_/CLK _6620_/D fanout446/X VGND VGND VPWR VPWR _6620_/Q sky130_fd_sc_hd__dfrtp_4
X_3832_ _3832_/A _3840_/B VGND VGND VPWR VPWR _3833_/B sky130_fd_sc_hd__nand2_1
X_6551_ _6648_/CLK _6551_/D _6426_/A VGND VGND VPWR VPWR _6551_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_192_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3763_ _6941_/Q _5362_/A _3509_/Y _6727_/Q _3762_/X VGND VGND VPWR VPWR _3769_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5502_ _5502_/A0 hold95/X _5505_/S VGND VGND VPWR VPWR _5502_/X sky130_fd_sc_hd__mux2_1
X_6482_ _6792_/CLK _6482_/D fanout442/X VGND VGND VPWR VPWR _6482_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_185_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3694_ _3694_/A _3694_/B _3694_/C _3694_/D VGND VGND VPWR VPWR _3704_/B sky130_fd_sc_hd__nor4_2
X_5433_ _5433_/A0 _5577_/A1 _5433_/S VGND VGND VPWR VPWR _7004_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput301 _3745_/Y VGND VGND VPWR VPWR reset sky130_fd_sc_hd__buf_12
Xoutput312 _7233_/X VGND VGND VPWR VPWR spimemio_flash_io3_di sky130_fd_sc_hd__buf_12
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput323 hold819/X VGND VGND VPWR VPWR hold205/A sky130_fd_sc_hd__buf_6
XFILLER_160_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput334 hold1338/X VGND VGND VPWR VPWR hold245/A sky130_fd_sc_hd__buf_6
X_5364_ hold780/X _5580_/A1 _5370_/S VGND VGND VPWR VPWR _6942_/D sky130_fd_sc_hd__mux2_1
Xoutput345 hold835/X VGND VGND VPWR VPWR hold259/A sky130_fd_sc_hd__buf_6
XFILLER_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7103_ _7103_/CLK _7103_/D fanout472/X VGND VGND VPWR VPWR _7103_/Q sky130_fd_sc_hd__dfrtp_2
X_4315_ hold97/X hold95/X _4315_/S VGND VGND VPWR VPWR hold98/A sky130_fd_sc_hd__mux2_1
XFILLER_99_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5295_ _5295_/A0 _5583_/A1 _5298_/S VGND VGND VPWR VPWR _5295_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7034_ _7035_/CLK _7034_/D fanout455/X VGND VGND VPWR VPWR _7034_/Q sky130_fd_sc_hd__dfrtp_4
X_4246_ _4246_/A0 _5556_/A1 _4249_/S VGND VGND VPWR VPWR _6672_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4177_ _4177_/A0 _5221_/A1 _4181_/S VGND VGND VPWR VPWR _4177_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6818_ _7111_/CLK _6818_/D fanout472/X VGND VGND VPWR VPWR _6818_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6749_ _6749_/CLK _6749_/D fanout440/X VGND VGND VPWR VPWR _6749_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4100_ _3737_/Y hold834/A _4106_/S VGND VGND VPWR VPWR _6554_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5080_ _5080_/A _5080_/B _5080_/C VGND VGND VPWR VPWR _5143_/A sky130_fd_sc_hd__and3_1
Xhold1709 _6797_/Q VGND VGND VPWR VPWR hold173/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4031_ hold215/X hold153/X _4056_/C VGND VGND VPWR VPWR _4031_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5982_ _6014_/A _6007_/C _6016_/C VGND VGND VPWR VPWR _5982_/X sky130_fd_sc_hd__and3_4
XFILLER_52_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4933_ _4374_/Y _5127_/A _4933_/C VGND VGND VPWR VPWR _5044_/C sky130_fd_sc_hd__and3b_1
XFILLER_178_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4864_ _5049_/B _4913_/A _4928_/C _4864_/D VGND VGND VPWR VPWR _4864_/X sky130_fd_sc_hd__and4_1
XFILLER_178_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_13 _3385_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_24 _3795_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6603_ _6794_/CLK _6603_/D fanout444/X VGND VGND VPWR VPWR _6603_/Q sky130_fd_sc_hd__dfrtp_4
X_3815_ _6657_/Q _3903_/A VGND VGND VPWR VPWR _3840_/B sky130_fd_sc_hd__nand2_2
XFILLER_193_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_35 _5678_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 _5990_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4795_ _4464_/Y _4570_/D _4713_/Y _4947_/A VGND VGND VPWR VPWR _4796_/C sky130_fd_sc_hd__o22a_1
XANTENNA_57 _6214_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6534_ _6747_/CLK _6534_/D fanout443/X VGND VGND VPWR VPWR _6534_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA_68 _6625_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3746_ _6981_/Q _5407_/A _4280_/A _6712_/Q VGND VGND VPWR VPWR _3746_/X sky130_fd_sc_hd__a22o_1
XANTENNA_79 input14/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6465_ _6656_/CLK _6465_/D _6415_/X VGND VGND VPWR VPWR _6465_/Q sky130_fd_sc_hd__dfrtp_4
X_3677_ _3676_/X _3677_/A1 _3739_/S VGND VGND VPWR VPWR _6776_/D sky130_fd_sc_hd__mux2_1
X_5416_ _5416_/A _5569_/B VGND VGND VPWR VPWR _5424_/S sky130_fd_sc_hd__and2_4
XFILLER_133_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6396_ _6399_/A _6423_/B VGND VGND VPWR VPWR _6396_/X sky130_fd_sc_hd__and2_1
XFILLER_88_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5347_ _5347_/A0 _5572_/A1 _5352_/S VGND VGND VPWR VPWR _5347_/X sky130_fd_sc_hd__mux2_1
Xoutput175 _3948_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[0] sky130_fd_sc_hd__buf_12
Xoutput186 _3947_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[1] sky130_fd_sc_hd__buf_12
Xoutput197 _3237_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[2] sky130_fd_sc_hd__buf_12
XFILLER_88_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5278_ _5278_/A0 _5503_/A1 _5280_/S VGND VGND VPWR VPWR _5278_/X sky130_fd_sc_hd__mux2_1
X_7017_ _7121_/CLK _7017_/D fanout468/X VGND VGND VPWR VPWR _7017_/Q sky130_fd_sc_hd__dfrtp_4
X_4229_ hold237/X _5518_/A1 _4239_/S VGND VGND VPWR VPWR _4229_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_824 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout380 hold20/X VGND VGND VPWR VPWR _5575_/A1 sky130_fd_sc_hd__buf_6
Xfanout391 _5249_/A1 VGND VGND VPWR VPWR _5555_/A1 sky130_fd_sc_hd__buf_12
XFILLER_93_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3600_ _6798_/Q _3319_/Y _3357_/Y _6482_/Q VGND VGND VPWR VPWR _3600_/X sky130_fd_sc_hd__a22o_2
XFILLER_174_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput11 mask_rev_in[16] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput22 mask_rev_in[26] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4580_ _4582_/A _4607_/B VGND VGND VPWR VPWR _4580_/Y sky130_fd_sc_hd__nand2_2
Xinput33 mask_rev_in[7] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput44 mgmt_gpio_in[17] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__clkbuf_2
Xinput55 mgmt_gpio_in[27] VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__clkbuf_4
X_3531_ _3553_/A _3531_/B VGND VGND VPWR VPWR _4322_/A sky130_fd_sc_hd__nor2_8
Xinput66 mgmt_gpio_in[37] VGND VGND VPWR VPWR _7233_/A sky130_fd_sc_hd__buf_4
Xinput77 ser_tx VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__clkbuf_2
Xhold806 hold806/A VGND VGND VPWR VPWR hold806/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold817 hold817/A VGND VGND VPWR VPWR hold817/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput88 spimemio_flash_io1_oeb VGND VGND VPWR VPWR _3962_/B sky130_fd_sc_hd__buf_4
Xhold828 hold828/A VGND VGND VPWR VPWR hold828/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput99 wb_adr_i[0] VGND VGND VPWR VPWR _4637_/B sky130_fd_sc_hd__buf_12
X_6250_ _6743_/Q _6014_/X _6244_/X _6249_/X VGND VGND VPWR VPWR _6255_/A sky130_fd_sc_hd__a211o_1
Xhold839 hold839/A VGND VGND VPWR VPWR hold839/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3462_ _3462_/A _3462_/B VGND VGND VPWR VPWR _3462_/Y sky130_fd_sc_hd__nand2_8
XFILLER_143_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5201_ hold686/X _5552_/A1 _5201_/S VGND VGND VPWR VPWR _5201_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6181_ _6979_/Q _5976_/B _5977_/X _7139_/Q _6180_/X VGND VGND VPWR VPWR _6181_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_124_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3393_ _7131_/Q _5569_/A _5236_/C input69/X VGND VGND VPWR VPWR _3393_/X sky130_fd_sc_hd__a22o_1
X_5132_ _4947_/B _4510_/B _4570_/A VGND VGND VPWR VPWR _5132_/X sky130_fd_sc_hd__a21o_1
Xhold2207 _6950_/Q VGND VGND VPWR VPWR hold684/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2218 _5310_/X VGND VGND VPWR VPWR _6894_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2229 hold723/X VGND VGND VPWR VPWR _5454_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1506 hold510/X VGND VGND VPWR VPWR _5523_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1517 hold209/X VGND VGND VPWR VPWR hold821/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5063_ _5063_/A _5063_/B _5063_/C _5063_/D VGND VGND VPWR VPWR _5155_/B sky130_fd_sc_hd__and4_1
Xhold1528 _5568_/X VGND VGND VPWR VPWR _7124_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1539 _6547_/Q VGND VGND VPWR VPWR hold830/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4014_ _4014_/A0 hold153/X _4047_/C VGND VGND VPWR VPWR _4014_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5965_ _6736_/Q _5656_/X _5679_/X _6593_/Q _5964_/X VGND VGND VPWR VPWR _5965_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_40_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4916_ _4969_/A _4652_/Y _4676_/Y _4633_/B VGND VGND VPWR VPWR _5047_/C sky130_fd_sc_hd__o22a_1
X_5896_ _6698_/Q _5672_/X _5679_/X _6590_/Q _5883_/X VGND VGND VPWR VPWR _5896_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_33_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4847_ _4638_/Y _4688_/B _5098_/A VGND VGND VPWR VPWR _4871_/A sky130_fd_sc_hd__o21a_1
XFILLER_166_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4778_ _4569_/B _4510_/B _4729_/A _4688_/A VGND VGND VPWR VPWR _4800_/B sky130_fd_sc_hd__o22a_1
XFILLER_5_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3729_ _6998_/Q _5425_/A _4268_/A _6703_/Q VGND VGND VPWR VPWR _3729_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6517_ _6522_/CLK _6517_/D fanout478/X VGND VGND VPWR VPWR _6517_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6448_ _6658_/CLK _6448_/D _6403_/X VGND VGND VPWR VPWR _6448_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_161_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6379_ _6684_/Q _6379_/A2 _6379_/B1 _6685_/Q VGND VGND VPWR VPWR _6379_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5750_ _5750_/A1 _3924_/Y _5647_/Y VGND VGND VPWR VPWR _5750_/X sky130_fd_sc_hd__o21ba_1
XFILLER_97_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4701_ _4701_/A _4701_/B VGND VGND VPWR VPWR _4826_/B sky130_fd_sc_hd__nor2_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5681_ _5689_/A _5684_/B _5689_/C VGND VGND VPWR VPWR _5681_/X sky130_fd_sc_hd__and3_4
X_4632_ _4594_/A _4463_/B _4568_/Y _4837_/B _4631_/X VGND VGND VPWR VPWR _4632_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_147_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4563_ _4615_/B _4693_/B VGND VGND VPWR VPWR _4922_/A sky130_fd_sc_hd__nand2_1
XFILLER_144_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold603 _5291_/X VGND VGND VPWR VPWR _6877_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold614 hold614/A VGND VGND VPWR VPWR hold614/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6302_ _6607_/Q _5982_/X _5992_/X _6710_/Q VGND VGND VPWR VPWR _6302_/X sky130_fd_sc_hd__a22o_1
X_3514_ _6913_/Q _5326_/A _5335_/A _6921_/Q _3513_/X VGND VGND VPWR VPWR _3515_/D
+ sky130_fd_sc_hd__a221o_1
Xhold625 hold625/A VGND VGND VPWR VPWR hold625/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4494_ _4652_/B _4560_/A VGND VGND VPWR VPWR _4840_/A sky130_fd_sc_hd__and2b_2
Xhold636 hold636/A VGND VGND VPWR VPWR hold636/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold647 hold647/A VGND VGND VPWR VPWR hold647/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold658 hold658/A VGND VGND VPWR VPWR hold658/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap366 _4579_/B VGND VGND VPWR VPWR _4598_/A sky130_fd_sc_hd__clkbuf_4
X_6233_ _6712_/Q _5973_/X _5988_/X _6569_/Q _6232_/X VGND VGND VPWR VPWR _6233_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold669 hold669/A VGND VGND VPWR VPWR hold669/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3445_ _7130_/Q _5569_/A _5353_/A _6938_/Q VGND VGND VPWR VPWR _3445_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2004 _7001_/Q VGND VGND VPWR VPWR hold542/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6164_ _6155_/X _6339_/B _6164_/C _6164_/D VGND VGND VPWR VPWR _6164_/X sky130_fd_sc_hd__and4b_2
XFILLER_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _7116_/Q _5551_/A _3339_/Y _6478_/Q VGND VGND VPWR VPWR _3376_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2015 _7080_/Q VGND VGND VPWR VPWR hold707/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2026 _7055_/Q VGND VGND VPWR VPWR hold337/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2037 _4074_/X VGND VGND VPWR VPWR _6532_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5115_ _5115_/A _5115_/B _5124_/C _5126_/C VGND VGND VPWR VPWR _5115_/X sky130_fd_sc_hd__and4_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2048 hold663/X VGND VGND VPWR VPWR _5381_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1303 _3978_/X VGND VGND VPWR VPWR hold152/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2059 _6632_/Q VGND VGND VPWR VPWR hold615/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1314 hold870/X VGND VGND VPWR VPWR hold246/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6095_ _7056_/Q _5990_/X _5996_/X _7048_/Q VGND VGND VPWR VPWR _6095_/X sky130_fd_sc_hd__a22o_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1325 _6535_/Q VGND VGND VPWR VPWR hold427/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1336 _7191_/Q VGND VGND VPWR VPWR hold871/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1347 hold271/X VGND VGND VPWR VPWR hold1347/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5046_ _5046_/A _5046_/B _5046_/C VGND VGND VPWR VPWR _5123_/B sky130_fd_sc_hd__and3_1
Xhold1358 hold190/X VGND VGND VPWR VPWR _5367_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1369 _6820_/Q VGND VGND VPWR VPWR hold248/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6997_ _7109_/CLK _6997_/D fanout452/X VGND VGND VPWR VPWR _6997_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_43_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5948_ _5969_/A1 _6342_/S _5946_/X _5947_/X VGND VGND VPWR VPWR _7171_/D sky130_fd_sc_hd__o22a_1
XFILLER_34_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5879_ _5879_/A _5879_/B _5879_/C _5879_/D VGND VGND VPWR VPWR _5879_/Y sky130_fd_sc_hd__nor4_1
XFILLER_21_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1870 hold578/X VGND VGND VPWR VPWR _4336_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1881 _7032_/Q VGND VGND VPWR VPWR hold509/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1892 _6759_/Q VGND VGND VPWR VPWR hold307/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3230_ _6920_/Q VGND VGND VPWR VPWR _3230_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6920_ _7123_/CLK _6920_/D fanout477/X VGND VGND VPWR VPWR _6920_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_63_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6851_ _7123_/CLK _6851_/D fanout479/X VGND VGND VPWR VPWR _6851_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_62_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5802_ _7002_/Q _5666_/X _5689_/X _7082_/Q VGND VGND VPWR VPWR _5802_/X sky130_fd_sc_hd__a22o_1
X_6782_ _6793_/CLK _6782_/D _3959_/B VGND VGND VPWR VPWR _6782_/Q sky130_fd_sc_hd__dfrtp_4
X_3994_ hold18/X hold875/X _3996_/S VGND VGND VPWR VPWR _3994_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5733_ _6999_/Q _5666_/X _5689_/X _7079_/Q _5732_/X VGND VGND VPWR VPWR _5733_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5664_ _5689_/A _5689_/B _5688_/C VGND VGND VPWR VPWR _5664_/X sky130_fd_sc_hd__and3_4
XFILLER_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_54_csclk _7093_/CLK VGND VGND VPWR VPWR _7084_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_129_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4615_ _4625_/A _4615_/B VGND VGND VPWR VPWR _5063_/B sky130_fd_sc_hd__nand2_2
X_5595_ _5595_/A0 _5593_/Y _5599_/D VGND VGND VPWR VPWR _7142_/D sky130_fd_sc_hd__mux2_1
Xhold400 _4061_/X VGND VGND VPWR VPWR _6521_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold411 hold411/A VGND VGND VPWR VPWR hold411/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4546_ _4569_/A _4601_/A _4543_/X _4544_/Y _4898_/A VGND VGND VPWR VPWR _4546_/X
+ sky130_fd_sc_hd__o2111a_1
Xhold422 hold422/A VGND VGND VPWR VPWR hold422/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold433 hold433/A VGND VGND VPWR VPWR hold433/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold444 _6537_/Q VGND VGND VPWR VPWR hold444/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold455 hold455/A VGND VGND VPWR VPWR hold455/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4477_ _4477_/A _4477_/B _4477_/C VGND VGND VPWR VPWR _4477_/Y sky130_fd_sc_hd__nand3_4
Xhold466 hold466/A VGND VGND VPWR VPWR hold466/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold477 hold477/A VGND VGND VPWR VPWR hold477/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold488 _5402_/X VGND VGND VPWR VPWR _6976_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3428_ _7172_/Q _6813_/Q _6815_/Q VGND VGND VPWR VPWR _3428_/X sky130_fd_sc_hd__mux2_4
Xclkbuf_leaf_69_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6794_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold499 hold499/A VGND VGND VPWR VPWR hold499/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6216_ _7179_/Q _3924_/Y _5647_/Y VGND VGND VPWR VPWR _6216_/X sky130_fd_sc_hd__o21ba_1
X_7196_ _7204_/CLK _7196_/D fanout484/X VGND VGND VPWR VPWR _7196_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_38_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6147_ _6994_/Q _6014_/X _6145_/X _6146_/X VGND VGND VPWR VPWR _6152_/A sky130_fd_sc_hd__a211o_1
X_3359_ _6908_/Q _5317_/A _5461_/A _7036_/Q VGND VGND VPWR VPWR _3359_/X sky130_fd_sc_hd__a22o_1
Xhold1100 _6955_/Q VGND VGND VPWR VPWR hold402/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1111 _5297_/X VGND VGND VPWR VPWR _6883_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 _5369_/X VGND VGND VPWR VPWR _6947_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1133 hold392/X VGND VGND VPWR VPWR _5306_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_100_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6078_ _6959_/Q _5992_/X _6012_/X _6999_/Q _6077_/X VGND VGND VPWR VPWR _6078_/X
+ sky130_fd_sc_hd__a221o_1
Xhold1144 _6931_/Q VGND VGND VPWR VPWR hold370/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1155 _7091_/Q VGND VGND VPWR VPWR hold380/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1166 _4118_/X VGND VGND VPWR VPWR _6570_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1177 hold93/X VGND VGND VPWR VPWR _3986_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5029_ _4417_/B _4648_/Y _4584_/Y VGND VGND VPWR VPWR _5029_/X sky130_fd_sc_hd__o21a_1
XFILLER_26_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1188 hold382/X VGND VGND VPWR VPWR _5288_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1199 hold459/X VGND VGND VPWR VPWR _5359_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_782 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2390 _6519_/Q VGND VGND VPWR VPWR hold2390/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4400_ _4575_/C _4594_/A VGND VGND VPWR VPWR _4454_/A sky130_fd_sc_hd__nand2_8
X_5380_ _5380_/A _5569_/B VGND VGND VPWR VPWR _5388_/S sky130_fd_sc_hd__and2_4
XFILLER_126_662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4331_ hold270/X _5581_/A1 _4333_/S VGND VGND VPWR VPWR _4331_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7050_ _7124_/CLK _7050_/D fanout459/X VGND VGND VPWR VPWR _7050_/Q sky130_fd_sc_hd__dfrtp_4
X_4262_ _4262_/A _5229_/C VGND VGND VPWR VPWR _4267_/S sky130_fd_sc_hd__and2_4
XFILLER_113_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6001_ _6015_/B _6018_/B _6019_/C _6019_/A VGND VGND VPWR VPWR _6001_/X sky130_fd_sc_hd__a22o_1
X_3213_ _7048_/Q VGND VGND VPWR VPWR _3213_/Y sky130_fd_sc_hd__clkinv_2
X_4193_ _4193_/A0 _5196_/A1 _4193_/S VGND VGND VPWR VPWR _6633_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6903_ _6903_/CLK hold3/X fanout460/X VGND VGND VPWR VPWR _6903_/Q sky130_fd_sc_hd__dfrtp_4
X_6834_ _7116_/CLK _6834_/D fanout457/X VGND VGND VPWR VPWR _6834_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6765_ _7183_/CLK _6765_/D _6346_/B VGND VGND VPWR VPWR _6765_/Q sky130_fd_sc_hd__dfrtp_1
X_3977_ _3977_/A _5229_/C VGND VGND VPWR VPWR _3987_/S sky130_fd_sc_hd__and2_2
XFILLER_10_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5716_ _6846_/Q _5842_/A2 _5682_/X _7038_/Q _5715_/X VGND VGND VPWR VPWR _5716_/X
+ sky130_fd_sc_hd__a221o_1
X_6696_ _6750_/CLK _6696_/D fanout446/X VGND VGND VPWR VPWR _6696_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5647_ _6490_/Q _5647_/B VGND VGND VPWR VPWR _5647_/Y sky130_fd_sc_hd__nor2_8
XFILLER_164_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5578_ hold33/X hold13/A VGND VGND VPWR VPWR _5586_/S sky130_fd_sc_hd__and2_4
Xhold230 hold230/A VGND VGND VPWR VPWR wb_dat_o[0] sky130_fd_sc_hd__buf_12
XFILLER_117_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold241 hold241/A VGND VGND VPWR VPWR hold241/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold252 hold252/A VGND VGND VPWR VPWR hold252/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4529_ _4396_/X _4529_/B _5151_/D _4529_/D VGND VGND VPWR VPWR _4529_/X sky130_fd_sc_hd__and4b_1
Xhold263 hold263/A VGND VGND VPWR VPWR hold839/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold274 hold274/A VGND VGND VPWR VPWR hold847/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold285 hold285/A VGND VGND VPWR VPWR hold861/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold296 hold296/A VGND VGND VPWR VPWR hold296/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7179_ _3950_/A1 _7179_/D fanout482/X VGND VGND VPWR VPWR _7179_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 _6785_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_114 _5503_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_125 _5872_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_136 hold153/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 hold27/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_158 _5670_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_169 _6599_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput9 mask_rev_in[14] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__buf_2
XFILLER_36_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3900_ _4395_/A _3900_/B _3900_/C _3900_/D VGND VGND VPWR VPWR _3921_/B sky130_fd_sc_hd__nand4b_4
XFILLER_51_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4880_ _5127_/A _4880_/B VGND VGND VPWR VPWR _4965_/C sky130_fd_sc_hd__and2_1
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3831_ _3830_/Y _3831_/B _3835_/S VGND VGND VPWR VPWR _3833_/A sky130_fd_sc_hd__and3b_1
XFILLER_177_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3762_ _7125_/Q _5569_/A _4268_/A _6702_/Q VGND VGND VPWR VPWR _3762_/X sky130_fd_sc_hd__a22o_1
X_6550_ _6750_/CLK _6550_/D fanout446/X VGND VGND VPWR VPWR _6550_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_9_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5501_ hold708/X _5582_/A1 _5505_/S VGND VGND VPWR VPWR _5501_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6481_ _6792_/CLK _6481_/D fanout442/X VGND VGND VPWR VPWR _6481_/Q sky130_fd_sc_hd__dfstp_4
X_3693_ _7102_/Q _3311_/Y _4140_/A _6590_/Q _3692_/X VGND VGND VPWR VPWR _3694_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_145_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5432_ _5432_/A0 _5585_/A1 _5433_/S VGND VGND VPWR VPWR _5432_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput302 _3970_/X VGND VGND VPWR VPWR ser_rx sky130_fd_sc_hd__buf_12
XFILLER_145_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput313 _7186_/Q VGND VGND VPWR VPWR wb_ack_o sky130_fd_sc_hd__buf_12
X_5363_ hold593/X _5561_/A1 _5370_/S VGND VGND VPWR VPWR _5363_/X sky130_fd_sc_hd__mux2_1
Xoutput324 hold821/X VGND VGND VPWR VPWR hold210/A sky130_fd_sc_hd__buf_6
XFILLER_114_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput335 hold1270/X VGND VGND VPWR VPWR hold212/A sky130_fd_sc_hd__buf_6
X_7102_ _7102_/CLK _7102_/D _6409_/A VGND VGND VPWR VPWR _7102_/Q sky130_fd_sc_hd__dfstp_2
X_4314_ _4314_/A0 _5303_/A1 _4315_/S VGND VGND VPWR VPWR _6740_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5294_ _5294_/A0 _5555_/A1 _5298_/S VGND VGND VPWR VPWR _5294_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4245_ _4245_/A0 _5582_/A1 _4249_/S VGND VGND VPWR VPWR _4245_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7033_ _7102_/CLK _7033_/D _6409_/A VGND VGND VPWR VPWR _7033_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4176_ _4176_/A _5229_/C VGND VGND VPWR VPWR _4181_/S sky130_fd_sc_hd__and2_4
XFILLER_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6817_ _6817_/CLK _6817_/D fanout445/X VGND VGND VPWR VPWR _6817_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6748_ _6757_/CLK _6748_/D fanout446/X VGND VGND VPWR VPWR _6748_/Q sky130_fd_sc_hd__dfrtp_4
Xwire429 _4649_/Y VGND VGND VPWR VPWR _4684_/A sky130_fd_sc_hd__buf_2
XFILLER_109_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6679_ _7152_/CLK _6679_/D _6346_/B VGND VGND VPWR VPWR _6679_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_152_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmgmt_gpio_14_buff_inst _3950_/X VGND VGND VPWR VPWR mgmt_gpio_out[14] sky130_fd_sc_hd__clkbuf_8
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4030_ _3343_/A wire438/X _4012_/X _4056_/C _5569_/B VGND VGND VPWR VPWR _4046_/S
+ sky130_fd_sc_hd__o221a_4
XFILLER_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5981_ _7153_/Q _7154_/Q VGND VGND VPWR VPWR _6016_/C sky130_fd_sc_hd__and2b_4
XFILLER_18_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4932_ _4925_/X _4931_/X _5115_/A VGND VGND VPWR VPWR _4932_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4863_ _4655_/A _4640_/Y _4655_/B _4704_/C VGND VGND VPWR VPWR _4864_/D sky130_fd_sc_hd__o31a_1
X_6602_ _6691_/CLK _6602_/D fanout444/X VGND VGND VPWR VPWR _6602_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_14 _3385_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_25 _5289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3814_ _3814_/A _3814_/B VGND VGND VPWR VPWR _6468_/D sky130_fd_sc_hd__xnor2_1
XFILLER_177_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_36 _5707_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4794_ _4729_/A _4712_/Y _4789_/X _4793_/X _5095_/A VGND VGND VPWR VPWR _4796_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_119_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_47 _5991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 _6295_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6533_ _6794_/CLK _6533_/D fanout444/X VGND VGND VPWR VPWR _6533_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA_69 _7096_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3745_ _3745_/A VGND VGND VPWR VPWR _3745_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6464_ _6656_/CLK _6464_/D _6414_/X VGND VGND VPWR VPWR _6464_/Q sky130_fd_sc_hd__dfrtp_4
X_3676_ _3739_/A1 _3675_/Y _3738_/S VGND VGND VPWR VPWR _3676_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5415_ _5415_/A0 _5559_/A1 _5415_/S VGND VGND VPWR VPWR _6988_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6395_ _6399_/A _6423_/B VGND VGND VPWR VPWR _6395_/X sky130_fd_sc_hd__and2_1
XFILLER_99_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5346_ _5346_/A0 _5571_/A1 _5352_/S VGND VGND VPWR VPWR _5346_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput176 _3230_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[10] sky130_fd_sc_hd__buf_12
Xoutput187 _3219_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[20] sky130_fd_sc_hd__buf_12
Xoutput198 _3209_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[30] sky130_fd_sc_hd__buf_12
XFILLER_99_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5277_ _5277_/A0 hold95/X _5280_/S VGND VGND VPWR VPWR _5277_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7016_ _7016_/CLK _7016_/D fanout475/X VGND VGND VPWR VPWR _7016_/Q sky130_fd_sc_hd__dfrtp_4
X_4228_ _4228_/A0 _4227_/X _4240_/S VGND VGND VPWR VPWR _6661_/D sky130_fd_sc_hd__mux2_1
XFILLER_46_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4159_ _4159_/A0 _5221_/A1 _4163_/S VGND VGND VPWR VPWR _6604_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_836 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout381 hold877/X VGND VGND VPWR VPWR hold878/A sky130_fd_sc_hd__buf_6
Xfanout392 _5267_/A1 VGND VGND VPWR VPWR _5249_/A1 sky130_fd_sc_hd__buf_8
XFILLER_47_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput12 mask_rev_in[17] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput23 mask_rev_in[27] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__buf_2
Xinput34 mask_rev_in[8] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput45 mgmt_gpio_in[18] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__buf_2
X_3530_ _3531_/B _3530_/B VGND VGND VPWR VPWR _4194_/A sky130_fd_sc_hd__nor2_8
Xinput56 mgmt_gpio_in[28] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__clkbuf_4
XFILLER_7_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold807 hold807/A VGND VGND VPWR VPWR hold807/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput67 mgmt_gpio_in[3] VGND VGND VPWR VPWR _3881_/C sky130_fd_sc_hd__buf_6
Xinput78 spi_csb VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__buf_4
XFILLER_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput89 spimemio_flash_io2_do VGND VGND VPWR VPWR input89/X sky130_fd_sc_hd__clkbuf_2
Xhold818 hold818/A VGND VGND VPWR VPWR hold818/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3461_ _3461_/A _3461_/B _3461_/C VGND VGND VPWR VPWR _3462_/B sky130_fd_sc_hd__and3_2
Xhold829 hold829/A VGND VGND VPWR VPWR hold829/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5200_ _5207_/A _5229_/B _5220_/C VGND VGND VPWR VPWR _5201_/S sky130_fd_sc_hd__and3_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3392_ _7185_/Q _6814_/Q _6815_/Q VGND VGND VPWR VPWR _3392_/X sky130_fd_sc_hd__mux2_8
X_6180_ _6931_/Q _5982_/X _6004_/X _6883_/Q VGND VGND VPWR VPWR _6180_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2208 _6589_/Q VGND VGND VPWR VPWR hold786/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5131_ _5131_/A _5131_/B _5131_/C VGND VGND VPWR VPWR _5134_/A sky130_fd_sc_hd__and3_1
Xhold2219 _6633_/Q VGND VGND VPWR VPWR hold465/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1507 _6612_/Q VGND VGND VPWR VPWR hold157/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5062_ _5062_/A VGND VGND VPWR VPWR _5135_/B sky130_fd_sc_hd__inv_2
Xhold1518 _6892_/Q VGND VGND VPWR VPWR hold504/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1529 _6805_/Q VGND VGND VPWR VPWR hold219/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4013_ _3648_/A _6432_/B _4012_/X _4047_/C _5569_/B VGND VGND VPWR VPWR _4029_/S
+ sky130_fd_sc_hd__o221a_4
XFILLER_65_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5964_ _6643_/Q _5655_/X _5663_/X _6633_/Q _5950_/Y VGND VGND VPWR VPWR _5964_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4915_ _5048_/A _4915_/B VGND VGND VPWR VPWR _5115_/B sky130_fd_sc_hd__nand2_1
XFILLER_178_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5895_ _6640_/Q _5655_/X _5656_/X _6733_/Q _5885_/Y VGND VGND VPWR VPWR _5895_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_33_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4846_ _4570_/C _4655_/A _4590_/Y _4691_/Y VGND VGND VPWR VPWR _4846_/X sky130_fd_sc_hd__o22a_1
XFILLER_193_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4777_ _4947_/A _4668_/Y _4531_/B VGND VGND VPWR VPWR _4777_/X sky130_fd_sc_hd__o21a_1
XFILLER_147_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6516_ _7138_/CLK hold7/X fanout480/X VGND VGND VPWR VPWR _6516_/Q sky130_fd_sc_hd__dfrtp_1
X_3728_ _6886_/Q _5299_/A _5497_/A _7062_/Q _3727_/X VGND VGND VPWR VPWR _3735_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_4_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6447_ _6656_/CLK _6447_/D _6402_/X VGND VGND VPWR VPWR _6447_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3659_ _7079_/Q _5515_/A hold67/A _7119_/Q _3658_/X VGND VGND VPWR VPWR _3664_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6378_ _6377_/X hold875/X _6384_/S VGND VGND VPWR VPWR _7200_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5329_ _5329_/A0 _5518_/A1 _5334_/S VGND VGND VPWR VPWR _6911_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4700_ _4718_/C _4751_/C VGND VGND VPWR VPWR _4701_/B sky130_fd_sc_hd__nand2_2
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ _5689_/A _5684_/B _5689_/C VGND VGND VPWR VPWR _5680_/X sky130_fd_sc_hd__and3b_4
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4631_ _4757_/A _4997_/A _4973_/C _4631_/D VGND VGND VPWR VPWR _4631_/X sky130_fd_sc_hd__and4_1
XFILLER_129_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4562_ _4562_/A _4693_/B VGND VGND VPWR VPWR _4894_/B sky130_fd_sc_hd__nand2_1
XFILLER_156_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6301_ _6755_/Q _5638_/X _6019_/X _6735_/Q _6300_/X VGND VGND VPWR VPWR _6304_/C
+ sky130_fd_sc_hd__a221o_1
Xhold604 hold604/A VGND VGND VPWR VPWR hold604/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold615 hold615/A VGND VGND VPWR VPWR hold615/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3513_ _7017_/Q _5443_/A _4212_/A _6653_/Q VGND VGND VPWR VPWR _3513_/X sky130_fd_sc_hd__a22o_1
Xhold626 hold626/A VGND VGND VPWR VPWR hold626/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4493_ _4649_/B _4639_/S VGND VGND VPWR VPWR _4652_/B sky130_fd_sc_hd__xnor2_2
Xhold637 hold637/A VGND VGND VPWR VPWR hold637/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold648 hold648/A VGND VGND VPWR VPWR hold648/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6232_ _6707_/Q _5992_/X _6012_/X _6747_/Q _6231_/X VGND VGND VPWR VPWR _6232_/X
+ sky130_fd_sc_hd__a221o_1
Xhold659 hold659/A VGND VGND VPWR VPWR hold659/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap367 _4579_/B VGND VGND VPWR VPWR _4473_/A sky130_fd_sc_hd__clkbuf_2
X_3444_ _3444_/A _3444_/B _3444_/C _3444_/D VGND VGND VPWR VPWR _3444_/Y sky130_fd_sc_hd__nor4_1
XFILLER_103_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3375_ _6892_/Q _5299_/A _5533_/A _7100_/Q _3374_/X VGND VGND VPWR VPWR _3384_/B
+ sky130_fd_sc_hd__a221o_2
X_6163_ _6163_/A _6163_/B _6163_/C _6163_/D VGND VGND VPWR VPWR _6164_/D sky130_fd_sc_hd__nor4_1
XFILLER_170_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2005 hold542/X VGND VGND VPWR VPWR _5430_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2016 hold707/X VGND VGND VPWR VPWR _5519_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2027 hold337/X VGND VGND VPWR VPWR _5491_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2038 _6733_/Q VGND VGND VPWR VPWR hold717/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _5114_/A _5114_/B _5114_/C VGND VGND VPWR VPWR _5126_/C sky130_fd_sc_hd__and3_1
XFILLER_57_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1304 hold152/X VGND VGND VPWR VPWR hold1304/X sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2049 _5381_/X VGND VGND VPWR VPWR _6957_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6094_ _6912_/Q _5991_/X _6018_/X _6968_/Q VGND VGND VPWR VPWR _6094_/X sky130_fd_sc_hd__a22o_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1315 hold246/X VGND VGND VPWR VPWR hold1315/X sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1326 _4078_/X VGND VGND VPWR VPWR hold428/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1337 hold871/X VGND VGND VPWR VPWR hold244/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1348 _7033_/Q VGND VGND VPWR VPWR hold187/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5045_ _4569_/B _4523_/Y _4583_/B _4688_/A VGND VGND VPWR VPWR _5046_/C sky130_fd_sc_hd__o22a_1
Xhold1359 _5367_/X VGND VGND VPWR VPWR _6945_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6996_ _7020_/CLK _6996_/D fanout458/X VGND VGND VPWR VPWR _6996_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5947_ _5947_/A1 _3924_/Y _5647_/Y VGND VGND VPWR VPWR _5947_/X sky130_fd_sc_hd__o21ba_1
XFILLER_159_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5878_ _6732_/Q _5656_/X _5663_/X _6629_/Q _5877_/X VGND VGND VPWR VPWR _5879_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4829_ _4454_/A _4719_/Y _4821_/X _4828_/X _4922_/B VGND VGND VPWR VPWR _4834_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_193_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1860 _6625_/Q VGND VGND VPWR VPWR hold569/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1871 _6848_/Q VGND VGND VPWR VPWR hold498/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_90_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1882 hold509/X VGND VGND VPWR VPWR _5465_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1893 _6772_/Q VGND VGND VPWR VPWR hold609/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_181_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6850_ _6850_/CLK _6850_/D fanout471/X VGND VGND VPWR VPWR _6850_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_62_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5801_ _7010_/Q _5686_/X _5796_/X _5800_/X VGND VGND VPWR VPWR _5801_/X sky130_fd_sc_hd__a211o_1
X_6781_ _6658_/CLK _6781_/D _6433_/X VGND VGND VPWR VPWR _6781_/Q sky130_fd_sc_hd__dfrtn_1
X_3993_ _3993_/A0 _5196_/A1 _3999_/S VGND VGND VPWR VPWR _6475_/D sky130_fd_sc_hd__mux2_1
X_5732_ _6991_/Q _5929_/B _5668_/X _7055_/Q _5731_/X VGND VGND VPWR VPWR _5732_/X
+ sky130_fd_sc_hd__a221o_1
X_5663_ _5689_/A _5684_/B _5688_/C VGND VGND VPWR VPWR _5663_/X sky130_fd_sc_hd__and3_4
X_4614_ _5073_/B _4614_/B _4614_/C _4614_/D VGND VGND VPWR VPWR _4614_/X sky130_fd_sc_hd__and4_1
XFILLER_175_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5594_ _5599_/D _5594_/B VGND VGND VPWR VPWR _5601_/A sky130_fd_sc_hd__nand2_1
XFILLER_175_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold401 hold401/A VGND VGND VPWR VPWR hold401/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4545_ _4625_/B _4724_/C VGND VGND VPWR VPWR _4898_/A sky130_fd_sc_hd__nand2_1
Xhold412 hold412/A VGND VGND VPWR VPWR hold412/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold423 hold423/A VGND VGND VPWR VPWR hold423/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold434 hold434/A VGND VGND VPWR VPWR hold434/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold445 hold445/A VGND VGND VPWR VPWR _6537_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold456 hold456/A VGND VGND VPWR VPWR hold456/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4476_ _4575_/C _4594_/A _4463_/B VGND VGND VPWR VPWR _4476_/X sky130_fd_sc_hd__a21o_2
Xhold467 hold467/A VGND VGND VPWR VPWR hold467/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold478 hold478/A VGND VGND VPWR VPWR hold478/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold489 hold489/A VGND VGND VPWR VPWR hold489/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6215_ _6844_/Q _6011_/Y _6214_/Y _6341_/S VGND VGND VPWR VPWR _6215_/X sky130_fd_sc_hd__o211a_2
XFILLER_132_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3427_ _3648_/B _3533_/B VGND VGND VPWR VPWR _3427_/Y sky130_fd_sc_hd__nor2_8
X_7195_ _7204_/CLK _7195_/D fanout484/X VGND VGND VPWR VPWR _7195_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6146_ _6906_/Q _5985_/X _5994_/X _7066_/Q _6144_/X VGND VGND VPWR VPWR _6146_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3358_ _7020_/Q _5443_/A _5506_/A _7076_/Q VGND VGND VPWR VPWR _3358_/X sky130_fd_sc_hd__a22o_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1101 hold402/X VGND VGND VPWR VPWR _5378_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1112 _7051_/Q VGND VGND VPWR VPWR hold371/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1123 _6438_/Q VGND VGND VPWR VPWR hold133/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1134 _5306_/X VGND VGND VPWR VPWR _6891_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_6077_ _6951_/Q _5997_/X _6004_/X _6879_/Q VGND VGND VPWR VPWR _6077_/X sky130_fd_sc_hd__a22o_1
XTAP_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3289_ _3322_/B _3430_/A VGND VGND VPWR VPWR _3764_/A sky130_fd_sc_hd__nand2_8
Xhold1145 hold370/X VGND VGND VPWR VPWR _5351_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1156 hold380/X VGND VGND VPWR VPWR _5531_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1167 _6728_/Q VGND VGND VPWR VPWR hold179/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5028_ _4417_/B _4688_/A _4800_/C _4898_/A VGND VGND VPWR VPWR _5148_/B sky130_fd_sc_hd__o211a_1
Xhold1178 _3986_/X VGND VGND VPWR VPWR hold107/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1189 _5288_/X VGND VGND VPWR VPWR _6875_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6979_ _7131_/CLK _6979_/D fanout469/X VGND VGND VPWR VPWR _6979_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_110_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold990 _5287_/X VGND VGND VPWR VPWR _6874_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_89_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2380 hold718/X VGND VGND VPWR VPWR _5565_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_64_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2391 _7129_/Q VGND VGND VPWR VPWR hold726/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1690 _7187_/Q VGND VGND VPWR VPWR hold848/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4330_ _4330_/A0 _5193_/A1 _4333_/S VGND VGND VPWR VPWR _4330_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4261_ _4261_/A0 _4339_/A1 _4261_/S VGND VGND VPWR VPWR _4261_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6000_ _5637_/A _6014_/A _6019_/C _5984_/X _5998_/X VGND VGND VPWR VPWR _6000_/X
+ sky130_fd_sc_hd__a311o_1
X_3212_ _7056_/Q VGND VGND VPWR VPWR _3212_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4192_ _4192_/A0 _5195_/A1 _4193_/S VGND VGND VPWR VPWR _6632_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6902_ _7127_/CLK _6902_/D fanout477/X VGND VGND VPWR VPWR _6902_/Q sky130_fd_sc_hd__dfstp_2
X_6833_ _6833_/CLK _6833_/D fanout454/X VGND VGND VPWR VPWR _6833_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6764_ _7183_/CLK _6764_/D _6346_/B VGND VGND VPWR VPWR _6764_/Q sky130_fd_sc_hd__dfrtp_1
X_3976_ _6434_/Q hold881/X _3996_/S VGND VGND VPWR VPWR _3976_/X sky130_fd_sc_hd__mux2_2
XFILLER_188_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5715_ _6934_/Q _5659_/X _5672_/X _6950_/Q VGND VGND VPWR VPWR _5715_/X sky130_fd_sc_hd__a22o_1
X_6695_ _6759_/CLK _6695_/D fanout449/X VGND VGND VPWR VPWR _6695_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5646_ _5646_/A1 _5643_/B _5645_/X VGND VGND VPWR VPWR _7159_/D sky130_fd_sc_hd__a21o_1
XFILLER_163_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5577_ _5577_/A0 _5577_/A1 _5577_/S VGND VGND VPWR VPWR _5577_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold220 hold220/A VGND VGND VPWR VPWR hold220/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_191_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4528_ _4947_/A _4426_/Y _4527_/X _4575_/C VGND VGND VPWR VPWR _4529_/D sky130_fd_sc_hd__o22a_1
Xhold231 hold231/A VGND VGND VPWR VPWR hold231/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold242 hold242/A VGND VGND VPWR VPWR hold831/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold253 hold943/X VGND VGND VPWR VPWR hold944/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold264 hold264/A VGND VGND VPWR VPWR wb_dat_o[17] sky130_fd_sc_hd__buf_12
XFILLER_49_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold275 hold275/A VGND VGND VPWR VPWR wb_dat_o[16] sky130_fd_sc_hd__buf_12
Xhold286 hold286/A VGND VGND VPWR VPWR wb_dat_o[5] sky130_fd_sc_hd__buf_12
XFILLER_78_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4459_ _4485_/B _4564_/C _4881_/A VGND VGND VPWR VPWR _4980_/A sky130_fd_sc_hd__and3_2
Xhold297 hold297/A VGND VGND VPWR VPWR _6707_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7178_ _3950_/A1 _7178_/D fanout482/X VGND VGND VPWR VPWR _7178_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6129_ _6129_/A _6129_/B _6129_/C _6129_/D VGND VGND VPWR VPWR _6139_/B sky130_fd_sc_hd__nor4_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_104 _6787_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_115 _5196_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 _6432_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_137 hold153/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_148 _3402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_159 _5678_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_53_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7035_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_17_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3830_ _6657_/Q _3834_/S VGND VGND VPWR VPWR _3830_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_68_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6809_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_32_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3761_ _7085_/Q _5524_/A _3391_/Y _7141_/Q _3760_/X VGND VGND VPWR VPWR _3769_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_186_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5500_ _5500_/A0 _5518_/A1 _5505_/S VGND VGND VPWR VPWR _5500_/X sky130_fd_sc_hd__mux2_1
X_6480_ _6792_/CLK _6480_/D fanout442/X VGND VGND VPWR VPWR _6480_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3692_ _6645_/Q _4206_/A _4194_/A _6635_/Q VGND VGND VPWR VPWR _3692_/X sky130_fd_sc_hd__a22o_1
XFILLER_185_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5431_ _5431_/A0 _5575_/A1 _5433_/S VGND VGND VPWR VPWR _5431_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput303 _5643_/A VGND VGND VPWR VPWR serial_clock sky130_fd_sc_hd__buf_12
Xoutput314 hold1291/X VGND VGND VPWR VPWR hold230/A sky130_fd_sc_hd__buf_6
XFILLER_160_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5362_ _5362_/A _5569_/B VGND VGND VPWR VPWR _5370_/S sky130_fd_sc_hd__and2_4
Xoutput325 hold1315/X VGND VGND VPWR VPWR hold247/A sky130_fd_sc_hd__buf_6
Xoutput336 hold1267/X VGND VGND VPWR VPWR hold233/A sky130_fd_sc_hd__buf_6
X_7101_ _7117_/CLK _7101_/D fanout457/X VGND VGND VPWR VPWR _7101_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_114_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4313_ hold183/X _5518_/A1 _4315_/S VGND VGND VPWR VPWR _6739_/D sky130_fd_sc_hd__mux2_1
X_5293_ _5293_/A0 _5572_/A1 _5298_/S VGND VGND VPWR VPWR _6879_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7032_ _7119_/CLK _7032_/D fanout472/X VGND VGND VPWR VPWR _7032_/Q sky130_fd_sc_hd__dfrtp_4
X_4244_ _4244_/A0 _5581_/A1 _4249_/S VGND VGND VPWR VPWR _6670_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4175_ _4175_/A0 hold95/X _4175_/S VGND VGND VPWR VPWR _4175_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6816_ _6816_/CLK _6816_/D _6409_/A VGND VGND VPWR VPWR _6816_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6747_ _6747_/CLK _6747_/D fanout439/X VGND VGND VPWR VPWR _6747_/Q sky130_fd_sc_hd__dfrtp_4
X_3959_ _6456_/Q _3959_/B VGND VGND VPWR VPWR _3959_/Y sky130_fd_sc_hd__nor2_2
XFILLER_51_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6678_ _7152_/CLK _6678_/D _6346_/B VGND VGND VPWR VPWR _6678_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_831 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5629_ _5629_/A1 _5631_/A _5628_/Y VGND VGND VPWR VPWR _7153_/D sky130_fd_sc_hd__a21oi_1
XFILLER_151_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5980_ _6017_/B _6018_/B _6007_/C VGND VGND VPWR VPWR _5980_/X sky130_fd_sc_hd__and3_4
X_4931_ _5123_/A _4931_/B _4931_/C _4931_/D VGND VGND VPWR VPWR _4931_/X sky130_fd_sc_hd__and4_1
XFILLER_64_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4862_ _4638_/Y _4713_/Y _4622_/C VGND VGND VPWR VPWR _4870_/B sky130_fd_sc_hd__o21a_1
XFILLER_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6601_ _6691_/CLK _6601_/D fanout443/X VGND VGND VPWR VPWR _6601_/Q sky130_fd_sc_hd__dfstp_2
X_3813_ _3811_/B _3813_/B VGND VGND VPWR VPWR _6469_/D sky130_fd_sc_hd__and2b_1
XANTENNA_15 _3385_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 _5505_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4793_ _4411_/Y _4712_/Y _4776_/Y _4792_/X _4531_/B VGND VGND VPWR VPWR _4793_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_193_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_37 _5685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_48 _5994_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6532_ _6691_/CLK _6532_/D fanout443/X VGND VGND VPWR VPWR _6532_/Q sky130_fd_sc_hd__dfrtp_4
X_3744_ _6457_/Q _6437_/Q _6808_/Q VGND VGND VPWR VPWR _3745_/A sky130_fd_sc_hd__nor3_1
XANTENNA_59 _6920_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6463_ _6656_/CLK _6463_/D _6413_/X VGND VGND VPWR VPWR _6463_/Q sky130_fd_sc_hd__dfrtp_4
X_3675_ _3675_/A _3675_/B _3675_/C VGND VGND VPWR VPWR _3675_/Y sky130_fd_sc_hd__nand3_4
XFILLER_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5414_ _5414_/A0 _5585_/A1 _5415_/S VGND VGND VPWR VPWR _6987_/D sky130_fd_sc_hd__mux2_1
X_6394_ _6399_/A _6423_/B VGND VGND VPWR VPWR _6394_/X sky130_fd_sc_hd__and2_1
XFILLER_133_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5345_ hold669/X _5561_/A1 _5352_/S VGND VGND VPWR VPWR _5345_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput177 _3229_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[11] sky130_fd_sc_hd__buf_12
XFILLER_142_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput188 _3218_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[21] sky130_fd_sc_hd__buf_12
XFILLER_114_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput199 _3208_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[31] sky130_fd_sc_hd__buf_12
X_5276_ _5276_/A0 _5303_/A1 _5280_/S VGND VGND VPWR VPWR _5276_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7015_ _7121_/CLK _7015_/D _6399_/A VGND VGND VPWR VPWR _7015_/Q sky130_fd_sc_hd__dfrtp_4
X_4227_ _5238_/A0 hold135/X _4239_/S VGND VGND VPWR VPWR _4227_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4158_ _4158_/A hold13/A VGND VGND VPWR VPWR _4163_/S sky130_fd_sc_hd__and2_4
XFILLER_110_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4089_ _3462_/Y hold824/A _4091_/S VGND VGND VPWR VPWR _6545_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout371 _4411_/Y VGND VGND VPWR VPWR _4947_/A sky130_fd_sc_hd__buf_12
XFILLER_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout382 hold95/X VGND VGND VPWR VPWR _5196_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_143_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout393 _4337_/A1 VGND VGND VPWR VPWR _5187_/A1 sky130_fd_sc_hd__buf_8
XFILLER_143_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput13 mask_rev_in[18] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__buf_2
XFILLER_128_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput24 mask_rev_in[28] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput35 mask_rev_in[9] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput46 mgmt_gpio_in[19] VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__buf_2
XFILLER_155_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput57 mgmt_gpio_in[29] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__clkbuf_2
Xinput68 mgmt_gpio_in[5] VGND VGND VPWR VPWR _3970_/A sky130_fd_sc_hd__buf_4
Xhold808 hold808/A VGND VGND VPWR VPWR hold808/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput79 spi_enabled VGND VGND VPWR VPWR _3971_/B sky130_fd_sc_hd__buf_6
Xhold819 hold819/A VGND VGND VPWR VPWR hold819/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3460_ _3460_/A _3460_/B _3460_/C _3460_/D VGND VGND VPWR VPWR _3461_/C sky130_fd_sc_hd__nor4_1
X_3391_ hold26/X _3516_/B VGND VGND VPWR VPWR _3391_/Y sky130_fd_sc_hd__nor2_8
XFILLER_124_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5130_ _5130_/A _5130_/B _5130_/C VGND VGND VPWR VPWR _5131_/C sky130_fd_sc_hd__and3_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2209 hold786/X VGND VGND VPWR VPWR _4141_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1508 hold157/X VGND VGND VPWR VPWR _4168_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5061_ _5061_/A _5061_/B VGND VGND VPWR VPWR _5062_/A sky130_fd_sc_hd__nand2_2
XFILLER_85_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1519 hold504/X VGND VGND VPWR VPWR _5307_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4012_ _6432_/B _4241_/A VGND VGND VPWR VPWR _4012_/X sky130_fd_sc_hd__and2b_4
XFILLER_93_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5963_ _6691_/Q _5659_/X _5687_/X _6603_/Q VGND VGND VPWR VPWR _5963_/X sky130_fd_sc_hd__a22o_1
X_4914_ _4633_/B _4688_/C _4871_/B _4898_/B VGND VGND VPWR VPWR _5046_/B sky130_fd_sc_hd__o211a_1
X_5894_ _6580_/Q _5688_/X _5887_/X _5888_/X _5893_/X VGND VGND VPWR VPWR _5894_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_80_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4845_ _4569_/C _4655_/A _4590_/Y _4688_/B VGND VGND VPWR VPWR _4845_/X sky130_fd_sc_hd__o22a_1
XFILLER_178_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4776_ _4776_/A _5081_/A VGND VGND VPWR VPWR _4776_/Y sky130_fd_sc_hd__nor2_1
XFILLER_165_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6515_ _7080_/CLK _6515_/D fanout480/X VGND VGND VPWR VPWR _6515_/Q sky130_fd_sc_hd__dfrtp_1
X_3727_ input72/X _4056_/C _4009_/A _6488_/Q VGND VGND VPWR VPWR _3727_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6446_ _6656_/CLK _6446_/D _6401_/X VGND VGND VPWR VPWR _6446_/Q sky130_fd_sc_hd__dfrtp_1
X_3658_ _6596_/Q _4146_/A _4268_/A _6704_/Q VGND VGND VPWR VPWR _3658_/X sky130_fd_sc_hd__a22o_2
X_6377_ _6686_/Q _6377_/A2 _6377_/B1 _6685_/Q _6376_/X VGND VGND VPWR VPWR _6377_/X
+ sky130_fd_sc_hd__a221o_1
X_3589_ _6792_/Q _3427_/Y _3562_/Y input95/X VGND VGND VPWR VPWR _3589_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5328_ hold692/X _5580_/A1 _5334_/S VGND VGND VPWR VPWR _6910_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5259_ _5259_/A0 _5583_/A1 _5262_/S VGND VGND VPWR VPWR _6849_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_726 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__1153_ clkbuf_0__1153_/X VGND VGND VPWR VPWR _6351_/A0 sky130_fd_sc_hd__clkbuf_16
XFILLER_184_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4630_ _4976_/A _5067_/B _4754_/D _4630_/D VGND VGND VPWR VPWR _4631_/D sky130_fd_sc_hd__and4b_1
XFILLER_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4561_ _4598_/B _4607_/B _4881_/B _3967_/A VGND VGND VPWR VPWR _4561_/X sky130_fd_sc_hd__a31o_1
XFILLER_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6300_ _6700_/Q _5997_/X _6017_/X _6772_/Q VGND VGND VPWR VPWR _6300_/X sky130_fd_sc_hd__a22o_1
X_3512_ _3530_/B _3533_/B VGND VGND VPWR VPWR _4212_/A sky130_fd_sc_hd__nor2_8
Xhold605 hold605/A VGND VGND VPWR VPWR hold605/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4492_ _4637_/B _4492_/B _4500_/B VGND VGND VPWR VPWR _4639_/S sky130_fd_sc_hd__and3_2
Xhold616 hold616/A VGND VGND VPWR VPWR hold616/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold627 hold627/A VGND VGND VPWR VPWR hold627/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold638 hold638/A VGND VGND VPWR VPWR hold638/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold649 hold649/A VGND VGND VPWR VPWR hold649/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6231_ _6697_/Q _5997_/X _6004_/X _6574_/Q VGND VGND VPWR VPWR _6231_/X sky130_fd_sc_hd__a22o_1
Xmax_cap357 _3530_/B VGND VGND VPWR VPWR _3535_/A sky130_fd_sc_hd__buf_12
XFILLER_116_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3443_ _6874_/Q _5281_/A _5461_/A _7034_/Q _3438_/X VGND VGND VPWR VPWR _3444_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _7138_/Q _5977_/X _5984_/X _7098_/Q _6161_/X VGND VGND VPWR VPWR _6163_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _7108_/Q _3311_/Y _5515_/A _7084_/Q _3360_/X VGND VGND VPWR VPWR _3374_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2006 _5430_/X VGND VGND VPWR VPWR _7001_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _5123_/C _5113_/B VGND VGND VPWR VPWR _5113_/Y sky130_fd_sc_hd__nand2_1
Xhold2017 _6910_/Q VGND VGND VPWR VPWR hold692/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2028 _5491_/X VGND VGND VPWR VPWR _7055_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2039 hold717/X VGND VGND VPWR VPWR _4306_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _6896_/Q _5989_/X _6013_/X _7080_/Q VGND VGND VPWR VPWR _6093_/X sky130_fd_sc_hd__a22o_1
Xhold1305 _4048_/X VGND VGND VPWR VPWR hold154/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1316 _6573_/Q VGND VGND VPWR VPWR hold142/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1327 _6884_/Q VGND VGND VPWR VPWR hold341/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _5044_/A _5044_/B _5044_/C VGND VGND VPWR VPWR _5086_/B sky130_fd_sc_hd__and3_1
Xhold1338 hold244/X VGND VGND VPWR VPWR hold1338/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1349 hold187/X VGND VGND VPWR VPWR _5466_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_66_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6995_ _7140_/CLK _6995_/D fanout469/X VGND VGND VPWR VPWR _6995_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5946_ _6528_/Q _5678_/Y _5940_/X _5945_/X _6341_/S VGND VGND VPWR VPWR _5946_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_179_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5877_ _6757_/Q _5664_/X _5679_/X _6589_/Q VGND VGND VPWR VPWR _5877_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4828_ _4384_/A _4675_/A _4633_/B _4825_/X _4827_/X VGND VGND VPWR VPWR _4828_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_193_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4759_ _5139_/A _4759_/B _4759_/C _4759_/D VGND VGND VPWR VPWR _4759_/X sky130_fd_sc_hd__and4_1
XFILLER_147_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6429_ _6432_/A _6433_/B VGND VGND VPWR VPWR _6429_/X sky130_fd_sc_hd__and2_1
XFILLER_108_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2540 _6463_/Q VGND VGND VPWR VPWR _3265_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1850 _6831_/Q VGND VGND VPWR VPWR hold237/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1861 hold569/X VGND VGND VPWR VPWR _4184_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1872 hold498/X VGND VGND VPWR VPWR _5258_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1883 _6744_/Q VGND VGND VPWR VPWR hold314/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1894 hold609/X VGND VGND VPWR VPWR _5173_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2 hold2/A VGND VGND VPWR VPWR hold2/X sky130_fd_sc_hd__buf_8
XFILLER_181_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5800_ _7058_/Q _5668_/X _5684_/X _6930_/Q VGND VGND VPWR VPWR _5800_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6780_ _3958_/A1 _6780_/D _6432_/X VGND VGND VPWR VPWR _6780_/Q sky130_fd_sc_hd__dfrtn_1
X_3992_ hold631/X _5195_/A1 _3999_/S VGND VGND VPWR VPWR _6474_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5731_ _6927_/Q _5684_/X _5686_/X _7007_/Q VGND VGND VPWR VPWR _5731_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5662_ _5689_/A _5684_/B _5688_/C VGND VGND VPWR VPWR _5662_/X sky130_fd_sc_hd__and3b_4
XFILLER_30_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4613_ _4570_/B _4523_/Y _4924_/A _5095_/B VGND VGND VPWR VPWR _4614_/D sky130_fd_sc_hd__o211a_1
XFILLER_129_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5593_ _7142_/Q _5594_/B VGND VGND VPWR VPWR _5593_/Y sky130_fd_sc_hd__nor2_1
XFILLER_175_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4544_ _4971_/A _4607_/B VGND VGND VPWR VPWR _4544_/Y sky130_fd_sc_hd__nand2_1
XFILLER_117_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold402 hold402/A VGND VGND VPWR VPWR hold402/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold413 hold413/A VGND VGND VPWR VPWR hold413/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold424 hold424/A VGND VGND VPWR VPWR hold424/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold435 hold435/A VGND VGND VPWR VPWR hold435/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold446 hold446/A VGND VGND VPWR VPWR hold446/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4475_ _4724_/C _4981_/A VGND VGND VPWR VPWR _5117_/A sky130_fd_sc_hd__nand2_2
Xhold457 hold457/A VGND VGND VPWR VPWR hold457/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold468 hold468/A VGND VGND VPWR VPWR hold468/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6214_ _6195_/X _6214_/B _6214_/C VGND VGND VPWR VPWR _6214_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_131_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold479 hold479/A VGND VGND VPWR VPWR hold479/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3426_ _3533_/B VGND VGND VPWR VPWR _5184_/B sky130_fd_sc_hd__clkinv_2
X_7194_ _7194_/CLK _7194_/D VGND VGND VPWR VPWR _7194_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6145_ _7058_/Q _5990_/X _5996_/X _7050_/Q VGND VGND VPWR VPWR _6145_/X sky130_fd_sc_hd__a22o_1
X_3357_ _3764_/B _3550_/B VGND VGND VPWR VPWR _3357_/Y sky130_fd_sc_hd__nor2_8
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1102 _5378_/X VGND VGND VPWR VPWR _6955_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1113 hold371/X VGND VGND VPWR VPWR _5486_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _6076_/A _6076_/B _6076_/C VGND VGND VPWR VPWR _6089_/C sky130_fd_sc_hd__nor3_1
Xhold1124 hold133/X VGND VGND VPWR VPWR _3980_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_3288_ _3429_/A hold66/X VGND VGND VPWR VPWR _3430_/A sky130_fd_sc_hd__and2_4
Xhold1135 _6914_/Q VGND VGND VPWR VPWR hold449/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1146 _5351_/X VGND VGND VPWR VPWR _6931_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1157 _5531_/X VGND VGND VPWR VPWR _7091_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5027_ _4947_/A _4995_/A _5034_/D _5034_/A _4509_/Y VGND VGND VPWR VPWR _5027_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_73_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1168 hold179/X VGND VGND VPWR VPWR _4300_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1179 hold107/X VGND VGND VPWR VPWR hold94/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6978_ _7084_/CLK _6978_/D fanout455/X VGND VGND VPWR VPWR _6978_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5929_ _6745_/Q _5929_/B VGND VGND VPWR VPWR _5929_/X sky130_fd_sc_hd__and2_1
XFILLER_70_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold980 _5386_/X VGND VGND VPWR VPWR _6962_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_89_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold991 _7044_/Q VGND VGND VPWR VPWR hold56/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_135_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2370 hold755/X VGND VGND VPWR VPWR _5429_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2381 _7021_/Q VGND VGND VPWR VPWR hold815/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_64_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2392 hold726/X VGND VGND VPWR VPWR _5574_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1680 hold734/X VGND VGND VPWR VPWR _4154_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1691 hold848/X VGND VGND VPWR VPWR hold191/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_189_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4260_ _4260_/A0 _5303_/A1 _4261_/S VGND VGND VPWR VPWR _4260_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3211_ _7064_/Q VGND VGND VPWR VPWR _3211_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4191_ hold587/X _5187_/A1 _4193_/S VGND VGND VPWR VPWR _6631_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6901_ _7077_/CLK _6901_/D fanout454/X VGND VGND VPWR VPWR _6901_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_47_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6832_ _6833_/CLK _6832_/D fanout457/X VGND VGND VPWR VPWR _6832_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6763_ _7183_/CLK _6763_/D _6346_/B VGND VGND VPWR VPWR _6763_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3975_ _6686_/Q _3975_/B VGND VGND VPWR VPWR _6677_/D sky130_fd_sc_hd__and2_1
X_5714_ _7030_/Q _5655_/X _5687_/X _6918_/Q VGND VGND VPWR VPWR _5714_/X sky130_fd_sc_hd__a22o_1
XFILLER_31_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6694_ _6750_/CLK _6694_/D fanout446/X VGND VGND VPWR VPWR _6694_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_191_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5645_ _7143_/Q _6492_/Q _5645_/C _7142_/Q VGND VGND VPWR VPWR _5645_/X sky130_fd_sc_hd__and4b_1
XFILLER_176_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5576_ _5576_/A0 _5576_/A1 _5577_/S VGND VGND VPWR VPWR _5576_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold210 hold210/A VGND VGND VPWR VPWR wb_dat_o[19] sky130_fd_sc_hd__buf_12
XFILLER_151_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4527_ _4462_/Y _4477_/Y _4466_/A _4463_/B VGND VGND VPWR VPWR _4527_/X sky130_fd_sc_hd__a211o_1
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold221 hold221/A VGND VGND VPWR VPWR hold221/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold232 hold232/A VGND VGND VPWR VPWR hold232/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold243 hold243/A VGND VGND VPWR VPWR wb_dat_o[23] sky130_fd_sc_hd__buf_12
XFILLER_132_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold254 hold254/A VGND VGND VPWR VPWR hold254/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold265 hold265/A VGND VGND VPWR VPWR hold841/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold276 hold276/A VGND VGND VPWR VPWR hold276/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4458_ _4598_/A _4881_/A VGND VGND VPWR VPWR _4491_/B sky130_fd_sc_hd__and2_4
XFILLER_49_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold287 hold287/A VGND VGND VPWR VPWR hold287/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold298 hold298/A VGND VGND VPWR VPWR hold298/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3409_ _7091_/Q _5524_/A _3347_/Y _7011_/Q _3408_/X VGND VGND VPWR VPWR _3409_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_120_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7177_ _3950_/A1 _7177_/D fanout468/X VGND VGND VPWR VPWR _7177_/Q sky130_fd_sc_hd__dfrtp_1
X_4389_ _4447_/B _4663_/D _4917_/A _4701_/A VGND VGND VPWR VPWR _4808_/A sky130_fd_sc_hd__nor4_4
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6128_ _6961_/Q _5992_/X _5999_/X _6865_/Q _6127_/X VGND VGND VPWR VPWR _6129_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6059_ _6974_/Q _5976_/B _5980_/X _6934_/Q VGND VGND VPWR VPWR _6059_/X sky130_fd_sc_hd__a22o_1
XTAP_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_105 _6485_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_116 _5556_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 _6432_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_138 _5407_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_149 _3438_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3760_ _7077_/Q _5515_/A _3336_/Y input20/X VGND VGND VPWR VPWR _3760_/X sky130_fd_sc_hd__a22o_1
XFILLER_32_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3691_ _6790_/Q _3427_/Y _4170_/A _6615_/Q _3690_/X VGND VGND VPWR VPWR _3694_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_158_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5430_ _5430_/A0 _5556_/A1 _5433_/S VGND VGND VPWR VPWR _5430_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput304 _3428_/X VGND VGND VPWR VPWR serial_data_1 sky130_fd_sc_hd__buf_12
X_5361_ _5361_/A0 _5559_/A1 _5361_/S VGND VGND VPWR VPWR _5361_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput315 hold833/X VGND VGND VPWR VPWR hold251/A sky130_fd_sc_hd__buf_6
Xoutput326 hold857/X VGND VGND VPWR VPWR hold199/A sky130_fd_sc_hd__buf_6
Xoutput337 hold1261/X VGND VGND VPWR VPWR hold207/A sky130_fd_sc_hd__buf_6
X_4312_ _4312_/A0 hold135/X _4315_/S VGND VGND VPWR VPWR _4312_/X sky130_fd_sc_hd__mux2_1
X_7100_ _7100_/CLK hold72/X fanout458/X VGND VGND VPWR VPWR _7100_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5292_ hold765/X _5580_/A1 _5298_/S VGND VGND VPWR VPWR _6878_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7031_ _7125_/CLK _7031_/D fanout454/X VGND VGND VPWR VPWR _7031_/Q sky130_fd_sc_hd__dfrtp_4
X_4243_ _4243_/A0 _5580_/A1 _4249_/S VGND VGND VPWR VPWR _4243_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4174_ _4174_/A0 _5303_/A1 _4175_/S VGND VGND VPWR VPWR _6617_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6815_ _7013_/CLK _6815_/D fanout452/X VGND VGND VPWR VPWR _6815_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_168_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6746_ _6750_/CLK _6746_/D fanout446/X VGND VGND VPWR VPWR _6746_/Q sky130_fd_sc_hd__dfrtp_4
X_3958_ input83/X _3958_/A1 _6456_/Q VGND VGND VPWR VPWR _3958_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3889_ _4720_/C _4649_/B VGND VGND VPWR VPWR _4394_/A sky130_fd_sc_hd__and2_1
XFILLER_136_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6677_ _7152_/CLK _6677_/D _6346_/B VGND VGND VPWR VPWR _6677_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5628_ _7153_/Q _5611_/Y _5631_/A VGND VGND VPWR VPWR _5628_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_164_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5559_ _5559_/A0 _5559_/A1 _5559_/S VGND VGND VPWR VPWR _5559_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7229_ _7229_/A VGND VGND VPWR VPWR _7229_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4930_ _4930_/A _5049_/C _4930_/C _4930_/D VGND VGND VPWR VPWR _4931_/D sky130_fd_sc_hd__and4_1
XFILLER_17_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4861_ _4569_/C _4655_/A _4590_/Y _4714_/Y VGND VGND VPWR VPWR _4871_/C sky130_fd_sc_hd__o22a_1
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6600_ _6817_/CLK _6600_/D fanout451/X VGND VGND VPWR VPWR _6600_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_177_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3812_ _3181_/Y _3814_/B _3879_/A VGND VGND VPWR VPWR _3813_/B sky130_fd_sc_hd__o21ai_1
XFILLER_177_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_16 _3385_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4792_ _4462_/Y _4464_/Y _4466_/A _4790_/X _4791_/X VGND VGND VPWR VPWR _4792_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_193_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_27 _5656_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_38 _5685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6531_ _6691_/CLK _6531_/D fanout442/X VGND VGND VPWR VPWR _6531_/Q sky130_fd_sc_hd__dfrtp_4
X_3743_ _6997_/Q _5425_/A _4092_/A _6548_/Q _3742_/X VGND VGND VPWR VPWR _3750_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA_49 _5997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3674_ _3674_/A _3674_/B _3674_/C _3674_/D VGND VGND VPWR VPWR _3675_/C sky130_fd_sc_hd__and4_2
X_6462_ _6656_/CLK _6462_/D _6412_/X VGND VGND VPWR VPWR _6462_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_146_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5413_ _5413_/A0 _5503_/A1 _5415_/S VGND VGND VPWR VPWR _6986_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6393_ _6409_/A _6423_/B VGND VGND VPWR VPWR _6393_/X sky130_fd_sc_hd__and2_1
XFILLER_173_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5344_ _5344_/A _5569_/B VGND VGND VPWR VPWR _5352_/S sky130_fd_sc_hd__and2_4
Xoutput178 _3228_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[12] sky130_fd_sc_hd__buf_12
Xoutput189 _3217_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[22] sky130_fd_sc_hd__buf_12
X_5275_ _5275_/A0 _5518_/A1 _5280_/S VGND VGND VPWR VPWR _5275_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4226_ _4226_/A0 _4225_/X _4240_/S VGND VGND VPWR VPWR _6660_/D sky130_fd_sc_hd__mux2_1
X_7014_ _7136_/CLK _7014_/D fanout475/X VGND VGND VPWR VPWR _7014_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4157_ _4157_/A0 _5196_/A1 _4157_/S VGND VGND VPWR VPWR _4157_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4088_ _6351_/A0 hold856/A _4091_/S VGND VGND VPWR VPWR _6544_/D sky130_fd_sc_hd__mux2_1
XFILLER_169_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6729_ _6729_/CLK _6729_/D fanout465/X VGND VGND VPWR VPWR _6729_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_165_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_52_csclk _7093_/CLK VGND VGND VPWR VPWR _6983_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_118_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_67_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6817_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_120_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout383 hold95/X VGND VGND VPWR VPWR _4339_/A1 sky130_fd_sc_hd__buf_4
XFILLER_120_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout394 hold2/X VGND VGND VPWR VPWR _4337_/A1 sky130_fd_sc_hd__buf_8
XFILLER_143_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput14 mask_rev_in[19] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__buf_2
Xinput25 mask_rev_in[29] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput36 mgmt_gpio_in[0] VGND VGND VPWR VPWR _3972_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_128_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput47 mgmt_gpio_in[1] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__buf_2
Xinput58 mgmt_gpio_in[2] VGND VGND VPWR VPWR wire1/A sky130_fd_sc_hd__buf_6
XFILLER_10_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput69 mgmt_gpio_in[6] VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold809 hold809/A VGND VGND VPWR VPWR hold809/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3390_ _3425_/A _3390_/B VGND VGND VPWR VPWR _3516_/B sky130_fd_sc_hd__nand2_8
XFILLER_124_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5060_ _5059_/X _5115_/A VGND VGND VPWR VPWR _5060_/X sky130_fd_sc_hd__and2b_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1509 _4168_/X VGND VGND VPWR VPWR hold158/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4011_ hold164/X hold135/X _4011_/S VGND VGND VPWR VPWR _4011_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5962_ _6638_/Q _5671_/X _5960_/X _5961_/X VGND VGND VPWR VPWR _5962_/X sky130_fd_sc_hd__a211o_1
XFILLER_52_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4913_ _4913_/A _4913_/B VGND VGND VPWR VPWR _5121_/B sky130_fd_sc_hd__and2_1
X_5893_ _6549_/Q _5673_/X _5890_/X _5892_/X VGND VGND VPWR VPWR _5893_/X sky130_fd_sc_hd__a211o_1
XFILLER_178_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4844_ _4569_/B _4655_/A _4590_/Y _4688_/A VGND VGND VPWR VPWR _4872_/A sky130_fd_sc_hd__o22a_1
XFILLER_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4775_ _4729_/A _4674_/Y _5063_/A VGND VGND VPWR VPWR _4796_/A sky130_fd_sc_hd__o21a_1
XFILLER_165_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6514_ _7080_/CLK hold48/X fanout480/X VGND VGND VPWR VPWR _6514_/Q sky130_fd_sc_hd__dfrtp_1
X_3726_ _3726_/A hold26/X VGND VGND VPWR VPWR _4009_/A sky130_fd_sc_hd__nor2_4
XFILLER_134_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6445_ _6656_/CLK _6445_/D _6400_/X VGND VGND VPWR VPWR _6445_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_174_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3657_ _7095_/Q _5533_/A _4274_/A _6709_/Q _3656_/X VGND VGND VPWR VPWR _3664_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_164_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6376_ _6684_/Q _6376_/A2 _6376_/B1 _4218_/Y VGND VGND VPWR VPWR _6376_/X sky130_fd_sc_hd__a22o_1
X_3588_ _7016_/Q _5443_/A _3336_/Y input23/X _3564_/X VGND VGND VPWR VPWR _3595_/A
+ sky130_fd_sc_hd__a221o_2
X_5327_ hold813/X _5552_/A1 _5334_/S VGND VGND VPWR VPWR _6909_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5258_ _5258_/A0 _5555_/A1 _5262_/S VGND VGND VPWR VPWR _6848_/D sky130_fd_sc_hd__mux2_1
XFILLER_75_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4209_ hold310/X _4337_/A1 _4211_/S VGND VGND VPWR VPWR _4209_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5189_ hold457/X _5196_/A1 _5190_/S VGND VGND VPWR VPWR _5189_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4560_ _4560_/A _4560_/B _4560_/C _4598_/C VGND VGND VPWR VPWR _4881_/B sky130_fd_sc_hd__and4_2
XFILLER_144_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3511_ _7129_/Q _5569_/A _5380_/A _6961_/Q _3510_/X VGND VGND VPWR VPWR _3515_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_156_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold606 hold606/A VGND VGND VPWR VPWR hold606/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4491_ _4598_/C _4491_/B VGND VGND VPWR VPWR _4491_/Y sky130_fd_sc_hd__nand2_8
Xhold617 hold617/A VGND VGND VPWR VPWR hold617/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold628 hold628/A VGND VGND VPWR VPWR hold628/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6230_ _6230_/A _6230_/B _6230_/C VGND VGND VPWR VPWR _6239_/C sky130_fd_sc_hd__nor3_2
X_3442_ _7002_/Q _5425_/A _5380_/A _6962_/Q _3441_/X VGND VGND VPWR VPWR _3444_/C
+ sky130_fd_sc_hd__a221o_1
Xhold639 hold639/A VGND VGND VPWR VPWR hold639/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap358 _3686_/B VGND VGND VPWR VPWR _3764_/B sky130_fd_sc_hd__buf_12
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3373_ _6844_/Q hold27/A _5236_/C _3973_/B _3372_/X VGND VGND VPWR VPWR _3384_/A
+ sky130_fd_sc_hd__a221o_2
X_6161_ _6930_/Q _5982_/X _5987_/X _7114_/Q VGND VGND VPWR VPWR _6161_/X sky130_fd_sc_hd__a22o_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2007 _7009_/Q VGND VGND VPWR VPWR hold533/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5112_ _5112_/A _5112_/B _5112_/C _5112_/D VGND VGND VPWR VPWR _5113_/B sky130_fd_sc_hd__and4_1
Xhold2018 _7110_/Q VGND VGND VPWR VPWR hold760/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2029 _6885_/Q VGND VGND VPWR VPWR hold783/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6092_ _6116_/A0 _6091_/X _6342_/S VGND VGND VPWR VPWR _6092_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1306 hold154/X VGND VGND VPWR VPWR _6509_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1317 hold142/X VGND VGND VPWR VPWR _4121_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5043_ _5043_/A _5043_/B VGND VGND VPWR VPWR _5043_/Y sky130_fd_sc_hd__nand2_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1328 hold341/X VGND VGND VPWR VPWR _5298_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1339 _6982_/Q VGND VGND VPWR VPWR hold636/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_66_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_wbbd_sck _7203_/Q VGND VGND VPWR VPWR clkbuf_0_wbbd_sck/X sky130_fd_sc_hd__clkbuf_16
X_6994_ _7084_/CLK _6994_/D fanout455/X VGND VGND VPWR VPWR _6994_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_25_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5945_ _6700_/Q _5672_/X _5941_/X _5943_/X _5944_/X VGND VGND VPWR VPWR _5945_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5876_ _6548_/Q _5673_/X _5682_/X _6450_/Q _5875_/X VGND VGND VPWR VPWR _5879_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4827_ _4947_/A _4701_/B _4812_/Y _4698_/Y _4928_/B VGND VGND VPWR VPWR _4827_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_138_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4758_ _4986_/C _4837_/B _4965_/B _4757_/X _4716_/Y VGND VGND VPWR VPWR _4759_/D
+ sky130_fd_sc_hd__a41o_1
XFILLER_193_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3709_ _7070_/Q _5506_/A _5515_/A _7078_/Q _3708_/X VGND VGND VPWR VPWR _3716_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4689_ _4710_/A _4719_/B VGND VGND VPWR VPWR _4689_/Y sky130_fd_sc_hd__nand2_1
XFILLER_162_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6428_ _6432_/A _6432_/B VGND VGND VPWR VPWR _6428_/X sky130_fd_sc_hd__and2_1
XFILLER_161_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6359_ _6685_/Q _6356_/Y _6357_/Y _6686_/Q _4836_/A VGND VGND VPWR VPWR _6359_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2530 _7147_/Q VGND VGND VPWR VPWR _5612_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_124_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_690 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1840 hold462/X VGND VGND VPWR VPWR _4032_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1851 hold237/X VGND VGND VPWR VPWR _5239_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1862 _4184_/X VGND VGND VPWR VPWR _6625_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1873 _6920_/Q VGND VGND VPWR VPWR hold468/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1884 _6648_/Q VGND VGND VPWR VPWR hold550/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1895 _5173_/X VGND VGND VPWR VPWR _6772_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold3 hold3/A VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_181_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3991_ hold574/X _5187_/A1 _3999_/S VGND VGND VPWR VPWR _6473_/D sky130_fd_sc_hd__mux2_1
X_5730_ _5750_/A1 _5729_/X _5730_/S VGND VGND VPWR VPWR _7161_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5661_ _7149_/Q _7148_/Q VGND VGND VPWR VPWR _5688_/C sky130_fd_sc_hd__and2b_4
XFILLER_31_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4612_ _4625_/A _4981_/A VGND VGND VPWR VPWR _5095_/B sky130_fd_sc_hd__nand2_1
XFILLER_176_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5592_ _6166_/S _3911_/B _3197_/Y VGND VGND VPWR VPWR _5594_/B sky130_fd_sc_hd__o21a_1
XFILLER_191_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4543_ _4464_/Y _4569_/C _4540_/X _5149_/A _4542_/Y VGND VGND VPWR VPWR _4543_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_116_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold403 hold403/A VGND VGND VPWR VPWR hold403/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold414 hold414/A VGND VGND VPWR VPWR hold414/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold425 hold425/A VGND VGND VPWR VPWR hold425/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold436 hold436/A VGND VGND VPWR VPWR hold436/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4474_ _4981_/A VGND VGND VPWR VPWR _4570_/B sky130_fd_sc_hd__inv_2
Xhold447 hold447/A VGND VGND VPWR VPWR hold447/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold458 hold458/A VGND VGND VPWR VPWR hold458/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold469 hold469/A VGND VGND VPWR VPWR hold469/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6213_ _6206_/X _6208_/X _6213_/C _6339_/B VGND VGND VPWR VPWR _6214_/C sky130_fd_sc_hd__and4bb_1
XFILLER_104_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3425_ _3425_/A _3430_/B VGND VGND VPWR VPWR _3533_/B sky130_fd_sc_hd__nand2_8
X_7193_ _7194_/CLK _7193_/D VGND VGND VPWR VPWR _7193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6144_ _6914_/Q _5991_/X _6018_/X _6970_/Q VGND VGND VPWR VPWR _6144_/X sky130_fd_sc_hd__a22o_1
X_3356_ _3563_/A _3550_/B VGND VGND VPWR VPWR _4239_/S sky130_fd_sc_hd__nor2_8
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1103 _6484_/Q VGND VGND VPWR VPWR hold431/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1114 _7019_/Q VGND VGND VPWR VPWR hold377/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3287_ _3563_/A _3354_/A VGND VGND VPWR VPWR _5569_/A sky130_fd_sc_hd__nor2_8
X_6075_ _7031_/Q _5986_/X _5998_/X _6887_/Q _6074_/X VGND VGND VPWR VPWR _6076_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_85_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1125 _3980_/X VGND VGND VPWR VPWR hold149/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_39_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1136 hold449/X VGND VGND VPWR VPWR _5332_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1147 _6813_/Q VGND VGND VPWR VPWR hold454/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5026_ _5150_/A _5026_/B _5026_/C VGND VGND VPWR VPWR _5034_/D sky130_fd_sc_hd__nand3_1
Xhold1158 _6923_/Q VGND VGND VPWR VPWR hold369/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1169 _4300_/X VGND VGND VPWR VPWR _6728_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_54_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6977_ _7119_/CLK _6977_/D fanout472/X VGND VGND VPWR VPWR _6977_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5928_ _3224_/Y _5872_/B _5677_/B VGND VGND VPWR VPWR _5928_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_179_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5859_ _7166_/Q _3924_/Y _5647_/Y VGND VGND VPWR VPWR _5859_/X sky130_fd_sc_hd__o21ba_1
XFILLER_166_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold970 hold970/A VGND VGND VPWR VPWR hold6/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold981 _6850_/Q VGND VGND VPWR VPWR hold981/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold992 hold56/X VGND VGND VPWR VPWR hold992/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2360 _6959_/Q VGND VGND VPWR VPWR hold624/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2371 _5429_/X VGND VGND VPWR VPWR _7000_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2382 hold815/X VGND VGND VPWR VPWR _5453_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2393 _5574_/X VGND VGND VPWR VPWR _7129_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1670 _7190_/Q VGND VGND VPWR VPWR hold854/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1681 _4154_/X VGND VGND VPWR VPWR _6600_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1692 _6709_/Q VGND VGND VPWR VPWR hold301/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3210_ _7072_/Q VGND VGND VPWR VPWR _3210_/Y sky130_fd_sc_hd__inv_2
X_4190_ _4190_/A0 _5186_/A1 _4193_/S VGND VGND VPWR VPWR _6630_/D sky130_fd_sc_hd__mux2_1
XFILLER_192_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6900_ _7124_/CLK _6900_/D fanout459/X VGND VGND VPWR VPWR _6900_/Q sky130_fd_sc_hd__dfrtp_4
X_6831_ _6833_/CLK _6831_/D fanout457/X VGND VGND VPWR VPWR _6831_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6762_ _7183_/CLK _6762_/D _6346_/B VGND VGND VPWR VPWR _6762_/Q sky130_fd_sc_hd__dfrtp_1
X_3974_ _6822_/Q _3974_/B VGND VGND VPWR VPWR _3974_/X sky130_fd_sc_hd__and2_4
X_5713_ _6894_/Q _5662_/X _5674_/X _6870_/Q _5712_/X VGND VGND VPWR VPWR _5718_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6693_ _6808_/CLK _6693_/D fanout440/X VGND VGND VPWR VPWR _6693_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_149_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5644_ _5644_/A1 _5643_/B _5643_/Y _6490_/Q VGND VGND VPWR VPWR _7158_/D sky130_fd_sc_hd__a22o_1
XFILLER_136_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5575_ hold965/X _5575_/A1 _5577_/S VGND VGND VPWR VPWR _5575_/X sky130_fd_sc_hd__mux2_1
Xhold200 hold200/A VGND VGND VPWR VPWR hold855/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold211 hold211/A VGND VGND VPWR VPWR hold211/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_191_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4526_ _5009_/A _5001_/A _4751_/B VGND VGND VPWR VPWR _4526_/X sky130_fd_sc_hd__and3_1
Xhold222 hold222/A VGND VGND VPWR VPWR hold222/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold233 hold233/A VGND VGND VPWR VPWR wb_dat_o[2] sky130_fd_sc_hd__buf_12
Xhold244 hold244/A VGND VGND VPWR VPWR hold244/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold255 hold255/A VGND VGND VPWR VPWR hold255/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold266 hold266/A VGND VGND VPWR VPWR wb_dat_o[8] sky130_fd_sc_hd__buf_12
X_4457_ _4457_/A _4469_/B _4457_/C VGND VGND VPWR VPWR _4881_/A sky130_fd_sc_hd__and3_4
XFILLER_171_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold277 hold277/A VGND VGND VPWR VPWR hold851/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold288 hold288/A VGND VGND VPWR VPWR hold863/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold299 hold299/A VGND VGND VPWR VPWR hold299/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3408_ _7083_/Q _5515_/A _5497_/A _7067_/Q VGND VGND VPWR VPWR _3408_/X sky130_fd_sc_hd__a22o_1
XFILLER_120_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7176_ _7204_/CLK _7176_/D fanout482/X VGND VGND VPWR VPWR _7176_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_172_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4388_ _4917_/A _4701_/A VGND VGND VPWR VPWR _4712_/A sky130_fd_sc_hd__nor2_8
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6127_ _6937_/Q _5980_/X _5982_/X _6929_/Q VGND VGND VPWR VPWR _6127_/X sky130_fd_sc_hd__a22o_1
X_3339_ _3764_/B _3563_/B VGND VGND VPWR VPWR _3339_/Y sky130_fd_sc_hd__nor2_8
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ _7062_/Q _5994_/X _5996_/X _7046_/Q _6057_/X VGND VGND VPWR VPWR _6058_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5009_ _5009_/A _5009_/B VGND VGND VPWR VPWR _5009_/Y sky130_fd_sc_hd__nor2_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 _5643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_117 _5303_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_128 _7186_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_139 _6794_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2190 _4327_/X VGND VGND VPWR VPWR _6751_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_64_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3690_ _6942_/Q _5362_/A _4286_/A _6718_/Q VGND VGND VPWR VPWR _3690_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput305 _3392_/X VGND VGND VPWR VPWR serial_data_2 sky130_fd_sc_hd__buf_12
X_5360_ _5360_/A0 _5576_/A1 _5361_/S VGND VGND VPWR VPWR _5360_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput316 hold827/X VGND VGND VPWR VPWR hold240/A sky130_fd_sc_hd__buf_6
Xoutput327 hold825/X VGND VGND VPWR VPWR hold224/A sky130_fd_sc_hd__buf_6
X_4311_ _4311_/A0 _5552_/A1 _4315_/S VGND VGND VPWR VPWR _6737_/D sky130_fd_sc_hd__mux2_1
Xoutput338 hold1285/X VGND VGND VPWR VPWR hold214/A sky130_fd_sc_hd__buf_6
X_5291_ hold602/X _5561_/A1 _5298_/S VGND VGND VPWR VPWR _5291_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7030_ _7113_/CLK _7030_/D fanout472/X VGND VGND VPWR VPWR _7030_/Q sky130_fd_sc_hd__dfstp_2
X_4242_ _4242_/A0 hold153/X _4249_/S VGND VGND VPWR VPWR _4242_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4173_ hold193/X _4337_/A1 _4175_/S VGND VGND VPWR VPWR _6616_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6814_ _7053_/CLK _6814_/D fanout452/X VGND VGND VPWR VPWR _6814_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6745_ _6757_/CLK _6745_/D fanout447/X VGND VGND VPWR VPWR _6745_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_177_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3957_ _6457_/Q _3959_/B VGND VGND VPWR VPWR _3957_/Y sky130_fd_sc_hd__nor2_2
XFILLER_192_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6676_ _7152_/CLK _6676_/D _6346_/B VGND VGND VPWR VPWR _6676_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_164_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3888_ _6455_/Q _6434_/Q _6423_/B VGND VGND VPWR VPWR _3975_/B sky130_fd_sc_hd__o21ai_2
X_5627_ _5647_/B _6019_/A _6017_/A _5605_/Y _5627_/B2 VGND VGND VPWR VPWR _7152_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_136_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5558_ _5558_/A0 _5576_/A1 _5559_/S VGND VGND VPWR VPWR _5558_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4509_ _4980_/A _4607_/B VGND VGND VPWR VPWR _4509_/Y sky130_fd_sc_hd__nand2_2
XFILLER_132_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5489_ hold807/X _5552_/A1 _5496_/S VGND VGND VPWR VPWR _5489_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7228_ _7228_/A VGND VGND VPWR VPWR _7228_/X sky130_fd_sc_hd__clkbuf_2
Xwire1 wire1/A VGND VGND VPWR VPWR wire1/X sky130_fd_sc_hd__buf_8
XFILLER_59_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7159_ _7186_/CLK _7159_/D fanout465/X VGND VGND VPWR VPWR _7159_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_747 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4860_ _4638_/Y _4683_/A _4683_/B _4586_/Y VGND VGND VPWR VPWR _4872_/C sky130_fd_sc_hd__o31a_1
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3811_ _3811_/A _3811_/B VGND VGND VPWR VPWR _6470_/D sky130_fd_sc_hd__xor2_1
X_4791_ _4791_/A _4791_/B _4791_/C _5034_/B VGND VGND VPWR VPWR _4791_/X sky130_fd_sc_hd__and4_1
XFILLER_159_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_17 _3385_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_28 _5656_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6530_ _6792_/CLK _6530_/D fanout442/X VGND VGND VPWR VPWR _6530_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_39 _5687_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3742_ _7053_/Q _5488_/A _4116_/A _6569_/Q VGND VGND VPWR VPWR _3742_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6461_ _6656_/CLK _6461_/D _6411_/X VGND VGND VPWR VPWR _6461_/Q sky130_fd_sc_hd__dfrtp_4
X_3673_ _3673_/A _3673_/B _3673_/C _3673_/D VGND VGND VPWR VPWR _3674_/D sky130_fd_sc_hd__nor4_1
XFILLER_118_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5412_ _5412_/A0 _5583_/A1 _5415_/S VGND VGND VPWR VPWR _6985_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6392_ _6426_/A _6432_/B VGND VGND VPWR VPWR _6392_/X sky130_fd_sc_hd__and2_1
XFILLER_114_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5343_ _5343_/A0 _5577_/A1 _5343_/S VGND VGND VPWR VPWR _5343_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput179 _3227_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[13] sky130_fd_sc_hd__buf_12
XFILLER_87_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5274_ _5274_/A0 _5499_/A1 _5280_/S VGND VGND VPWR VPWR _5274_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7013_ _7013_/CLK _7013_/D fanout453/X VGND VGND VPWR VPWR _7013_/Q sky130_fd_sc_hd__dfstp_2
X_4225_ _5237_/A0 _5552_/A1 _4239_/S VGND VGND VPWR VPWR _4225_/X sky130_fd_sc_hd__mux2_1
X_4156_ _4156_/A0 _5195_/A1 _4157_/S VGND VGND VPWR VPWR _4156_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4087_ _3616_/Y hold820/A _4091_/S VGND VGND VPWR VPWR _6543_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4989_ _5150_/B _4989_/B VGND VGND VPWR VPWR _4995_/B sky130_fd_sc_hd__nor2_4
XFILLER_11_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6728_ _6731_/CLK _6728_/D fanout465/X VGND VGND VPWR VPWR _6728_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_183_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6659_ _7152_/CLK _6659_/D _6346_/B VGND VGND VPWR VPWR _6659_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout373 hold6/X VGND VGND VPWR VPWR _5559_/A1 sky130_fd_sc_hd__clkbuf_16
Xfanout384 hold94/X VGND VGND VPWR VPWR hold95/A sky130_fd_sc_hd__buf_4
XFILLER_101_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout395 hold2/X VGND VGND VPWR VPWR _5518_/A1 sky130_fd_sc_hd__buf_12
XFILLER_59_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput15 mask_rev_in[1] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput26 mask_rev_in[2] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput37 mgmt_gpio_in[10] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__buf_2
Xinput48 mgmt_gpio_in[20] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__buf_2
XFILLER_128_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput59 mgmt_gpio_in[30] VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__clkbuf_4
XFILLER_143_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4010_ hold668/X _5552_/A1 _4011_/S VGND VGND VPWR VPWR _6487_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5961_ _6751_/Q _5666_/X _5689_/X _6628_/Q VGND VGND VPWR VPWR _5961_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4912_ _4640_/Y _4648_/Y _4679_/Y _4564_/Y _4658_/B VGND VGND VPWR VPWR _4913_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_45_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5892_ _6610_/Q _5660_/X _5669_/X _6650_/Q _5891_/X VGND VGND VPWR VPWR _5892_/X
+ sky130_fd_sc_hd__a221o_1
X_4843_ _4500_/Y _4652_/Y _4930_/A VGND VGND VPWR VPWR _5126_/A sky130_fd_sc_hd__o21a_1
XFILLER_178_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4774_ _4947_/A _4688_/B _4536_/Y VGND VGND VPWR VPWR _4774_/X sky130_fd_sc_hd__o21a_1
XFILLER_165_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6513_ _7016_/CLK _6513_/D fanout475/X VGND VGND VPWR VPWR _6513_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3725_ _3725_/A _3725_/B _3725_/C _3725_/D VGND VGND VPWR VPWR _3736_/C sky130_fd_sc_hd__nor4_1
XFILLER_158_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6444_ _3940_/A1 _6444_/D _6399_/X VGND VGND VPWR VPWR hold4/A sky130_fd_sc_hd__dfrtp_1
X_3656_ _7047_/Q _5479_/A _4077_/A _6537_/Q VGND VGND VPWR VPWR _3656_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6375_ _6374_/X _6375_/A1 _6384_/S VGND VGND VPWR VPWR _7199_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3587_ _3587_/A _3587_/B _3587_/C _3587_/D VGND VGND VPWR VPWR _3616_/C sky130_fd_sc_hd__nor4_2
XFILLER_114_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5326_ _5326_/A _5551_/B VGND VGND VPWR VPWR _5334_/S sky130_fd_sc_hd__and2_4
XFILLER_115_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5257_ _5257_/A0 _5572_/A1 _5262_/S VGND VGND VPWR VPWR _6847_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4208_ _4208_/A0 _5193_/A1 _4211_/S VGND VGND VPWR VPWR _4208_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5188_ _5188_/A0 _5195_/A1 _5190_/S VGND VGND VPWR VPWR _5188_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4139_ _4139_/A0 _4339_/A1 _4139_/S VGND VGND VPWR VPWR _6588_/D sky130_fd_sc_hd__mux2_1
XFILLER_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3510_ _7105_/Q _3311_/Y _3509_/Y _6731_/Q VGND VGND VPWR VPWR _3510_/X sky130_fd_sc_hd__a22o_1
XFILLER_128_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4490_ _4598_/C _4491_/B VGND VGND VPWR VPWR _4628_/A sky130_fd_sc_hd__and2_2
Xhold607 hold607/A VGND VGND VPWR VPWR hold607/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold618 hold618/A VGND VGND VPWR VPWR hold618/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold629 hold629/A VGND VGND VPWR VPWR hold629/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3441_ _6914_/Q _5326_/A _3427_/Y _6794_/Q VGND VGND VPWR VPWR _3441_/X sky130_fd_sc_hd__a22o_1
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap359 _3431_/A VGND VGND VPWR VPWR _3563_/A sky130_fd_sc_hd__buf_12
XFILLER_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6160_ _6866_/Q _5999_/X _6019_/X _6986_/Q _6143_/X VGND VGND VPWR VPWR _6163_/C
+ sky130_fd_sc_hd__a221o_1
X_3372_ _6486_/Q _3357_/Y _3369_/X _3371_/X VGND VGND VPWR VPWR _3372_/X sky130_fd_sc_hd__a211o_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5111_ _4990_/B _4995_/A _4699_/Y _4924_/C _4924_/A VGND VGND VPWR VPWR _5112_/D
+ sky130_fd_sc_hd__o2111a_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2008 hold533/X VGND VGND VPWR VPWR _5439_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_151_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2019 _6592_/Q VGND VGND VPWR VPWR hold601/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _7174_/Q _6090_/X _6166_/S VGND VGND VPWR VPWR _6091_/X sky130_fd_sc_hd__mux2_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1307 _7222_/A VGND VGND VPWR VPWR hold162/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1318 _4121_/X VGND VGND VPWR VPWR _6573_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5042_ _5042_/A _5149_/B _5086_/A _5042_/D VGND VGND VPWR VPWR _5043_/B sky130_fd_sc_hd__and4_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1329 _5298_/X VGND VGND VPWR VPWR _6884_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_38_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6993_ _7008_/CLK _6993_/D fanout472/X VGND VGND VPWR VPWR _6993_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_51_csclk _7093_/CLK VGND VGND VPWR VPWR _7132_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_81_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5944_ _6597_/Q _5670_/X _5685_/X _6772_/Q _5927_/X VGND VGND VPWR VPWR _5944_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_40_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5875_ _6747_/Q _5666_/X _5685_/X _6769_/Q VGND VGND VPWR VPWR _5875_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4826_ _4826_/A _4826_/B VGND VGND VPWR VPWR _4928_/B sky130_fd_sc_hd__nand2_1
XFILLER_119_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4757_ _4757_/A _4920_/B _4757_/C _4757_/D VGND VGND VPWR VPWR _4757_/X sky130_fd_sc_hd__and4_1
X_3708_ _7046_/Q _5479_/A _5236_/C input47/X VGND VGND VPWR VPWR _3708_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4688_ _4688_/A _4688_/B _4688_/C VGND VGND VPWR VPWR _4688_/X sky130_fd_sc_hd__and3_1
XFILLER_107_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6427_ _6432_/A _6432_/B VGND VGND VPWR VPWR _6427_/X sky130_fd_sc_hd__and2_1
XFILLER_134_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3639_ input22/X _3336_/Y _4188_/A _6631_/Q VGND VGND VPWR VPWR _3639_/X sky130_fd_sc_hd__a22o_1
XFILLER_162_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6358_ _6358_/A _6358_/B VGND VGND VPWR VPWR _6358_/Y sky130_fd_sc_hd__nand2_2
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5309_ hold793/X _5570_/A1 _5316_/S VGND VGND VPWR VPWR _5309_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6289_ _6270_/X _6289_/B _6289_/C VGND VGND VPWR VPWR _6289_/Y sky130_fd_sc_hd__nand3b_2
XFILLER_88_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2520 _5606_/X VGND VGND VPWR VPWR _7146_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2531 _7152_/Q VGND VGND VPWR VPWR _5627_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1830 _6660_/Q VGND VGND VPWR VPWR hold801/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1841 _4032_/X VGND VGND VPWR VPWR hold463/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1852 _6626_/Q VGND VGND VPWR VPWR hold305/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1863 _6619_/Q VGND VGND VPWR VPWR hold647/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1874 hold468/X VGND VGND VPWR VPWR _5339_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1885 hold550/X VGND VGND VPWR VPWR _4211_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_90_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1896 _6714_/Q VGND VGND VPWR VPWR hold290/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_19_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7111_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_140_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold4 hold4/A VGND VGND VPWR VPWR hold4/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xnet399_2 _3940_/A1 VGND VGND VPWR VPWR _3954_/B sky130_fd_sc_hd__inv_2
X_3990_ hold525/X _5193_/A1 _3999_/S VGND VGND VPWR VPWR _6472_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5660_ _5686_/A _5676_/B _5686_/B VGND VGND VPWR VPWR _5660_/X sky130_fd_sc_hd__and3_4
XFILLER_88_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4611_ _4611_/A _4693_/B VGND VGND VPWR VPWR _4924_/A sky130_fd_sc_hd__nand2_2
X_5591_ _5599_/D VGND VGND VPWR VPWR _5591_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4542_ _4971_/A _4972_/A VGND VGND VPWR VPWR _4542_/Y sky130_fd_sc_hd__nand2_1
XFILLER_190_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold404 hold404/A VGND VGND VPWR VPWR hold404/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold415 hold415/A VGND VGND VPWR VPWR hold415/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold426 hold426/A VGND VGND VPWR VPWR hold426/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4473_ _4473_/A _4598_/B _4564_/C VGND VGND VPWR VPWR _4981_/A sky130_fd_sc_hd__and3_4
Xhold437 hold437/A VGND VGND VPWR VPWR hold437/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold448 _4051_/X VGND VGND VPWR VPWR _6512_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold459 hold459/A VGND VGND VPWR VPWR hold459/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6212_ _7044_/Q _6016_/X _6209_/X _6211_/X VGND VGND VPWR VPWR _6213_/C sky130_fd_sc_hd__a211oi_1
X_3424_ _3423_/X _3424_/A1 _3739_/S VGND VGND VPWR VPWR _6780_/D sky130_fd_sc_hd__mux2_1
X_7192_ _7194_/CLK _7192_/D VGND VGND VPWR VPWR _7192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6143_ _7090_/Q _5638_/X _6015_/X _7018_/Q VGND VGND VPWR VPWR _6143_/X sky130_fd_sc_hd__a22o_1
XFILLER_112_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3355_ _3355_/A _3430_/B VGND VGND VPWR VPWR _3355_/Y sky130_fd_sc_hd__nand2_8
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _6975_/Q _5976_/B _5993_/X _7007_/Q VGND VGND VPWR VPWR _6074_/X sky130_fd_sc_hd__a22o_1
XFILLER_100_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0__1153_ _3558_/Y VGND VGND VPWR VPWR clkbuf_0__1153_/X sky130_fd_sc_hd__clkbuf_16
Xhold1104 _6987_/Q VGND VGND VPWR VPWR hold401/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_3286_ _3309_/A _3322_/B VGND VGND VPWR VPWR _3354_/A sky130_fd_sc_hd__nand2_8
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1115 hold377/X VGND VGND VPWR VPWR _5450_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1126 hold149/X VGND VGND VPWR VPWR hold134/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1137 _5332_/X VGND VGND VPWR VPWR _6914_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5025_ _5015_/X _5024_/Y _5139_/A _5140_/A VGND VGND VPWR VPWR _5025_/X sky130_fd_sc_hd__o211a_1
Xhold1148 hold454/X VGND VGND VPWR VPWR _5215_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1159 hold369/X VGND VGND VPWR VPWR _5342_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_66_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6976_ _7140_/CLK _6976_/D fanout471/X VGND VGND VPWR VPWR _6976_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5927_ _6538_/Q _5651_/X _5688_/X _6582_/Q VGND VGND VPWR VPWR _5927_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5858_ _6844_/Q _5678_/Y _5849_/X _5857_/X _6341_/S VGND VGND VPWR VPWR _5858_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4809_ _4637_/C _4637_/D _4719_/Y _4691_/Y _4583_/B VGND VGND VPWR VPWR _4818_/A
+ sky130_fd_sc_hd__o32a_1
X_5789_ _6937_/Q _5659_/X _5663_/X _7025_/Q _5788_/X VGND VGND VPWR VPWR _5792_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold960 _3997_/X VGND VGND VPWR VPWR hold960/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_134_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold971 _4064_/X VGND VGND VPWR VPWR hold15/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold982 hold982/A VGND VGND VPWR VPWR hold982/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold993 _5478_/X VGND VGND VPWR VPWR hold57/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_122_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2350 _5232_/X VGND VGND VPWR VPWR _6825_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2361 hold624/X VGND VGND VPWR VPWR _5383_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_48_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2372 _7041_/Q VGND VGND VPWR VPWR hold713/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2383 _5453_/X VGND VGND VPWR VPWR _7021_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2394 _7025_/Q VGND VGND VPWR VPWR hold738/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1660 hold592/X VGND VGND VPWR VPWR _4271_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1671 hold854/X VGND VGND VPWR VPWR hold200/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1682 _7062_/Q VGND VGND VPWR VPWR hold467/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1693 _6919_/Q VGND VGND VPWR VPWR hold159/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_151_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6830_ _7053_/CLK _6830_/D fanout454/X VGND VGND VPWR VPWR _6830_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_51_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6761_ _6761_/CLK _6761_/D fanout449/X VGND VGND VPWR VPWR _6761_/Q sky130_fd_sc_hd__dfrtp_4
X_3973_ _6821_/Q _3973_/B VGND VGND VPWR VPWR _3973_/X sky130_fd_sc_hd__and2_4
XFILLER_90_494 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5712_ _7062_/Q _5671_/X _5689_/X _7078_/Q VGND VGND VPWR VPWR _5712_/X sky130_fd_sc_hd__a22o_1
XFILLER_149_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6692_ _6742_/CLK _6692_/D fanout440/X VGND VGND VPWR VPWR _6692_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5643_ _5643_/A _5643_/B VGND VGND VPWR VPWR _5643_/Y sky130_fd_sc_hd__nor2_1
XFILLER_163_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5574_ _5574_/A0 _5583_/A1 _5577_/S VGND VGND VPWR VPWR _5574_/X sky130_fd_sc_hd__mux2_1
Xhold201 hold201/A VGND VGND VPWR VPWR wb_dat_o[27] sky130_fd_sc_hd__buf_12
X_4525_ _4625_/A _5033_/A VGND VGND VPWR VPWR _5067_/A sky130_fd_sc_hd__nand2_2
Xhold212 hold212/A VGND VGND VPWR VPWR wb_dat_o[29] sky130_fd_sc_hd__buf_12
Xhold223 hold223/A VGND VGND VPWR VPWR hold825/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold234 hold234/A VGND VGND VPWR VPWR hold234/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold245 hold245/A VGND VGND VPWR VPWR wb_dat_o[28] sky130_fd_sc_hd__buf_12
XFILLER_144_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold256 hold256/A VGND VGND VPWR VPWR hold256/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4456_ _4450_/A _4450_/B _4451_/A VGND VGND VPWR VPWR _4564_/C sky130_fd_sc_hd__o21a_4
XFILLER_172_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold267 hold267/A VGND VGND VPWR VPWR hold843/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold278 hold278/A VGND VGND VPWR VPWR wb_dat_o[7] sky130_fd_sc_hd__buf_12
XFILLER_171_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold289 hold289/A VGND VGND VPWR VPWR wb_dat_o[6] sky130_fd_sc_hd__buf_12
X_3407_ _6867_/Q _5272_/A _5344_/A _6931_/Q VGND VGND VPWR VPWR _3407_/X sky130_fd_sc_hd__a22o_1
X_7175_ _7204_/CLK _7175_/D fanout482/X VGND VGND VPWR VPWR _7175_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4387_ _4921_/A _4886_/A VGND VGND VPWR VPWR _4387_/Y sky130_fd_sc_hd__nor2_1
XFILLER_86_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6126_ _7121_/Q _5978_/X _6015_/X _7017_/Q _6125_/X VGND VGND VPWR VPWR _6129_/C
+ sky130_fd_sc_hd__a221o_1
X_3338_ _3338_/A _3563_/A VGND VGND VPWR VPWR hold67/A sky130_fd_sc_hd__nor2_8
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6057_ _6854_/Q _5983_/X _5998_/X _6886_/Q VGND VGND VPWR VPWR _6057_/X sky130_fd_sc_hd__a22o_1
XTAP_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3269_ _3268_/X hold909/X _3996_/S VGND VGND VPWR VPWR _3269_/X sky130_fd_sc_hd__mux2_4
XTAP_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5008_ _4683_/A _5007_/Y _4999_/D VGND VGND VPWR VPWR _5022_/A sky130_fd_sc_hd__o21a_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 wire350/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 _5303_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_129 _3950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6959_ _7137_/CLK _6959_/D fanout476/X VGND VGND VPWR VPWR _6959_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_10_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold790 hold790/A VGND VGND VPWR VPWR hold790/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2180 _6784_/Q VGND VGND VPWR VPWR hold791/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_162_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2191 _6593_/Q VGND VGND VPWR VPWR hold450/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1490 _4279_/X VGND VGND VPWR VPWR hold108/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_0__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _3958_/A1
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput306 _3953_/X VGND VGND VPWR VPWR serial_load sky130_fd_sc_hd__buf_12
Xoutput317 hold859/X VGND VGND VPWR VPWR hold282/A sky130_fd_sc_hd__buf_6
X_4310_ _4310_/A _5551_/B VGND VGND VPWR VPWR _4315_/S sky130_fd_sc_hd__and2_2
Xoutput328 hold823/X VGND VGND VPWR VPWR hold218/A sky130_fd_sc_hd__buf_6
XFILLER_153_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput339 hold1297/X VGND VGND VPWR VPWR hold227/A sky130_fd_sc_hd__buf_6
X_5290_ _5290_/A hold13/A VGND VGND VPWR VPWR _5298_/S sky130_fd_sc_hd__and2_4
XFILLER_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4241_ _4241_/A hold13/A VGND VGND VPWR VPWR _4249_/S sky130_fd_sc_hd__and2_4
XFILLER_68_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4172_ _4172_/A0 _5186_/A1 _4175_/S VGND VGND VPWR VPWR _6615_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6813_ _7053_/CLK _6813_/D fanout452/X VGND VGND VPWR VPWR _6813_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_169_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3956_ input84/X _3881_/C _6457_/Q VGND VGND VPWR VPWR _3956_/X sky130_fd_sc_hd__mux2_4
X_6744_ _6757_/CLK _6744_/D fanout447/X VGND VGND VPWR VPWR _6744_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_177_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6675_ _7080_/CLK hold17/X fanout480/X VGND VGND VPWR VPWR _7229_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3887_ _6455_/Q _6434_/Q _6423_/B VGND VGND VPWR VPWR _3969_/B sky130_fd_sc_hd__o21a_4
X_5626_ _7152_/Q _7151_/Q VGND VGND VPWR VPWR _6017_/A sky130_fd_sc_hd__and2b_4
XFILLER_136_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5557_ hold917/X hold20/X _5559_/S VGND VGND VPWR VPWR _5557_/X sky130_fd_sc_hd__mux2_1
X_4508_ _4625_/A _4508_/B VGND VGND VPWR VPWR _5136_/A sky130_fd_sc_hd__nand2_2
XFILLER_172_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5488_ _5488_/A _5551_/B VGND VGND VPWR VPWR _5496_/S sky130_fd_sc_hd__and2_4
XFILLER_104_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7227_ _7227_/A VGND VGND VPWR VPWR _7227_/X sky130_fd_sc_hd__clkbuf_2
X_4439_ _4701_/A _4808_/B VGND VGND VPWR VPWR _4469_/B sky130_fd_sc_hd__xnor2_4
XFILLER_104_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7158_ _7186_/CLK _7158_/D fanout466/X VGND VGND VPWR VPWR _7158_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6109_ _7088_/Q _5638_/X _6015_/X _7016_/Q VGND VGND VPWR VPWR _6109_/X sky130_fd_sc_hd__a22o_1
XFILLER_100_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7089_ _7121_/CLK _7089_/D _6399_/A VGND VGND VPWR VPWR _7089_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_74_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3810_ _6470_/Q _6469_/Q _6468_/Q VGND VGND VPWR VPWR _3904_/A sky130_fd_sc_hd__and3_4
X_4790_ _4411_/Y _4662_/Y _4782_/X VGND VGND VPWR VPWR _4790_/X sky130_fd_sc_hd__o21ba_1
XFILLER_20_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_18 _3396_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3741_ _6901_/Q _5317_/A _4140_/A _6589_/Q _3740_/X VGND VGND VPWR VPWR _3750_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA_29 _5659_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6460_ _6656_/CLK _6460_/D _6410_/X VGND VGND VPWR VPWR _6460_/Q sky130_fd_sc_hd__dfrtp_4
X_3672_ _6481_/Q _3357_/Y _4170_/A _6616_/Q _3671_/X VGND VGND VPWR VPWR _3673_/D
+ sky130_fd_sc_hd__a221o_1
X_5411_ hold638/X _5582_/A1 _5415_/S VGND VGND VPWR VPWR _6984_/D sky130_fd_sc_hd__mux2_1
X_6391_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6391_/X sky130_fd_sc_hd__and2_1
X_5342_ _5342_/A0 _5576_/A1 _5343_/S VGND VGND VPWR VPWR _5342_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5273_ hold782/X _5570_/A1 _5280_/S VGND VGND VPWR VPWR _5273_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7012_ _7132_/CLK _7012_/D fanout459/X VGND VGND VPWR VPWR _7012_/Q sky130_fd_sc_hd__dfrtp_4
X_4224_ _3550_/B _6432_/B _4012_/X _5236_/C _5551_/B VGND VGND VPWR VPWR _4240_/S
+ sky130_fd_sc_hd__o221a_4
XFILLER_141_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4155_ hold241/X _4337_/A1 _4157_/S VGND VGND VPWR VPWR _4155_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4086_ _3675_/Y hold818/A _4091_/S VGND VGND VPWR VPWR _6542_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4988_ _4988_/A _5009_/B VGND VGND VPWR VPWR _5021_/B sky130_fd_sc_hd__nand2_1
XFILLER_168_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6727_ _6727_/CLK _6727_/D fanout450/X VGND VGND VPWR VPWR _6727_/Q sky130_fd_sc_hd__dfrtp_2
X_3939_ _6503_/Q wire1/A _6459_/Q VGND VGND VPWR VPWR _3939_/X sky130_fd_sc_hd__mux2_2
XFILLER_137_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6658_ _6658_/CLK _6658_/D _6425_/X VGND VGND VPWR VPWR _6658_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_137_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5609_ _7147_/Q _7146_/Q VGND VGND VPWR VPWR _5684_/B sky130_fd_sc_hd__and2_4
X_6589_ _6747_/CLK _6589_/D fanout443/X VGND VGND VPWR VPWR _6589_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout374 hold6/X VGND VGND VPWR VPWR _5577_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_143_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout385 _5556_/A1 VGND VGND VPWR VPWR _5583_/A1 sky130_fd_sc_hd__buf_6
Xfanout396 _5581_/A1 VGND VGND VPWR VPWR _5572_/A1 sky130_fd_sc_hd__buf_12
XFILLER_74_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput16 mask_rev_in[20] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__buf_2
XFILLER_168_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput27 mask_rev_in[30] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput38 mgmt_gpio_in[11] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__clkbuf_4
Xinput49 mgmt_gpio_in[21] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__buf_2
XFILLER_182_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5960_ _6746_/Q _5929_/B _5668_/X _6648_/Q _5949_/X VGND VGND VPWR VPWR _5960_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4911_ _4633_/B _4688_/B _4845_/X _4901_/B VGND VGND VPWR VPWR _5107_/A sky130_fd_sc_hd__o211a_1
X_5891_ _6570_/Q _5674_/X _5680_/X _6708_/Q VGND VGND VPWR VPWR _5891_/X sky130_fd_sc_hd__a22o_1
X_4842_ _4590_/Y _4676_/Y _4628_/Y VGND VGND VPWR VPWR _4930_/A sky130_fd_sc_hd__o21a_1
XFILLER_178_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4773_ _4729_/A _4688_/C _4542_/Y VGND VGND VPWR VPWR _4800_/A sky130_fd_sc_hd__o21a_1
X_3724_ _6934_/Q _5353_/A _4152_/A _6600_/Q _3723_/X VGND VGND VPWR VPWR _3725_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6512_ _7080_/CLK _6512_/D fanout480/X VGND VGND VPWR VPWR _6512_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3655_ _3655_/A _3655_/B _3655_/C _3655_/D VGND VGND VPWR VPWR _3674_/B sky130_fd_sc_hd__nor4_1
X_6443_ _3940_/A1 _6443_/D _6398_/X VGND VGND VPWR VPWR hold76/A sky130_fd_sc_hd__dfrtp_1
XFILLER_162_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6374_ _6686_/Q _6374_/A2 _6374_/B1 _6685_/Q _6373_/X VGND VGND VPWR VPWR _6374_/X
+ sky130_fd_sc_hd__a221o_1
X_3586_ _6960_/Q _5380_/A _3431_/Y input64/X _3585_/X VGND VGND VPWR VPWR _3587_/D
+ sky130_fd_sc_hd__a221o_2
X_5325_ _5325_/A0 _5577_/A1 _5325_/S VGND VGND VPWR VPWR _5325_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5256_ hold771/X _5580_/A1 _5262_/S VGND VGND VPWR VPWR _6846_/D sky130_fd_sc_hd__mux2_1
X_4207_ _4207_/A0 _5221_/A1 _4211_/S VGND VGND VPWR VPWR _4207_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5187_ _5187_/A0 _5187_/A1 _5190_/S VGND VGND VPWR VPWR _5187_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4138_ _4138_/A0 _5303_/A1 _4139_/S VGND VGND VPWR VPWR _4138_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4069_ hold262/X _5249_/A1 _4070_/S VGND VGND VPWR VPWR _6528_/D sky130_fd_sc_hd__mux2_1
XFILLER_24_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold608 hold608/A VGND VGND VPWR VPWR hold608/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3440_ _7026_/Q _5452_/A _5407_/A _6986_/Q _3437_/X VGND VGND VPWR VPWR _3444_/B
+ sky130_fd_sc_hd__a221o_1
Xhold619 hold619/A VGND VGND VPWR VPWR hold619/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3371_ _7132_/Q _5569_/A _5326_/A _6916_/Q _3370_/X VGND VGND VPWR VPWR _3371_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5110_ _5110_/A _5110_/B VGND VGND VPWR VPWR _5110_/Y sky130_fd_sc_hd__nand2_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2009 _6511_/Q VGND VGND VPWR VPWR hold120/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6090_ _6839_/Q _6011_/Y _6089_/X VGND VGND VPWR VPWR _6090_/X sky130_fd_sc_hd__o21ba_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _5041_/A _5148_/B _5162_/B VGND VGND VPWR VPWR _5042_/D sky130_fd_sc_hd__and3_1
Xhold1308 hold162/X VGND VGND VPWR VPWR _4242_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1319 _6984_/Q VGND VGND VPWR VPWR hold638/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_38_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6992_ _7123_/CLK _6992_/D fanout478/X VGND VGND VPWR VPWR _6992_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_92_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5943_ _6735_/Q _5656_/X _5679_/X _6592_/Q _5942_/X VGND VGND VPWR VPWR _5943_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5874_ _6594_/Q _5670_/X _5671_/X _6634_/Q _5873_/X VGND VGND VPWR VPWR _5879_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_33_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4825_ _4822_/Y _4825_/B _4825_/C _4924_/B VGND VGND VPWR VPWR _4825_/X sky130_fd_sc_hd__and4b_1
XFILLER_138_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4756_ _5009_/B _4732_/B _4811_/B VGND VGND VPWR VPWR _4757_/D sky130_fd_sc_hd__o21ai_1
X_3707_ input15/X _3307_/Y _3389_/Y _3706_/X VGND VGND VPWR VPWR _3707_/X sky130_fd_sc_hd__a211o_1
XFILLER_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4687_ _4712_/A _4691_/B VGND VGND VPWR VPWR _4688_/C sky130_fd_sc_hd__nand2_8
XFILLER_107_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3638_ _7031_/Q _5461_/A _5169_/A _6771_/Q _3637_/X VGND VGND VPWR VPWR _3645_/A
+ sky130_fd_sc_hd__a221o_1
X_6426_ _6426_/A _6432_/B VGND VGND VPWR VPWR _6426_/X sky130_fd_sc_hd__and2_1
XFILLER_161_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6357_ _6357_/A _6358_/A VGND VGND VPWR VPWR _6357_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3569_ _6952_/Q _5371_/A _5308_/A _6896_/Q _3561_/X VGND VGND VPWR VPWR _3569_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5308_ _5308_/A _5569_/B VGND VGND VPWR VPWR _5316_/S sky130_fd_sc_hd__and2_4
X_6288_ _6281_/X _6283_/X _6288_/C _6339_/B VGND VGND VPWR VPWR _6289_/C sky130_fd_sc_hd__and4bb_2
XFILLER_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2510 _7141_/Q VGND VGND VPWR VPWR _5588_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2521 _7142_/Q VGND VGND VPWR VPWR _5595_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_48_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2532 _6819_/Q VGND VGND VPWR VPWR hold273/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5239_ _5239_/A0 _5518_/A1 _5244_/S VGND VGND VPWR VPWR _5239_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1820 hold255/X VGND VGND VPWR VPWR _5500_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1831 hold801/X VGND VGND VPWR VPWR _4226_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1842 _6628_/Q VGND VGND VPWR VPWR hold515/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1853 _4185_/X VGND VGND VPWR VPWR _6626_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_124_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1864 hold647/X VGND VGND VPWR VPWR _4177_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1875 _6967_/Q VGND VGND VPWR VPWR hold225/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1886 _4211_/X VGND VGND VPWR VPWR _6648_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1897 hold290/X VGND VGND VPWR VPWR _4283_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_16_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold5 hold5/A VGND VGND VPWR VPWR hold5/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4610_ _4610_/A _4611_/A VGND VGND VPWR VPWR _4614_/C sky130_fd_sc_hd__nand2_1
XFILLER_175_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5590_ _6490_/Q _6492_/Q _6491_/Q _3924_/Y VGND VGND VPWR VPWR _5599_/D sky130_fd_sc_hd__o31a_4
XFILLER_175_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4541_ _4971_/A _4724_/C VGND VGND VPWR VPWR _5149_/A sky130_fd_sc_hd__nand2_2
XFILLER_191_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold405 _6503_/Q VGND VGND VPWR VPWR hold405/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold416 hold416/A VGND VGND VPWR VPWR _6834_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4472_ _4564_/C _4486_/B VGND VGND VPWR VPWR _4510_/A sky130_fd_sc_hd__nand2_4
XFILLER_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold427 hold427/A VGND VGND VPWR VPWR hold427/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold438 hold438/A VGND VGND VPWR VPWR hold438/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold449 hold449/A VGND VGND VPWR VPWR hold449/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6211_ _7140_/Q _5977_/X _5985_/X _6908_/Q _6210_/X VGND VGND VPWR VPWR _6211_/X
+ sky130_fd_sc_hd__a221o_1
X_3423_ _3464_/A1 _3422_/Y _3857_/B VGND VGND VPWR VPWR _3423_/X sky130_fd_sc_hd__mux2_1
X_7191_ _7194_/CLK _7191_/D VGND VGND VPWR VPWR _7191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6142_ _6142_/A1 _6342_/S _6140_/X _6141_/X VGND VGND VPWR VPWR _7177_/D sky130_fd_sc_hd__o22a_1
X_3354_ _3354_/A _3487_/A VGND VGND VPWR VPWR _5353_/A sky130_fd_sc_hd__nor2_8
XFILLER_124_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_607 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _7023_/Q _5971_/X _6007_/X _6847_/Q _6068_/X VGND VGND VPWR VPWR _6076_/B
+ sky130_fd_sc_hd__a221o_1
X_3285_ _3305_/B _3285_/B VGND VGND VPWR VPWR _3322_/B sky130_fd_sc_hd__and2b_4
Xhold1105 hold401/X VGND VGND VPWR VPWR _5414_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1116 _5450_/X VGND VGND VPWR VPWR _7019_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1127 hold134/X VGND VGND VPWR VPWR hold1127/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5024_ _5139_/B _5024_/B VGND VGND VPWR VPWR _5024_/Y sky130_fd_sc_hd__nand2_1
Xhold1138 _6708_/Q VGND VGND VPWR VPWR hold155/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1149 _7067_/Q VGND VGND VPWR VPWR hold385/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_54_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6975_ _7047_/CLK _6975_/D fanout459/X VGND VGND VPWR VPWR _6975_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5926_ _5947_/A1 _6342_/S _5924_/X _5925_/X VGND VGND VPWR VPWR _5926_/X sky130_fd_sc_hd__o22a_1
XFILLER_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5857_ _6868_/Q _5673_/X _5850_/X _5851_/X _5856_/X VGND VGND VPWR VPWR _5857_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_139_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4808_ _4808_/A _4808_/B VGND VGND VPWR VPWR _4832_/B sky130_fd_sc_hd__nand2_1
XFILLER_186_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5788_ _7017_/Q _5664_/X _5681_/X _7089_/Q VGND VGND VPWR VPWR _5788_/X sky130_fd_sc_hd__a22o_1
X_4739_ _5011_/A _4712_/Y _4727_/Y _4823_/C _4738_/Y VGND VGND VPWR VPWR _4739_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_5_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6409_ _6409_/A _6423_/B VGND VGND VPWR VPWR _6409_/X sky130_fd_sc_hd__and2_1
XFILLER_150_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold950 _5235_/X VGND VGND VPWR VPWR hold92/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold961 _6906_/Q VGND VGND VPWR VPWR hold961/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_150_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold972 hold15/X VGND VGND VPWR VPWR _6524_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold983 _6930_/Q VGND VGND VPWR VPWR hold983/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_1_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold994 _6954_/Q VGND VGND VPWR VPWR hold994/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2340 _7038_/Q VGND VGND VPWR VPWR hold759/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2351 _6897_/Q VGND VGND VPWR VPWR hold693/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2362 _5383_/X VGND VGND VPWR VPWR _6959_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2373 hold713/X VGND VGND VPWR VPWR _5475_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_185_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2384 _7128_/Q VGND VGND VPWR VPWR hold770/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1650 _5227_/X VGND VGND VPWR VPWR _6821_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2395 hold738/X VGND VGND VPWR VPWR _5457_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1661 _4271_/X VGND VGND VPWR VPWR _6704_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1672 _6548_/Q VGND VGND VPWR VPWR hold676/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1683 hold467/X VGND VGND VPWR VPWR _5499_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1694 hold159/X VGND VGND VPWR VPWR _5338_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_50_csclk _7093_/CLK VGND VGND VPWR VPWR _7124_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_99_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6760_ _6760_/CLK _6760_/D _6433_/A VGND VGND VPWR VPWR _6760_/Q sky130_fd_sc_hd__dfrtp_4
X_3972_ _3972_/A input1/X VGND VGND VPWR VPWR _3972_/X sky130_fd_sc_hd__and2_2
XFILLER_62_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5711_ _6982_/Q _5656_/X _5663_/X _7022_/Q _5710_/X VGND VGND VPWR VPWR _5718_/A
+ sky130_fd_sc_hd__a221o_1
X_6691_ _6691_/CLK _6691_/D fanout445/X VGND VGND VPWR VPWR _6691_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_149_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5642_ _5589_/Y _5604_/Y _5641_/Y _6492_/Q VGND VGND VPWR VPWR _5643_/B sky130_fd_sc_hd__a22o_2
XFILLER_176_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5573_ _5573_/A0 _5582_/A1 _5577_/S VGND VGND VPWR VPWR _5573_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_780 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold202 hold202/A VGND VGND VPWR VPWR hold202/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4524_ _4596_/A _5048_/A VGND VGND VPWR VPWR _5114_/A sky130_fd_sc_hd__nand2_2
XFILLER_156_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold213 hold213/A VGND VGND VPWR VPWR hold213/X sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_18_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7113_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold224 hold224/A VGND VGND VPWR VPWR wb_dat_o[21] sky130_fd_sc_hd__buf_12
Xhold235 hold235/A VGND VGND VPWR VPWR hold829/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold246 hold246/A VGND VGND VPWR VPWR hold246/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4455_ _4590_/B _4488_/B VGND VGND VPWR VPWR _4947_/B sky130_fd_sc_hd__nand2_4
Xhold257 hold257/A VGND VGND VPWR VPWR hold257/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold268 hold268/A VGND VGND VPWR VPWR wb_dat_o[15] sky130_fd_sc_hd__buf_12
XFILLER_132_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold279 hold279/A VGND VGND VPWR VPWR hold279/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3406_ _3406_/A _3406_/B VGND VGND VPWR VPWR _3422_/A sky130_fd_sc_hd__nor2_2
X_4386_ _5011_/A _4578_/A VGND VGND VPWR VPWR _4886_/A sky130_fd_sc_hd__nor2_2
X_7174_ _3950_/A1 _7174_/D fanout482/X VGND VGND VPWR VPWR _7174_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3337_ _3535_/A _3563_/B VGND VGND VPWR VPWR _5533_/A sky130_fd_sc_hd__nor2_8
XFILLER_86_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6125_ _6921_/Q _5995_/X _5997_/X _6953_/Q VGND VGND VPWR VPWR _6125_/X sky130_fd_sc_hd__a22o_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3268_ _6461_/Q _6460_/Q _6657_/Q VGND VGND VPWR VPWR _3268_/X sky130_fd_sc_hd__mux2_1
X_6056_ _7102_/Q _6008_/X _6018_/X _6966_/Q _6055_/X VGND VGND VPWR VPWR _6056_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5007_ _5009_/B _4735_/B _4677_/B _4733_/X VGND VGND VPWR VPWR _5007_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_39_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3199_ _6658_/Q VGND VGND VPWR VPWR _3199_/Y sky130_fd_sc_hd__inv_2
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_108 _6339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_119 _5187_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6958_ _7136_/CLK _6958_/D fanout476/X VGND VGND VPWR VPWR _6958_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_41_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5909_ _6636_/Q _5671_/X _5906_/X _5907_/X _5908_/X VGND VGND VPWR VPWR _5909_/X
+ sky130_fd_sc_hd__a2111o_1
X_6889_ _7103_/CLK _6889_/D fanout472/X VGND VGND VPWR VPWR _6889_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_139_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold780 hold780/A VGND VGND VPWR VPWR hold780/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold791 hold791/A VGND VGND VPWR VPWR hold791/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2170 _4040_/X VGND VGND VPWR VPWR _6505_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2181 hold791/X VGND VGND VPWR VPWR _5179_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_36_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2192 hold450/X VGND VGND VPWR VPWR _4145_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_18_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1480 hold492/X VGND VGND VPWR VPWR _5325_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1491 _6924_/Q VGND VGND VPWR VPWR hold477/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput307 _3952_/X VGND VGND VPWR VPWR serial_resetn sky130_fd_sc_hd__buf_12
Xoutput318 hold837/X VGND VGND VPWR VPWR hold261/A sky130_fd_sc_hd__buf_6
XFILLER_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput329 hold831/X VGND VGND VPWR VPWR hold243/A sky130_fd_sc_hd__buf_6
XFILLER_126_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4240_ _4240_/A0 _4239_/X _4240_/S VGND VGND VPWR VPWR _6667_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4171_ _4171_/A0 _5221_/A1 _4175_/S VGND VGND VPWR VPWR _6614_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6812_ _7053_/CLK _6812_/D fanout454/X VGND VGND VPWR VPWR _6812_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_36_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6743_ _6750_/CLK _6743_/D fanout446/X VGND VGND VPWR VPWR _6743_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_149_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3955_ _3996_/S _3955_/A2 _6423_/B _3954_/Y VGND VGND VPWR VPWR _3955_/X sky130_fd_sc_hd__a22o_2
XFILLER_50_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6674_ _7080_/CLK _6674_/D fanout480/X VGND VGND VPWR VPWR _7228_/A sky130_fd_sc_hd__dfrtp_1
X_3886_ _7158_/Q _6810_/Q _6815_/Q VGND VGND VPWR VPWR _5643_/A sky130_fd_sc_hd__mux2_8
XFILLER_192_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5625_ _7152_/Q _7151_/Q _6491_/Q VGND VGND VPWR VPWR _5631_/A sky130_fd_sc_hd__and3_1
XFILLER_164_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5556_ _5556_/A0 _5556_/A1 _5559_/S VGND VGND VPWR VPWR _7113_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4507_ _4508_/B VGND VGND VPWR VPWR _4507_/Y sky130_fd_sc_hd__inv_2
X_5487_ _5487_/A0 _5577_/A1 _5487_/S VGND VGND VPWR VPWR _7052_/D sky130_fd_sc_hd__mux2_1
XFILLER_104_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7226_ _7226_/A VGND VGND VPWR VPWR _7226_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_160_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4438_ _4485_/B VGND VGND VPWR VPWR _4438_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7157_ _7186_/CLK _7157_/D fanout457/X VGND VGND VPWR VPWR _7157_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4369_ _4955_/A _4513_/B VGND VGND VPWR VPWR _4596_/A sky130_fd_sc_hd__and2_4
XFILLER_58_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6108_ _6936_/Q _5980_/X _6017_/X _7072_/Q _6093_/X VGND VGND VPWR VPWR _6113_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7088_ _7126_/CLK _7088_/D fanout480/X VGND VGND VPWR VPWR _7088_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_18_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6039_ _6039_/A _6039_/B _6039_/C _6039_/D VGND VGND VPWR VPWR _6040_/B sky130_fd_sc_hd__nor4_2
XFILLER_100_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_19 _3422_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3740_ _6853_/Q _5263_/A _4122_/A _6574_/Q VGND VGND VPWR VPWR _3740_/X sky130_fd_sc_hd__a22o_1
XFILLER_41_690 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3671_ input37/X _3293_/Y _4140_/A _6591_/Q VGND VGND VPWR VPWR _3671_/X sky130_fd_sc_hd__a22o_1
X_5410_ _5410_/A0 _5518_/A1 _5415_/S VGND VGND VPWR VPWR _6983_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6390_ _6414_/A _6433_/B VGND VGND VPWR VPWR _6390_/X sky130_fd_sc_hd__and2_1
XFILLER_126_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5341_ _5341_/A0 _5503_/A1 _5343_/S VGND VGND VPWR VPWR _5341_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5272_ _5272_/A _5551_/B VGND VGND VPWR VPWR _5280_/S sky130_fd_sc_hd__and2_4
XFILLER_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7011_ _7140_/CLK _7011_/D fanout469/X VGND VGND VPWR VPWR _7011_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4223_ _3184_/Y _3996_/S _6680_/D _5139_/A _4222_/Y VGND VGND VPWR VPWR _6659_/D
+ sky130_fd_sc_hd__a2111o_1
X_4154_ _4154_/A0 _5186_/A1 _4157_/S VGND VGND VPWR VPWR _4154_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4085_ _3737_/Y hold838/A _4091_/S VGND VGND VPWR VPWR _6541_/D sky130_fd_sc_hd__mux2_1
XFILLER_36_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4987_ _4384_/A _4990_/B _4683_/B _4823_/A VGND VGND VPWR VPWR _5083_/B sky130_fd_sc_hd__o31a_1
XFILLER_149_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6726_ _6817_/CLK _6726_/D fanout445/X VGND VGND VPWR VPWR _6726_/Q sky130_fd_sc_hd__dfrtp_4
X_3938_ _6826_/Q input81/X _3971_/B VGND VGND VPWR VPWR _3938_/X sky130_fd_sc_hd__mux2_8
XFILLER_177_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6657_ _6658_/CLK _6657_/D _6424_/X VGND VGND VPWR VPWR _6657_/Q sky130_fd_sc_hd__dfrtp_4
X_3869_ _3869_/A _3869_/B VGND VGND VPWR VPWR _3869_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_192_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5608_ _6491_/Q _5679_/B VGND VGND VPWR VPWR _5613_/B sky130_fd_sc_hd__nand2_1
X_6588_ _6588_/CLK _6588_/D fanout447/X VGND VGND VPWR VPWR _6588_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_3_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5539_ hold947/X hold20/X _5541_/S VGND VGND VPWR VPWR _5539_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7209_ _7209_/A VGND VGND VPWR VPWR _7209_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_160_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout364 _5730_/S VGND VGND VPWR VPWR _6342_/S sky130_fd_sc_hd__buf_12
XFILLER_101_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout375 hold969/X VGND VGND VPWR VPWR hold970/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout386 _5538_/A1 VGND VGND VPWR VPWR _5556_/A1 sky130_fd_sc_hd__buf_8
Xfanout397 hold2/X VGND VGND VPWR VPWR _5581_/A1 sky130_fd_sc_hd__buf_12
XFILLER_100_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput17 mask_rev_in[21] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput28 mask_rev_in[31] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput39 mgmt_gpio_in[12] VGND VGND VPWR VPWR _3974_/B sky130_fd_sc_hd__buf_4
XFILLER_6_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4910_ _4655_/A _4640_/Y _4655_/B _4704_/C _4791_/A VGND VGND VPWR VPWR _5049_/C
+ sky130_fd_sc_hd__o311a_1
XTAP_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5890_ _6753_/Q _5681_/X _5889_/X VGND VGND VPWR VPWR _5890_/X sky130_fd_sc_hd__a21o_1
XFILLER_61_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4841_ _4917_/D _4915_/B VGND VGND VPWR VPWR _5108_/C sky130_fd_sc_hd__nand2_1
XFILLER_61_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4772_ _5136_/A _4973_/C VGND VGND VPWR VPWR _4959_/B sky130_fd_sc_hd__nand2_1
XFILLER_193_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6511_ _7138_/CLK _6511_/D fanout480/X VGND VGND VPWR VPWR _6511_/Q sky130_fd_sc_hd__dfrtp_1
X_3723_ _6990_/Q _5416_/A _5326_/A _6910_/Q VGND VGND VPWR VPWR _3723_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6442_ _3940_/A1 _6442_/D _6397_/X VGND VGND VPWR VPWR hold18/A sky130_fd_sc_hd__dfrtp_1
XFILLER_173_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3654_ _7039_/Q _5470_/A _4122_/A _6576_/Q _3653_/X VGND VGND VPWR VPWR _3655_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6373_ _6684_/Q _6373_/A2 _6373_/B1 _4218_/Y VGND VGND VPWR VPWR _6373_/X sky130_fd_sc_hd__a22o_1
X_3585_ _6572_/Q _4116_/A _4158_/A _6607_/Q VGND VGND VPWR VPWR _3585_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5324_ _5324_/A0 _5576_/A1 _5325_/S VGND VGND VPWR VPWR _5324_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5255_ hold666/X _5561_/A1 _5262_/S VGND VGND VPWR VPWR _6845_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4206_ _4206_/A _5229_/C VGND VGND VPWR VPWR _4211_/S sky130_fd_sc_hd__and2_4
XFILLER_29_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5186_ _5186_/A0 _5186_/A1 _5190_/S VGND VGND VPWR VPWR _5186_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4137_ hold577/X _5187_/A1 _4139_/S VGND VGND VPWR VPWR _4137_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4068_ _4068_/A0 _5581_/A1 _4070_/S VGND VGND VPWR VPWR _6527_/D sky130_fd_sc_hd__mux2_1
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6709_ _6729_/CLK _6709_/D fanout465/X VGND VGND VPWR VPWR _6709_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_137_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold609 hold609/A VGND VGND VPWR VPWR hold609/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3370_ input42/X _4056_/C _5524_/A _7092_/Q VGND VGND VPWR VPWR _3370_/X sky130_fd_sc_hd__a22o_1
XFILLER_170_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5040_ _4454_/A _4463_/B _4570_/D _4954_/D _5039_/Y VGND VGND VPWR VPWR _5162_/B
+ sky130_fd_sc_hd__o311a_1
Xhold1309 _4242_/X VGND VGND VPWR VPWR hold163/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6991_ _7131_/CLK _6991_/D fanout469/X VGND VGND VPWR VPWR _6991_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5942_ _6642_/Q _5655_/X _5663_/X _6632_/Q _5928_/Y VGND VGND VPWR VPWR _5942_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5873_ _6742_/Q _5929_/B _5678_/B _5872_/Y VGND VGND VPWR VPWR _5873_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4824_ _4995_/A _4698_/Y _4583_/B VGND VGND VPWR VPWR _4825_/C sky130_fd_sc_hd__a21o_1
XFILLER_21_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4755_ _4976_/A _4755_/B _4755_/C _4997_/A VGND VGND VPWR VPWR _4757_/C sky130_fd_sc_hd__and4b_1
XFILLER_193_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3706_ _6974_/Q _5398_/A _4116_/A _6570_/Q _3705_/X VGND VGND VPWR VPWR _3706_/X
+ sky130_fd_sc_hd__a221o_2
X_4686_ _4712_/A _4714_/B _4713_/C VGND VGND VPWR VPWR _4686_/X sky130_fd_sc_hd__and3_1
XFILLER_162_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6425_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6425_/X sky130_fd_sc_hd__and2_1
X_3637_ _6967_/Q _5389_/A _5497_/A _7063_/Q VGND VGND VPWR VPWR _3637_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6356_ _6358_/A _6356_/B VGND VGND VPWR VPWR _6356_/Y sky130_fd_sc_hd__nand2_1
XFILLER_1_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3568_ _6602_/Q _4152_/A _4256_/A _6695_/Q VGND VGND VPWR VPWR _3568_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5307_ _5307_/A0 _5577_/A1 _5307_/S VGND VGND VPWR VPWR _5307_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6287_ _6452_/Q _6016_/X _6284_/X _6286_/X VGND VGND VPWR VPWR _6288_/C sky130_fd_sc_hd__a211oi_2
XFILLER_88_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3499_ _3499_/A _3499_/B _3499_/C _3499_/D VGND VGND VPWR VPWR _3558_/B sky130_fd_sc_hd__nor4_2
Xhold2500 _7153_/Q VGND VGND VPWR VPWR _5629_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2511 _6468_/Q VGND VGND VPWR VPWR _3814_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2522 _7186_/Q VGND VGND VPWR VPWR _6345_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2533 _6814_/Q VGND VGND VPWR VPWR hold115/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5238_ _5238_/A0 hold135/X _5244_/S VGND VGND VPWR VPWR _5238_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1810 _6752_/Q VGND VGND VPWR VPWR hold643/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1821 _5500_/X VGND VGND VPWR VPWR _7063_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1832 _6912_/Q VGND VGND VPWR VPWR hold456/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5169_ _5169_/A _5229_/C VGND VGND VPWR VPWR _5174_/S sky130_fd_sc_hd__and2_2
XFILLER_68_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1843 hold515/X VGND VGND VPWR VPWR _4187_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1854 _6552_/Q VGND VGND VPWR VPWR hold530/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1865 _4177_/X VGND VGND VPWR VPWR _6619_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1876 hold225/X VGND VGND VPWR VPWR _5392_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_83_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1887 _6773_/Q VGND VGND VPWR VPWR hold461/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1898 _4283_/X VGND VGND VPWR VPWR _6714_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold6 hold6/A VGND VGND VPWR VPWR hold6/X sky130_fd_sc_hd__buf_12
XFILLER_75_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4540_ _4601_/A _4569_/C _4537_/X _4894_/A _4539_/Y VGND VGND VPWR VPWR _4540_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_144_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold406 hold406/A VGND VGND VPWR VPWR hold406/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4471_ _4485_/B _4564_/C _4568_/A VGND VGND VPWR VPWR _4611_/A sky130_fd_sc_hd__and3_4
XFILLER_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold417 hold417/A VGND VGND VPWR VPWR hold417/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold428 hold428/A VGND VGND VPWR VPWR _6535_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6210_ _6996_/Q _6014_/X _6017_/X _7076_/Q VGND VGND VPWR VPWR _6210_/X sky130_fd_sc_hd__a22o_1
Xhold439 _7214_/A VGND VGND VPWR VPWR hold439/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3422_ _3422_/A _3422_/B _3422_/C VGND VGND VPWR VPWR _3422_/Y sky130_fd_sc_hd__nand3_4
X_7190_ _7194_/CLK _7190_/D VGND VGND VPWR VPWR _7190_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6141_ _6141_/A1 _3924_/Y _5647_/Y VGND VGND VPWR VPWR _6141_/X sky130_fd_sc_hd__o21ba_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _3353_/A hold26/X VGND VGND VPWR VPWR hold27/A sky130_fd_sc_hd__nor2_8
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6072_ _6991_/Q _6014_/X _6070_/X _6071_/X VGND VGND VPWR VPWR _6076_/A sky130_fd_sc_hd__a211o_1
XFILLER_85_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ hold89/X hold53/A VGND VGND VPWR VPWR _3431_/A sky130_fd_sc_hd__nand2_8
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1106 _6867_/Q VGND VGND VPWR VPWR hold363/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1117 _7066_/Q VGND VGND VPWR VPWR hold438/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1128 _4160_/X VGND VGND VPWR VPWR _6605_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5023_ _5023_/A _5083_/C _5023_/C _5023_/D VGND VGND VPWR VPWR _5024_/B sky130_fd_sc_hd__and4_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1139 hold155/X VGND VGND VPWR VPWR _4276_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_38_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6974_ _7133_/CLK _6974_/D fanout472/X VGND VGND VPWR VPWR _6974_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5925_ _6490_/Q _7169_/Q _5649_/Y VGND VGND VPWR VPWR _5925_/X sky130_fd_sc_hd__a21o_1
X_5856_ _6892_/Q _5688_/X _5852_/X _5853_/X _5855_/X VGND VGND VPWR VPWR _5856_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_21_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4807_ _4947_/A _4590_/Y _4370_/Y VGND VGND VPWR VPWR _5114_/B sky130_fd_sc_hd__a21o_2
XFILLER_21_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5787_ _6929_/Q _5684_/X _5689_/X _7081_/Q _5786_/X VGND VGND VPWR VPWR _5792_/B
+ sky130_fd_sc_hd__a221o_1
X_4738_ _5009_/A _4738_/B _5150_/C VGND VGND VPWR VPWR _4738_/Y sky130_fd_sc_hd__nand3_1
XFILLER_135_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4669_ _4638_/Y _4995_/A _4668_/Y _4583_/B VGND VGND VPWR VPWR _4669_/X sky130_fd_sc_hd__o22a_1
XFILLER_79_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6408_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6408_/X sky130_fd_sc_hd__and2_1
XFILLER_162_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold940 _6522_/Q VGND VGND VPWR VPWR hold60/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold951 _6915_/Q VGND VGND VPWR VPWR hold951/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold962 hold962/A VGND VGND VPWR VPWR hold962/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_134_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold973 _6516_/Q VGND VGND VPWR VPWR hold973/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold984 hold984/A VGND VGND VPWR VPWR hold984/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_6339_ _6330_/X _6339_/B _6339_/C _6339_/D VGND VGND VPWR VPWR _6339_/X sky130_fd_sc_hd__and4b_1
Xhold995 hold995/A VGND VGND VPWR VPWR hold995/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_131_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2330 _6998_/Q VGND VGND VPWR VPWR hold753/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2341 _7039_/Q VGND VGND VPWR VPWR hold607/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2352 hold693/X VGND VGND VPWR VPWR _5313_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2363 _7086_/Q VGND VGND VPWR VPWR hold769/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2374 _7093_/Q VGND VGND VPWR VPWR hold802/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1640 _6567_/Q VGND VGND VPWR VPWR hold862/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2385 hold770/X VGND VGND VPWR VPWR _5573_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1651 _6857_/Q VGND VGND VPWR VPWR hold99/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2396 _5457_/X VGND VGND VPWR VPWR _7025_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1662 _6691_/Q VGND VGND VPWR VPWR hold479/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1673 hold676/X VGND VGND VPWR VPWR _4093_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1684 _5499_/X VGND VGND VPWR VPWR _7062_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1695 _7012_/Q VGND VGND VPWR VPWR hold553/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_151_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3971_ _3971_/A _3971_/B VGND VGND VPWR VPWR _3971_/X sky130_fd_sc_hd__and2_2
XFILLER_189_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5710_ _6998_/Q _5666_/X _5673_/X _6862_/Q VGND VGND VPWR VPWR _5710_/X sky130_fd_sc_hd__a22o_1
X_6690_ _6691_/CLK _6690_/D fanout450/X VGND VGND VPWR VPWR _6690_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5641_ _5645_/C _5641_/B VGND VGND VPWR VPWR _5641_/Y sky130_fd_sc_hd__nand2_1
XFILLER_191_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5572_ _5572_/A0 _5572_/A1 _5577_/S VGND VGND VPWR VPWR _5572_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4523_ _4523_/A _4595_/B VGND VGND VPWR VPWR _4523_/Y sky130_fd_sc_hd__nand2_8
XFILLER_8_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold203 hold203/A VGND VGND VPWR VPWR hold203/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold214 hold214/A VGND VGND VPWR VPWR wb_dat_o[31] sky130_fd_sc_hd__buf_12
Xhold225 hold225/A VGND VGND VPWR VPWR hold225/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold236 hold236/A VGND VGND VPWR VPWR wb_dat_o[14] sky130_fd_sc_hd__buf_12
XFILLER_132_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4454_ _4454_/A _4463_/B VGND VGND VPWR VPWR _4724_/C sky130_fd_sc_hd__nor2_8
Xhold247 hold247/A VGND VGND VPWR VPWR wb_dat_o[1] sky130_fd_sc_hd__buf_12
Xhold258 hold258/A VGND VGND VPWR VPWR hold835/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold269 hold269/A VGND VGND VPWR VPWR hold269/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3405_ _3391_/Y _3392_/X _3402_/X _3403_/X _3404_/X VGND VGND VPWR VPWR _3406_/B
+ sky130_fd_sc_hd__a2111o_1
X_7173_ _7203_/CLK _7173_/D fanout468/X VGND VGND VPWR VPWR _7173_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4385_ _5001_/A _4751_/B VGND VGND VPWR VPWR _4578_/A sky130_fd_sc_hd__nand2_2
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6124_ _6857_/Q _5983_/X _5993_/X _7009_/Q _6123_/X VGND VGND VPWR VPWR _6129_/B
+ sky130_fd_sc_hd__a221o_1
X_3336_ _3338_/A _3686_/B VGND VGND VPWR VPWR _3336_/Y sky130_fd_sc_hd__nor2_8
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _6862_/Q _5999_/X _6007_/X _6846_/Q VGND VGND VPWR VPWR _6055_/X sky130_fd_sc_hd__a22o_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _3267_/A hold66/X VGND VGND VPWR VPWR _3355_/A sky130_fd_sc_hd__and2_4
XFILLER_39_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _5139_/A _5140_/A VGND VGND VPWR VPWR _5006_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3198_ _6491_/Q VGND VGND VPWR VPWR _5647_/B sky130_fd_sc_hd__clkinv_4
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_109 _6339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6957_ _7018_/CLK _6957_/D fanout460/X VGND VGND VPWR VPWR _6957_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_41_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5908_ _6749_/Q _5666_/X _5689_/X _6626_/Q VGND VGND VPWR VPWR _5908_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6888_ _7131_/CLK _6888_/D fanout469/X VGND VGND VPWR VPWR _6888_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5839_ _3243_/Y _5872_/B _5677_/B VGND VGND VPWR VPWR _5839_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_10_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold770 hold770/A VGND VGND VPWR VPWR hold770/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold781 hold781/A VGND VGND VPWR VPWR hold781/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold792 hold792/A VGND VGND VPWR VPWR hold792/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2160 _6576_/Q VGND VGND VPWR VPWR hold567/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_77_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2171 _6510_/Q VGND VGND VPWR VPWR hold744/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_162_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2182 _6785_/Q VGND VGND VPWR VPWR hold730/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2193 _6788_/Q VGND VGND VPWR VPWR hold490/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1470 _4027_/X VGND VGND VPWR VPWR _6499_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1481 _5325_/X VGND VGND VPWR VPWR _6908_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1492 hold477/X VGND VGND VPWR VPWR _5343_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput308 _3971_/X VGND VGND VPWR VPWR spi_sdi sky130_fd_sc_hd__buf_12
XFILLER_126_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput319 hold829/X VGND VGND VPWR VPWR hold236/A sky130_fd_sc_hd__buf_6
XFILLER_99_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4170_ _4170_/A _5229_/C VGND VGND VPWR VPWR _4175_/S sky130_fd_sc_hd__and2_4
XFILLER_68_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6811_ _7013_/CLK _6811_/D fanout452/X VGND VGND VPWR VPWR _6811_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6742_ _6742_/CLK _6742_/D fanout439/X VGND VGND VPWR VPWR _6742_/Q sky130_fd_sc_hd__dfrtp_4
X_3954_ _3996_/S _3954_/B VGND VGND VPWR VPWR _3954_/Y sky130_fd_sc_hd__nor2_2
XFILLER_149_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6673_ _7016_/CLK hold21/X fanout480/X VGND VGND VPWR VPWR _7227_/A sky130_fd_sc_hd__dfrtp_1
X_3885_ _6449_/Q _3885_/A2 _6656_/Q _3904_/A VGND VGND VPWR VPWR _6434_/D sky130_fd_sc_hd__o211a_1
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5624_ _7152_/Q _7151_/Q VGND VGND VPWR VPWR _6014_/A sky130_fd_sc_hd__and2_4
XFILLER_176_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5555_ _5555_/A0 _5555_/A1 _5559_/S VGND VGND VPWR VPWR _7112_/D sky130_fd_sc_hd__mux2_1
XFILLER_191_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4506_ _4506_/A _4840_/A _4917_/B _4917_/C VGND VGND VPWR VPWR _4508_/B sky130_fd_sc_hd__and4_2
X_5486_ _5486_/A0 _5576_/A1 _5487_/S VGND VGND VPWR VPWR _7051_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7225_ _7225_/A VGND VGND VPWR VPWR _7225_/X sky130_fd_sc_hd__clkbuf_2
X_4437_ _4560_/B _4560_/C _4341_/X _4394_/Y VGND VGND VPWR VPWR _4437_/Y sky130_fd_sc_hd__a211oi_1
X_7156_ _3950_/A1 _7156_/D fanout468/X VGND VGND VPWR VPWR _7156_/Q sky130_fd_sc_hd__dfrtp_4
X_4368_ _4368_/A _4368_/B VGND VGND VPWR VPWR _4513_/B sky130_fd_sc_hd__nor2_4
XFILLER_101_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6107_ _7120_/Q _5978_/X _5995_/X _6920_/Q _6106_/X VGND VGND VPWR VPWR _6113_/A
+ sky130_fd_sc_hd__a221o_1
X_3319_ _3764_/B _3549_/B VGND VGND VPWR VPWR _3319_/Y sky130_fd_sc_hd__nor2_8
XFILLER_112_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7087_ _7121_/CLK _7087_/D _6399_/A VGND VGND VPWR VPWR _7087_/Q sky130_fd_sc_hd__dfrtp_4
X_4299_ _4299_/A0 _5221_/A1 _4303_/S VGND VGND VPWR VPWR _6727_/D sky130_fd_sc_hd__mux2_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6038_ _6909_/Q _5991_/X _5993_/X _7005_/Q _6037_/X VGND VGND VPWR VPWR _6039_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_64_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _6810_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_127_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_17_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7102_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3670_ _6847_/Q hold40/A hold27/A _6839_/Q _3669_/X VGND VGND VPWR VPWR _3673_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_9_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5340_ _5340_/A0 _5583_/A1 _5343_/S VGND VGND VPWR VPWR _6921_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5271_ _5271_/A0 _5577_/A1 _5271_/S VGND VGND VPWR VPWR _5271_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7010_ _7084_/CLK _7010_/D fanout456/X VGND VGND VPWR VPWR _7010_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_102_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4222_ _6677_/Q _4222_/B _4222_/C VGND VGND VPWR VPWR _4222_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_68_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4153_ _4153_/A0 _5221_/A1 _4157_/S VGND VGND VPWR VPWR _4153_/X sky130_fd_sc_hd__mux2_1
X_4084_ _3803_/Y hold846/A _4091_/S VGND VGND VPWR VPWR _6540_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4986_ _4716_/Y _5127_/B _4986_/C VGND VGND VPWR VPWR _5005_/B sky130_fd_sc_hd__and3b_1
XFILLER_149_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6725_ _6810_/CLK _6725_/D fanout457/X VGND VGND VPWR VPWR _6725_/Q sky130_fd_sc_hd__dfrtp_4
X_3937_ _6824_/Q input78/X _3971_/B VGND VGND VPWR VPWR _3937_/X sky130_fd_sc_hd__mux2_8
XFILLER_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6656_ _6656_/CLK _6656_/D _6423_/X VGND VGND VPWR VPWR _6656_/Q sky130_fd_sc_hd__dfrtp_4
X_3868_ _6446_/Q _3868_/B VGND VGND VPWR VPWR _3869_/B sky130_fd_sc_hd__nor2_1
XFILLER_165_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5607_ _7147_/Q _7146_/Q VGND VGND VPWR VPWR _5679_/B sky130_fd_sc_hd__nor2_8
X_6587_ _6757_/CLK _6587_/D fanout447/X VGND VGND VPWR VPWR _6587_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_180_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3799_ _6722_/Q _4292_/A _4310_/A _6737_/Q VGND VGND VPWR VPWR _3799_/X sky130_fd_sc_hd__a22o_1
XFILLER_152_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5538_ _5538_/A0 _5538_/A1 _5541_/S VGND VGND VPWR VPWR _7097_/D sky130_fd_sc_hd__mux2_1
XFILLER_192_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5469_ _5469_/A0 _5559_/A1 _5469_/S VGND VGND VPWR VPWR _7036_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7208_ _7208_/A VGND VGND VPWR VPWR _7208_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7139_ _7139_/CLK _7139_/D fanout478/X VGND VGND VPWR VPWR _7139_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout376 hold78/X VGND VGND VPWR VPWR _5585_/A1 sky130_fd_sc_hd__buf_8
XFILLER_74_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout387 hold1180/X VGND VGND VPWR VPWR _5538_/A1 sky130_fd_sc_hd__clkbuf_16
Xfanout398 _5193_/A1 VGND VGND VPWR VPWR _5186_/A1 sky130_fd_sc_hd__buf_8
XFILLER_100_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput18 mask_rev_in[22] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput29 mask_rev_in[3] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_812 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4840_ _4840_/A _4917_/B _4857_/C VGND VGND VPWR VPWR _4915_/B sky130_fd_sc_hd__and3_1
XFILLER_61_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4771_ _4719_/A _4590_/B _4719_/B _4981_/A _4607_/B VGND VGND VPWR VPWR _4771_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_14_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6510_ _6523_/CLK _6510_/D fanout480/X VGND VGND VPWR VPWR _6510_/Q sky130_fd_sc_hd__dfrtp_1
X_3722_ _7014_/Q _5443_/A _3648_/Y _6819_/Q _3721_/X VGND VGND VPWR VPWR _3725_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6441_ _3940_/A1 _6441_/D _6396_/X VGND VGND VPWR VPWR _6441_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3653_ input13/X _3310_/Y _3562_/Y input97/X VGND VGND VPWR VPWR _3653_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6372_ _6371_/X _6372_/A1 _6384_/S VGND VGND VPWR VPWR _7198_/D sky130_fd_sc_hd__mux2_1
X_3584_ input55/X _4241_/A _4286_/A _6720_/Q _3566_/X VGND VGND VPWR VPWR _3587_/C
+ sky130_fd_sc_hd__a221o_1
X_5323_ hold962/X _5575_/A1 _5325_/S VGND VGND VPWR VPWR _5323_/X sky130_fd_sc_hd__mux2_1
X_5254_ hold40/X _5569_/B VGND VGND VPWR VPWR _5262_/S sky130_fd_sc_hd__and2_4
X_4205_ _4205_/A0 _5196_/A1 _4205_/S VGND VGND VPWR VPWR _6643_/D sky130_fd_sc_hd__mux2_1
X_5185_ _5185_/A0 _5208_/A1 _5190_/S VGND VGND VPWR VPWR _5185_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_6_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_6_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4136_ _4136_/A0 _5186_/A1 _4139_/S VGND VGND VPWR VPWR _4136_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4067_ _4067_/A0 _5544_/A1 _4070_/S VGND VGND VPWR VPWR _4067_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4969_ _4969_/A _4969_/B VGND VGND VPWR VPWR _5001_/B sky130_fd_sc_hd__nand2_1
XFILLER_184_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6708_ _6760_/CLK _6708_/D _6433_/A VGND VGND VPWR VPWR _6708_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_149_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6639_ _6793_/CLK _6639_/D fanout443/X VGND VGND VPWR VPWR _6639_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6990_ _7123_/CLK _6990_/D fanout477/X VGND VGND VPWR VPWR _6990_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_81_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5941_ _6690_/Q _5659_/X _5687_/X _6602_/Q VGND VGND VPWR VPWR _5941_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5872_ _6717_/Q _5872_/B VGND VGND VPWR VPWR _5872_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4823_ _4823_/A _5083_/A _4823_/C VGND VGND VPWR VPWR _4825_/B sky130_fd_sc_hd__and3_1
XFILLER_179_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4754_ _4722_/X _4754_/B _5083_/A _4754_/D VGND VGND VPWR VPWR _4755_/B sky130_fd_sc_hd__and4b_1
X_3705_ _7110_/Q _5551_/A _5407_/A _6982_/Q VGND VGND VPWR VPWR _3705_/X sky130_fd_sc_hd__a22o_1
X_4685_ _4717_/B _4691_/B VGND VGND VPWR VPWR _4688_/B sky130_fd_sc_hd__nand2_8
XFILLER_146_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3636_ _3636_/A _3636_/B _3636_/C _3636_/D VGND VGND VPWR VPWR _3636_/Y sky130_fd_sc_hd__nor4_1
X_6424_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6424_/X sky130_fd_sc_hd__and2_1
XFILLER_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6355_ _6358_/A _6355_/A2 _6682_/Q VGND VGND VPWR VPWR _6355_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_115_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3567_ _6888_/Q _5299_/A _4128_/A _6582_/Q VGND VGND VPWR VPWR _3567_/X sky130_fd_sc_hd__a22o_1
X_5306_ _5306_/A0 _5576_/A1 _5307_/S VGND VGND VPWR VPWR _5306_/X sky130_fd_sc_hd__mux2_1
X_6286_ _6581_/Q _5998_/X _6004_/X _6576_/Q _6285_/X VGND VGND VPWR VPWR _6286_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3498_ _6613_/Q _4164_/A _4328_/A _6756_/Q _3495_/X VGND VGND VPWR VPWR _3499_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2501 _6434_/Q VGND VGND VPWR VPWR _3885_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5237_ _5237_/A0 _5552_/A1 _5244_/S VGND VGND VPWR VPWR _5237_/X sky130_fd_sc_hd__mux2_1
Xhold2512 _7148_/Q VGND VGND VPWR VPWR _5614_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2523 _6457_/Q VGND VGND VPWR VPWR _3853_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2534 _6653_/Q VGND VGND VPWR VPWR hold116/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1800 _6549_/Q VGND VGND VPWR VPWR hold564/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1811 hold643/X VGND VGND VPWR VPWR _4329_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1822 _6911_/Q VGND VGND VPWR VPWR hold256/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5168_ _5137_/X _5162_/Y _5167_/X _5159_/Y VGND VGND VPWR VPWR _6768_/D sky130_fd_sc_hd__a211o_1
XFILLER_57_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1833 hold456/X VGND VGND VPWR VPWR _5330_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1844 _4187_/X VGND VGND VPWR VPWR _6628_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1855 hold530/X VGND VGND VPWR VPWR _4097_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4119_ hold294/X _5581_/A1 _4121_/S VGND VGND VPWR VPWR _4119_/X sky130_fd_sc_hd__mux2_1
Xhold1866 _6944_/Q VGND VGND VPWR VPWR hold471/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1877 _7208_/A VGND VGND VPWR VPWR hold464/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_83_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5099_ _4611_/A _4981_/B _5095_/Y _4897_/B VGND VGND VPWR VPWR _5099_/X sky130_fd_sc_hd__a211o_1
Xhold1888 hold461/X VGND VGND VPWR VPWR _5174_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1899 _6968_/Q VGND VGND VPWR VPWR hold491/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold7 hold7/A VGND VGND VPWR VPWR hold7/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4470_ _4485_/B _4568_/A VGND VGND VPWR VPWR _4486_/B sky130_fd_sc_hd__and2_2
XFILLER_171_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold407 hold407/A VGND VGND VPWR VPWR hold407/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold418 hold418/A VGND VGND VPWR VPWR hold418/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold429 hold429/A VGND VGND VPWR VPWR hold429/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3421_ _3421_/A _3421_/B _3421_/C _3421_/D VGND VGND VPWR VPWR _3422_/C sky130_fd_sc_hd__nor4_4
XFILLER_109_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6140_ _6841_/Q _6011_/Y _6139_/Y _6341_/S VGND VGND VPWR VPWR _6140_/X sky130_fd_sc_hd__o211a_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3352_ hold52/A hold25/X VGND VGND VPWR VPWR _3648_/B sky130_fd_sc_hd__nand2_8
XFILLER_171_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _6903_/Q _5985_/X _5994_/X _7063_/Q _6069_/X VGND VGND VPWR VPWR _6071_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ hold89/X hold53/X VGND VGND VPWR VPWR hold90/A sky130_fd_sc_hd__and2_2
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1107 hold363/X VGND VGND VPWR VPWR _5279_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5022_ _5022_/A _5080_/B _5022_/C _5140_/B VGND VGND VPWR VPWR _5023_/D sky130_fd_sc_hd__and4_1
Xhold1118 hold438/X VGND VGND VPWR VPWR _5503_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1129 _6794_/Q VGND VGND VPWR VPWR hold437/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_39_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6973_ _7125_/CLK _6973_/D fanout454/X VGND VGND VPWR VPWR _6973_/Q sky130_fd_sc_hd__dfstp_2
X_5924_ _6527_/Q _5678_/Y _5914_/X _5923_/X _6341_/S VGND VGND VPWR VPWR _5924_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5855_ _7068_/Q _5671_/X _5854_/X VGND VGND VPWR VPWR _5855_/X sky130_fd_sc_hd__a21o_1
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4806_ _4933_/C _5044_/A _4805_/X _4374_/Y VGND VGND VPWR VPWR _4906_/A sky130_fd_sc_hd__a31o_1
X_5786_ _6993_/Q _5929_/B _5678_/B _5785_/Y VGND VGND VPWR VPWR _5786_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4737_ _4718_/X _4733_/X _4734_/Y _4738_/B VGND VGND VPWR VPWR _4737_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_119_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4668_ _4712_/A _4712_/B _4672_/B VGND VGND VPWR VPWR _4668_/Y sky130_fd_sc_hd__nand3_4
XFILLER_134_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6407_ _6426_/A _6432_/B VGND VGND VPWR VPWR _6407_/X sky130_fd_sc_hd__and2_1
X_3619_ _6959_/Q _5380_/A _4280_/A _6714_/Q VGND VGND VPWR VPWR _3619_/X sky130_fd_sc_hd__a22o_1
Xhold930 _7122_/Q VGND VGND VPWR VPWR hold930/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_134_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4599_ _4625_/A _5048_/A _4981_/A VGND VGND VPWR VPWR _5112_/A sky130_fd_sc_hd__o21ai_1
Xhold941 hold60/X VGND VGND VPWR VPWR hold941/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold952 _5333_/X VGND VGND VPWR VPWR hold79/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_162_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold963 _5323_/X VGND VGND VPWR VPWR _6906_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold974 hold974/A VGND VGND VPWR VPWR hold974/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_6338_ _6338_/A _6338_/B _6338_/C _6338_/D VGND VGND VPWR VPWR _6339_/D sky130_fd_sc_hd__nor4_1
Xhold985 _5350_/X VGND VGND VPWR VPWR _6930_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold996 _5377_/X VGND VGND VPWR VPWR _6954_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6269_ _6621_/Q _5993_/X _6018_/X _6719_/Q _6268_/X VGND VGND VPWR VPWR _6269_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2320 _6718_/Q VGND VGND VPWR VPWR hold768/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2331 _5427_/X VGND VGND VPWR VPWR _6998_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2342 hold607/X VGND VGND VPWR VPWR _5473_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2353 _5313_/X VGND VGND VPWR VPWR _6897_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2364 _5526_/X VGND VGND VPWR VPWR _7086_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1630 _6742_/Q VGND VGND VPWR VPWR hold677/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2375 _6847_/Q VGND VGND VPWR VPWR hold633/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1641 hold862/X VGND VGND VPWR VPWR hold288/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_151_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2386 _5573_/X VGND VGND VPWR VPWR _7128_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1652 _6690_/Q VGND VGND VPWR VPWR hold627/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2397 _6849_/Q VGND VGND VPWR VPWR hold724/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1663 hold479/X VGND VGND VPWR VPWR _4255_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1674 _6582_/Q VGND VGND VPWR VPWR hold625/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1685 _7079_/Q VGND VGND VPWR VPWR hold184/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1696 hold553/X VGND VGND VPWR VPWR _5442_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3970_ _3970_/A _3970_/B VGND VGND VPWR VPWR _3970_/X sky130_fd_sc_hd__and2_2
XFILLER_50_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5640_ _5640_/A1 _5638_/X _5639_/Y _7156_/Q VGND VGND VPWR VPWR _5640_/X sky130_fd_sc_hd__a22o_1
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5571_ _5571_/A0 _5571_/A1 _5577_/S VGND VGND VPWR VPWR _5571_/X sky130_fd_sc_hd__mux2_1
X_4522_ _4594_/A _4522_/B VGND VGND VPWR VPWR _5048_/A sky130_fd_sc_hd__nor2_4
XFILLER_129_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold204 hold204/A VGND VGND VPWR VPWR hold819/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold215 hold215/A VGND VGND VPWR VPWR hold215/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold226 hold226/A VGND VGND VPWR VPWR hold226/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4453_ _4483_/B _4598_/C VGND VGND VPWR VPWR _4569_/B sky130_fd_sc_hd__nand2_4
Xhold237 hold237/A VGND VGND VPWR VPWR hold237/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold248 hold248/A VGND VGND VPWR VPWR hold248/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3404_ input18/X _3310_/Y _4241_/A input59/X _3394_/X VGND VGND VPWR VPWR _3404_/X
+ sky130_fd_sc_hd__a221o_1
Xhold259 hold259/A VGND VGND VPWR VPWR wb_dat_o[9] sky130_fd_sc_hd__buf_12
XFILLER_144_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7172_ _7186_/CLK _7172_/D fanout465/X VGND VGND VPWR VPWR _7172_/Q sky130_fd_sc_hd__dfrtp_4
X_4384_ _4384_/A _4675_/A VGND VGND VPWR VPWR _4988_/A sky130_fd_sc_hd__nor2_4
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6123_ _7129_/Q _5973_/X _6014_/X _6993_/Q VGND VGND VPWR VPWR _6123_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3335_ _3487_/A _3726_/A VGND VGND VPWR VPWR _5326_/A sky130_fd_sc_hd__nor2_8
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6054_ _6054_/A _6054_/B _6054_/C _6054_/D VGND VGND VPWR VPWR _6064_/B sky130_fd_sc_hd__nor4_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3266_ _3265_/X hold889/X _3996_/S VGND VGND VPWR VPWR _3266_/X sky130_fd_sc_hd__mux2_4
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _5114_/B _5005_/B _5124_/C VGND VGND VPWR VPWR _5140_/A sky130_fd_sc_hd__and3_1
XFILLER_100_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3197_ _6492_/Q VGND VGND VPWR VPWR _3197_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6956_ _7130_/CLK hold46/X fanout458/X VGND VGND VPWR VPWR _6956_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5907_ _6744_/Q _5929_/B _5686_/X _6621_/Q VGND VGND VPWR VPWR _5907_/X sky130_fd_sc_hd__a22o_1
X_6887_ _7109_/CLK _6887_/D fanout452/X VGND VGND VPWR VPWR _6887_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5838_ _5838_/A0 _5837_/X _6342_/S VGND VGND VPWR VPWR _5838_/X sky130_fd_sc_hd__mux2_1
X_5769_ _7024_/Q _5663_/X _5673_/X _6864_/Q _5768_/X VGND VGND VPWR VPWR _5770_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_30_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold760 hold760/A VGND VGND VPWR VPWR hold760/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold771 hold771/A VGND VGND VPWR VPWR hold771/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold782 hold782/A VGND VGND VPWR VPWR hold782/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold793 hold793/A VGND VGND VPWR VPWR hold793/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2150 _6966_/Q VGND VGND VPWR VPWR hold777/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2161 hold567/X VGND VGND VPWR VPWR _4125_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_162_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2172 hold744/X VGND VGND VPWR VPWR _4049_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2183 hold730/X VGND VGND VPWR VPWR _5180_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2194 hold490/X VGND VGND VPWR VPWR _5183_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1460 _5460_/X VGND VGND VPWR VPWR _7028_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1471 _6980_/Q VGND VGND VPWR VPWR hold507/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_18_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1482 _6551_/Q VGND VGND VPWR VPWR hold340/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1493 _5343_/X VGND VGND VPWR VPWR _6924_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput309 _3965_/X VGND VGND VPWR VPWR spimemio_flash_io0_di sky130_fd_sc_hd__buf_12
XFILLER_181_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6810_ _6810_/CLK _6810_/D fanout453/X VGND VGND VPWR VPWR _6810_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6741_ _6822_/CLK hold98/X fanout453/X VGND VGND VPWR VPWR _6741_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3953_ _7159_/Q _6811_/Q _6815_/Q VGND VGND VPWR VPWR _3953_/X sky130_fd_sc_hd__mux2_4
XFILLER_32_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6672_ _7016_/CLK _6672_/D fanout476/X VGND VGND VPWR VPWR _7226_/A sky130_fd_sc_hd__dfrtp_1
X_3884_ wire1/X _3853_/S _3883_/X _3927_/A1 VGND VGND VPWR VPWR _6435_/D sky130_fd_sc_hd__a22o_1
XFILLER_31_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5623_ _5623_/A VGND VGND VPWR VPWR _7151_/D sky130_fd_sc_hd__inv_2
XFILLER_164_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5554_ _5554_/A0 _5572_/A1 _5559_/S VGND VGND VPWR VPWR _7111_/D sky130_fd_sc_hd__mux2_1
XFILLER_191_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4505_ _4643_/D _4643_/C VGND VGND VPWR VPWR _4917_/C sky130_fd_sc_hd__and2_1
X_5485_ _5485_/A0 _5575_/A1 _5487_/S VGND VGND VPWR VPWR _7050_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7224_ _7224_/A VGND VGND VPWR VPWR _7224_/X sky130_fd_sc_hd__clkbuf_2
X_4436_ _4492_/B _4500_/B _4649_/B VGND VGND VPWR VPWR _4560_/C sky130_fd_sc_hd__a21o_1
XFILLER_104_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4367_ _4420_/A _4420_/C _4461_/B VGND VGND VPWR VPWR _4368_/B sky130_fd_sc_hd__a21bo_2
X_7155_ _7204_/CLK _7155_/D fanout468/X VGND VGND VPWR VPWR _7155_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_59_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3318_ _3355_/A _3390_/B VGND VGND VPWR VPWR _3549_/B sky130_fd_sc_hd__nand2_8
X_6106_ _7104_/Q _6008_/X _6016_/X _7040_/Q VGND VGND VPWR VPWR _6106_/X sky130_fd_sc_hd__a22o_1
X_7086_ _7105_/CLK _7086_/D fanout473/X VGND VGND VPWR VPWR _7086_/Q sky130_fd_sc_hd__dfstp_2
X_4298_ hold90/X _5184_/B _5229_/C VGND VGND VPWR VPWR _4303_/S sky130_fd_sc_hd__and3_4
XFILLER_86_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6037_ _6933_/Q _5980_/X _5990_/X _7053_/Q VGND VGND VPWR VPWR _6037_/X sky130_fd_sc_hd__a22o_1
X_3249_ _3248_/X hold903/X _3996_/S VGND VGND VPWR VPWR _3249_/X sky130_fd_sc_hd__mux2_8
XFILLER_86_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6939_ _7140_/CLK _6939_/D fanout471/X VGND VGND VPWR VPWR _6939_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_csclk _3955_/X VGND VGND VPWR VPWR clkbuf_0_csclk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_151_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold590 hold590/A VGND VGND VPWR VPWR hold590/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1290 hold868/X VGND VGND VPWR VPWR hold229/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5270_ hold356/X _5576_/A1 _5271_/S VGND VGND VPWR VPWR _5270_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4221_ _6678_/Q _6679_/Q _6681_/Q VGND VGND VPWR VPWR _4222_/C sky130_fd_sc_hd__nor3_1
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4152_ _4152_/A _5229_/C VGND VGND VPWR VPWR _4157_/S sky130_fd_sc_hd__and2_4
XFILLER_68_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4083_ _6681_/Q _6346_/B VGND VGND VPWR VPWR _4091_/S sky130_fd_sc_hd__nand2_8
XFILLER_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4985_ _5135_/A _5061_/B _4985_/C _4985_/D VGND VGND VPWR VPWR _4985_/Y sky130_fd_sc_hd__nand4_1
XFILLER_168_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6724_ _6817_/CLK _6724_/D fanout453/X VGND VGND VPWR VPWR _6724_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_20_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3936_ _6823_/Q input80/X _3971_/B VGND VGND VPWR VPWR _3936_/X sky130_fd_sc_hd__mux2_8
XFILLER_177_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_2_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_2_0_csclk/X sky130_fd_sc_hd__clkbuf_8
X_6655_ _6658_/CLK _6655_/D _6422_/X VGND VGND VPWR VPWR _6655_/Q sky130_fd_sc_hd__dfrtp_1
X_3867_ _3867_/A1 _3866_/A _3866_/Y _6446_/Q VGND VGND VPWR VPWR _3867_/X sky130_fd_sc_hd__o22a_1
XFILLER_191_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5606_ _6491_/Q _5604_/Y _5606_/S VGND VGND VPWR VPWR _5606_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6586_ _6742_/CLK _6586_/D fanout439/X VGND VGND VPWR VPWR _6586_/Q sky130_fd_sc_hd__dfstp_2
X_3798_ _6933_/Q _5353_/A _4239_/S _3972_/A _3797_/X VGND VGND VPWR VPWR _3801_/C
+ sky130_fd_sc_hd__a221o_1
X_5537_ _5537_/A0 _5582_/A1 _5541_/S VGND VGND VPWR VPWR _7096_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5468_ hold936/X hold78/X _5469_/S VGND VGND VPWR VPWR _5468_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7207_ _7207_/A VGND VGND VPWR VPWR _7207_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4419_ _4955_/A _4955_/B _4936_/B VGND VGND VPWR VPWR _4948_/A sky130_fd_sc_hd__and3_2
X_5399_ hold657/X _5570_/A1 _5406_/S VGND VGND VPWR VPWR _6973_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7138_ _7138_/CLK _7138_/D fanout479/X VGND VGND VPWR VPWR _7138_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_113_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout377 hold78/X VGND VGND VPWR VPWR _5576_/A1 sky130_fd_sc_hd__buf_6
XFILLER_143_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout388 _5303_/A1 VGND VGND VPWR VPWR _5195_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7069_ _7109_/CLK _7069_/D fanout457/X VGND VGND VPWR VPWR _7069_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout399 hold135/X VGND VGND VPWR VPWR _5193_/A1 sky130_fd_sc_hd__buf_8
XFILLER_101_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput19 mask_rev_in[23] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__clkbuf_2
XFILLER_183_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4770_ _4770_/A _4770_/B VGND VGND VPWR VPWR _5138_/C sky130_fd_sc_hd__and2_1
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3721_ _6862_/Q _5272_/A _4241_/A input53/X VGND VGND VPWR VPWR _3721_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6440_ _3940_/A1 _6440_/D _6395_/X VGND VGND VPWR VPWR _6440_/Q sky130_fd_sc_hd__dfrtp_1
X_3652_ _6641_/Q _4200_/A _4322_/A _6749_/Q _3651_/X VGND VGND VPWR VPWR _3655_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_174_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6371_ _6684_/Q _6371_/A2 _6371_/B1 _4218_/Y _6370_/X VGND VGND VPWR VPWR _6371_/X
+ sky130_fd_sc_hd__a221o_1
X_3583_ _6904_/Q _5317_/A _5290_/A _6880_/Q _3567_/X VGND VGND VPWR VPWR _3587_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5322_ _5322_/A0 _5583_/A1 _5325_/S VGND VGND VPWR VPWR _6905_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_851 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5253_ _5253_/A0 hold6/X _5253_/S VGND VGND VPWR VPWR _5253_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4204_ _4204_/A0 _5195_/A1 _4205_/S VGND VGND VPWR VPWR _6642_/D sky130_fd_sc_hd__mux2_1
X_5184_ _5226_/B _5184_/B _5220_/C VGND VGND VPWR VPWR _5190_/S sky130_fd_sc_hd__and3_4
XFILLER_96_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4135_ _4135_/A0 _5208_/A1 _4139_/S VGND VGND VPWR VPWR _6584_/D sky130_fd_sc_hd__mux2_1
XFILLER_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_63_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _6822_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_83_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4066_ hold302/X hold153/X _4070_/S VGND VGND VPWR VPWR _4066_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4968_ _4981_/B VGND VGND VPWR VPWR _4968_/Y sky130_fd_sc_hd__inv_2
X_6707_ _6760_/CLK _6707_/D _6433_/A VGND VGND VPWR VPWR _6707_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_177_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3919_ _6686_/Q _3969_/B _3919_/B1 VGND VGND VPWR VPWR _6686_/D sky130_fd_sc_hd__a21o_1
XFILLER_149_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4899_ _5034_/A _5100_/C VGND VGND VPWR VPWR _5073_/C sky130_fd_sc_hd__and2_1
X_6638_ _6750_/CLK _6638_/D fanout446/X VGND VGND VPWR VPWR _6638_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_164_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6569_ _6729_/CLK _6569_/D fanout465/X VGND VGND VPWR VPWR _6569_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_152_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_16_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _6945_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_121_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5940_ _6755_/Q _5681_/X _5935_/X _5936_/X _5939_/X VGND VGND VPWR VPWR _5940_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5871_ _6639_/Q _5655_/X _5662_/X _6584_/Q _5870_/X VGND VGND VPWR VPWR _5879_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4822_ _4729_/A _4698_/Y _4689_/Y VGND VGND VPWR VPWR _4822_/Y sky130_fd_sc_hd__o21ai_1
X_4753_ _4752_/X _4753_/B _5138_/B _4770_/B VGND VGND VPWR VPWR _4754_/B sky130_fd_sc_hd__and4b_1
XFILLER_147_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3704_ _3704_/A _3704_/B _3704_/C VGND VGND VPWR VPWR _3737_/A sky130_fd_sc_hd__and3_1
XFILLER_186_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4684_ _4684_/A _4722_/C VGND VGND VPWR VPWR _4688_/A sky130_fd_sc_hd__nand2_8
X_6423_ _6433_/A _6423_/B VGND VGND VPWR VPWR _6423_/X sky130_fd_sc_hd__and2_1
X_3635_ _6951_/Q _5371_/A _5317_/A _6903_/Q _3634_/X VGND VGND VPWR VPWR _3636_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6354_ _3385_/Y hold866/A _6354_/S VGND VGND VPWR VPWR _7194_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3566_ _7112_/Q _5551_/A _4280_/A _6715_/Q VGND VGND VPWR VPWR _3566_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5305_ _5305_/A0 _5503_/A1 _5307_/S VGND VGND VPWR VPWR _5305_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6285_ _6606_/Q _5982_/X _6005_/X _6694_/Q VGND VGND VPWR VPWR _6285_/X sky130_fd_sc_hd__a22o_1
X_3497_ _3530_/B _3648_/A VGND VGND VPWR VPWR _4328_/A sky130_fd_sc_hd__nor2_8
XFILLER_103_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2502 _6460_/Q VGND VGND VPWR VPWR _3846_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5236_ _6432_/B _5407_/B _5236_/C VGND VGND VPWR VPWR _5244_/S sky130_fd_sc_hd__and3b_4
Xhold2513 hold22/A VGND VGND VPWR VPWR _5147_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2524 _6455_/Q VGND VGND VPWR VPWR _3856_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_124_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2535 _7138_/Q VGND VGND VPWR VPWR hold42/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1801 hold564/X VGND VGND VPWR VPWR _4094_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1812 _4329_/X VGND VGND VPWR VPWR _6752_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1823 hold256/X VGND VGND VPWR VPWR _5329_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5167_ hold110/A _4836_/A _5135_/X _5156_/Y _5166_/X VGND VGND VPWR VPWR _5167_/X
+ sky130_fd_sc_hd__a221o_1
Xhold1834 _6770_/Q VGND VGND VPWR VPWR hold543/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1845 _6701_/Q VGND VGND VPWR VPWR hold534/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1856 _6609_/Q VGND VGND VPWR VPWR hold650/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_110_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4118_ _4118_/A0 _5544_/A1 _4121_/S VGND VGND VPWR VPWR _4118_/X sky130_fd_sc_hd__mux2_1
Xhold1867 hold471/X VGND VGND VPWR VPWR _5366_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5098_ _5098_/A _5098_/B _5098_/C VGND VGND VPWR VPWR _5131_/B sky130_fd_sc_hd__and3_1
Xhold1878 hold464/X VGND VGND VPWR VPWR _4232_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1889 _5174_/X VGND VGND VPWR VPWR _6773_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_83_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4049_ _4049_/A0 _5571_/A1 _4055_/S VGND VGND VPWR VPWR _4049_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold8 hold8/A VGND VGND VPWR VPWR hold8/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire350 _5879_/Y VGND VGND VPWR VPWR wire350/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire372 _4218_/Y VGND VGND VPWR VPWR _4220_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_128_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold408 hold408/A VGND VGND VPWR VPWR hold408/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold419 hold419/A VGND VGND VPWR VPWR hold419/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3420_ _7019_/Q _5443_/A _3315_/Y input9/X _3419_/X VGND VGND VPWR VPWR _3421_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_171_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3351_ hold52/X hold25/X VGND VGND VPWR VPWR _5226_/B sky130_fd_sc_hd__and2_4
XFILLER_140_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3282_ _3333_/A _3338_/A VGND VGND VPWR VPWR _5272_/A sky130_fd_sc_hd__nor2_8
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _7055_/Q _5990_/X _5996_/X _7047_/Q VGND VGND VPWR VPWR _6070_/X sky130_fd_sc_hd__a22o_1
XFILLER_98_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1108 _5279_/X VGND VGND VPWR VPWR _6867_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5021_ _5021_/A _5021_/B _5021_/C VGND VGND VPWR VPWR _5140_/B sky130_fd_sc_hd__and3_1
XFILLER_39_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1119 _5503_/X VGND VGND VPWR VPWR _7066_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6972_ _7084_/CLK _6972_/D fanout455/X VGND VGND VPWR VPWR _6972_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_80_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5923_ _6591_/Q _5679_/X _5915_/X _5917_/X _5922_/X VGND VGND VPWR VPWR _5923_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_22_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5854_ _7004_/Q _5666_/X _5689_/X _7084_/Q VGND VGND VPWR VPWR _5854_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4805_ _4959_/B _4805_/B _5032_/A _5089_/A VGND VGND VPWR VPWR _4805_/X sky130_fd_sc_hd__and4b_1
XFILLER_167_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5785_ _6969_/Q _5872_/B VGND VGND VPWR VPWR _5785_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4736_ _4955_/D _5150_/C VGND VGND VPWR VPWR _4736_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4667_ _4590_/B _4662_/Y _4995_/A _4638_/B VGND VGND VPWR VPWR _4667_/X sky130_fd_sc_hd__o22a_1
XFILLER_119_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6406_ _6426_/A _6432_/B VGND VGND VPWR VPWR _6406_/X sky130_fd_sc_hd__and2_1
X_3618_ _3617_/X _3618_/A1 _3739_/S VGND VGND VPWR VPWR _6777_/D sky130_fd_sc_hd__mux2_1
Xhold920 _5296_/X VGND VGND VPWR VPWR hold55/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_134_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold931 _5566_/X VGND VGND VPWR VPWR hold68/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4598_ _4598_/A _4598_/B _4598_/C _4607_/B VGND VGND VPWR VPWR _5102_/A sky130_fd_sc_hd__nand4_2
XFILLER_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold942 _4062_/X VGND VGND VPWR VPWR hold61/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold953 _7107_/Q VGND VGND VPWR VPWR hold84/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold964 _7130_/Q VGND VGND VPWR VPWR hold964/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_6337_ _6608_/Q _5982_/X _5987_/X _6731_/Q _6319_/X VGND VGND VPWR VPWR _6338_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3549_ _3553_/A _3549_/B VGND VGND VPWR VPWR _3977_/A sky130_fd_sc_hd__nor2_4
Xhold975 _4055_/X VGND VGND VPWR VPWR hold7/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold986 _6964_/Q VGND VGND VPWR VPWR hold43/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold997 _6852_/Q VGND VGND VPWR VPWR hold997/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6268_ _6591_/Q _5985_/X _6012_/X _6749_/Q VGND VGND VPWR VPWR _6268_/X sky130_fd_sc_hd__a22o_1
Xhold2310 _6951_/Q VGND VGND VPWR VPWR hold560/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2321 hold768/X VGND VGND VPWR VPWR _4288_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2332 hold2390/X VGND VGND VPWR VPWR hold540/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2343 _6901_/Q VGND VGND VPWR VPWR hold785/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5219_ hold13/X _5219_/B VGND VGND VPWR VPWR _6816_/D sky130_fd_sc_hd__and2_1
XFILLER_29_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6199_ _6940_/Q _5980_/X _6019_/X _6988_/Q _6198_/X VGND VGND VPWR VPWR _6204_/B
+ sky130_fd_sc_hd__a221o_1
Xhold2354 _6918_/Q VGND VGND VPWR VPWR hold766/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2365 _6520_/Q VGND VGND VPWR VPWR hold704/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1620 _4137_/X VGND VGND VPWR VPWR _6586_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1631 hold677/X VGND VGND VPWR VPWR _4317_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2376 hold633/X VGND VGND VPWR VPWR _5257_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1642 _6812_/Q VGND VGND VPWR VPWR hold228/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2387 _6942_/Q VGND VGND VPWR VPWR hold780/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1653 hold627/X VGND VGND VPWR VPWR _4254_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2398 hold724/X VGND VGND VPWR VPWR _5259_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1664 _4255_/X VGND VGND VPWR VPWR _6691_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1675 hold625/X VGND VGND VPWR VPWR _4132_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1686 hold184/X VGND VGND VPWR VPWR _5518_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_151_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1697 _7188_/Q VGND VGND VPWR VPWR hold844/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5570_ hold787/X _5570_/A1 _5577_/S VGND VGND VPWR VPWR _5570_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4521_ _4596_/A _4917_/D VGND VGND VPWR VPWR _5127_/A sky130_fd_sc_hd__nand2_2
XFILLER_184_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold205 hold205/A VGND VGND VPWR VPWR wb_dat_o[18] sky130_fd_sc_hd__buf_12
X_4452_ _4483_/B _4598_/C VGND VGND VPWR VPWR _4625_/B sky130_fd_sc_hd__and2_1
Xhold216 _4057_/X VGND VGND VPWR VPWR _6517_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold227 hold227/A VGND VGND VPWR VPWR wb_dat_o[3] sky130_fd_sc_hd__buf_12
XFILLER_116_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold238 _5239_/X VGND VGND VPWR VPWR _6831_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold249 hold249/A VGND VGND VPWR VPWR _6820_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3403_ _6979_/Q _5398_/A _3339_/Y _6477_/Q _3393_/X VGND VGND VPWR VPWR _3403_/X
+ sky130_fd_sc_hd__a221o_1
X_7171_ _7186_/CLK _7171_/D fanout466/X VGND VGND VPWR VPWR _7171_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4383_ _4717_/A _4713_/A VGND VGND VPWR VPWR _4675_/A sky130_fd_sc_hd__nand2_2
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6122_ _7137_/Q _5977_/X _6017_/X _7073_/Q _6121_/X VGND VGND VPWR VPWR _6129_/A
+ sky130_fd_sc_hd__a221o_1
X_3334_ _3349_/A _3563_/B VGND VGND VPWR VPWR _5461_/A sky130_fd_sc_hd__nor2_8
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _7118_/Q _5978_/X _6014_/X _6990_/Q _6052_/X VGND VGND VPWR VPWR _6054_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ _3265_/A0 _6462_/Q _6657_/Q VGND VGND VPWR VPWR _3265_/X sky130_fd_sc_hd__mux2_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5004_ _4932_/Y _4964_/X _5003_/X _5139_/A hold37/A VGND VGND VPWR VPWR _6764_/D
+ sky130_fd_sc_hd__o32a_1
X_3196_ _5611_/A VGND VGND VPWR VPWR _5610_/A sky130_fd_sc_hd__clkinv_2
XFILLER_54_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6955_ _7123_/CLK _6955_/D fanout479/X VGND VGND VPWR VPWR _6955_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5906_ _6646_/Q _5668_/X _5684_/X _6606_/Q VGND VGND VPWR VPWR _5906_/X sky130_fd_sc_hd__a22o_1
X_6886_ _7131_/CLK _6886_/D fanout469/X VGND VGND VPWR VPWR _6886_/Q sky130_fd_sc_hd__dfstp_2
X_5837_ _7165_/Q _5836_/X _6341_/S VGND VGND VPWR VPWR _5837_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5768_ _6944_/Q _5658_/X _5687_/X _6920_/Q VGND VGND VPWR VPWR _5768_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4719_ _4719_/A _4719_/B VGND VGND VPWR VPWR _4719_/Y sky130_fd_sc_hd__nand2_1
X_5699_ _6853_/Q _5651_/X _5668_/X _7053_/Q _5698_/X VGND VGND VPWR VPWR _5699_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_175_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold750 hold750/A VGND VGND VPWR VPWR hold750/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold761 hold761/A VGND VGND VPWR VPWR hold761/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold772 hold772/A VGND VGND VPWR VPWR hold772/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold783 hold783/A VGND VGND VPWR VPWR hold783/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold794 hold794/A VGND VGND VPWR VPWR hold794/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2140 _6799_/Q VGND VGND VPWR VPWR hold443/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2151 _7218_/A VGND VGND VPWR VPWR hold610/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2162 _4125_/X VGND VGND VPWR VPWR _6576_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2173 _6722_/Q VGND VGND VPWR VPWR hold812/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_92_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2184 _6786_/Q VGND VGND VPWR VPWR hold588/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_18_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2195 _6749_/Q VGND VGND VPWR VPWR hold621/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1450 _5271_/X VGND VGND VPWR VPWR _6860_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1461 _6488_/Q VGND VGND VPWR VPWR hold164/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1472 hold507/X VGND VGND VPWR VPWR _5406_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1483 _4096_/X VGND VGND VPWR VPWR _6551_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1494 _6569_/Q VGND VGND VPWR VPWR hold316/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6740_ _7013_/CLK _6740_/D fanout453/X VGND VGND VPWR VPWR _6740_/Q sky130_fd_sc_hd__dfrtp_4
X_3952_ _7157_/Q _6812_/Q _6815_/Q VGND VGND VPWR VPWR _3952_/X sky130_fd_sc_hd__mux2_2
XFILLER_189_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6671_ _7016_/CLK _6671_/D fanout476/X VGND VGND VPWR VPWR _7225_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_188_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3883_ _6468_/Q _6437_/Q _3852_/B VGND VGND VPWR VPWR _3883_/X sky130_fd_sc_hd__a21o_1
XFILLER_31_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5622_ _5604_/Y _5640_/A1 _7151_/Q VGND VGND VPWR VPWR _5623_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5553_ hold760/X _5571_/A1 _5559_/S VGND VGND VPWR VPWR _7110_/D sky130_fd_sc_hd__mux2_1
XFILLER_191_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4504_ _4506_/A _4643_/D VGND VGND VPWR VPWR _4504_/X sky130_fd_sc_hd__and2_1
XFILLER_144_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5484_ _5484_/A0 hold95/X _5487_/S VGND VGND VPWR VPWR _7049_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7223_ _7223_/A VGND VGND VPWR VPWR _7223_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4435_ _4649_/B _4492_/B _4500_/B VGND VGND VPWR VPWR _4560_/B sky130_fd_sc_hd__nand3_2
XFILLER_99_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7154_ _7204_/CLK _7154_/D fanout468/X VGND VGND VPWR VPWR _7154_/Q sky130_fd_sc_hd__dfrtp_4
X_4366_ _4701_/A _4365_/B _4917_/A VGND VGND VPWR VPWR _4420_/C sky130_fd_sc_hd__a21o_1
XFILLER_113_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6105_ _7128_/Q _5973_/X _5988_/X _6872_/Q _6104_/X VGND VGND VPWR VPWR _6105_/X
+ sky130_fd_sc_hd__a221o_1
X_3317_ _3355_/A _3390_/B VGND VGND VPWR VPWR _5220_/B sky130_fd_sc_hd__and2_2
XFILLER_101_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7085_ _7117_/CLK _7085_/D fanout456/X VGND VGND VPWR VPWR _7085_/Q sky130_fd_sc_hd__dfstp_2
X_4297_ _4297_/A0 _5196_/A1 _4297_/S VGND VGND VPWR VPWR _6726_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _7133_/Q _5977_/X _5998_/X _6885_/Q _6035_/X VGND VGND VPWR VPWR _6039_/C
+ sky130_fd_sc_hd__a221o_1
X_3248_ _3265_/A0 _6657_/Q _3247_/Y VGND VGND VPWR VPWR _3248_/X sky130_fd_sc_hd__a21bo_1
XFILLER_27_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6938_ _7124_/CLK _6938_/D fanout459/X VGND VGND VPWR VPWR _6938_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6869_ _7077_/CLK _6869_/D fanout456/X VGND VGND VPWR VPWR _6869_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_22_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold580 hold580/A VGND VGND VPWR VPWR hold580/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold591 hold591/A VGND VGND VPWR VPWR hold591/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1280 _5234_/X VGND VGND VPWR VPWR _6827_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_18_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1291 hold229/X VGND VGND VPWR VPWR hold1291/X sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4220_ _6682_/Q _4220_/B VGND VGND VPWR VPWR _5139_/A sky130_fd_sc_hd__nand2b_4
XFILLER_99_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4151_ _4151_/A0 _5196_/A1 _4151_/S VGND VGND VPWR VPWR _6598_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4082_ hold516/X _4339_/A1 _4082_/S VGND VGND VPWR VPWR _4082_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4984_ _5069_/A _4984_/B _4984_/C VGND VGND VPWR VPWR _4985_/D sky130_fd_sc_hd__and3_1
XFILLER_23_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6723_ _6817_/CLK _6723_/D fanout451/X VGND VGND VPWR VPWR _6723_/Q sky130_fd_sc_hd__dfrtp_2
X_3935_ _3204_/Y input82/X _3971_/B VGND VGND VPWR VPWR _3935_/X sky130_fd_sc_hd__mux2_8
XFILLER_149_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6654_ _6658_/CLK _6654_/D _6421_/X VGND VGND VPWR VPWR _6654_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_149_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3866_ _3866_/A _3869_/A VGND VGND VPWR VPWR _3866_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5605_ _5610_/A _5647_/B VGND VGND VPWR VPWR _5605_/Y sky130_fd_sc_hd__nand2_1
XFILLER_164_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6585_ _6742_/CLK _6585_/D fanout439/X VGND VGND VPWR VPWR _6585_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_176_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3797_ _6789_/Q _3427_/Y _5169_/A _6769_/Q VGND VGND VPWR VPWR _3797_/X sky130_fd_sc_hd__a22o_1
XFILLER_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5536_ _5536_/A0 _5572_/A1 _5541_/S VGND VGND VPWR VPWR _7095_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5467_ _5467_/A0 _5503_/A1 _5469_/S VGND VGND VPWR VPWR _7034_/D sky130_fd_sc_hd__mux2_1
X_7206_ _7206_/A VGND VGND VPWR VPWR _7206_/X sky130_fd_sc_hd__clkbuf_2
X_4418_ _4917_/A _4461_/B VGND VGND VPWR VPWR _4936_/B sky130_fd_sc_hd__nor2_1
X_5398_ _5398_/A _5407_/B VGND VGND VPWR VPWR _5406_/S sky130_fd_sc_hd__and2_4
XFILLER_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7137_ _7137_/CLK _7137_/D fanout473/X VGND VGND VPWR VPWR _7137_/Q sky130_fd_sc_hd__dfrtp_4
X_4349_ _4575_/C _4637_/D VGND VGND VPWR VPWR _4718_/A sky130_fd_sc_hd__nand2_8
XFILLER_86_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout356 _6011_/Y VGND VGND VPWR VPWR _6339_/B sky130_fd_sc_hd__buf_12
XFILLER_47_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout378 hold899/X VGND VGND VPWR VPWR hold900/A sky130_fd_sc_hd__buf_6
X_7068_ _7084_/CLK _7068_/D fanout455/X VGND VGND VPWR VPWR _7068_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout389 _5267_/A1 VGND VGND VPWR VPWR _5303_/A1 sky130_fd_sc_hd__buf_12
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6019_ _6019_/A _6019_/B _6019_/C VGND VGND VPWR VPWR _6019_/X sky130_fd_sc_hd__and3_4
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3720_ _6958_/Q _5380_/A _4182_/A _6625_/Q _3719_/X VGND VGND VPWR VPWR _3725_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_147_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3651_ _6887_/Q _5299_/A _4316_/A _6744_/Q VGND VGND VPWR VPWR _3651_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6370_ _6686_/Q _6370_/A2 _6370_/B1 _6685_/Q VGND VGND VPWR VPWR _6370_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3582_ _6690_/Q _4250_/A _4262_/A _6700_/Q _3581_/X VGND VGND VPWR VPWR _3587_/A
+ sky130_fd_sc_hd__a221o_2
X_5321_ _5321_/A0 _5555_/A1 _5325_/S VGND VGND VPWR VPWR _6904_/D sky130_fd_sc_hd__mux2_1
XFILLER_154_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5252_ _5252_/A0 _5585_/A1 _5253_/S VGND VGND VPWR VPWR _6843_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4203_ hold583/X _5187_/A1 _4205_/S VGND VGND VPWR VPWR _6641_/D sky130_fd_sc_hd__mux2_1
X_5183_ _5183_/A0 _5196_/A1 _5183_/S VGND VGND VPWR VPWR _6788_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4134_ _4134_/A _5229_/C VGND VGND VPWR VPWR _4139_/S sky130_fd_sc_hd__and2_4
XFILLER_68_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4065_ _4065_/A hold13/A VGND VGND VPWR VPWR _4070_/S sky130_fd_sc_hd__and2_2
XFILLER_36_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4967_ _4595_/B _4476_/X _4522_/B VGND VGND VPWR VPWR _4981_/B sky130_fd_sc_hd__o21ai_4
X_6706_ _7013_/CLK _6706_/D fanout452/X VGND VGND VPWR VPWR _6706_/Q sky130_fd_sc_hd__dfstp_2
X_3918_ _3918_/A1 _3969_/B _3918_/B1 VGND VGND VPWR VPWR _6685_/D sky130_fd_sc_hd__a21o_1
X_4898_ _4898_/A _4898_/B VGND VGND VPWR VPWR _4902_/A sky130_fd_sc_hd__and2_1
XFILLER_177_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6637_ _6761_/CLK _6637_/D _6426_/A VGND VGND VPWR VPWR _6637_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3849_ _6654_/Q _3904_/A VGND VGND VPWR VPWR _3850_/S sky130_fd_sc_hd__nand2_2
XFILLER_137_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6568_ _6568_/CLK _6568_/D VGND VGND VPWR VPWR _6568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5519_ _5519_/A0 _5582_/A1 _5523_/S VGND VGND VPWR VPWR _7080_/D sky130_fd_sc_hd__mux2_1
X_6499_ _7016_/CLK _6499_/D fanout475/X VGND VGND VPWR VPWR _7220_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_133_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5870_ _6530_/Q _5653_/X _5689_/X _6624_/Q VGND VGND VPWR VPWR _5870_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4821_ _4676_/Y _4688_/A _4691_/Y _4812_/Y VGND VGND VPWR VPWR _4821_/X sky130_fd_sc_hd__a31o_1
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4752_ _4804_/A _4683_/Y _4750_/X _4751_/X VGND VGND VPWR VPWR _4752_/X sky130_fd_sc_hd__a211o_1
XFILLER_21_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3703_ _3703_/A _3703_/B _3703_/C _3703_/D VGND VGND VPWR VPWR _3704_/C sky130_fd_sc_hd__nor4_1
XFILLER_174_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4683_ _4683_/A _4683_/B VGND VGND VPWR VPWR _4683_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6422_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6422_/X sky130_fd_sc_hd__and2_1
X_3634_ _6651_/Q _4212_/A _4176_/A _6621_/Q VGND VGND VPWR VPWR _3634_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6353_ _3422_/Y hold864/A _6354_/S VGND VGND VPWR VPWR _7193_/D sky130_fd_sc_hd__mux2_1
X_3565_ _6856_/Q _5263_/A _4092_/A _6551_/Q VGND VGND VPWR VPWR _3565_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5304_ _5304_/A0 _5556_/A1 _5307_/S VGND VGND VPWR VPWR _6889_/D sky130_fd_sc_hd__mux2_1
X_6284_ _6689_/Q _5980_/X _6008_/X _6739_/Q VGND VGND VPWR VPWR _6284_/X sky130_fd_sc_hd__a22o_1
XFILLER_88_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3496_ _3550_/A _3549_/B VGND VGND VPWR VPWR _4164_/A sky130_fd_sc_hd__nor2_8
XFILLER_130_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5235_ hold949/X hold20/X hold91/X VGND VGND VPWR VPWR _5235_/X sky130_fd_sc_hd__mux2_1
Xhold2503 _3844_/X VGND VGND VPWR VPWR _6461_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2514 _7154_/Q VGND VGND VPWR VPWR _5633_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2525 _6491_/Q VGND VGND VPWR VPWR _5640_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2536 _7011_/Q VGND VGND VPWR VPWR hold360/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1802 _6936_/Q VGND VGND VPWR VPWR hold460/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1813 _6635_/Q VGND VGND VPWR VPWR hold586/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5166_ _5145_/Y _5165_/Y _5140_/X VGND VGND VPWR VPWR _5166_/X sky130_fd_sc_hd__o21a_1
Xhold1824 _6771_/Q VGND VGND VPWR VPWR hold561/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1835 hold543/X VGND VGND VPWR VPWR _5171_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1846 hold534/X VGND VGND VPWR VPWR _4267_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4117_ _4117_/A0 hold153/X _4121_/S VGND VGND VPWR VPWR _4117_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1857 hold650/X VGND VGND VPWR VPWR _4165_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1868 _5366_/X VGND VGND VPWR VPWR _6944_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5097_ _4569_/C _4968_/Y _4542_/Y VGND VGND VPWR VPWR _5098_/C sky130_fd_sc_hd__o21a_1
Xhold1879 _6969_/Q VGND VGND VPWR VPWR hold425/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4048_ hold874/X hold153/X _4055_/S VGND VGND VPWR VPWR _4048_/X sky130_fd_sc_hd__mux2_1
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5999_ _6014_/A _6019_/C _6007_/C VGND VGND VPWR VPWR _5999_/X sky130_fd_sc_hd__and3_4
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput290 _6482_/Q VGND VGND VPWR VPWR pll_trim[3] sky130_fd_sc_hd__buf_12
XFILLER_58_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold9 hold9/A VGND VGND VPWR VPWR hold9/X sky130_fd_sc_hd__buf_8
XFILLER_181_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_62_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7013_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_144_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold409 hold409/A VGND VGND VPWR VPWR hold409/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3350_ _3354_/A _3535_/A VGND VGND VPWR VPWR _5497_/A sky130_fd_sc_hd__nor2_8
XFILLER_124_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ hold31/X _3309_/A VGND VGND VPWR VPWR _3338_/A sky130_fd_sc_hd__nand2_8
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _4993_/A _4727_/A _5001_/A VGND VGND VPWR VPWR _5021_/C sky130_fd_sc_hd__o21ai_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1109 _6883_/Q VGND VGND VPWR VPWR hold410/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_38_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6971_ _7091_/CLK _6971_/D fanout471/X VGND VGND VPWR VPWR _6971_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5922_ _6586_/Q _5662_/X _5919_/X _5921_/X VGND VGND VPWR VPWR _5922_/X sky130_fd_sc_hd__a211o_1
XFILLER_34_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5853_ _6996_/Q _5929_/B _5686_/X _7012_/Q VGND VGND VPWR VPWR _5853_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_15_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7121_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_179_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4804_ _4804_/A _4948_/A VGND VGND VPWR VPWR _5032_/A sky130_fd_sc_hd__nand2_1
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5784_ _6857_/Q _5651_/X _5685_/X _7073_/Q _5783_/X VGND VGND VPWR VPWR _5792_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4735_ _4955_/D _4735_/B VGND VGND VPWR VPWR _4735_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4666_ _4666_/A _5026_/C VGND VGND VPWR VPWR _4995_/A sky130_fd_sc_hd__nand2_8
XFILLER_175_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6405_ _6414_/A _6433_/B VGND VGND VPWR VPWR _6405_/X sky130_fd_sc_hd__and2_1
X_3617_ _3677_/A1 _3616_/Y _3738_/S VGND VGND VPWR VPWR _3617_/X sky130_fd_sc_hd__mux2_1
Xhold910 _3269_/X VGND VGND VPWR VPWR _3272_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_190_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold921 _6946_/Q VGND VGND VPWR VPWR hold80/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4597_ _5033_/A _4724_/C VGND VGND VPWR VPWR _5067_/B sky130_fd_sc_hd__nand2_1
Xhold932 _7219_/A VGND VGND VPWR VPWR hold932/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_134_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold943 _6506_/Q VGND VGND VPWR VPWR hold943/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_6336_ _6552_/Q _5999_/X _6019_/X _6736_/Q _6335_/X VGND VGND VPWR VPWR _6338_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold954 _6762_/Q VGND VGND VPWR VPWR hold29/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_3548_ _6905_/Q _5317_/A _5470_/A _7041_/Q _3547_/X VGND VGND VPWR VPWR _3556_/B
+ sky130_fd_sc_hd__a221o_2
Xhold965 hold965/A VGND VGND VPWR VPWR hold965/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_103_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold976 _7140_/Q VGND VGND VPWR VPWR hold976/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold987 _5388_/X VGND VGND VPWR VPWR hold44/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold998 _5262_/X VGND VGND VPWR VPWR hold41/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6267_ _6291_/A2 _6266_/X _6342_/S VGND VGND VPWR VPWR _6267_/X sky130_fd_sc_hd__mux2_1
Xhold2300 _6578_/Q VGND VGND VPWR VPWR hold575/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3479_ _3550_/A _3516_/B VGND VGND VPWR VPWR _4158_/A sky130_fd_sc_hd__nor2_8
Xhold2311 hold560/X VGND VGND VPWR VPWR _5374_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2322 _6480_/Q VGND VGND VPWR VPWR hold737/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5218_ hold420/X hold153/X _5218_/S VGND VGND VPWR VPWR _5218_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2333 _4035_/X VGND VGND VPWR VPWR _4036_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2344 _6989_/Q VGND VGND VPWR VPWR hold792/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6198_ _6900_/Q _5989_/X _6013_/X _7084_/Q VGND VGND VPWR VPWR _6198_/X sky130_fd_sc_hd__a22o_1
XFILLER_57_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1610 _5397_/X VGND VGND VPWR VPWR _6972_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2355 _6846_/Q VGND VGND VPWR VPWR hold771/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1621 _7224_/A VGND VGND VPWR VPWR hold127/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2366 hold704/X VGND VGND VPWR VPWR _4060_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1632 _7132_/Q VGND VGND VPWR VPWR hold544/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2377 _6727_/Q VGND VGND VPWR VPWR hold800/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5149_ _5149_/A _5149_/B _5149_/C _5149_/D VGND VGND VPWR VPWR _5152_/A sky130_fd_sc_hd__and4_1
Xhold1643 hold228/X VGND VGND VPWR VPWR _5214_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2388 _6518_/Q VGND VGND VPWR VPWR hold742/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1654 _4254_/X VGND VGND VPWR VPWR _6690_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_151_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2399 _7073_/Q VGND VGND VPWR VPWR hold716/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1665 _7226_/A VGND VGND VPWR VPWR hold359/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_151_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1676 _6624_/Q VGND VGND VPWR VPWR hold630/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1687 _6603_/Q VGND VGND VPWR VPWR hold485/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1698 hold844/X VGND VGND VPWR VPWR hold188/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_71_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4520_ _4523_/A _4638_/B VGND VGND VPWR VPWR _4655_/A sky130_fd_sc_hd__nand2_8
XFILLER_157_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold206 hold206/A VGND VGND VPWR VPWR hold206/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4451_ _4451_/A _4451_/B VGND VGND VPWR VPWR _4598_/C sky130_fd_sc_hd__and2_4
XFILLER_171_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold217 hold217/A VGND VGND VPWR VPWR hold823/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold228 hold228/A VGND VGND VPWR VPWR hold228/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold239 hold239/A VGND VGND VPWR VPWR hold827/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3402_ _6883_/Q _5290_/A _3399_/X _3401_/X VGND VGND VPWR VPWR _3402_/X sky130_fd_sc_hd__a211o_1
X_7170_ _7183_/CLK _7170_/D fanout466/X VGND VGND VPWR VPWR _7170_/Q sky130_fd_sc_hd__dfrtp_1
X_4382_ _4717_/A _4713_/A VGND VGND VPWR VPWR _4751_/B sky130_fd_sc_hd__and2_4
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6121_ _7033_/Q _5986_/X _5988_/X _6873_/Q VGND VGND VPWR VPWR _6121_/X sky130_fd_sc_hd__a22o_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _3333_/A _3354_/A VGND VGND VPWR VPWR _5281_/A sky130_fd_sc_hd__nor2_8
XFILLER_124_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6052_ _6894_/Q _5989_/X _6015_/X _7014_/Q VGND VGND VPWR VPWR _6052_/X sky130_fd_sc_hd__a22o_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ _3267_/A VGND VGND VPWR VPWR _3429_/A sky130_fd_sc_hd__inv_2
XFILLER_105_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _5061_/A _4985_/Y _5005_/B _5002_/Y _4836_/A VGND VGND VPWR VPWR _5003_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3195_ _6490_/Q VGND VGND VPWR VPWR _6166_/S sky130_fd_sc_hd__clkinv_4
XFILLER_94_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6954_ _7130_/CLK _6954_/D fanout458/X VGND VGND VPWR VPWR _6954_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5905_ _3201_/Y _5872_/B _5677_/B VGND VGND VPWR VPWR _5905_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_179_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6885_ _7125_/CLK _6885_/D fanout454/X VGND VGND VPWR VPWR _6885_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_50_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5836_ _5826_/Y _5835_/Y _6843_/Q _5678_/Y VGND VGND VPWR VPWR _5836_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_167_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5767_ _6896_/Q _5662_/X _5684_/X _6928_/Q _5766_/X VGND VGND VPWR VPWR _5770_/C
+ sky130_fd_sc_hd__a221o_1
X_4718_ _4718_/A _4719_/A _4718_/C VGND VGND VPWR VPWR _4718_/X sky130_fd_sc_hd__and3_1
XFILLER_5_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5698_ _7029_/Q _5655_/X _5678_/B _6965_/Q _5707_/B VGND VGND VPWR VPWR _5698_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_108_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4649_ _4720_/C _4649_/B _4649_/C _4649_/D VGND VGND VPWR VPWR _4649_/Y sky130_fd_sc_hd__nor4_2
XFILLER_135_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold740 hold740/A VGND VGND VPWR VPWR hold740/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold751 hold751/A VGND VGND VPWR VPWR hold751/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold762 hold762/A VGND VGND VPWR VPWR hold762/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold773 hold773/A VGND VGND VPWR VPWR hold773/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold784 hold784/A VGND VGND VPWR VPWR hold784/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6319_ _6706_/Q _5977_/X _5984_/X _6618_/Q VGND VGND VPWR VPWR _6319_/X sky130_fd_sc_hd__a22o_1
Xhold795 hold795/A VGND VGND VPWR VPWR hold795/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2130 _6735_/Q VGND VGND VPWR VPWR hold648/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_103_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2141 _7057_/Q VGND VGND VPWR VPWR hold719/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2152 hold610/X VGND VGND VPWR VPWR _4023_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2163 _6937_/Q VGND VGND VPWR VPWR hold763/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2174 hold812/X VGND VGND VPWR VPWR _4293_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_92_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1440 _4270_/X VGND VGND VPWR VPWR _6703_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2185 _6748_/Q VGND VGND VPWR VPWR hold568/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1451 _6650_/Q VGND VGND VPWR VPWR _4214_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2196 hold621/X VGND VGND VPWR VPWR _4325_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1462 _4011_/X VGND VGND VPWR VPWR _6488_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1473 _6536_/Q VGND VGND VPWR VPWR hold547/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_176_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1484 _6525_/Q VGND VGND VPWR VPWR hold302/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1495 hold316/X VGND VGND VPWR VPWR _4117_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3951_ _6506_/Q input93/X _6820_/Q VGND VGND VPWR VPWR _3951_/X sky130_fd_sc_hd__mux2_4
XFILLER_189_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6670_ _7016_/CLK _6670_/D fanout476/X VGND VGND VPWR VPWR _7224_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_91_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3882_ _6409_/A _6423_/B VGND VGND VPWR VPWR _3882_/X sky130_fd_sc_hd__and2_1
XFILLER_176_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5621_ _5621_/A VGND VGND VPWR VPWR _7150_/D sky130_fd_sc_hd__inv_2
XFILLER_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5552_ hold809/X _5552_/A1 _5559_/S VGND VGND VPWR VPWR _7109_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4503_ _4637_/B _4808_/B _4701_/A VGND VGND VPWR VPWR _4643_/C sky130_fd_sc_hd__a21o_1
XFILLER_117_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5483_ _5483_/A0 _5555_/A1 _5487_/S VGND VGND VPWR VPWR _7048_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7222_ _7222_/A VGND VGND VPWR VPWR _7222_/X sky130_fd_sc_hd__clkbuf_2
X_4434_ _4447_/B _4663_/D _4682_/A _4808_/B VGND VGND VPWR VPWR _4500_/B sky130_fd_sc_hd__and4_4
XFILLER_117_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7153_ _7204_/CLK _7153_/D fanout468/X VGND VGND VPWR VPWR _7153_/Q sky130_fd_sc_hd__dfrtp_4
X_4365_ _4701_/A _4365_/B VGND VGND VPWR VPWR _4461_/B sky130_fd_sc_hd__xnor2_4
XFILLER_59_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6104_ _6960_/Q _5992_/X _6012_/X _7000_/Q _6103_/X VGND VGND VPWR VPWR _6104_/X
+ sky130_fd_sc_hd__a221o_1
X_3316_ hold32/X _3535_/A VGND VGND VPWR VPWR _5506_/A sky130_fd_sc_hd__nor2_8
X_7084_ _7084_/CLK _7084_/D fanout456/X VGND VGND VPWR VPWR _7084_/Q sky130_fd_sc_hd__dfrtp_4
X_4296_ _4296_/A0 _5303_/A1 _4297_/S VGND VGND VPWR VPWR _4296_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6035_ _7109_/Q _5987_/X _5997_/X _6949_/Q VGND VGND VPWR VPWR _6035_/X sky130_fd_sc_hd__a22o_1
X_3247_ _6464_/Q _3862_/A VGND VGND VPWR VPWR _3247_/Y sky130_fd_sc_hd__nand2_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6937_ _7135_/CLK _6937_/D fanout473/X VGND VGND VPWR VPWR _6937_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6868_ _7130_/CLK _6868_/D fanout458/X VGND VGND VPWR VPWR _6868_/Q sky130_fd_sc_hd__dfrtp_4
X_5819_ _6915_/Q _5670_/X _5682_/X _7043_/Q _5818_/X VGND VGND VPWR VPWR _5826_/A
+ sky130_fd_sc_hd__a221o_1
X_6799_ _6809_/CLK _6799_/D fanout444/X VGND VGND VPWR VPWR _6799_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_167_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold570 hold570/A VGND VGND VPWR VPWR hold570/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold581 hold581/A VGND VGND VPWR VPWR hold581/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold592 hold592/A VGND VGND VPWR VPWR hold592/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1270 hold211/X VGND VGND VPWR VPWR hold1270/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1281 _7018_/Q VGND VGND VPWR VPWR hold531/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1292 _6731_/Q VGND VGND VPWR VPWR hold129/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_18_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4150_ _4150_/A0 _5195_/A1 _4151_/S VGND VGND VPWR VPWR _6597_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4081_ hold328/X _5303_/A1 _4082_/S VGND VGND VPWR VPWR _4081_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4983_ _5103_/B _4983_/B _4983_/C VGND VGND VPWR VPWR _4984_/C sky130_fd_sc_hd__and3_1
XFILLER_23_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6722_ _6822_/CLK _6722_/D fanout451/X VGND VGND VPWR VPWR _6722_/Q sky130_fd_sc_hd__dfrtp_2
X_3934_ _3203_/Y input90/X _3934_/S VGND VGND VPWR VPWR _3934_/X sky130_fd_sc_hd__mux2_4
X_6653_ _6711_/CLK _6653_/D _6414_/A VGND VGND VPWR VPWR _6653_/Q sky130_fd_sc_hd__dfrtp_4
X_3865_ _3870_/A _3870_/B VGND VGND VPWR VPWR _3869_/A sky130_fd_sc_hd__nor2_2
XFILLER_137_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5604_ _6489_/Q _6491_/Q VGND VGND VPWR VPWR _5604_/Y sky130_fd_sc_hd__nor2_1
X_3796_ _6795_/Q _3319_/Y _5299_/A _6885_/Q _3795_/X VGND VGND VPWR VPWR _3801_/B
+ sky130_fd_sc_hd__a221o_1
X_6584_ _6747_/CLK _6584_/D fanout450/X VGND VGND VPWR VPWR _6584_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_191_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5535_ hold222/X _5544_/A1 _5541_/S VGND VGND VPWR VPWR _7094_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5466_ _5466_/A0 _5538_/A1 _5469_/S VGND VGND VPWR VPWR _7033_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4417_ _4947_/A _4417_/B VGND VGND VPWR VPWR _5150_/B sky130_fd_sc_hd__nand2_4
XFILLER_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5397_ _5397_/A0 _5559_/A1 _5397_/S VGND VGND VPWR VPWR _5397_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4348_ _4575_/C _4637_/D VGND VGND VPWR VPWR _4576_/A sky130_fd_sc_hd__and2_4
X_7136_ _7136_/CLK _7136_/D fanout475/X VGND VGND VPWR VPWR _7136_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_86_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7067_ _7091_/CLK _7067_/D fanout472/X VGND VGND VPWR VPWR _7067_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout379 hold20/X VGND VGND VPWR VPWR _5503_/A1 sky130_fd_sc_hd__clkbuf_16
X_4279_ _4279_/A0 _5538_/A1 _4279_/S VGND VGND VPWR VPWR _4279_/X sky130_fd_sc_hd__mux2_1
X_6018_ _6019_/B _6018_/B _6019_/C VGND VGND VPWR VPWR _6018_/X sky130_fd_sc_hd__and3_4
XFILLER_27_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3650_ _7087_/Q _5524_/A _4065_/A _6527_/Q _3649_/X VGND VGND VPWR VPWR _3655_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_159_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3581_ _6848_/Q hold40/A _4077_/A _6538_/Q VGND VGND VPWR VPWR _3581_/X sky130_fd_sc_hd__a22o_1
X_5320_ _5320_/A0 _5320_/A1 _5325_/S VGND VGND VPWR VPWR _5320_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5251_ hold64/X hold20/X _5253_/S VGND VGND VPWR VPWR _5251_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4202_ _4202_/A0 _5186_/A1 _4205_/S VGND VGND VPWR VPWR _6640_/D sky130_fd_sc_hd__mux2_1
X_5182_ _5182_/A0 _5195_/A1 _5183_/S VGND VGND VPWR VPWR _6787_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4133_ _4133_/A0 _4339_/A1 _4133_/S VGND VGND VPWR VPWR _6583_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4064_ _6524_/Q hold6/X hold14/X VGND VGND VPWR VPWR _4064_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4966_ _4581_/X _4969_/B _4878_/Y _4491_/Y _4628_/Y VGND VGND VPWR VPWR _5074_/B
+ sky130_fd_sc_hd__o221a_1
X_6705_ _7013_/CLK _6705_/D fanout453/X VGND VGND VPWR VPWR _6705_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_177_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3917_ _3917_/A1 _3969_/B _3917_/B1 VGND VGND VPWR VPWR _6684_/D sky130_fd_sc_hd__a21o_1
X_4897_ _4921_/B _4897_/B VGND VGND VPWR VPWR _4903_/C sky130_fd_sc_hd__nor2_1
XFILLER_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6636_ _6759_/CLK _6636_/D _6426_/A VGND VGND VPWR VPWR _6636_/Q sky130_fd_sc_hd__dfstp_2
X_3848_ _6470_/Q _6468_/Q _6654_/Q VGND VGND VPWR VPWR _3880_/S sky130_fd_sc_hd__and3_1
XFILLER_137_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3779_ _6817_/Q hold90/A _5220_/B _4194_/A _6634_/Q VGND VGND VPWR VPWR _3779_/X
+ sky130_fd_sc_hd__a32o_1
X_6567_ _6568_/CLK _6567_/D VGND VGND VPWR VPWR _6567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5518_ _5518_/A0 _5518_/A1 _5523_/S VGND VGND VPWR VPWR _7079_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6498_ _7016_/CLK _6498_/D fanout475/X VGND VGND VPWR VPWR _7219_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_145_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5449_ _5449_/A0 _5575_/A1 _5451_/S VGND VGND VPWR VPWR _7018_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7119_ _7119_/CLK _7119_/D fanout470/X VGND VGND VPWR VPWR _7119_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _6385_/A3 sky130_fd_sc_hd__clkbuf_16
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4820_ _4820_/A _4820_/B _4820_/C VGND VGND VPWR VPWR _4834_/A sky130_fd_sc_hd__and3_1
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4751_ _5009_/A _4751_/B _4751_/C VGND VGND VPWR VPWR _4751_/X sky130_fd_sc_hd__and3_1
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3702_ _7022_/Q _5452_/A hold67/A _7118_/Q _3701_/X VGND VGND VPWR VPWR _3703_/D
+ sky130_fd_sc_hd__a221o_2
X_4682_ _4682_/A _4717_/A VGND VGND VPWR VPWR _4683_/B sky130_fd_sc_hd__nand2_2
XFILLER_146_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3633_ _6975_/Q _5398_/A _5281_/A _6871_/Q _3632_/X VGND VGND VPWR VPWR _3636_/C
+ sky130_fd_sc_hd__a221o_1
X_6421_ _6432_/A _6433_/B VGND VGND VPWR VPWR _6421_/X sky130_fd_sc_hd__and2_1
XFILLER_135_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3564_ _7088_/Q _5524_/A _4170_/A _6617_/Q VGND VGND VPWR VPWR _3564_/X sky130_fd_sc_hd__a22o_1
X_6352_ _3462_/Y hold865/A _6354_/S VGND VGND VPWR VPWR _7192_/D sky130_fd_sc_hd__mux2_1
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5303_ _5303_/A0 _5303_/A1 _5307_/S VGND VGND VPWR VPWR _5303_/X sky130_fd_sc_hd__mux2_1
X_6283_ _6611_/Q _5976_/B _5984_/X _6616_/Q _6282_/X VGND VGND VPWR VPWR _6283_/X
+ sky130_fd_sc_hd__a221o_1
X_3495_ _7081_/Q _5515_/A _3391_/Y _6810_/Q VGND VGND VPWR VPWR _3495_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5234_ _5234_/A0 _5538_/A1 hold91/X VGND VGND VPWR VPWR _5234_/X sky130_fd_sc_hd__mux2_1
Xhold2504 _6456_/Q VGND VGND VPWR VPWR _3854_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2515 _6492_/Q VGND VGND VPWR VPWR _3916_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2526 _5640_/X VGND VGND VPWR VPWR _7156_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2537 _6842_/Q VGND VGND VPWR VPWR hold64/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5165_ _5015_/X _5165_/B _5165_/C VGND VGND VPWR VPWR _5165_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1803 hold460/X VGND VGND VPWR VPWR _5357_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1814 hold586/X VGND VGND VPWR VPWR _4196_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1825 hold561/X VGND VGND VPWR VPWR _5172_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1836 _5171_/X VGND VGND VPWR VPWR _6770_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4116_ _4116_/A hold13/A VGND VGND VPWR VPWR _4121_/S sky130_fd_sc_hd__and2_2
XFILLER_83_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1847 _6896_/Q VGND VGND VPWR VPWR hold484/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5096_ _4611_/A _4981_/B _5095_/Y _4897_/B VGND VGND VPWR VPWR _5156_/B sky130_fd_sc_hd__a211oi_2
Xhold1858 _6822_/Q VGND VGND VPWR VPWR _5228_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1869 _6758_/Q VGND VGND VPWR VPWR hold578/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_110_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4047_ _6432_/B hold13/A _4047_/C VGND VGND VPWR VPWR _4055_/S sky130_fd_sc_hd__and3b_4
XFILLER_37_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5998_ _6019_/A _6015_/B _6007_/C VGND VGND VPWR VPWR _5998_/X sky130_fd_sc_hd__and3_4
XFILLER_169_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4949_ _5067_/A _5023_/A VGND VGND VPWR VPWR _4949_/Y sky130_fd_sc_hd__nand2_1
XFILLER_184_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6619_ _6750_/CLK _6619_/D fanout446/X VGND VGND VPWR VPWR _6619_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_193_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput280 _6797_/Q VGND VGND VPWR VPWR pll_trim[18] sky130_fd_sc_hd__buf_12
Xoutput291 _6483_/Q VGND VGND VPWR VPWR pll_trim[4] sky130_fd_sc_hd__buf_12
XFILLER_181_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3280_ _3429_/A hold66/X VGND VGND VPWR VPWR _3309_/A sky130_fd_sc_hd__nor2_8
XFILLER_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6970_ _7116_/CLK _6970_/D fanout457/X VGND VGND VPWR VPWR _6970_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5921_ _6537_/Q _5651_/X _5688_/X _6581_/Q _5920_/X VGND VGND VPWR VPWR _5921_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_81_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5852_ _7060_/Q _5668_/X _5684_/X _6932_/Q VGND VGND VPWR VPWR _5852_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4803_ _5108_/B _5138_/C _4803_/C _4803_/D VGND VGND VPWR VPWR _4805_/B sky130_fd_sc_hd__and4_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5783_ _7009_/Q _5686_/X _5688_/X _6889_/Q VGND VGND VPWR VPWR _5783_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4734_ _5011_/A _4664_/Y _4584_/Y VGND VGND VPWR VPWR _4734_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4665_ _4738_/B _5026_/C VGND VGND VPWR VPWR _4730_/B sky130_fd_sc_hd__and2_1
XFILLER_175_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6404_ _6414_/A _6433_/B VGND VGND VPWR VPWR _6404_/X sky130_fd_sc_hd__and2_1
X_3616_ _3573_/X _3616_/B _3616_/C _3616_/D VGND VGND VPWR VPWR _3616_/Y sky130_fd_sc_hd__nand4b_4
XFILLER_128_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold900 hold900/A VGND VGND VPWR VPWR hold78/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold911 _3285_/B VGND VGND VPWR VPWR _3305_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold922 hold80/X VGND VGND VPWR VPWR hold922/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4596_ _4596_/A _4934_/B VGND VGND VPWR VPWR _4880_/B sky130_fd_sc_hd__nand2_1
Xhold933 hold933/A VGND VGND VPWR VPWR hold933/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_6335_ _6756_/Q _5638_/X _6015_/X _6761_/Q VGND VGND VPWR VPWR _6335_/X sky130_fd_sc_hd__a22o_1
Xhold944 hold944/A VGND VGND VPWR VPWR hold944/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_89_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold955 hold29/X VGND VGND VPWR VPWR hold955/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_3547_ _3940_/A1 _5236_/C _3431_/Y _7232_/A VGND VGND VPWR VPWR _3547_/X sky130_fd_sc_hd__a22o_2
Xhold966 _5575_/X VGND VGND VPWR VPWR _7130_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_89_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold977 _5586_/X VGND VGND VPWR VPWR hold34/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold988 _6874_/Q VGND VGND VPWR VPWR hold988/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_3478_ _6857_/Q _5263_/A _4310_/A _6741_/Q VGND VGND VPWR VPWR _3478_/X sky130_fd_sc_hd__a22o_1
Xhold999 _7002_/Q VGND VGND VPWR VPWR hold999/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_6266_ _7181_/Q _6265_/X _6341_/S VGND VGND VPWR VPWR _6266_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2301 hold575/X VGND VGND VPWR VPWR _4127_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2312 _6481_/Q VGND VGND VPWR VPWR hold579/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5217_ hold143/X hold135/X _5217_/S VGND VGND VPWR VPWR _5217_/X sky130_fd_sc_hd__mux2_1
Xhold2323 _6640_/Q VGND VGND VPWR VPWR hold736/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2334 _4036_/X VGND VGND VPWR VPWR hold406/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6197_ _7132_/Q _5973_/X _5998_/X _6892_/Q _6196_/X VGND VGND VPWR VPWR _6204_/A
+ sky130_fd_sc_hd__a221o_1
Xhold1600 _5266_/X VGND VGND VPWR VPWR hold145/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2345 _5417_/X VGND VGND VPWR VPWR _6989_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1611 _6581_/Q VGND VGND VPWR VPWR hold562/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2356 _6893_/Q VGND VGND VPWR VPWR hold793/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1622 hold127/X VGND VGND VPWR VPWR _4244_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2367 _7095_/Q VGND VGND VPWR VPWR hold623/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1633 hold544/X VGND VGND VPWR VPWR _5577_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2378 hold800/X VGND VGND VPWR VPWR _4299_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5148_ _5148_/A _5148_/B _5148_/C VGND VGND VPWR VPWR _5149_/D sky130_fd_sc_hd__and3_1
Xhold1644 _6699_/Q VGND VGND VPWR VPWR hold584/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2389 hold742/X VGND VGND VPWR VPWR _4058_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1655 _6601_/Q VGND VGND VPWR VPWR hold241/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1666 hold359/X VGND VGND VPWR VPWR _4246_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1677 hold630/X VGND VGND VPWR VPWR _4183_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5079_ _4688_/B _4995_/B _5009_/Y _4688_/C VGND VGND VPWR VPWR _5080_/C sky130_fd_sc_hd__o22a_1
Xhold1688 hold485/X VGND VGND VPWR VPWR _4157_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1699 _6804_/Q VGND VGND VPWR VPWR hold699/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_71_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4450_ _4450_/A _4450_/B VGND VGND VPWR VPWR _4451_/B sky130_fd_sc_hd__nor2_1
Xhold207 hold207/A VGND VGND VPWR VPWR wb_dat_o[30] sky130_fd_sc_hd__buf_12
XFILLER_116_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold218 hold218/A VGND VGND VPWR VPWR wb_dat_o[22] sky130_fd_sc_hd__buf_12
XFILLER_144_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold229 hold229/A VGND VGND VPWR VPWR hold229/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3401_ _6907_/Q _5317_/A _5488_/A _7059_/Q _3400_/X VGND VGND VPWR VPWR _3401_/X
+ sky130_fd_sc_hd__a221o_1
X_4381_ _4701_/A _4917_/A VGND VGND VPWR VPWR _4713_/A sky130_fd_sc_hd__and2b_4
XFILLER_125_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3332_ _3333_/A _3764_/A VGND VGND VPWR VPWR _5299_/A sky130_fd_sc_hd__nor2_8
X_6120_ _6977_/Q _5976_/B _6008_/X _7105_/Q _6119_/X VGND VGND VPWR VPWR _6120_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_171_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ _3262_/X _3263_/A1 _3996_/S VGND VGND VPWR VPWR _3263_/X sky130_fd_sc_hd__mux2_1
X_6051_ _7022_/Q _5971_/X _5987_/X _7110_/Q _6050_/X VGND VGND VPWR VPWR _6054_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _5114_/B _5002_/B _5124_/C VGND VGND VPWR VPWR _5002_/Y sky130_fd_sc_hd__nand3_1
X_3194_ _7155_/Q VGND VGND VPWR VPWR _5637_/A sky130_fd_sc_hd__clkinv_4
XFILLER_94_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6953_ _7105_/CLK _6953_/D fanout473/X VGND VGND VPWR VPWR _6953_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5904_ _5904_/A1 _6342_/S _5902_/X _5903_/X VGND VGND VPWR VPWR _7169_/D sky130_fd_sc_hd__o22a_1
XFILLER_50_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6884_ _7130_/CLK _6884_/D fanout458/X VGND VGND VPWR VPWR _6884_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5835_ _5835_/A _5835_/B _5835_/C _5835_/D VGND VGND VPWR VPWR _5835_/Y sky130_fd_sc_hd__nor4_2
XFILLER_179_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5766_ _6848_/Q _5842_/A2 _5656_/X _6984_/Q VGND VGND VPWR VPWR _5766_/X sky130_fd_sc_hd__a22o_1
X_4717_ _4717_/A _4717_/B _4732_/B VGND VGND VPWR VPWR _4727_/A sky130_fd_sc_hd__and3_2
XFILLER_175_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5697_ _6925_/Q _5684_/X _5694_/X _5696_/X VGND VGND VPWR VPWR _5697_/X sky130_fd_sc_hd__a211o_1
XFILLER_108_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4648_ _4682_/A _4712_/B VGND VGND VPWR VPWR _4648_/Y sky130_fd_sc_hd__nand2_2
XFILLER_135_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold730 hold730/A VGND VGND VPWR VPWR hold730/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold741 hold741/A VGND VGND VPWR VPWR hold741/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_146_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4579_ _4751_/B _4579_/B _4693_/B VGND VGND VPWR VPWR _4889_/B sky130_fd_sc_hd__nand3_2
Xhold752 hold752/A VGND VGND VPWR VPWR hold752/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold763 hold763/A VGND VGND VPWR VPWR hold763/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6318_ _6593_/Q _5985_/X _5994_/X _6638_/Q VGND VGND VPWR VPWR _6318_/X sky130_fd_sc_hd__a22o_1
Xhold774 hold774/A VGND VGND VPWR VPWR hold774/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold785 hold785/A VGND VGND VPWR VPWR hold785/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold796 hold796/A VGND VGND VPWR VPWR hold796/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6249_ _6590_/Q _5985_/X _5994_/X _6635_/Q _6243_/X VGND VGND VPWR VPWR _6249_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_77_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2120 hold740/X VGND VGND VPWR VPWR _5520_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2131 hold648/X VGND VGND VPWR VPWR _4308_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2142 hold719/X VGND VGND VPWR VPWR _5493_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2153 _4023_/X VGND VGND VPWR VPWR _6497_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2164 hold763/X VGND VGND VPWR VPWR _5358_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1430 hold332/X VGND VGND VPWR VPWR _4138_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2175 _6913_/Q VGND VGND VPWR VPWR hold762/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1441 _7060_/Q VGND VGND VPWR VPWR hold414/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2186 hold568/X VGND VGND VPWR VPWR _4324_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2197 _4325_/X VGND VGND VPWR VPWR _6749_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1452 _4214_/X VGND VGND VPWR VPWR hold150/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1463 _6756_/Q VGND VGND VPWR VPWR _4333_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1474 hold547/X VGND VGND VPWR VPWR _4079_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_61_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7053_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1485 _6900_/Q VGND VGND VPWR VPWR hold478/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1496 _4117_/X VGND VGND VPWR VPWR hold317/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_76_csclk _6727_/CLK VGND VGND VPWR VPWR _6808_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_14_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7134_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_122_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_csclk _6850_/CLK VGND VGND VPWR VPWR _7080_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold90 hold90/A VGND VGND VPWR VPWR hold90/X sky130_fd_sc_hd__clkdlybuf4s25_2
XFILLER_91_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3950_ _6507_/Q _3950_/A1 _6818_/Q VGND VGND VPWR VPWR _3950_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3881_ _6817_/Q _6864_/Q _3881_/C VGND VGND VPWR VPWR _3881_/Y sky130_fd_sc_hd__nor3_4
XFILLER_149_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5620_ _5619_/Y _5686_/A _5620_/S VGND VGND VPWR VPWR _5621_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5551_ _5551_/A _5551_/B VGND VGND VPWR VPWR _5559_/S sky130_fd_sc_hd__and2_4
XFILLER_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4502_ _4498_/X _4499_/Y _4500_/Y _4501_/X VGND VGND VPWR VPWR _4917_/B sky130_fd_sc_hd__a2bb2oi_2
XFILLER_8_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5482_ _5482_/A0 hold2/X _5487_/S VGND VGND VPWR VPWR _5482_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7221_ _7221_/A VGND VGND VPWR VPWR _7221_/X sky130_fd_sc_hd__clkbuf_2
X_4433_ _4663_/D _4451_/A VGND VGND VPWR VPWR _4486_/A sky130_fd_sc_hd__nor2_8
XFILLER_144_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7152_ _7152_/CLK _7152_/D _6399_/A VGND VGND VPWR VPWR _7152_/Q sky130_fd_sc_hd__dfstp_4
X_4364_ _4360_/A _4360_/B _4362_/B _4362_/A VGND VGND VPWR VPWR _4368_/A sky130_fd_sc_hd__a22o_4
XFILLER_116_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6103_ _6952_/Q _5997_/X _6004_/X _6880_/Q VGND VGND VPWR VPWR _6103_/X sky130_fd_sc_hd__a22o_1
X_3315_ _3354_/A _3686_/B VGND VGND VPWR VPWR _3315_/Y sky130_fd_sc_hd__nor2_8
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4295_ hold591/X _5187_/A1 _4297_/S VGND VGND VPWR VPWR _6724_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7083_ _7091_/CLK _7083_/D fanout481/X VGND VGND VPWR VPWR _7083_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_140_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6034_ _7117_/Q _5978_/X _5992_/X _6957_/Q _6033_/X VGND VGND VPWR VPWR _6039_/B
+ sky130_fd_sc_hd__a221o_1
X_3246_ _6470_/Q _6469_/Q _6468_/Q VGND VGND VPWR VPWR _3738_/S sky130_fd_sc_hd__nor3_4
XFILLER_100_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6936_ _7091_/CLK _6936_/D fanout471/X VGND VGND VPWR VPWR _6936_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6867_ _7140_/CLK _6867_/D fanout469/X VGND VGND VPWR VPWR _6867_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5818_ _7003_/Q _5666_/X _5674_/X _6875_/Q VGND VGND VPWR VPWR _5818_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6798_ _6809_/CLK _6798_/D fanout444/X VGND VGND VPWR VPWR _6798_/Q sky130_fd_sc_hd__dfstp_2
X_5749_ _6839_/Q _5678_/Y _5740_/X _5748_/X _6341_/S VGND VGND VPWR VPWR _5749_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold560 hold560/A VGND VGND VPWR VPWR hold560/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold571 hold571/A VGND VGND VPWR VPWR hold571/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold582 hold582/A VGND VGND VPWR VPWR hold582/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold593 hold593/A VGND VGND VPWR VPWR hold593/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_173_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1260 hold864/X VGND VGND VPWR VPWR hold206/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1271 _6866_/Q VGND VGND VPWR VPWR hold527/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1282 hold531/X VGND VGND VPWR VPWR _5449_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1293 hold129/X VGND VGND VPWR VPWR _4303_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__1153_ clkbuf_0__1153_/X VGND VGND VPWR VPWR _4112_/A0 sky130_fd_sc_hd__clkbuf_16
XFILLER_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4080_ hold444/X _5187_/A1 _4082_/S VGND VGND VPWR VPWR _4080_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4982_ _4569_/B _4570_/A _4570_/B _4570_/D _4968_/Y VGND VGND VPWR VPWR _4983_/C
+ sky130_fd_sc_hd__a41o_1
X_6721_ _6788_/CLK _6721_/D fanout439/X VGND VGND VPWR VPWR _6721_/Q sky130_fd_sc_hd__dfrtp_4
X_3933_ _3202_/Y input92/X _3934_/S VGND VGND VPWR VPWR _3933_/X sky130_fd_sc_hd__mux2_4
XFILLER_189_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_824 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6652_ _6711_/CLK _6652_/D _6432_/A VGND VGND VPWR VPWR _6652_/Q sky130_fd_sc_hd__dfrtp_4
X_3864_ _3904_/A _3863_/Y _3866_/A VGND VGND VPWR VPWR _3870_/B sky130_fd_sc_hd__a21oi_1
XFILLER_176_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5603_ _3193_/Y _5601_/B _5602_/Y VGND VGND VPWR VPWR _7145_/D sky130_fd_sc_hd__a21oi_1
XFILLER_164_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6583_ _6757_/CLK _6583_/D fanout447/X VGND VGND VPWR VPWR _6583_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_118_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3795_ input43/X _4047_/C _4241_/A input52/X VGND VGND VPWR VPWR _3795_/X sky130_fd_sc_hd__a22o_4
X_5534_ hold802/X _5561_/A1 _5541_/S VGND VGND VPWR VPWR _7093_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5465_ _5465_/A0 _5555_/A1 _5469_/S VGND VGND VPWR VPWR _7032_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7204_ _7204_/CLK _7204_/D fanout484/X VGND VGND VPWR VPWR _7204_/Q sky130_fd_sc_hd__dfrtp_1
X_4416_ _4719_/A _4595_/B VGND VGND VPWR VPWR _4417_/B sky130_fd_sc_hd__nand2_8
XFILLER_99_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5396_ _5396_/A0 _5576_/A1 _5397_/S VGND VGND VPWR VPWR _5396_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7135_ _7135_/CLK _7135_/D fanout474/X VGND VGND VPWR VPWR _7135_/Q sky130_fd_sc_hd__dfrtp_4
X_4347_ _4917_/A _4701_/A VGND VGND VPWR VPWR _4682_/A sky130_fd_sc_hd__and2_4
XFILLER_98_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7066_ _7116_/CLK _7066_/D fanout455/X VGND VGND VPWR VPWR _7066_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4278_ _4278_/A0 _5249_/A1 _4279_/S VGND VGND VPWR VPWR _4278_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6017_ _6017_/A _6017_/B _6019_/B VGND VGND VPWR VPWR _6017_/X sky130_fd_sc_hd__and3_4
XFILLER_100_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3229_ _6928_/Q VGND VGND VPWR VPWR _3229_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _3955_/A2 sky130_fd_sc_hd__clkbuf_16
XFILLER_54_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6919_ _7100_/CLK _6919_/D fanout458/X VGND VGND VPWR VPWR _6919_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold390 hold390/A VGND VGND VPWR VPWR hold390/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1090 _4248_/X VGND VGND VPWR VPWR _6674_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_46_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3580_ _3580_/A _3580_/B _3580_/C _3580_/D VGND VGND VPWR VPWR _3616_/B sky130_fd_sc_hd__nor4_4
XFILLER_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_748 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5250_ _5250_/A0 _5538_/A1 _5253_/S VGND VGND VPWR VPWR _6841_/D sky130_fd_sc_hd__mux2_1
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4201_ _4201_/A0 _5208_/A1 _4205_/S VGND VGND VPWR VPWR _6639_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5181_ hold588/X _5187_/A1 _5183_/S VGND VGND VPWR VPWR _6786_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4132_ _4132_/A0 _5195_/A1 _4133_/S VGND VGND VPWR VPWR _6582_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4063_ _4063_/A0 _5585_/A1 hold14/X VGND VGND VPWR VPWR _4063_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4965_ _4561_/X _4965_/B _4965_/C VGND VGND VPWR VPWR _5061_/A sky130_fd_sc_hd__and3b_1
X_6704_ _6817_/CLK _6704_/D fanout445/X VGND VGND VPWR VPWR _6704_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3916_ _6490_/Q _3909_/X _3912_/B _3915_/Y _3916_/B2 VGND VGND VPWR VPWR _3916_/X
+ sky130_fd_sc_hd__a32o_1
X_4896_ _5117_/A _4924_/A VGND VGND VPWR VPWR _4897_/B sky130_fd_sc_hd__nand2_2
X_6635_ _6750_/CLK _6635_/D fanout446/X VGND VGND VPWR VPWR _6635_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3847_ _6654_/Q _3847_/B VGND VGND VPWR VPWR _3852_/B sky130_fd_sc_hd__nand2_1
XFILLER_149_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6566_ _6568_/CLK _6566_/D VGND VGND VPWR VPWR _6566_/Q sky130_fd_sc_hd__dfxtp_1
X_3778_ _7061_/Q _5497_/A _3539_/Y _6530_/Q _3777_/X VGND VGND VPWR VPWR _3783_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5517_ hold694/X _5580_/A1 _5523_/S VGND VGND VPWR VPWR _7078_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6497_ _7016_/CLK _6497_/D fanout475/X VGND VGND VPWR VPWR _7218_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5448_ _5448_/A0 _5538_/A1 _5451_/S VGND VGND VPWR VPWR _5448_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5379_ _5379_/A0 hold6/X _5379_/S VGND VGND VPWR VPWR _5379_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7118_ _7126_/CLK _7118_/D fanout477/X VGND VGND VPWR VPWR _7118_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_87_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7049_ _7065_/CLK _7049_/D fanout460/X VGND VGND VPWR VPWR _7049_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_47_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4750_ _4637_/C _4719_/A _4683_/Y _4749_/X VGND VGND VPWR VPWR _4750_/X sky130_fd_sc_hd__a31o_1
XFILLER_33_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3701_ input44/X _3330_/Y _5263_/A _6854_/Q VGND VGND VPWR VPWR _3701_/X sky130_fd_sc_hd__a22o_1
X_4681_ _4682_/A _4717_/A VGND VGND VPWR VPWR _4722_/C sky130_fd_sc_hd__and2_2
XFILLER_146_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6420_ _6426_/A _6432_/B VGND VGND VPWR VPWR _6420_/X sky130_fd_sc_hd__and2_1
XFILLER_147_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3632_ _6863_/Q _5272_/A _3319_/Y _6797_/Q VGND VGND VPWR VPWR _3632_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6351_ _6351_/A0 hold871/A _6354_/S VGND VGND VPWR VPWR _7191_/D sky130_fd_sc_hd__mux2_1
X_3563_ _3563_/A _3563_/B VGND VGND VPWR VPWR _5202_/A sky130_fd_sc_hd__nor2_4
XFILLER_155_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5302_ _5302_/A0 _5518_/A1 _5307_/S VGND VGND VPWR VPWR _6887_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6282_ _6537_/Q _5983_/X _5986_/X _6641_/Q VGND VGND VPWR VPWR _6282_/X sky130_fd_sc_hd__a22o_1
X_3494_ input30/X _3307_/Y _4200_/A _6643_/Q _3493_/X VGND VGND VPWR VPWR _3499_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5233_ _5233_/A0 _5249_/A1 hold91/X VGND VGND VPWR VPWR _5233_/X sky130_fd_sc_hd__mux2_1
Xhold2505 _6437_/Q VGND VGND VPWR VPWR _3880_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2516 _3916_/X VGND VGND VPWR VPWR _6492_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2527 _6462_/Q VGND VGND VPWR VPWR _3840_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2538 _6605_/Q VGND VGND VPWR VPWR hold167/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5164_ _5011_/A _4691_/Y _4818_/A _5163_/X VGND VGND VPWR VPWR _5165_/C sky130_fd_sc_hd__o211a_1
Xhold1804 _5357_/X VGND VGND VPWR VPWR _6936_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1815 _4196_/X VGND VGND VPWR VPWR _6635_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1826 _5172_/X VGND VGND VPWR VPWR _6771_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_4115_ _3385_/Y hold850/A _4115_/S VGND VGND VPWR VPWR _6568_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1837 _6550_/Q VGND VGND VPWR VPWR hold295/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1848 hold484/X VGND VGND VPWR VPWR _5312_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5095_ _5095_/A _5095_/B VGND VGND VPWR VPWR _5095_/Y sky130_fd_sc_hd__nand2_1
Xhold1859 _5228_/X VGND VGND VPWR VPWR hold136/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4046_ hold338/X _4045_/X _4046_/S VGND VGND VPWR VPWR _4046_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5997_ _6019_/A _6017_/B _6007_/C VGND VGND VPWR VPWR _5997_/X sky130_fd_sc_hd__and3_4
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4948_ _4948_/A _5033_/B VGND VGND VPWR VPWR _5136_/B sky130_fd_sc_hd__nand2_1
XFILLER_177_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4879_ _4510_/A _4564_/Y _4569_/X _4570_/X _4878_/Y VGND VGND VPWR VPWR _4879_/X
+ sky130_fd_sc_hd__a41o_1
X_6618_ _6822_/CLK hold96/X fanout451/X VGND VGND VPWR VPWR _6618_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6549_ _6750_/CLK _6549_/D fanout446/X VGND VGND VPWR VPWR _6549_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput270 _6791_/Q VGND VGND VPWR VPWR pll_sel[2] sky130_fd_sc_hd__buf_12
XFILLER_133_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput281 _6798_/Q VGND VGND VPWR VPWR pll_trim[19] sky130_fd_sc_hd__buf_12
Xoutput292 _6484_/Q VGND VGND VPWR VPWR pll_trim[5] sky130_fd_sc_hd__buf_12
XFILLER_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5920_ _6596_/Q _5670_/X _5685_/X _6771_/Q VGND VGND VPWR VPWR _5920_/X sky130_fd_sc_hd__a22o_1
XFILLER_19_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5851_ _6964_/Q _5680_/X _5681_/X _7092_/Q VGND VGND VPWR VPWR _5851_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4802_ _5090_/C _4802_/B _4802_/C VGND VGND VPWR VPWR _4803_/D sky130_fd_sc_hd__and3_1
X_5782_ _5782_/A _5782_/B _5782_/C VGND VGND VPWR VPWR _5782_/Y sky130_fd_sc_hd__nor3_1
X_4733_ _4808_/A _4607_/B _4727_/A VGND VGND VPWR VPWR _4733_/X sky130_fd_sc_hd__a21o_1
XFILLER_175_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4664_ _5026_/C VGND VGND VPWR VPWR _4664_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6403_ _6432_/A _6433_/B VGND VGND VPWR VPWR _6403_/X sky130_fd_sc_hd__and2_1
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3615_ _3615_/A _3615_/B _3615_/C VGND VGND VPWR VPWR _3616_/D sky130_fd_sc_hd__and3_1
XFILLER_116_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold901 _5198_/X VGND VGND VPWR VPWR _6801_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_4595_ _4638_/A _4595_/B VGND VGND VPWR VPWR _4633_/B sky130_fd_sc_hd__nand2_8
Xhold912 _3308_/X VGND VGND VPWR VPWR _3430_/B sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_116_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold923 _5368_/X VGND VGND VPWR VPWR hold81/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold934 _4025_/X VGND VGND VPWR VPWR _6498_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_6334_ _6588_/Q _5989_/X _6013_/X _6628_/Q _6333_/X VGND VGND VPWR VPWR _6338_/B
+ sky130_fd_sc_hd__a221o_1
X_3546_ _6873_/Q _5281_/A _3347_/Y _7009_/Q _3545_/X VGND VGND VPWR VPWR _3556_/A
+ sky130_fd_sc_hd__a221o_1
Xhold945 _4042_/X VGND VGND VPWR VPWR _6506_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold956 _3271_/X VGND VGND VPWR VPWR hold30/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_115_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold967 _7202_/Q VGND VGND VPWR VPWR hold967/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold978 _6962_/Q VGND VGND VPWR VPWR hold978/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_89_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold989 hold989/A VGND VGND VPWR VPWR hold989/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_6265_ _6526_/Q _6339_/B _6264_/X VGND VGND VPWR VPWR _6265_/X sky130_fd_sc_hd__o21ba_1
X_3477_ _3535_/A _3549_/B VGND VGND VPWR VPWR _4310_/A sky130_fd_sc_hd__nor2_4
Xhold2302 _4127_/X VGND VGND VPWR VPWR _6578_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5216_ hold115/X hold78/X _5217_/S VGND VGND VPWR VPWR _5216_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2313 _6871_/Q VGND VGND VPWR VPWR hold582/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2324 hold736/X VGND VGND VPWR VPWR _4202_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6196_ _6884_/Q _6004_/X _6008_/X _7108_/Q VGND VGND VPWR VPWR _6196_/X sky130_fd_sc_hd__a22o_1
Xhold2335 hold406/X VGND VGND VPWR VPWR _6503_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2346 _6997_/Q VGND VGND VPWR VPWR hold797/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1601 _6754_/Q VGND VGND VPWR VPWR hold270/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1612 hold562/X VGND VGND VPWR VPWR _4131_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2357 _5309_/X VGND VGND VPWR VPWR _6893_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1623 _6584_/Q VGND VGND VPWR VPWR hold673/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5147_ _5147_/A1 _4836_/A _5134_/Y _5135_/X _5128_/Y VGND VGND VPWR VPWR _5147_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2368 hold623/X VGND VGND VPWR VPWR _5536_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1634 _5577_/X VGND VGND VPWR VPWR _7132_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2379 _7121_/Q VGND VGND VPWR VPWR hold718/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1645 _6602_/Q VGND VGND VPWR VPWR hold622/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1656 _4155_/X VGND VGND VPWR VPWR _6601_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1667 _6599_/Q VGND VGND VPWR VPWR hold629/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1678 _4183_/X VGND VGND VPWR VPWR _6624_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5078_ hold65/A _4836_/A _5025_/X _5077_/X VGND VGND VPWR VPWR _6765_/D sky130_fd_sc_hd__a211o_1
XFILLER_38_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1689 _4157_/X VGND VGND VPWR VPWR _6603_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_4029_ _4029_/A0 _4028_/X _4029_/S VGND VGND VPWR VPWR _4029_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold208 hold208/A VGND VGND VPWR VPWR hold208/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold219 hold219/A VGND VGND VPWR VPWR hold219/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3400_ input50/X _4047_/C hold27/A _6843_/Q VGND VGND VPWR VPWR _3400_/X sky130_fd_sc_hd__a22o_1
XFILLER_171_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4380_ _5009_/A _4811_/B VGND VGND VPWR VPWR _4921_/A sky130_fd_sc_hd__and2_1
XFILLER_125_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3331_ _3333_/A _3470_/A VGND VGND VPWR VPWR _5263_/A sky130_fd_sc_hd__nor2_8
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _7126_/Q _5973_/X _5988_/X _6870_/Q VGND VGND VPWR VPWR _6050_/X sky130_fd_sc_hd__a22o_1
XFILLER_140_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _6462_/Q _6461_/Q _6657_/Q VGND VGND VPWR VPWR _3262_/X sky130_fd_sc_hd__mux2_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5001_ _5001_/A _5001_/B VGND VGND VPWR VPWR _5124_/C sky130_fd_sc_hd__nand2_2
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3193_ _3193_/A VGND VGND VPWR VPWR _3193_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6952_ _7139_/CLK _6952_/D fanout478/X VGND VGND VPWR VPWR _6952_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5903_ _5903_/A1 _3924_/Y _5647_/Y VGND VGND VPWR VPWR _5903_/X sky130_fd_sc_hd__o21ba_1
XFILLER_50_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6883_ _7139_/CLK _6883_/D fanout478/X VGND VGND VPWR VPWR _6883_/Q sky130_fd_sc_hd__dfrtp_4
X_5834_ _6947_/Q _5658_/X _5673_/X _6867_/Q _5833_/X VGND VGND VPWR VPWR _5835_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5765_ _6976_/Q _5660_/X _5689_/X _7080_/Q _5764_/X VGND VGND VPWR VPWR _5770_/B
+ sky130_fd_sc_hd__a221o_1
X_4716_ _4384_/A _4658_/A _4638_/Y _4220_/B VGND VGND VPWR VPWR _4716_/Y sky130_fd_sc_hd__o31ai_4
X_5696_ _6869_/Q _5674_/X _5679_/X _6901_/Q _5695_/X VGND VGND VPWR VPWR _5696_/X
+ sky130_fd_sc_hd__a221o_1
X_4647_ _4682_/A _4712_/B VGND VGND VPWR VPWR _4735_/B sky130_fd_sc_hd__and2_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold720 hold720/A VGND VGND VPWR VPWR hold720/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold731 hold731/A VGND VGND VPWR VPWR hold731/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4578_ _4578_/A _4583_/B VGND VGND VPWR VPWR _4976_/A sky130_fd_sc_hd__nor2_4
Xhold742 hold742/A VGND VGND VPWR VPWR hold742/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold753 hold753/A VGND VGND VPWR VPWR hold753/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6317_ _6341_/A0 _6342_/S _6315_/X _6316_/X VGND VGND VPWR VPWR _7184_/D sky130_fd_sc_hd__o22a_1
Xhold764 hold764/A VGND VGND VPWR VPWR hold764/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3529_ _3529_/A _3529_/B _3529_/C _3529_/D VGND VGND VPWR VPWR _3557_/B sky130_fd_sc_hd__nor4_1
XFILLER_131_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold775 hold775/A VGND VGND VPWR VPWR hold775/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold786 hold786/A VGND VGND VPWR VPWR hold786/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold797 hold797/A VGND VGND VPWR VPWR hold797/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6248_ _6703_/Q _5977_/X _5984_/X _6615_/Q _6247_/X VGND VGND VPWR VPWR _6263_/B
+ sky130_fd_sc_hd__a221o_1
Xhold2110 _6791_/Q VGND VGND VPWR VPWR hold573/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2121 _7014_/Q VGND VGND VPWR VPWR hold761/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2132 _6512_/Q VGND VGND VPWR VPWR hold447/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_131_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2143 _5493_/X VGND VGND VPWR VPWR _7057_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2154 _6472_/Q VGND VGND VPWR VPWR hold525/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6179_ _6179_/A _6179_/B _6179_/C _6179_/D VGND VGND VPWR VPWR _6189_/B sky130_fd_sc_hd__nor4_2
Xhold1420 _6515_/Q VGND VGND VPWR VPWR hold383/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2165 _6574_/Q VGND VGND VPWR VPWR hold790/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1431 _4138_/X VGND VGND VPWR VPWR _6587_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2176 hold762/X VGND VGND VPWR VPWR _5331_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1442 hold414/X VGND VGND VPWR VPWR _5496_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2187 _4324_/X VGND VGND VPWR VPWR _6748_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1453 _6979_/Q VGND VGND VPWR VPWR hold374/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2198 _6999_/Q VGND VGND VPWR VPWR hold511/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1464 _4333_/X VGND VGND VPWR VPWR hold113/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1475 _4079_/X VGND VGND VPWR VPWR hold548/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1486 hold478/X VGND VGND VPWR VPWR _5316_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1497 _6710_/Q VGND VGND VPWR VPWR hold165/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold80 hold80/A VGND VGND VPWR VPWR hold80/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold91 hold91/A VGND VGND VPWR VPWR hold91/X sky130_fd_sc_hd__clkbuf_8
XFILLER_35_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3880_ _3880_/A0 _3879_/X _3880_/S VGND VGND VPWR VPWR _6437_/D sky130_fd_sc_hd__mux2_1
XFILLER_188_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5550_ _5550_/A0 _5577_/A1 _5550_/S VGND VGND VPWR VPWR _7108_/D sky130_fd_sc_hd__mux2_1
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4501_ _4637_/B _4498_/B _4663_/D VGND VGND VPWR VPWR _4501_/X sky130_fd_sc_hd__a21o_1
X_5481_ hold502/X _5499_/A1 _5487_/S VGND VGND VPWR VPWR _7046_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7220_ _7220_/A VGND VGND VPWR VPWR _7220_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4432_ _4447_/B _4457_/A VGND VGND VPWR VPWR _4451_/A sky130_fd_sc_hd__xor2_4
XFILLER_6_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7151_ _7152_/CLK _7151_/D _6399_/A VGND VGND VPWR VPWR _7151_/Q sky130_fd_sc_hd__dfstp_4
X_4363_ _4465_/B _4363_/B VGND VGND VPWR VPWR _4955_/B sky130_fd_sc_hd__and2_1
XFILLER_98_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6102_ _6102_/A _6102_/B _6102_/C VGND VGND VPWR VPWR _6114_/C sky130_fd_sc_hd__nor3_1
X_3314_ _3343_/A _3535_/A VGND VGND VPWR VPWR _5524_/A sky130_fd_sc_hd__nor2_8
X_7082_ _7124_/CLK _7082_/D fanout460/X VGND VGND VPWR VPWR _7082_/Q sky130_fd_sc_hd__dfrtp_4
X_4294_ _4294_/A0 _5186_/A1 _4297_/S VGND VGND VPWR VPWR _6723_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6033_ _7029_/Q _5986_/X _5996_/X _7045_/Q VGND VGND VPWR VPWR _6033_/X sky130_fd_sc_hd__a22o_1
XFILLER_101_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3245_ _4917_/A VGND VGND VPWR VPWR _4506_/A sky130_fd_sc_hd__clkinv_4
XFILLER_140_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6935_ _7035_/CLK _6935_/D fanout456/X VGND VGND VPWR VPWR _6935_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_25_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6866_ _7084_/CLK _6866_/D fanout455/X VGND VGND VPWR VPWR _6866_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_148_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5817_ _5817_/A1 _6342_/S _5815_/X _5816_/X VGND VGND VPWR VPWR _7165_/D sky130_fd_sc_hd__o22a_1
X_6797_ _6822_/CLK _6797_/D fanout451/X VGND VGND VPWR VPWR _6797_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_167_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5748_ _6887_/Q _5688_/X _5741_/X _5744_/X _5747_/X VGND VGND VPWR VPWR _5748_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_176_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5679_ _5689_/A _5679_/B _5687_/C VGND VGND VPWR VPWR _5679_/X sky130_fd_sc_hd__and3b_4
XFILLER_191_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold550 hold550/A VGND VGND VPWR VPWR hold550/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold561 hold561/A VGND VGND VPWR VPWR hold561/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold572 hold572/A VGND VGND VPWR VPWR hold572/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold583 hold583/A VGND VGND VPWR VPWR hold583/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold594 _5363_/X VGND VGND VPWR VPWR _6941_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1250 _6529_/Q VGND VGND VPWR VPWR hold122/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_18_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1261 hold206/X VGND VGND VPWR VPWR hold1261/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1272 hold527/X VGND VGND VPWR VPWR _5278_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1283 _7194_/Q VGND VGND VPWR VPWR hold866/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1294 _4303_/X VGND VGND VPWR VPWR _6731_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_727 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput170 wb_we_i VGND VGND VPWR VPWR _6358_/A sky130_fd_sc_hd__buf_2
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4981_ _4981_/A _4981_/B VGND VGND VPWR VPWR _5063_/D sky130_fd_sc_hd__nand2_1
XFILLER_51_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3932_ _6827_/Q input89/X _3934_/S VGND VGND VPWR VPWR _3932_/X sky130_fd_sc_hd__mux2_8
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6720_ _6750_/CLK _6720_/D fanout447/X VGND VGND VPWR VPWR _6720_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_16_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6651_ _6760_/CLK _6651_/D _6433_/A VGND VGND VPWR VPWR _6651_/Q sky130_fd_sc_hd__dfstp_2
X_3863_ _3863_/A _3878_/S VGND VGND VPWR VPWR _3863_/Y sky130_fd_sc_hd__nor2_1
XFILLER_176_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5602_ _3193_/Y _5601_/B _5601_/A VGND VGND VPWR VPWR _5602_/Y sky130_fd_sc_hd__o21ai_1
X_6582_ _6691_/CLK _6582_/D fanout450/X VGND VGND VPWR VPWR _6582_/Q sky130_fd_sc_hd__dfrtp_4
X_3794_ _7069_/Q _5506_/A _4256_/A _6692_/Q _3793_/X VGND VGND VPWR VPWR _3801_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5533_ _5533_/A _5569_/B VGND VGND VPWR VPWR _5541_/S sky130_fd_sc_hd__and2_4
XFILLER_157_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5464_ _5464_/A0 _5518_/A1 _5469_/S VGND VGND VPWR VPWR _7031_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_60_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7109_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_117_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7203_ _7203_/CLK _7203_/D _6346_/B VGND VGND VPWR VPWR _7203_/Q sky130_fd_sc_hd__dfrtp_2
X_4415_ _4594_/A _4415_/B VGND VGND VPWR VPWR _5026_/B sky130_fd_sc_hd__nor2_4
XFILLER_172_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5395_ _5395_/A0 _5503_/A1 _5397_/S VGND VGND VPWR VPWR _5395_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7134_ _7134_/CLK _7134_/D fanout468/X VGND VGND VPWR VPWR _7134_/Q sky130_fd_sc_hd__dfstp_4
X_4346_ _4346_/A _4346_/B _4346_/C VGND VGND VPWR VPWR _4492_/B sky130_fd_sc_hd__and3_4
XFILLER_59_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_75_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6749_/CLK sky130_fd_sc_hd__clkbuf_16
X_7065_ _7065_/CLK _7065_/D fanout460/X VGND VGND VPWR VPWR _7065_/Q sky130_fd_sc_hd__dfrtp_4
X_4277_ hold301/X _5581_/A1 _4279_/S VGND VGND VPWR VPWR _6709_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6016_ _6017_/A _6019_/B _6016_/C VGND VGND VPWR VPWR _6016_/X sky130_fd_sc_hd__and3_4
X_3228_ _6936_/Q VGND VGND VPWR VPWR _3228_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6918_ _7137_/CLK _6918_/D fanout476/X VGND VGND VPWR VPWR _6918_/Q sky130_fd_sc_hd__dfstp_2
Xclkbuf_leaf_13_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7097_/CLK sky130_fd_sc_hd__clkbuf_16
X_6849_ _7121_/CLK _6849_/D fanout473/X VGND VGND VPWR VPWR _6849_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length369 _5653_/X VGND VGND VPWR VPWR _5842_/A2 sky130_fd_sc_hd__buf_8
Xclkbuf_leaf_28_csclk _6850_/CLK VGND VGND VPWR VPWR _7138_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_164_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold380 hold380/A VGND VGND VPWR VPWR hold380/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold391 hold391/A VGND VGND VPWR VPWR hold391/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1080 hold435/X VGND VGND VPWR VPWR _5395_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_46_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1091 _7131_/Q VGND VGND VPWR VPWR hold378/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_788 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4200_ _4200_/A _5220_/C VGND VGND VPWR VPWR _4205_/S sky130_fd_sc_hd__and2_2
X_5180_ _5180_/A0 _5186_/A1 _5183_/S VGND VGND VPWR VPWR _6785_/D sky130_fd_sc_hd__mux2_1
XFILLER_123_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4131_ _4131_/A0 _5187_/A1 _4133_/S VGND VGND VPWR VPWR _4131_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4062_ hold941/X hold20/X hold14/X VGND VGND VPWR VPWR _4062_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4964_ _4963_/X _5044_/C VGND VGND VPWR VPWR _4964_/X sky130_fd_sc_hd__and2b_1
XFILLER_52_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6703_ _6822_/CLK _6703_/D fanout453/X VGND VGND VPWR VPWR _6703_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_189_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3915_ _7142_/Q _7143_/Q _5645_/C VGND VGND VPWR VPWR _3915_/Y sky130_fd_sc_hd__nand3b_2
X_4895_ _5136_/A _4997_/A VGND VGND VPWR VPWR _4921_/B sky130_fd_sc_hd__nand2_1
XFILLER_32_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_780 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6634_ _6749_/CLK _6634_/D fanout439/X VGND VGND VPWR VPWR _6634_/Q sky130_fd_sc_hd__dfrtp_4
X_3846_ _3845_/X _3846_/A1 _3846_/S VGND VGND VPWR VPWR _6460_/D sky130_fd_sc_hd__mux2_1
XFILLER_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3777_ _6784_/Q _5178_/A _4200_/A _6639_/Q VGND VGND VPWR VPWR _3777_/X sky130_fd_sc_hd__a22o_1
X_6565_ _6568_/CLK _6565_/D VGND VGND VPWR VPWR _6565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5516_ hold637/X _5561_/A1 _5523_/S VGND VGND VPWR VPWR _7077_/D sky130_fd_sc_hd__mux2_1
X_6496_ _6523_/CLK _6496_/D fanout481/X VGND VGND VPWR VPWR _7217_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_161_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5447_ _5447_/A0 _5582_/A1 _5451_/S VGND VGND VPWR VPWR _7016_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5378_ _5378_/A0 _5585_/A1 _5379_/S VGND VGND VPWR VPWR _5378_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7117_ _7117_/CLK _7117_/D fanout457/X VGND VGND VPWR VPWR _7117_/Q sky130_fd_sc_hd__dfstp_1
X_4329_ _4329_/A0 _5221_/A1 _4333_/S VGND VGND VPWR VPWR _4329_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7048_ _7133_/CLK _7048_/D fanout470/X VGND VGND VPWR VPWR _7048_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_75_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3700_ _7126_/Q _5569_/A hold27/A _6838_/Q _3699_/X VGND VGND VPWR VPWR _3703_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_41_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4680_ _4590_/Y _4674_/Y _4679_/Y _4668_/Y _4678_/X VGND VGND VPWR VPWR _4703_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_187_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3631_ _6999_/Q _5425_/A _3311_/Y _7103_/Q _3630_/X VGND VGND VPWR VPWR _3636_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6350_ _3616_/Y hold854/A _6354_/S VGND VGND VPWR VPWR _7190_/D sky130_fd_sc_hd__mux2_1
X_3562_ _3764_/A _3648_/B VGND VGND VPWR VPWR _3562_/Y sky130_fd_sc_hd__nor2_4
X_5301_ hold481/X _5499_/A1 _5307_/S VGND VGND VPWR VPWR _6886_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6281_ _6724_/Q _5978_/X _5992_/X _6709_/Q _6280_/X VGND VGND VPWR VPWR _6281_/X
+ sky130_fd_sc_hd__a221o_1
X_3493_ _3974_/B _3293_/Y _4280_/A _6716_/Q VGND VGND VPWR VPWR _3493_/X sky130_fd_sc_hd__a22o_1
X_5232_ _5232_/A0 _5572_/A1 hold91/X VGND VGND VPWR VPWR _5232_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2506 _7158_/Q VGND VGND VPWR VPWR _5644_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2517 _7172_/Q VGND VGND VPWR VPWR _5970_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5163_ _4590_/Y _4691_/Y _4995_/B _4674_/Y VGND VGND VPWR VPWR _5163_/X sky130_fd_sc_hd__o22a_1
Xhold2528 _6491_/Q VGND VGND VPWR VPWR _5610_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2539 _7160_/Q VGND VGND VPWR VPWR _5729_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1805 _7209_/A VGND VGND VPWR VPWR hold353/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1816 _6621_/Q VGND VGND VPWR VPWR hold306/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4114_ _3422_/Y hold862/A _4115_/S VGND VGND VPWR VPWR _6567_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1827 _6928_/Q VGND VGND VPWR VPWR hold495/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5094_ _3187_/Y _5139_/A _5085_/X _5093_/X VGND VGND VPWR VPWR _5119_/A sky130_fd_sc_hd__o211a_1
XFILLER_56_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1838 hold295/X VGND VGND VPWR VPWR _4095_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1849 _5312_/X VGND VGND VPWR VPWR _6896_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_83_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4045_ _4045_/A0 hold6/X _4056_/C VGND VGND VPWR VPWR _4045_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5996_ _6019_/A _6019_/B _6016_/C VGND VGND VPWR VPWR _5996_/X sky130_fd_sc_hd__and3_4
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4947_ _4947_/A _4947_/B VGND VGND VPWR VPWR _5033_/B sky130_fd_sc_hd__nand2_2
XFILLER_178_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4878_ _4934_/B _5048_/A VGND VGND VPWR VPWR _4878_/Y sky130_fd_sc_hd__nor2_1
XFILLER_165_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6617_ _6810_/CLK _6617_/D fanout452/X VGND VGND VPWR VPWR _6617_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_193_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3829_ _3829_/A1 _3835_/S _3827_/Y _3828_/X VGND VGND VPWR VPWR _6466_/D sky130_fd_sc_hd__o22a_1
XFILLER_119_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6548_ _6747_/CLK _6548_/D fanout439/X VGND VGND VPWR VPWR _6548_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_145_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6479_ _6793_/CLK _6479_/D fanout442/X VGND VGND VPWR VPWR _6479_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_161_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput260 _6803_/Q VGND VGND VPWR VPWR pll_bypass sky130_fd_sc_hd__buf_12
XFILLER_0_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput271 _6479_/Q VGND VGND VPWR VPWR pll_trim[0] sky130_fd_sc_hd__buf_12
Xoutput282 _6480_/Q VGND VGND VPWR VPWR pll_trim[1] sky130_fd_sc_hd__buf_12
Xoutput293 _6485_/Q VGND VGND VPWR VPWR pll_trim[6] sky130_fd_sc_hd__buf_12
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5850_ _6948_/Q _5658_/X _5664_/X _7020_/Q VGND VGND VPWR VPWR _5850_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4801_ _5011_/A _4729_/A _4514_/B VGND VGND VPWR VPWR _4802_/C sky130_fd_sc_hd__a21o_1
XFILLER_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5781_ _6905_/Q _5679_/X _5778_/X _5780_/X VGND VGND VPWR VPWR _5782_/C sky130_fd_sc_hd__a211o_1
X_4732_ _4988_/A _4732_/B VGND VGND VPWR VPWR _4755_/C sky130_fd_sc_hd__nand2_1
XFILLER_30_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4663_ _4447_/B _4917_/A _4701_/A _4663_/D VGND VGND VPWR VPWR _5026_/C sky130_fd_sc_hd__and4bb_4
XFILLER_174_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3614_ _3614_/A _3614_/B _3614_/C _3614_/D VGND VGND VPWR VPWR _3615_/C sky130_fd_sc_hd__nor4_1
X_6402_ _6414_/A _6423_/B VGND VGND VPWR VPWR _6402_/X sky130_fd_sc_hd__and2_1
XFILLER_147_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4594_ _4594_/A _4990_/B VGND VGND VPWR VPWR _4826_/A sky130_fd_sc_hd__nor2_4
Xhold902 _6766_/Q VGND VGND VPWR VPWR hold51/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_190_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold913 _3355_/Y VGND VGND VPWR VPWR _3550_/B sky130_fd_sc_hd__buf_12
Xhold924 _6514_/Q VGND VGND VPWR VPWR hold47/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6333_ _6691_/Q _5980_/X _6017_/X _6773_/Q VGND VGND VPWR VPWR _6333_/X sky130_fd_sc_hd__a22o_1
X_3545_ _7121_/Q hold67/A _4134_/A _6588_/Q VGND VGND VPWR VPWR _3545_/X sky130_fd_sc_hd__a22o_1
XFILLER_190_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold935 _7035_/Q VGND VGND VPWR VPWR hold935/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold946 _7098_/Q VGND VGND VPWR VPWR hold82/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold957 hold30/X VGND VGND VPWR VPWR _3305_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold968 _3998_/X VGND VGND VPWR VPWR hold5/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6264_ _6258_/X _6339_/B _6264_/C _6264_/D VGND VGND VPWR VPWR _6264_/X sky130_fd_sc_hd__and4b_1
XFILLER_103_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold979 hold979/A VGND VGND VPWR VPWR hold979/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_3476_ _7025_/Q _5452_/A _4206_/A _6648_/Q _3474_/X VGND VGND VPWR VPWR _3481_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5215_ _5215_/A0 _5503_/A1 _5217_/S VGND VGND VPWR VPWR _6813_/D sky130_fd_sc_hd__mux2_1
Xhold2303 _7127_/Q VGND VGND VPWR VPWR hold552/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6195_ _6924_/Q _5995_/X _6018_/X _6972_/Q _6194_/X VGND VGND VPWR VPWR _6195_/X
+ sky130_fd_sc_hd__a221o_1
Xhold2314 hold582/X VGND VGND VPWR VPWR _5284_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2325 _6479_/Q VGND VGND VPWR VPWR hold796/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2336 _7125_/Q VGND VGND VPWR VPWR hold787/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2347 _5426_/X VGND VGND VPWR VPWR _6997_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1602 _4331_/X VGND VGND VPWR VPWR _6754_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5146_ _5143_/Y _5145_/Y _5140_/X VGND VGND VPWR VPWR _5146_/X sky130_fd_sc_hd__o21a_1
Xhold2358 _6958_/Q VGND VGND VPWR VPWR hold764/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1613 _4131_/X VGND VGND VPWR VPWR _6581_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2369 _7000_/Q VGND VGND VPWR VPWR hold755/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1624 hold673/X VGND VGND VPWR VPWR _4135_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1635 _6688_/Q VGND VGND VPWR VPWR hold725/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1646 hold622/X VGND VGND VPWR VPWR _4156_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1657 _6614_/Q VGND VGND VPWR VPWR hold626/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5077_ _5043_/Y _5086_/B _5060_/X _5076_/Y VGND VGND VPWR VPWR _5077_/X sky130_fd_sc_hd__a211o_1
Xhold1668 hold629/X VGND VGND VPWR VPWR _4153_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1679 _6600_/Q VGND VGND VPWR VPWR hold734/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4028_ hold973/X hold6/X _4047_/C VGND VGND VPWR VPWR _4028_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5979_ _7155_/Q _7156_/Q VGND VGND VPWR VPWR _6007_/C sky130_fd_sc_hd__nor2_8
XFILLER_178_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold209 hold209/A VGND VGND VPWR VPWR hold209/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3330_ _3431_/A _3648_/A VGND VGND VPWR VPWR _3330_/Y sky130_fd_sc_hd__nor2_4
XFILLER_98_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ hold52/X _3261_/B VGND VGND VPWR VPWR _3501_/A sky130_fd_sc_hd__nand2b_4
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _5000_/A _5000_/B VGND VGND VPWR VPWR _5002_/B sky130_fd_sc_hd__and2_1
XFILLER_39_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3192_ _6654_/Q VGND VGND VPWR VPWR _3903_/A sky130_fd_sc_hd__inv_4
XFILLER_39_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6951_ _7119_/CLK _6951_/D fanout472/X VGND VGND VPWR VPWR _6951_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5902_ _6526_/Q _5678_/Y _5894_/X _5901_/X _6341_/S VGND VGND VPWR VPWR _5902_/X
+ sky130_fd_sc_hd__o221a_1
X_6882_ _7140_/CLK hold55/X fanout469/X VGND VGND VPWR VPWR _6882_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5833_ _7019_/Q _5664_/X _5686_/X _7011_/Q VGND VGND VPWR VPWR _5833_/X sky130_fd_sc_hd__a22o_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5764_ _7000_/Q _5666_/X _5678_/B _5763_/Y VGND VGND VPWR VPWR _5764_/X sky130_fd_sc_hd__a22o_1
X_4715_ _4651_/X _4709_/X _4636_/X VGND VGND VPWR VPWR _4759_/C sky130_fd_sc_hd__a21o_1
XFILLER_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5695_ _6941_/Q _5658_/X _5669_/X _7045_/Q VGND VGND VPWR VPWR _5695_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4646_ _4917_/A _4712_/B VGND VGND VPWR VPWR _4718_/C sky130_fd_sc_hd__and2_1
XFILLER_190_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold710 hold710/A VGND VGND VPWR VPWR hold710/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold721 hold721/A VGND VGND VPWR VPWR hold721/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4577_ _4811_/B _4710_/A VGND VGND VPWR VPWR _4997_/A sky130_fd_sc_hd__nand2_2
Xhold732 hold732/A VGND VGND VPWR VPWR hold732/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold743 _4058_/X VGND VGND VPWR VPWR _6518_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6316_ _6316_/A1 _3924_/Y _5647_/Y VGND VGND VPWR VPWR _6316_/X sky130_fd_sc_hd__o21ba_1
Xhold754 hold754/A VGND VGND VPWR VPWR hold754/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3528_ _6977_/Q _5398_/A _5299_/A _6889_/Q _3527_/X VGND VGND VPWR VPWR _3529_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_104_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold765 hold765/A VGND VGND VPWR VPWR hold765/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold776 hold776/A VGND VGND VPWR VPWR hold776/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold787 hold787/A VGND VGND VPWR VPWR hold787/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold798 hold798/A VGND VGND VPWR VPWR hold798/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6247_ _6605_/Q _5982_/X _5987_/X _6728_/Q VGND VGND VPWR VPWR _6247_/X sky130_fd_sc_hd__a22o_1
X_3459_ _6946_/Q _5362_/A _5290_/A _6882_/Q _3432_/X VGND VGND VPWR VPWR _3460_/D
+ sky130_fd_sc_hd__a221o_1
Xhold2100 _6881_/Q VGND VGND VPWR VPWR hold721/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2111 hold573/X VGND VGND VPWR VPWR _5187_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2122 _7216_/A VGND VGND VPWR VPWR hold417/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2133 hold447/X VGND VGND VPWR VPWR _4051_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2144 _7056_/Q VGND VGND VPWR VPWR hold767/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6178_ _6947_/Q _6005_/X _6015_/X _7019_/Q _6177_/X VGND VGND VPWR VPWR _6179_/D
+ sky130_fd_sc_hd__a221o_1
Xhold1410 _4063_/X VGND VGND VPWR VPWR hold398/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2155 _6796_/Q VGND VGND VPWR VPWR hold529/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1421 hold383/X VGND VGND VPWR VPWR _4054_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2166 hold790/X VGND VGND VPWR VPWR _4123_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1432 _7036_/Q VGND VGND VPWR VPWR hold423/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2177 _6577_/Q VGND VGND VPWR VPWR hold662/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1443 _5496_/X VGND VGND VPWR VPWR _7060_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2188 _6751_/Q VGND VGND VPWR VPWR hold526/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5129_ _4569_/B _4968_/Y _4586_/Y _4550_/Y VGND VGND VPWR VPWR _5130_/C sky130_fd_sc_hd__o211a_1
Xhold1454 _7006_/Q VGND VGND VPWR VPWR hold141/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2199 hold511/X VGND VGND VPWR VPWR _5428_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1465 _7116_/Q VGND VGND VPWR VPWR hold424/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1476 _6712_/Q VGND VGND VPWR VPWR hold319/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1487 _5316_/X VGND VGND VPWR VPWR _6900_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1498 hold165/X VGND VGND VPWR VPWR _4278_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold70 hold70/A VGND VGND VPWR VPWR hold70/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold81 hold81/A VGND VGND VPWR VPWR hold81/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold92 hold92/A VGND VGND VPWR VPWR hold92/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_817 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4500_ _4637_/B _4500_/B VGND VGND VPWR VPWR _4500_/Y sky130_fd_sc_hd__nand2_4
X_5480_ hold788/X _5570_/A1 _5487_/S VGND VGND VPWR VPWR _7045_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4431_ _4447_/B _4682_/A _4808_/B VGND VGND VPWR VPWR _4498_/B sky130_fd_sc_hd__and3_1
XANTENNA_1 _6475_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4362_ _4362_/A _4362_/B VGND VGND VPWR VPWR _4363_/B sky130_fd_sc_hd__nand2_1
X_7150_ _7204_/CLK _7150_/D fanout468/X VGND VGND VPWR VPWR _7150_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_99_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3313_ hold52/X _3313_/B VGND VGND VPWR VPWR _3530_/B sky130_fd_sc_hd__nand2_8
XFILLER_98_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6101_ _7032_/Q _5986_/X _5998_/X _6888_/Q _6100_/X VGND VGND VPWR VPWR _6102_/C
+ sky130_fd_sc_hd__a221o_1
X_7081_ _7137_/CLK _7081_/D fanout476/X VGND VGND VPWR VPWR _7081_/Q sky130_fd_sc_hd__dfrtp_4
X_4293_ _4293_/A0 _5552_/A1 _4297_/S VGND VGND VPWR VPWR _6722_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6032_ _7125_/Q _5973_/X _5988_/X _6869_/Q _6031_/X VGND VGND VPWR VPWR _6032_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_98_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3244_ _4637_/D VGND VGND VPWR VPWR _4594_/A sky130_fd_sc_hd__inv_6
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6934_ _7127_/CLK _6934_/D fanout477/X VGND VGND VPWR VPWR _6934_/Q sky130_fd_sc_hd__dfstp_2
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6865_ _7013_/CLK _6865_/D fanout452/X VGND VGND VPWR VPWR _6865_/Q sky130_fd_sc_hd__dfrtp_4
X_5816_ _5816_/A1 _3924_/Y _5647_/Y VGND VGND VPWR VPWR _5816_/X sky130_fd_sc_hd__o21ba_1
XFILLER_179_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6796_ _6809_/CLK _6796_/D fanout444/X VGND VGND VPWR VPWR _6796_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_10_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5747_ _7087_/Q _5681_/X _5745_/X _5746_/X VGND VGND VPWR VPWR _5747_/X sky130_fd_sc_hd__a211o_1
XFILLER_148_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5678_ _5686_/A _5678_/B VGND VGND VPWR VPWR _5678_/Y sky130_fd_sc_hd__nand2b_4
XFILLER_175_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4629_ _4522_/B _4491_/Y _5102_/A _4602_/Y _4627_/X VGND VGND VPWR VPWR _4630_/D
+ sky130_fd_sc_hd__o2111a_1
Xhold540 hold540/A VGND VGND VPWR VPWR hold540/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold551 hold551/A VGND VGND VPWR VPWR hold551/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold562 hold562/A VGND VGND VPWR VPWR hold562/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold573 hold573/A VGND VGND VPWR VPWR hold573/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_173_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold584 hold584/A VGND VGND VPWR VPWR hold584/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold595 hold595/A VGND VGND VPWR VPWR hold595/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1240 hold38/X VGND VGND VPWR VPWR _3267_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1251 _7074_/Q VGND VGND VPWR VPWR hold506/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_58_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1262 _6730_/Q VGND VGND VPWR VPWR hold208/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1273 _5278_/X VGND VGND VPWR VPWR _6866_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1284 hold866/X VGND VGND VPWR VPWR hold213/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1295 _6564_/Q VGND VGND VPWR VPWR hold867/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput160 wb_dat_i[6] VGND VGND VPWR VPWR _6380_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4980_ _4980_/A _4981_/B VGND VGND VPWR VPWR _5100_/B sky130_fd_sc_hd__nand2_1
XFILLER_63_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3931_ _6828_/Q input91/X _3934_/S VGND VGND VPWR VPWR _3931_/X sky130_fd_sc_hd__mux2_8
XFILLER_177_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6650_ _6760_/CLK _6650_/D _6433_/A VGND VGND VPWR VPWR _6650_/Q sky130_fd_sc_hd__dfrtp_4
X_3862_ _3862_/A _6656_/Q _3903_/A VGND VGND VPWR VPWR _3878_/S sky130_fd_sc_hd__nand3_4
X_5601_ _5601_/A _5601_/B _5601_/C VGND VGND VPWR VPWR _7144_/D sky130_fd_sc_hd__and3_1
XFILLER_176_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6581_ _6747_/CLK _6581_/D fanout450/X VGND VGND VPWR VPWR _6581_/Q sky130_fd_sc_hd__dfstp_2
X_3793_ _7093_/Q _5533_/A _4134_/A _6584_/Q VGND VGND VPWR VPWR _3793_/X sky130_fd_sc_hd__a22o_1
XFILLER_191_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5532_ hold35/X hold6/X _5532_/S VGND VGND VPWR VPWR _5532_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_9_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _6816_/CLK sky130_fd_sc_hd__clkbuf_16
X_5463_ hold604/X _5499_/A1 _5469_/S VGND VGND VPWR VPWR _7030_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7202_ _7204_/CLK _7202_/D fanout484/X VGND VGND VPWR VPWR _7202_/Q sky130_fd_sc_hd__dfrtp_1
X_4414_ _4575_/C _4637_/D VGND VGND VPWR VPWR _4595_/B sky130_fd_sc_hd__and2b_4
XFILLER_172_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5394_ _5394_/A0 _5556_/A1 _5397_/S VGND VGND VPWR VPWR _6969_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7133_ _7133_/CLK _7133_/D fanout471/X VGND VGND VPWR VPWR _7133_/Q sky130_fd_sc_hd__dfstp_4
X_4345_ _4345_/A _4345_/B _4345_/C _4345_/D VGND VGND VPWR VPWR _4346_/C sky130_fd_sc_hd__and4_1
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4276_ _4276_/A0 _5544_/A1 _4279_/S VGND VGND VPWR VPWR _4276_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7064_ _7138_/CLK _7064_/D fanout477/X VGND VGND VPWR VPWR _7064_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3227_ _6944_/Q VGND VGND VPWR VPWR _3227_/Y sky130_fd_sc_hd__inv_2
X_6015_ _6019_/A _6015_/B _6019_/B VGND VGND VPWR VPWR _6015_/X sky130_fd_sc_hd__and3_4
XFILLER_86_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6917_ _7117_/CLK _6917_/D fanout456/X VGND VGND VPWR VPWR _6917_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_54_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6848_ _7008_/CLK _6848_/D fanout477/X VGND VGND VPWR VPWR _6848_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6779_ _6658_/CLK _6779_/D _6431_/X VGND VGND VPWR VPWR _6779_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_183_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold370 hold370/A VGND VGND VPWR VPWR hold370/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold381 hold999/X VGND VGND VPWR VPWR hold381/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold392 hold392/A VGND VGND VPWR VPWR hold392/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1070 hold404/X VGND VGND VPWR VPWR _5540_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1081 _5395_/X VGND VGND VPWR VPWR _6970_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1092 hold378/X VGND VGND VPWR VPWR _5576_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4130_ _4130_/A0 _5186_/A1 _4133_/S VGND VGND VPWR VPWR _6580_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4061_ _4061_/A0 _5556_/A1 hold14/X VGND VGND VPWR VPWR _4061_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4963_ _4963_/A _5148_/A _4963_/C VGND VGND VPWR VPWR _4963_/X sky130_fd_sc_hd__and3_1
X_6702_ _7013_/CLK _6702_/D fanout452/X VGND VGND VPWR VPWR _6702_/Q sky130_fd_sc_hd__dfrtp_4
X_3914_ _7144_/Q _7145_/Q VGND VGND VPWR VPWR _5645_/C sky130_fd_sc_hd__nor2_2
X_4894_ _4894_/A _4894_/B VGND VGND VPWR VPWR _4903_/B sky130_fd_sc_hd__and2_1
XFILLER_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6633_ _6742_/CLK _6633_/D fanout439/X VGND VGND VPWR VPWR _6633_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3845_ _3182_/Y wire1/X _6657_/Q VGND VGND VPWR VPWR _3845_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6564_ _6568_/CLK _6564_/D VGND VGND VPWR VPWR _6564_/Q sky130_fd_sc_hd__dfxtp_1
X_3776_ _6624_/Q _4182_/A _5175_/A _6782_/Q _3775_/X VGND VGND VPWR VPWR _3783_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5515_ _5515_/A _5551_/B VGND VGND VPWR VPWR _5523_/S sky130_fd_sc_hd__and2_4
XFILLER_145_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6495_ _6523_/CLK _6495_/D fanout480/X VGND VGND VPWR VPWR _7216_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_145_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5446_ _5446_/A0 _5581_/A1 _5451_/S VGND VGND VPWR VPWR _7015_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5377_ hold995/X _5503_/A1 _5379_/S VGND VGND VPWR VPWR _5377_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7116_ _7116_/CLK _7116_/D fanout454/X VGND VGND VPWR VPWR _7116_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4328_ _4328_/A hold13/A VGND VGND VPWR VPWR _4333_/S sky130_fd_sc_hd__and2_4
XFILLER_141_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7047_ _7047_/CLK hold75/X fanout459/X VGND VGND VPWR VPWR _7047_/Q sky130_fd_sc_hd__dfrtp_4
X_4259_ _4259_/A0 _4337_/A1 _4261_/S VGND VGND VPWR VPWR _4259_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_74_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6788_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_147_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3630_ _3303_/X _5184_/B _3427_/Y _6791_/Q _3389_/Y VGND VGND VPWR VPWR _3630_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_139_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3561_ _6928_/Q _5344_/A _5353_/A _6936_/Q VGND VGND VPWR VPWR _3561_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5300_ hold783/X _5570_/A1 _5307_/S VGND VGND VPWR VPWR _6885_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6280_ _6631_/Q _5971_/X _6017_/X _6771_/Q VGND VGND VPWR VPWR _6280_/X sky130_fd_sc_hd__a22o_1
X_3492_ _3563_/A _3531_/B VGND VGND VPWR VPWR _4280_/A sky130_fd_sc_hd__nor2_4
XFILLER_154_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5231_ _5231_/A0 _5544_/A1 hold91/X VGND VGND VPWR VPWR _5231_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2507 _7185_/Q VGND VGND VPWR VPWR _6342_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2518 _7143_/Q VGND VGND VPWR VPWR _5598_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5162_ _5162_/A _5162_/B _5162_/C VGND VGND VPWR VPWR _5162_/Y sky130_fd_sc_hd__nand3_1
Xhold2529 _5635_/Y VGND VGND VPWR VPWR _5636_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xclkbuf_leaf_12_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _6826_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_69_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1806 hold353/X VGND VGND VPWR VPWR _4234_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4113_ _3462_/Y hold860/A _4115_/S VGND VGND VPWR VPWR _6566_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1817 hold306/X VGND VGND VPWR VPWR _4179_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5093_ _5088_/X _5136_/C _5092_/X _5086_/Y VGND VGND VPWR VPWR _5093_/X sky130_fd_sc_hd__a31o_1
XFILLER_57_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1828 hold495/X VGND VGND VPWR VPWR _5348_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1839 _6501_/Q VGND VGND VPWR VPWR hold462/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4044_ _4044_/A0 _4043_/X _4046_/S VGND VGND VPWR VPWR _4044_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_27_csclk _6850_/CLK VGND VGND VPWR VPWR _7127_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_37_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5995_ _6019_/A _6007_/C _6016_/C VGND VGND VPWR VPWR _5995_/X sky130_fd_sc_hd__and3_4
XFILLER_52_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4946_ _4368_/B _4407_/Y _4935_/X _4800_/A VGND VGND VPWR VPWR _5041_/A sky130_fd_sc_hd__o31a_1
XFILLER_193_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4877_ _5127_/A _4965_/B _5044_/B _4876_/X _4636_/X VGND VGND VPWR VPWR _4906_/C
+ sky130_fd_sc_hd__a41o_1
XFILLER_137_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6616_ _6809_/CLK _6616_/D fanout444/X VGND VGND VPWR VPWR _6616_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_138_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3828_ _3832_/A _6657_/Q _3846_/S VGND VGND VPWR VPWR _3828_/X sky130_fd_sc_hd__a21o_1
XFILLER_137_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6547_ _7194_/CLK _6547_/D VGND VGND VPWR VPWR _6547_/Q sky130_fd_sc_hd__dfxtp_1
X_3759_ _3759_/A _3759_/B _3759_/C _3759_/D VGND VGND VPWR VPWR _3770_/B sky130_fd_sc_hd__nor4_1
X_6478_ _6822_/CLK _6478_/D fanout451/X VGND VGND VPWR VPWR _6478_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_118_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5429_ _5429_/A0 _5582_/A1 _5433_/S VGND VGND VPWR VPWR _5429_/X sky130_fd_sc_hd__mux2_1
Xoutput250 _3957_/Y VGND VGND VPWR VPWR pad_flash_csb_oeb sky130_fd_sc_hd__buf_12
Xoutput261 _6783_/Q VGND VGND VPWR VPWR pll_dco_ena sky130_fd_sc_hd__buf_12
Xoutput272 _6473_/Q VGND VGND VPWR VPWR pll_trim[10] sky130_fd_sc_hd__buf_12
Xoutput283 _6799_/Q VGND VGND VPWR VPWR pll_trim[20] sky130_fd_sc_hd__buf_12
XFILLER_160_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput294 _6486_/Q VGND VGND VPWR VPWR pll_trim[7] sky130_fd_sc_hd__buf_12
XFILLER_181_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire355 _6204_/Y VGND VGND VPWR VPWR _6214_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4800_ _4800_/A _4800_/B _4800_/C _4800_/D VGND VGND VPWR VPWR _4803_/C sky130_fd_sc_hd__and4_1
XFILLER_34_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5780_ _6985_/Q _5656_/X _5680_/X _6961_/Q _5779_/X VGND VGND VPWR VPWR _5780_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_159_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ _4731_/A _4993_/B VGND VGND VPWR VPWR _4753_/B sky130_fd_sc_hd__nand2_1
XFILLER_187_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4662_ _4738_/B _5150_/C VGND VGND VPWR VPWR _4662_/Y sky130_fd_sc_hd__nand2_2
XFILLER_119_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6401_ _6414_/A _6423_/B VGND VGND VPWR VPWR _6401_/X sky130_fd_sc_hd__and2_1
X_3613_ _7080_/Q _5515_/A _4334_/A _6760_/Q _3612_/X VGND VGND VPWR VPWR _3614_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_116_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4593_ _4637_/C _4638_/A VGND VGND VPWR VPWR _4990_/B sky130_fd_sc_hd__nand2b_4
XFILLER_128_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold903 hold51/X VGND VGND VPWR VPWR hold903/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold914 _3357_/Y VGND VGND VPWR VPWR _4000_/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6332_ _6726_/Q _5978_/X _5995_/X _6603_/Q _6331_/X VGND VGND VPWR VPWR _6338_/A
+ sky130_fd_sc_hd__a221o_1
Xhold925 hold47/X VGND VGND VPWR VPWR hold925/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_3544_ hold54/X _3648_/A VGND VGND VPWR VPWR _4134_/A sky130_fd_sc_hd__nor2_8
Xhold936 hold936/A VGND VGND VPWR VPWR hold936/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_116_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold947 hold82/X VGND VGND VPWR VPWR hold947/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold958 _3353_/A VGND VGND VPWR VPWR _3563_/B sky130_fd_sc_hd__clkdlybuf4s50_2
X_6263_ _6263_/A _6263_/B _6263_/C _6263_/D VGND VGND VPWR VPWR _6264_/D sky130_fd_sc_hd__nor4_2
XFILLER_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold969 hold5/X VGND VGND VPWR VPWR hold969/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_3475_ _3530_/B _3516_/B VGND VGND VPWR VPWR _4206_/A sky130_fd_sc_hd__nor2_8
XFILLER_103_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5214_ _5214_/A0 _5518_/A1 _5217_/S VGND VGND VPWR VPWR _6812_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6194_ _7060_/Q _5990_/X _5991_/X _6916_/Q _6193_/X VGND VGND VPWR VPWR _6194_/X
+ sky130_fd_sc_hd__a221o_1
Xhold2304 hold552/X VGND VGND VPWR VPWR _5572_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2315 _5284_/X VGND VGND VPWR VPWR _6871_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2326 _6927_/Q VGND VGND VPWR VPWR hold570/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2337 _5570_/X VGND VGND VPWR VPWR _7125_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2348 _7230_/A VGND VGND VPWR VPWR hold612/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1603 _6554_/Q VGND VGND VPWR VPWR hold834/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5145_ _4683_/A _5144_/X _5022_/A VGND VGND VPWR VPWR _5145_/Y sky130_fd_sc_hd__o21ai_2
Xhold1614 _6687_/Q VGND VGND VPWR VPWR hold608/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2359 _5382_/X VGND VGND VPWR VPWR _6958_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1625 _6524_/Q VGND VGND VPWR VPWR _4045_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1636 hold725/X VGND VGND VPWR VPWR _4252_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1647 _4156_/X VGND VGND VPWR VPWR _6602_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1658 hold626/X VGND VGND VPWR VPWR _4171_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5076_ _5066_/X _5074_/X _5062_/A VGND VGND VPWR VPWR _5076_/Y sky130_fd_sc_hd__a21oi_1
Xhold1669 _4153_/X VGND VGND VPWR VPWR _6599_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4027_ _4027_/A0 _4026_/X _4029_/S VGND VGND VPWR VPWR _4027_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5978_ _6008_/A _6014_/A _6019_/C VGND VGND VPWR VPWR _5978_/X sky130_fd_sc_hd__and3_4
X_4929_ _5126_/B _4929_/B _5112_/B VGND VGND VPWR VPWR _4930_/D sky130_fd_sc_hd__and3_1
XFILLER_178_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmgmt_gpio_9_buff_inst _3940_/X VGND VGND VPWR VPWR mgmt_gpio_out[9] sky130_fd_sc_hd__clkbuf_8
XFILLER_134_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _3302_/A hold88/X _3260_/C VGND VGND VPWR VPWR _3260_/X sky130_fd_sc_hd__and3_2
XFILLER_140_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3191_ _6685_/Q VGND VGND VPWR VPWR _3969_/A sky130_fd_sc_hd__inv_2
XFILLER_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6950_ _7126_/CLK _6950_/D fanout474/X VGND VGND VPWR VPWR _6950_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_47_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5901_ _6630_/Q _5663_/X _5895_/X _5896_/X _5900_/X VGND VGND VPWR VPWR _5901_/X
+ sky130_fd_sc_hd__a2111o_2
X_6881_ _7137_/CLK _6881_/D fanout473/X VGND VGND VPWR VPWR _6881_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5832_ _6939_/Q _5659_/X _5663_/X _7027_/Q _5831_/X VGND VGND VPWR VPWR _5835_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5763_ _5763_/A _5872_/B VGND VGND VPWR VPWR _5763_/Y sky130_fd_sc_hd__nand2_1
XFILLER_148_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4714_ _4717_/B _4714_/B _4751_/C VGND VGND VPWR VPWR _4714_/Y sky130_fd_sc_hd__nand3_4
XFILLER_187_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5694_ _6933_/Q _5659_/X _5693_/X VGND VGND VPWR VPWR _5694_/X sky130_fd_sc_hd__a21o_1
XFILLER_147_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4645_ _4447_/B _4663_/D VGND VGND VPWR VPWR _4712_/B sky130_fd_sc_hd__and2b_4
XFILLER_148_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold700 hold700/A VGND VGND VPWR VPWR hold700/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4576_ _4576_/A _4638_/A VGND VGND VPWR VPWR _4583_/B sky130_fd_sc_hd__nand2_8
Xhold711 hold711/A VGND VGND VPWR VPWR hold711/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap430 _4649_/Y VGND VGND VPWR VPWR _4672_/B sky130_fd_sc_hd__buf_2
Xhold722 hold722/A VGND VGND VPWR VPWR hold722/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold733 hold733/A VGND VGND VPWR VPWR hold733/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6315_ _6528_/Q _6339_/B _6314_/Y _6341_/S VGND VGND VPWR VPWR _6315_/X sky130_fd_sc_hd__o211a_1
Xhold744 hold744/A VGND VGND VPWR VPWR hold744/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3527_ input16/X _3310_/Y _4065_/A _6529_/Q VGND VGND VPWR VPWR _3527_/X sky130_fd_sc_hd__a22o_1
Xhold755 hold755/A VGND VGND VPWR VPWR hold755/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold766 hold766/A VGND VGND VPWR VPWR hold766/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold777 hold777/A VGND VGND VPWR VPWR hold777/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold788 hold788/A VGND VGND VPWR VPWR hold788/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold799 hold799/A VGND VGND VPWR VPWR hold799/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6246_ _6549_/Q _5999_/X _6019_/X _6733_/Q _6245_/X VGND VGND VPWR VPWR _6263_/A
+ sky130_fd_sc_hd__a221o_1
X_3458_ input40/X _4056_/C _5317_/A _6906_/Q _3457_/X VGND VGND VPWR VPWR _3460_/C
+ sky130_fd_sc_hd__a221o_1
Xhold2101 hold721/X VGND VGND VPWR VPWR _5295_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2112 _5187_/X VGND VGND VPWR VPWR _6791_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2123 hold417/X VGND VGND VPWR VPWR _4019_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6177_ _7083_/Q _6013_/X _6017_/X _7075_/Q VGND VGND VPWR VPWR _6177_/X sky130_fd_sc_hd__a22o_1
Xhold2134 _7134_/Q VGND VGND VPWR VPWR hold775/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_3389_ _3686_/B _3470_/A VGND VGND VPWR VPWR _3389_/Y sky130_fd_sc_hd__nor2_4
Xhold1400 hold413/X VGND VGND VPWR VPWR _5415_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2145 hold767/X VGND VGND VPWR VPWR _5492_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2156 _7217_/A VGND VGND VPWR VPWR hold655/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1411 _6695_/Q VGND VGND VPWR VPWR hold322/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1422 _4054_/X VGND VGND VPWR VPWR hold384/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2167 _4123_/X VGND VGND VPWR VPWR _6574_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1433 hold423/X VGND VGND VPWR VPWR _5469_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5128_ _5121_/X _5123_/X _5127_/X VGND VGND VPWR VPWR _5128_/Y sky130_fd_sc_hd__a21boi_1
Xhold2178 hold662/X VGND VGND VPWR VPWR _4126_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2189 hold526/X VGND VGND VPWR VPWR _4327_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1444 _6707_/Q VGND VGND VPWR VPWR hold296/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1455 _5436_/X VGND VGND VPWR VPWR _7006_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1466 hold424/X VGND VGND VPWR VPWR _5559_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_55_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1477 hold319/X VGND VGND VPWR VPWR _4281_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1488 _6981_/Q VGND VGND VPWR VPWR hold664/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5059_ _5123_/B _5059_/B _5059_/C VGND VGND VPWR VPWR _5059_/X sky130_fd_sc_hd__and3_1
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1499 _4278_/X VGND VGND VPWR VPWR hold166/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold60 hold60/A VGND VGND VPWR VPWR hold60/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold71 hold71/A VGND VGND VPWR VPWR hold71/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold82 hold82/A VGND VGND VPWR VPWR hold82/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold93 hold93/A VGND VGND VPWR VPWR hold93/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4430_ _4682_/A _4808_/B VGND VGND VPWR VPWR _4457_/A sky130_fd_sc_hd__nand2_4
XANTENNA_2 _3239_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4361_ _4447_/B _4682_/A _4365_/B _4663_/D VGND VGND VPWR VPWR _4362_/B sky130_fd_sc_hd__a31o_1
XFILLER_125_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6100_ _6976_/Q _5976_/B _5993_/X _7008_/Q VGND VGND VPWR VPWR _6100_/X sky130_fd_sc_hd__a22o_1
X_3312_ _3349_/A _3764_/A VGND VGND VPWR VPWR _5443_/A sky130_fd_sc_hd__nor2_8
X_7080_ _7080_/CLK _7080_/D fanout480/X VGND VGND VPWR VPWR _7080_/Q sky130_fd_sc_hd__dfrtp_4
X_4292_ _4292_/A _5220_/C VGND VGND VPWR VPWR _4297_/S sky130_fd_sc_hd__and2_2
XFILLER_140_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6031_ _7021_/Q _5971_/X _5994_/X _7061_/Q _6030_/X VGND VGND VPWR VPWR _6031_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_58_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3243_ _6972_/Q VGND VGND VPWR VPWR _3243_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6933_ _7125_/CLK _6933_/D fanout454/X VGND VGND VPWR VPWR _6933_/Q sky130_fd_sc_hd__dfstp_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6864_ _7020_/CLK _6864_/D fanout458/X VGND VGND VPWR VPWR _6864_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5815_ _6842_/Q _5678_/Y _5808_/X _5814_/X _6341_/S VGND VGND VPWR VPWR _5815_/X
+ sky130_fd_sc_hd__o221a_2
X_6795_ _6822_/CLK _6795_/D fanout451/X VGND VGND VPWR VPWR _6795_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_50_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5746_ _6863_/Q _5673_/X _5680_/X _6959_/Q VGND VGND VPWR VPWR _5746_/X sky130_fd_sc_hd__a22o_1
XFILLER_182_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5677_ _5872_/B _5677_/B VGND VGND VPWR VPWR _5707_/B sky130_fd_sc_hd__nor2_8
XFILLER_108_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4628_ _4628_/A _4917_/D VGND VGND VPWR VPWR _4628_/Y sky130_fd_sc_hd__nand2_1
Xhold530 hold530/A VGND VGND VPWR VPWR hold530/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4559_ _4598_/B _4598_/C VGND VGND VPWR VPWR _4601_/B sky130_fd_sc_hd__nand2_1
Xhold541 _4059_/X VGND VGND VPWR VPWR _6519_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold552 hold552/A VGND VGND VPWR VPWR hold552/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold563 hold563/A VGND VGND VPWR VPWR hold563/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold574 hold574/A VGND VGND VPWR VPWR hold574/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_173_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold585 hold585/A VGND VGND VPWR VPWR hold585/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_173_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold596 _3989_/X VGND VGND VPWR VPWR _6471_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6229_ _6639_/Q _5986_/X _5998_/X _6579_/Q _6228_/X VGND VGND VPWR VPWR _6230_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1230 hold503/X VGND VGND VPWR VPWR _5530_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1241 _3328_/X VGND VGND VPWR VPWR _5222_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_100_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1252 hold506/X VGND VGND VPWR VPWR _5512_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1263 hold208/X VGND VGND VPWR VPWR _4302_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1274 _7102_/Q VGND VGND VPWR VPWR hold284/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1285 hold213/X VGND VGND VPWR VPWR hold1285/X sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1296 hold867/X VGND VGND VPWR VPWR hold226/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput150 wb_dat_i[26] VGND VGND VPWR VPWR _6367_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput161 wb_dat_i[7] VGND VGND VPWR VPWR _6383_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3930_ _6656_/Q _3929_/Y _3739_/S VGND VGND VPWR VPWR _6436_/D sky130_fd_sc_hd__o21a_1
XFILLER_17_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3861_ _3879_/A _6468_/Q _3903_/A _3738_/S _3847_/B VGND VGND VPWR VPWR _3868_/B
+ sky130_fd_sc_hd__a2111oi_4
XFILLER_189_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5600_ _7142_/Q _7143_/Q _5599_/D _7144_/Q VGND VGND VPWR VPWR _5601_/C sky130_fd_sc_hd__a31o_1
X_6580_ _6808_/CLK _6580_/D fanout439/X VGND VGND VPWR VPWR _6580_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_82_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3792_ _3792_/A _3792_/B _3792_/C _3792_/D VGND VGND VPWR VPWR _3802_/C sky130_fd_sc_hd__nor4_1
XFILLER_158_851 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5531_ _5531_/A0 _5576_/A1 _5532_/S VGND VGND VPWR VPWR _5531_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5462_ hold795/X _5552_/A1 _5469_/S VGND VGND VPWR VPWR _7029_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7201_ _7204_/CLK _7201_/D fanout484/X VGND VGND VPWR VPWR _7201_/Q sky130_fd_sc_hd__dfrtp_1
X_4413_ _4804_/A VGND VGND VPWR VPWR _4415_/B sky130_fd_sc_hd__clkinv_2
XFILLER_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5393_ _5393_/A0 _5555_/A1 _5397_/S VGND VGND VPWR VPWR _6968_/D sky130_fd_sc_hd__mux2_1
X_7132_ _7132_/CLK _7132_/D fanout459/X VGND VGND VPWR VPWR _7132_/Q sky130_fd_sc_hd__dfrtp_4
X_4344_ _4344_/A _4344_/B _4344_/C _4344_/D VGND VGND VPWR VPWR _4346_/B sky130_fd_sc_hd__and4_1
X_7063_ _7077_/CLK _7063_/D fanout456/X VGND VGND VPWR VPWR _7063_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4275_ hold296/X hold153/X _4279_/S VGND VGND VPWR VPWR _4275_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6014_ _6014_/A _6019_/B _6019_/C VGND VGND VPWR VPWR _6014_/X sky130_fd_sc_hd__and3_4
X_3226_ _6952_/Q VGND VGND VPWR VPWR _3226_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6916_ _7084_/CLK _6916_/D fanout455/X VGND VGND VPWR VPWR _6916_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_70_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6847_ _7111_/CLK _6847_/D fanout472/X VGND VGND VPWR VPWR _6847_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6778_ _6658_/CLK _6778_/D _6430_/X VGND VGND VPWR VPWR _6778_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_139_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5729_ _5729_/A0 _5728_/X _6341_/S VGND VGND VPWR VPWR _5729_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold360 hold360/A VGND VGND VPWR VPWR hold360/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold371 hold371/A VGND VGND VPWR VPWR hold371/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold382 hold382/A VGND VGND VPWR VPWR hold382/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold393 hold994/X VGND VGND VPWR VPWR hold995/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1060 hold87/X VGND VGND VPWR VPWR _3255_/B sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1071 _6851_/Q VGND VGND VPWR VPWR hold390/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1082 _6995_/Q VGND VGND VPWR VPWR hold361/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1093 _5576_/X VGND VGND VPWR VPWR _7131_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_200 _5678_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4060_ _4060_/A0 _5582_/A1 hold14/X VGND VGND VPWR VPWR _4060_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4962_ _5162_/A _4962_/B _4962_/C VGND VGND VPWR VPWR _4963_/C sky130_fd_sc_hd__and3_1
XFILLER_51_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6701_ _6759_/CLK _6701_/D fanout447/X VGND VGND VPWR VPWR _6701_/Q sky130_fd_sc_hd__dfrtp_4
X_3913_ _6816_/Q _5611_/A _3912_/X _6490_/Q VGND VGND VPWR VPWR _6491_/D sky130_fd_sc_hd__a22o_1
XFILLER_32_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4893_ _4893_/A _4922_/A VGND VGND VPWR VPWR _5155_/A sky130_fd_sc_hd__and2_1
XFILLER_149_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6632_ _6742_/CLK _6632_/D fanout440/X VGND VGND VPWR VPWR _6632_/Q sky130_fd_sc_hd__dfrtp_4
X_3844_ _3846_/A1 _3843_/Y _3842_/X VGND VGND VPWR VPWR _3844_/X sky130_fd_sc_hd__a21o_1
XFILLER_192_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6563_ _6568_/CLK _6563_/D VGND VGND VPWR VPWR _6563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3775_ _6877_/Q _5290_/A _3648_/Y _6820_/Q VGND VGND VPWR VPWR _3775_/X sky130_fd_sc_hd__a22o_2
XFILLER_164_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5514_ _5514_/A0 _5577_/A1 _5514_/S VGND VGND VPWR VPWR _7076_/D sky130_fd_sc_hd__mux2_1
XFILLER_192_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6494_ _6523_/CLK _6494_/D fanout480/X VGND VGND VPWR VPWR _7215_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_173_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5445_ hold761/X _5580_/A1 _5451_/S VGND VGND VPWR VPWR _7014_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5376_ _5376_/A0 _5583_/A1 _5379_/S VGND VGND VPWR VPWR _6953_/D sky130_fd_sc_hd__mux2_1
XFILLER_154_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7115_ _7140_/CLK _7115_/D fanout470/X VGND VGND VPWR VPWR _7115_/Q sky130_fd_sc_hd__dfrtp_4
X_4327_ _4327_/A0 _4339_/A1 _4327_/S VGND VGND VPWR VPWR _4327_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7046_ _7131_/CLK _7046_/D fanout470/X VGND VGND VPWR VPWR _7046_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_47_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4258_ _4258_/A0 _5193_/A1 _4261_/S VGND VGND VPWR VPWR _4258_/X sky130_fd_sc_hd__mux2_1
X_3209_ _7080_/Q VGND VGND VPWR VPWR _3209_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4189_ _4189_/A0 _5208_/A1 _4193_/S VGND VGND VPWR VPWR _6629_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold190 hold190/A VGND VGND VPWR VPWR hold190/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_8_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _6731_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_160_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3560_ _3559_/X _6778_/Q _3739_/S VGND VGND VPWR VPWR _6778_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3491_ _3553_/A _3550_/B VGND VGND VPWR VPWR _4200_/A sky130_fd_sc_hd__nor2_4
XFILLER_154_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5230_ _5230_/A0 hold153/X hold91/X VGND VGND VPWR VPWR _5230_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5161_ _4417_/B _4698_/Y _4788_/X _5117_/X _5160_/X VGND VGND VPWR VPWR _5162_/C
+ sky130_fd_sc_hd__o2111a_1
Xhold2508 _6448_/Q VGND VGND VPWR VPWR _3860_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2519 _7146_/Q VGND VGND VPWR VPWR _5606_/S sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4112_ _4112_/A0 hold872/A _4115_/S VGND VGND VPWR VPWR _6565_/D sky130_fd_sc_hd__mux2_1
XFILLER_111_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1807 _6620_/Q VGND VGND VPWR VPWR hold565/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1818 _4179_/X VGND VGND VPWR VPWR _6621_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5092_ _5149_/B _5137_/B _5092_/C VGND VGND VPWR VPWR _5092_/X sky130_fd_sc_hd__and3_1
XFILLER_96_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1829 _5348_/X VGND VGND VPWR VPWR _6928_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4043_ hold397/X _5585_/A1 _4056_/C VGND VGND VPWR VPWR _4043_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5994_ _6017_/B _6019_/B _6018_/B VGND VGND VPWR VPWR _5994_/X sky130_fd_sc_hd__and3_4
XFILLER_24_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4945_ _4368_/A _4477_/Y _4729_/A _4550_/Y _4944_/X VGND VGND VPWR VPWR _5090_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_52_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4876_ _4522_/B _4507_/Y _5108_/C _5089_/B _4875_/X VGND VGND VPWR VPWR _4876_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_177_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6615_ _6794_/CLK _6615_/D fanout444/X VGND VGND VPWR VPWR _6615_/Q sky130_fd_sc_hd__dfrtp_4
X_3827_ _6657_/Q _3827_/B _3827_/C VGND VGND VPWR VPWR _3827_/Y sky130_fd_sc_hd__nor3_1
XFILLER_193_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6546_ _7194_/CLK _6546_/D VGND VGND VPWR VPWR _6546_/Q sky130_fd_sc_hd__dfxtp_1
X_3758_ _7013_/Q _5443_/A _4146_/A _6594_/Q _3757_/X VGND VGND VPWR VPWR _3759_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_824 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6477_ _6822_/CLK _6477_/D fanout451/X VGND VGND VPWR VPWR _6477_/Q sky130_fd_sc_hd__dfstp_4
X_3689_ _6753_/Q _4328_/A _4077_/A _6536_/Q _3688_/X VGND VGND VPWR VPWR _3694_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5428_ _5428_/A0 _5572_/A1 _5433_/S VGND VGND VPWR VPWR _5428_/X sky130_fd_sc_hd__mux2_1
Xoutput240 _3932_/X VGND VGND VPWR VPWR mgmt_gpio_out[36] sky130_fd_sc_hd__buf_12
XFILLER_133_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput251 _3964_/X VGND VGND VPWR VPWR pad_flash_io0_do sky130_fd_sc_hd__buf_12
Xoutput262 _6784_/Q VGND VGND VPWR VPWR pll_div[0] sky130_fd_sc_hd__buf_12
XFILLER_0_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput273 _6474_/Q VGND VGND VPWR VPWR pll_trim[11] sky130_fd_sc_hd__buf_12
XFILLER_114_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput284 _6800_/Q VGND VGND VPWR VPWR pll_trim[21] sky130_fd_sc_hd__buf_12
X_5359_ _5359_/A0 _5575_/A1 _5361_/S VGND VGND VPWR VPWR _5359_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput295 _6471_/Q VGND VGND VPWR VPWR pll_trim[8] sky130_fd_sc_hd__buf_12
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7029_ _7109_/CLK _7029_/D fanout453/X VGND VGND VPWR VPWR _7029_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_114_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4730_ _4955_/D _4730_/B VGND VGND VPWR VPWR _4823_/C sky130_fd_sc_hd__nand2_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4661_ _5150_/C VGND VGND VPWR VPWR _4661_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6400_ _6414_/A _6433_/B VGND VGND VPWR VPWR _6400_/X sky130_fd_sc_hd__and2_1
XFILLER_174_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3612_ _7128_/Q _5569_/A _4140_/A _6592_/Q _3611_/X VGND VGND VPWR VPWR _3612_/X
+ sky130_fd_sc_hd__a221o_1
X_4592_ _4575_/C _4638_/A VGND VGND VPWR VPWR _4989_/B sky130_fd_sc_hd__and2b_2
XFILLER_116_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6331_ _6741_/Q _6008_/X _6016_/X _6454_/Q VGND VGND VPWR VPWR _6331_/X sky130_fd_sc_hd__a22o_1
Xhold904 _3249_/X VGND VGND VPWR VPWR hold52/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_116_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3543_ _3543_/A _3543_/B _3543_/C VGND VGND VPWR VPWR _3557_/C sky130_fd_sc_hd__nor3_2
XFILLER_127_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold915 _4007_/X VGND VGND VPWR VPWR _6485_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold926 _4053_/X VGND VGND VPWR VPWR hold48/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold937 _5468_/X VGND VGND VPWR VPWR _7035_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold948 _5539_/X VGND VGND VPWR VPWR hold83/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold959 _3339_/Y VGND VGND VPWR VPWR _3988_/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6262_ _6585_/Q _5989_/X _6013_/X _6625_/Q _6261_/X VGND VGND VPWR VPWR _6263_/D
+ sky130_fd_sc_hd__a221o_1
X_3474_ _6849_/Q hold40/A _4116_/A _6573_/Q VGND VGND VPWR VPWR _3474_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5213_ _5213_/A0 _5303_/A1 _5217_/S VGND VGND VPWR VPWR _6811_/D sky130_fd_sc_hd__mux2_1
XFILLER_103_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6193_ _7028_/Q _5971_/X _5987_/X _7116_/Q VGND VGND VPWR VPWR _6193_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2305 _5572_/X VGND VGND VPWR VPWR _7127_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2316 _7101_/Q VGND VGND VPWR VPWR hold817/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2327 hold570/X VGND VGND VPWR VPWR _5347_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5144_ _4648_/Y _4995_/B _5011_/X _4661_/Y _4735_/Y VGND VGND VPWR VPWR _5144_/X
+ sky130_fd_sc_hd__o221a_1
Xhold2338 _6639_/Q VGND VGND VPWR VPWR hold799/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2349 hold612/X VGND VGND VPWR VPWR _5232_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1604 hold834/X VGND VGND VPWR VPWR hold258/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1615 hold608/X VGND VGND VPWR VPWR _4251_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1626 _4046_/X VGND VGND VPWR VPWR hold339/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1637 _4252_/X VGND VGND VPWR VPWR _6688_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5075_ _4402_/Y _4947_/B _4510_/B _4510_/A VGND VGND VPWR VPWR _5100_/D sky130_fd_sc_hd__a31o_1
Xhold1648 _6821_/Q VGND VGND VPWR VPWR hold691/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1659 _6704_/Q VGND VGND VPWR VPWR hold592/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4026_ _4054_/A0 _5585_/A1 _4047_/C VGND VGND VPWR VPWR _4026_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5977_ _6015_/B _6008_/A _6017_/A VGND VGND VPWR VPWR _5977_/X sky130_fd_sc_hd__and3_4
XFILLER_52_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4928_ _5100_/C _4928_/B _4928_/C VGND VGND VPWR VPWR _5112_/B sky130_fd_sc_hd__and3_1
XFILLER_21_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4859_ _4701_/A _4638_/Y _4701_/B _5073_/B VGND VGND VPWR VPWR _4859_/X sky130_fd_sc_hd__o31a_1
XFILLER_165_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6529_ _6731_/CLK _6529_/D fanout465/X VGND VGND VPWR VPWR _6529_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_118_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_73_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6793_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_11_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _6760_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_26_csclk _6850_/CLK VGND VGND VPWR VPWR _7126_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_171_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3190_ _6684_/Q VGND VGND VPWR VPWR _3967_/A sky130_fd_sc_hd__clkinv_2
XFILLER_182_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5900_ _6585_/Q _5662_/X _5897_/X _5898_/X _5899_/X VGND VGND VPWR VPWR _5900_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_81_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6880_ _7140_/CLK _6880_/D fanout469/X VGND VGND VPWR VPWR _6880_/Q sky130_fd_sc_hd__dfrtp_4
X_5831_ _6851_/Q _5842_/A2 _5662_/X _6899_/Q VGND VGND VPWR VPWR _5831_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5762_ _6912_/Q _5670_/X _5674_/X _6872_/Q _5761_/X VGND VGND VPWR VPWR _5770_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4713_ _4713_/A _4714_/B _4713_/C VGND VGND VPWR VPWR _4713_/Y sky130_fd_sc_hd__nand3_4
X_5693_ _6877_/Q _5667_/X _5688_/X _6885_/Q VGND VGND VPWR VPWR _5693_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4644_ _4732_/B _5048_/B VGND VGND VPWR VPWR _5121_/A sky130_fd_sc_hd__nand2_1
XFILLER_190_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4575_ _4637_/A _4637_/B _4575_/C _4637_/D VGND VGND VPWR VPWR _4710_/A sky130_fd_sc_hd__and4bb_4
Xhold701 hold701/A VGND VGND VPWR VPWR hold701/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold712 hold712/A VGND VGND VPWR VPWR hold712/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold723 hold723/A VGND VGND VPWR VPWR hold723/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold734 hold734/A VGND VGND VPWR VPWR hold734/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3526_ hold26/X _3550_/B VGND VGND VPWR VPWR _4065_/A sky130_fd_sc_hd__nor2_4
X_6314_ _6295_/X _6314_/B _6314_/C VGND VGND VPWR VPWR _6314_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_89_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold745 _4049_/X VGND VGND VPWR VPWR _6510_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold756 hold756/A VGND VGND VPWR VPWR hold756/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold767 hold767/A VGND VGND VPWR VPWR hold767/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold778 hold778/A VGND VGND VPWR VPWR hold778/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6245_ _6753_/Q _5638_/X _6015_/X _6758_/Q VGND VGND VPWR VPWR _6245_/X sky130_fd_sc_hd__a22o_1
Xhold789 hold789/A VGND VGND VPWR VPWR hold789/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3457_ hold49/A _3311_/Y _5551_/A _7114_/Q VGND VGND VPWR VPWR _3457_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2102 _5295_/X VGND VGND VPWR VPWR _6881_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2113 _6917_/Q VGND VGND VPWR VPWR hold678/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2124 _4019_/X VGND VGND VPWR VPWR _6495_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_6176_ _7115_/Q _5987_/X _5993_/X _7011_/Q _6175_/X VGND VGND VPWR VPWR _6179_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2135 _6747_/Q VGND VGND VPWR VPWR hold789/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_3388_ _3387_/X _3388_/A1 _3739_/S VGND VGND VPWR VPWR _6781_/D sky130_fd_sc_hd__mux2_1
Xhold1401 _6647_/Q VGND VGND VPWR VPWR hold325/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2146 _5492_/X VGND VGND VPWR VPWR _7056_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2157 hold655/X VGND VGND VPWR VPWR _4021_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1412 hold322/X VGND VGND VPWR VPWR _4260_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5127_ _5127_/A _5127_/B _5127_/C _5127_/D VGND VGND VPWR VPWR _5127_/X sky130_fd_sc_hd__and4_1
Xhold1423 _6834_/Q VGND VGND VPWR VPWR hold415/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2168 _7213_/A VGND VGND VPWR VPWR hold635/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1434 _6486_/Q VGND VGND VPWR VPWR hold395/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2179 _4126_/X VGND VGND VPWR VPWR _6577_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_183_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1445 _4275_/X VGND VGND VPWR VPWR hold297/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1456 _6815_/Q VGND VGND VPWR VPWR hold143/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1467 _5559_/X VGND VGND VPWR VPWR _7116_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5058_ _5108_/B _5110_/A _5058_/C _5058_/D VGND VGND VPWR VPWR _5059_/C sky130_fd_sc_hd__and4_1
XFILLER_55_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1478 _4281_/X VGND VGND VPWR VPWR hold320/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1489 _6711_/Q VGND VGND VPWR VPWR _4279_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4009_ _4009_/A _5551_/B VGND VGND VPWR VPWR _4011_/S sky130_fd_sc_hd__and2_1
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold50 hold50/A VGND VGND VPWR VPWR hold50/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold61 hold61/A VGND VGND VPWR VPWR hold61/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold72 hold72/A VGND VGND VPWR VPWR hold72/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold83 hold83/A VGND VGND VPWR VPWR hold83/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold94 hold94/A VGND VGND VPWR VPWR hold94/X sky130_fd_sc_hd__clkbuf_4
Xhold1990 _6618_/Q VGND VGND VPWR VPWR _4175_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_3 _5344_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4360_ _4360_/A _4360_/B VGND VGND VPWR VPWR _4465_/B sky130_fd_sc_hd__nand2_2
XFILLER_98_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3311_ _3563_/A _3726_/A VGND VGND VPWR VPWR _3311_/Y sky130_fd_sc_hd__nor2_8
XFILLER_4_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4291_ _4291_/A0 _5196_/A1 _4291_/S VGND VGND VPWR VPWR _6721_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6030_ _6925_/Q _5982_/X _6014_/X _6989_/Q VGND VGND VPWR VPWR _6030_/X sky130_fd_sc_hd__a22o_1
XFILLER_112_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3242_ _6970_/Q VGND VGND VPWR VPWR _3242_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6932_ _7130_/CLK _6932_/D fanout458/X VGND VGND VPWR VPWR _6932_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6863_ _6941_/CLK _6863_/D fanout460/X VGND VGND VPWR VPWR _6863_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_34_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5814_ _7026_/Q _5663_/X _5809_/X _5811_/X _5813_/X VGND VGND VPWR VPWR _5814_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6794_ _6794_/CLK _6794_/D fanout444/X VGND VGND VPWR VPWR _6794_/Q sky130_fd_sc_hd__dfrtp_4
X_5745_ _6943_/Q _5658_/X _5664_/X _7015_/Q VGND VGND VPWR VPWR _5745_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5676_ _5679_/B _5676_/B VGND VGND VPWR VPWR _5677_/B sky130_fd_sc_hd__nand2_8
XFILLER_135_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4627_ _4522_/B _4569_/B _4889_/B _4586_/Y _4626_/X VGND VGND VPWR VPWR _4627_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_135_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold520 hold520/A VGND VGND VPWR VPWR hold520/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold531 hold531/A VGND VGND VPWR VPWR hold531/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4558_ _4767_/A _5114_/A _4556_/X _4557_/X _4374_/Y VGND VGND VPWR VPWR _4558_/X
+ sky130_fd_sc_hd__a41o_1
Xhold542 hold542/A VGND VGND VPWR VPWR hold542/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold553 hold553/A VGND VGND VPWR VPWR hold553/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold564 hold564/A VGND VGND VPWR VPWR hold564/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold575 hold575/A VGND VGND VPWR VPWR hold575/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3509_ _3563_/A _3533_/B VGND VGND VPWR VPWR _3509_/Y sky130_fd_sc_hd__nor2_4
XFILLER_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold586 hold586/A VGND VGND VPWR VPWR hold586/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4489_ _4981_/A _4972_/A VGND VGND VPWR VPWR _5095_/A sky130_fd_sc_hd__nand2_2
Xhold597 hold597/A VGND VGND VPWR VPWR hold597/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6228_ _6609_/Q _5976_/B _5993_/X _6619_/Q VGND VGND VPWR VPWR _6228_/X sky130_fd_sc_hd__a22o_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _6898_/Q _5989_/X _6013_/X _7082_/Q _6158_/X VGND VGND VPWR VPWR _6163_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_66_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1220 _6608_/Q VGND VGND VPWR VPWR hold119/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1231 _5530_/X VGND VGND VPWR VPWR _7090_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1242 _5225_/S VGND VGND VPWR VPWR _5224_/S sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1253 _6607_/Q VGND VGND VPWR VPWR hold195/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1264 _4302_/X VGND VGND VPWR VPWR _6730_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1275 _6755_/Q VGND VGND VPWR VPWR hold186/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_122_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1286 _6716_/Q VGND VGND VPWR VPWR hold128/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1297 hold226/X VGND VGND VPWR VPWR hold1297/X sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput140 wb_dat_i[17] VGND VGND VPWR VPWR _6364_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_95_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput151 wb_dat_i[27] VGND VGND VPWR VPWR _6370_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput162 wb_dat_i[8] VGND VGND VPWR VPWR _6361_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3860_ _3860_/A0 wire1/X _3860_/S VGND VGND VPWR VPWR _6448_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3791_ _6450_/Q _3977_/A _4286_/A _6717_/Q _3790_/X VGND VGND VPWR VPWR _3792_/D
+ sky130_fd_sc_hd__a221o_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5530_ _5530_/A0 _5575_/A1 _5532_/S VGND VGND VPWR VPWR _5530_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5461_ _5461_/A _5551_/B VGND VGND VPWR VPWR _5469_/S sky130_fd_sc_hd__and2_4
XFILLER_118_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4412_ _4575_/C _4719_/A VGND VGND VPWR VPWR _4804_/A sky130_fd_sc_hd__and2b_2
X_7200_ _7204_/CLK _7200_/D fanout484/X VGND VGND VPWR VPWR _7200_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_160_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5392_ _5392_/A0 _5518_/A1 _5397_/S VGND VGND VPWR VPWR _6967_/D sky130_fd_sc_hd__mux2_1
XFILLER_126_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4343_ _4343_/A _4343_/B _4343_/C _4343_/D VGND VGND VPWR VPWR _4346_/A sky130_fd_sc_hd__and4_1
X_7131_ _7131_/CLK _7131_/D fanout469/X VGND VGND VPWR VPWR _7131_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7062_ _7140_/CLK _7062_/D fanout471/X VGND VGND VPWR VPWR _7062_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_86_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4274_ _4274_/A hold13/A VGND VGND VPWR VPWR _4279_/S sky130_fd_sc_hd__and2_4
XFILLER_140_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6013_ _6019_/A _6017_/B _6019_/B VGND VGND VPWR VPWR _6013_/X sky130_fd_sc_hd__and3_4
X_3225_ _6960_/Q VGND VGND VPWR VPWR _3225_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6915_ _7139_/CLK hold79/X fanout478/X VGND VGND VPWR VPWR _6915_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6846_ _7136_/CLK _6846_/D fanout476/X VGND VGND VPWR VPWR _6846_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_50_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6777_ _6658_/CLK _6777_/D _6429_/X VGND VGND VPWR VPWR _6777_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_149_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3989_ hold595/X _5221_/A1 _3999_/S VGND VGND VPWR VPWR _3989_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5728_ _5718_/Y _5727_/Y _6838_/Q _5678_/Y VGND VGND VPWR VPWR _5728_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5659_ _5686_/A _5679_/B _5689_/C VGND VGND VPWR VPWR _5659_/X sky130_fd_sc_hd__and3b_4
XFILLER_164_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold350 hold350/A VGND VGND VPWR VPWR hold350/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold361 hold361/A VGND VGND VPWR VPWR hold361/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold372 hold372/A VGND VGND VPWR VPWR hold372/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold383 hold383/A VGND VGND VPWR VPWR hold383/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold394 hold394/A VGND VGND VPWR VPWR hold394/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1050 _6476_/Q VGND VGND VPWR VPWR hold411/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1061 _3255_/Y VGND VGND VPWR VPWR hold88/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1072 hold390/X VGND VGND VPWR VPWR _5261_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1083 hold361/X VGND VGND VPWR VPWR _5423_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_133_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1094 _7139_/Q VGND VGND VPWR VPWR hold403/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_201 _5689_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4961_ _5151_/C _4961_/B _5042_/A _4961_/D VGND VGND VPWR VPWR _4962_/C sky130_fd_sc_hd__and4_1
X_6700_ _6757_/CLK _6700_/D fanout447/X VGND VGND VPWR VPWR _6700_/Q sky130_fd_sc_hd__dfrtp_4
X_3912_ _3909_/X _3912_/B VGND VGND VPWR VPWR _3912_/X sky130_fd_sc_hd__and2b_1
X_4892_ _4892_/A _4892_/B _4892_/C _4892_/D VGND VGND VPWR VPWR _4892_/X sky130_fd_sc_hd__and4_1
XFILLER_189_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6631_ _6792_/CLK _6631_/D fanout442/X VGND VGND VPWR VPWR _6631_/Q sky130_fd_sc_hd__dfstp_2
X_3843_ _6461_/Q _3840_/B _3846_/S VGND VGND VPWR VPWR _3843_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_149_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3774_ _7109_/Q _5551_/A _3486_/Y _3772_/X _3773_/X VGND VGND VPWR VPWR _3774_/X
+ sky130_fd_sc_hd__a2111o_1
X_6562_ _6568_/CLK _6562_/D VGND VGND VPWR VPWR _6562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5513_ _5513_/A0 _5585_/A1 _5514_/S VGND VGND VPWR VPWR _5513_/X sky130_fd_sc_hd__mux2_1
X_6493_ _6523_/CLK _6493_/D fanout480/X VGND VGND VPWR VPWR _7214_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_173_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5444_ hold778/X _5570_/A1 _5451_/S VGND VGND VPWR VPWR _7013_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5375_ _5375_/A0 _5582_/A1 _5379_/S VGND VGND VPWR VPWR _6952_/D sky130_fd_sc_hd__mux2_1
X_7114_ _7140_/CLK hold59/X fanout470/X VGND VGND VPWR VPWR _7114_/Q sky130_fd_sc_hd__dfrtp_2
X_4326_ _4326_/A0 _5303_/A1 _4327_/S VGND VGND VPWR VPWR _4326_/X sky130_fd_sc_hd__mux2_1
X_4257_ _4257_/A0 _5208_/A1 _4261_/S VGND VGND VPWR VPWR _4257_/X sky130_fd_sc_hd__mux2_1
X_7045_ _7077_/CLK _7045_/D fanout456/X VGND VGND VPWR VPWR _7045_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_59_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3208_ _7088_/Q VGND VGND VPWR VPWR _3208_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4188_ _4188_/A _5220_/C VGND VGND VPWR VPWR _4193_/S sky130_fd_sc_hd__and2_4
XFILLER_28_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6829_ _7053_/CLK _6829_/D fanout452/X VGND VGND VPWR VPWR _6829_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_183_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold180 hold932/X VGND VGND VPWR VPWR hold933/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold191 hold191/A VGND VGND VPWR VPWR hold849/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3490_ _6969_/Q _5389_/A _3389_/Y _3486_/Y _3489_/X VGND VGND VPWR VPWR _3499_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_185_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5160_ _4417_/B _4691_/Y _4785_/X _5152_/B _4893_/A VGND VGND VPWR VPWR _5160_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2509 _7159_/Q VGND VGND VPWR VPWR _5646_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4111_ _3616_/Y hold867/A _4115_/S VGND VGND VPWR VPWR _6564_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5091_ _4417_/B _4688_/C _4779_/X _4954_/A _5149_/A VGND VGND VPWR VPWR _5092_/C
+ sky130_fd_sc_hd__o2111a_1
Xhold1808 hold565/X VGND VGND VPWR VPWR _4178_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1819 _7063_/Q VGND VGND VPWR VPWR hold255/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4042_ hold944/X _4041_/X _4046_/S VGND VGND VPWR VPWR _4042_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5993_ _6015_/B _6017_/A _6019_/B VGND VGND VPWR VPWR _5993_/X sky130_fd_sc_hd__and3_4
X_4944_ _4601_/A _4491_/Y _4514_/B _4947_/A VGND VGND VPWR VPWR _4944_/X sky130_fd_sc_hd__o22a_1
XFILLER_177_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4875_ _5124_/B _4930_/A _4875_/C _4875_/D VGND VGND VPWR VPWR _4875_/X sky130_fd_sc_hd__and4_1
XFILLER_177_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6614_ _6817_/CLK _6614_/D fanout444/X VGND VGND VPWR VPWR _6614_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3826_ hold86/A _3826_/B VGND VGND VPWR VPWR _3827_/C sky130_fd_sc_hd__nor2_1
XFILLER_193_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6545_ _7194_/CLK _6545_/D VGND VGND VPWR VPWR _6545_/Q sky130_fd_sc_hd__dfxtp_1
X_3757_ input4/X _3307_/Y _3339_/Y _6471_/Q VGND VGND VPWR VPWR _3757_/X sky130_fd_sc_hd__a22o_1
XFILLER_180_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6476_ _6822_/CLK _6476_/D fanout451/X VGND VGND VPWR VPWR _6476_/Q sky130_fd_sc_hd__dfstp_2
X_3688_ _6688_/Q _4250_/A _4092_/A _6549_/Q VGND VGND VPWR VPWR _3688_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput230 _7225_/X VGND VGND VPWR VPWR mgmt_gpio_out[27] sky130_fd_sc_hd__buf_12
X_5427_ hold753/X _5580_/A1 _5433_/S VGND VGND VPWR VPWR _5427_/X sky130_fd_sc_hd__mux2_1
Xoutput241 _3931_/X VGND VGND VPWR VPWR mgmt_gpio_out[37] sky130_fd_sc_hd__buf_12
Xoutput252 _3961_/A VGND VGND VPWR VPWR pad_flash_io0_ieb sky130_fd_sc_hd__buf_12
Xoutput263 _6785_/Q VGND VGND VPWR VPWR pll_div[1] sky130_fd_sc_hd__buf_12
XFILLER_121_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput274 _6475_/Q VGND VGND VPWR VPWR pll_trim[12] sky130_fd_sc_hd__buf_12
Xoutput285 _6801_/Q VGND VGND VPWR VPWR pll_trim[22] sky130_fd_sc_hd__buf_12
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5358_ _5358_/A0 _5583_/A1 _5361_/S VGND VGND VPWR VPWR _6937_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput296 _6472_/Q VGND VGND VPWR VPWR pll_trim[9] sky130_fd_sc_hd__buf_12
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4309_ _4309_/A0 _5196_/A1 _4309_/S VGND VGND VPWR VPWR _6736_/D sky130_fd_sc_hd__mux2_1
X_5289_ _5289_/A0 _5559_/A1 _5289_/S VGND VGND VPWR VPWR _5289_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7028_ _7116_/CLK _7028_/D fanout455/X VGND VGND VPWR VPWR _7028_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_75_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire346 _3735_/Y VGND VGND VPWR VPWR _3736_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_139_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire368 _4437_/Y VGND VGND VPWR VPWR _4579_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_137_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4660_ _4713_/A _4712_/B VGND VGND VPWR VPWR _5150_/C sky130_fd_sc_hd__and2_4
XFILLER_119_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3611_ _3881_/C _5236_/C _4268_/A _6705_/Q VGND VGND VPWR VPWR _3611_/X sky130_fd_sc_hd__a22o_1
X_4591_ _4596_/A _5009_/B VGND VGND VPWR VPWR _4837_/B sky130_fd_sc_hd__nand2_2
X_6330_ _6716_/Q _5973_/X _5988_/X _6573_/Q _6329_/X VGND VGND VPWR VPWR _6330_/X
+ sky130_fd_sc_hd__a221o_1
X_3542_ _7065_/Q _5497_/A _3539_/Y _6534_/Q _3541_/X VGND VGND VPWR VPWR _3543_/C
+ sky130_fd_sc_hd__a221o_1
Xhold905 _3648_/B VGND VGND VPWR VPWR hold26/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_115_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold916 _7114_/Q VGND VGND VPWR VPWR hold58/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold927 _6835_/Q VGND VGND VPWR VPWR hold927/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold938 _7042_/Q VGND VGND VPWR VPWR hold69/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold949 _6828_/Q VGND VGND VPWR VPWR hold949/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_6_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6261_ _6688_/Q _5980_/X _6017_/X _6770_/Q VGND VGND VPWR VPWR _6261_/X sky130_fd_sc_hd__a22o_1
X_3473_ hold54/X _3531_/B VGND VGND VPWR VPWR _4116_/A sky130_fd_sc_hd__nor2_4
X_5212_ _5212_/A0 hold95/X _5217_/S VGND VGND VPWR VPWR _6810_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6192_ _6192_/A1 _5730_/S _6190_/X _6191_/X VGND VGND VPWR VPWR _7179_/D sky130_fd_sc_hd__o22a_1
Xhold2306 _6502_/Q VGND VGND VPWR VPWR hold811/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2317 _6902_/Q VGND VGND VPWR VPWR hold773/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2328 _5347_/X VGND VGND VPWR VPWR _6927_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5143_ _5143_/A _5143_/B VGND VGND VPWR VPWR _5143_/Y sky130_fd_sc_hd__nand2_1
Xhold2339 hold799/X VGND VGND VPWR VPWR _4201_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1605 _6585_/Q VGND VGND VPWR VPWR hold680/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1616 _4251_/X VGND VGND VPWR VPWR _6687_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1627 _6692_/Q VGND VGND VPWR VPWR hold685/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5074_ _5103_/A _5074_/B _5074_/C _5156_/A VGND VGND VPWR VPWR _5074_/X sky130_fd_sc_hd__and4_1
Xhold1638 _6606_/Q VGND VGND VPWR VPWR hold203/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1649 hold691/X VGND VGND VPWR VPWR _5227_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4025_ hold933/X _4024_/X _4029_/S VGND VGND VPWR VPWR _4025_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5976_ _6973_/Q _5976_/B VGND VGND VPWR VPWR _5976_/X sky130_fd_sc_hd__and2_1
XFILLER_40_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4927_ _4633_/B _4688_/B _4845_/X _5121_/B _4901_/B VGND VGND VPWR VPWR _4931_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_33_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4858_ _4705_/Y _4857_/Y _4640_/Y VGND VGND VPWR VPWR _4928_/C sky130_fd_sc_hd__a21o_1
XFILLER_193_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3809_ _6470_/Q _6469_/Q VGND VGND VPWR VPWR _3847_/B sky130_fd_sc_hd__and2_2
XFILLER_119_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4789_ _4464_/Y _4570_/B _4674_/Y _4947_/A VGND VGND VPWR VPWR _4789_/X sky130_fd_sc_hd__o22a_1
XFILLER_4_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6528_ _6816_/CLK _6528_/D _6409_/A VGND VGND VPWR VPWR _6528_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_119_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_7_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _6729_/CLK sky130_fd_sc_hd__clkbuf_16
X_6459_ _6656_/CLK _6459_/D _6409_/X VGND VGND VPWR VPWR _6459_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5830_ _6931_/Q _5684_/X _5689_/X _7083_/Q _5829_/X VGND VGND VPWR VPWR _5835_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5761_ _7064_/Q _5671_/X _5672_/X _6952_/Q VGND VGND VPWR VPWR _5761_/X sky130_fd_sc_hd__a22o_1
XFILLER_188_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4712_ _4712_/A _4712_/B _4712_/C VGND VGND VPWR VPWR _4712_/Y sky130_fd_sc_hd__nand3_4
XFILLER_175_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5692_ _7061_/Q _5671_/X _5685_/X _7069_/Q _5691_/X VGND VGND VPWR VPWR _5692_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_187_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4643_ _4506_/A _4642_/Y _4643_/C _4643_/D VGND VGND VPWR VPWR _5048_/B sky130_fd_sc_hd__and4bb_2
XFILLER_190_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4574_ _4575_/C _4638_/A VGND VGND VPWR VPWR _5011_/B sky130_fd_sc_hd__nand2_4
Xhold702 hold702/A VGND VGND VPWR VPWR hold702/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold713 hold713/A VGND VGND VPWR VPWR hold713/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6313_ _6306_/X _6308_/X _6313_/C _6339_/B VGND VGND VPWR VPWR _6314_/C sky130_fd_sc_hd__and4bb_1
XFILLER_115_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold724 hold724/A VGND VGND VPWR VPWR hold724/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap432 _4582_/A VGND VGND VPWR VPWR _4724_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_190_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold735 hold735/A VGND VGND VPWR VPWR hold735/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3525_ _6993_/Q _5416_/A _5308_/A _6897_/Q _3524_/X VGND VGND VPWR VPWR _3529_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_116_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold746 hold746/A VGND VGND VPWR VPWR hold746/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold757 hold757/A VGND VGND VPWR VPWR hold757/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold768 hold768/A VGND VGND VPWR VPWR hold768/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold779 hold779/A VGND VGND VPWR VPWR hold779/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6244_ _6645_/Q _5990_/X _5996_/X _6650_/Q VGND VGND VPWR VPWR _6244_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3456_ _6858_/Q _5263_/A _5335_/A _6922_/Q _3455_/X VGND VGND VPWR VPWR _3460_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2103 _7111_/Q VGND VGND VPWR VPWR hold632/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2114 _6877_/Q VGND VGND VPWR VPWR hold602/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_3387_ _3424_/A1 _3385_/Y _3857_/B VGND VGND VPWR VPWR _3387_/X sky130_fd_sc_hd__mux2_1
X_6175_ _6859_/Q _5983_/X _5988_/X _6875_/Q VGND VGND VPWR VPWR _6175_/X sky130_fd_sc_hd__a22o_1
Xhold2125 _6795_/Q VGND VGND VPWR VPWR hold779/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2136 hold789/X VGND VGND VPWR VPWR _4323_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2147 _6575_/Q VGND VGND VPWR VPWR hold715/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1402 hold325/X VGND VGND VPWR VPWR _4210_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2158 _4021_/X VGND VGND VPWR VPWR _6496_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1413 _4260_/X VGND VGND VPWR VPWR _6695_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5126_ _5126_/A _5126_/B _5126_/C VGND VGND VPWR VPWR _5127_/D sky130_fd_sc_hd__and3_1
Xhold1424 hold415/X VGND VGND VPWR VPWR _5242_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2169 hold635/X VGND VGND VPWR VPWR _4040_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1435 _6738_/Q VGND VGND VPWR VPWR hold137/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1446 _7133_/Q VGND VGND VPWR VPWR hold292/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1457 _5217_/X VGND VGND VPWR VPWR _6815_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1468 _7220_/A VGND VGND VPWR VPWR hold616/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5057_ _4384_/A _4969_/A _5115_/B _4930_/C _5114_/C VGND VGND VPWR VPWR _5058_/D
+ sky130_fd_sc_hd__o2111a_1
Xhold1479 _6908_/Q VGND VGND VPWR VPWR hold492/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_55_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4008_ hold395/X _5559_/A1 _4008_/S VGND VGND VPWR VPWR _6486_/D sky130_fd_sc_hd__mux2_1
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5959_ _6552_/Q _5673_/X _5954_/X _5955_/X _5958_/X VGND VGND VPWR VPWR _5959_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_179_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold40 hold40/A VGND VGND VPWR VPWR hold40/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold51 hold51/A VGND VGND VPWR VPWR hold51/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold62 hold62/A VGND VGND VPWR VPWR hold62/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold73 hold73/A VGND VGND VPWR VPWR hold73/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold84 hold84/A VGND VGND VPWR VPWR hold84/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold95 hold95/A VGND VGND VPWR VPWR hold95/X sky130_fd_sc_hd__buf_12
XFILLER_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1980 hold590/X VGND VGND VPWR VPWR _4139_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1991 _4175_/X VGND VGND VPWR VPWR hold96/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_90_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_4 _3311_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3310_ _3764_/B _3531_/B VGND VGND VPWR VPWR _3310_/Y sky130_fd_sc_hd__nor2_8
X_4290_ _4290_/A0 _5303_/A1 _4291_/S VGND VGND VPWR VPWR _4290_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3241_ _6721_/Q VGND VGND VPWR VPWR _3241_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6931_ _7091_/CLK _6931_/D fanout471/X VGND VGND VPWR VPWR _6931_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6862_ _7008_/CLK _6862_/D fanout474/X VGND VGND VPWR VPWR _6862_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5813_ _6858_/Q _5651_/X _5688_/X _6890_/Q _5812_/X VGND VGND VPWR VPWR _5813_/X
+ sky130_fd_sc_hd__a221o_1
X_6793_ _6793_/CLK _6793_/D fanout442/X VGND VGND VPWR VPWR _6793_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_50_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5744_ _6895_/Q _5662_/X _5742_/X _5743_/X VGND VGND VPWR VPWR _5744_/X sky130_fd_sc_hd__a211o_1
XFILLER_148_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5675_ _5679_/B _5676_/B VGND VGND VPWR VPWR _5678_/B sky130_fd_sc_hd__and2_4
Xclkbuf_leaf_72_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6747_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_135_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4626_ _4522_/B _4569_/A _4898_/B _4624_/X _4625_/Y VGND VGND VPWR VPWR _4626_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_163_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold510 hold510/A VGND VGND VPWR VPWR hold510/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold521 hold521/A VGND VGND VPWR VPWR hold521/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4557_ _4384_/A _4658_/A _4417_/B _5127_/A VGND VGND VPWR VPWR _4557_/X sky130_fd_sc_hd__o31a_1
Xhold532 hold532/A VGND VGND VPWR VPWR hold532/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold543 hold543/A VGND VGND VPWR VPWR hold543/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold554 hold554/A VGND VGND VPWR VPWR hold554/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold565 hold565/A VGND VGND VPWR VPWR hold565/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3508_ _7097_/Q _5533_/A _4182_/A _6628_/Q _3506_/X VGND VGND VPWR VPWR _3515_/B
+ sky130_fd_sc_hd__a221o_1
Xhold576 hold576/A VGND VGND VPWR VPWR hold576/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4488_ _4595_/B _4488_/B VGND VGND VPWR VPWR _4510_/B sky130_fd_sc_hd__nand2_4
Xhold587 hold587/A VGND VGND VPWR VPWR hold587/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold598 hold598/A VGND VGND VPWR VPWR hold598/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6227_ _6629_/Q _5971_/X _6007_/X _6530_/Q _6226_/X VGND VGND VPWR VPWR _6230_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_104_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3439_ _7018_/Q _5443_/A _3319_/Y _6800_/Q _3433_/X VGND VGND VPWR VPWR _3444_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_58_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _6938_/Q _5980_/X _6017_/X _7074_/Q VGND VGND VPWR VPWR _6158_/X sky130_fd_sc_hd__a22o_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1210 hold254/X VGND VGND VPWR VPWR _4067_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1221 hold119/X VGND VGND VPWR VPWR _4163_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xclkbuf_leaf_10_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _6711_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_66_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1232 _7017_/Q VGND VGND VPWR VPWR hold123/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1243 _5224_/X VGND VGND VPWR VPWR _6819_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5109_ _4500_/Y _4640_/Y _4919_/C _5125_/B _4757_/A VGND VGND VPWR VPWR _5110_/B
+ sky130_fd_sc_hd__o2111a_1
X_6089_ _6079_/X _6339_/B _6089_/C _6089_/D VGND VGND VPWR VPWR _6089_/X sky130_fd_sc_hd__and4b_1
Xhold1254 hold195/X VGND VGND VPWR VPWR _4162_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1265 _6563_/Q VGND VGND VPWR VPWR hold869/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1276 hold186/X VGND VGND VPWR VPWR _4332_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1287 hold128/X VGND VGND VPWR VPWR _4285_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1298 _6826_/Q VGND VGND VPWR VPWR hold221/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_csclk _6850_/CLK VGND VGND VPWR VPWR _7016_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_53_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput130 wb_adr_i[9] VGND VGND VPWR VPWR _4345_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput141 wb_dat_i[18] VGND VGND VPWR VPWR _6368_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput152 wb_dat_i[28] VGND VGND VPWR VPWR _6374_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput163 wb_dat_i[9] VGND VGND VPWR VPWR _6365_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3790_ _6629_/Q _4188_/A _4262_/A _6697_/Q VGND VGND VPWR VPWR _3790_/X sky130_fd_sc_hd__a22o_1
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5460_ _5460_/A0 _5559_/A1 _5460_/S VGND VGND VPWR VPWR _5460_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4411_ _4719_/A _4590_/B VGND VGND VPWR VPWR _4411_/Y sky130_fd_sc_hd__nand2_4
XFILLER_126_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5391_ hold777/X _5580_/A1 _5397_/S VGND VGND VPWR VPWR _6966_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7130_ _7130_/CLK _7130_/D fanout460/X VGND VGND VPWR VPWR _7130_/Q sky130_fd_sc_hd__dfrtp_2
X_4342_ _4720_/C _4395_/A VGND VGND VPWR VPWR _4560_/A sky130_fd_sc_hd__nor2_4
XFILLER_113_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7061_ _7109_/CLK _7061_/D fanout453/X VGND VGND VPWR VPWR _7061_/Q sky130_fd_sc_hd__dfstp_2
X_4273_ _4273_/A0 hold95/X _4273_/S VGND VGND VPWR VPWR _4273_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6012_ _6015_/B _6019_/B _6018_/B VGND VGND VPWR VPWR _6012_/X sky130_fd_sc_hd__and3_4
X_3224_ _6720_/Q VGND VGND VPWR VPWR _3224_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
.ends

