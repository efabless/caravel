magic
tech sky130A
timestamp 1637698310
<< fillblock >>
rect 186540 7419 197809 9621
use font_53  font_53_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598768855
transform 1 0 187474 0 1 7963
box 0 0 540 1260
use font_61  font_61_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598775307
transform 1 0 188192 0 1 7967
box 0 0 540 900
use font_69  font_69_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598776260
transform 1 0 188908 0 1 7967
box 0 0 360 1260
use font_6C  font_6C_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598776550
transform 1 0 189441 0 1 7971
box 0 0 180 1260
use font_69  font_69_1
timestamp 1598776260
transform 1 0 189798 0 1 7971
box 0 0 360 1260
use font_6E  font_6E_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598776997
transform 1 0 190337 0 1 7971
box 0 0 540 900
use font_67  font_67_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598776042
transform 1 0 191057 0 1 7971
box 0 -360 540 900
use font_54  font_54_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598768910
transform 1 0 192288 0 1 7971
box 0 0 540 1260
use font_68  font_68_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598776130
transform 1 0 193003 0 1 7965
box 0 0 540 1260
use font_65  font_65_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598775915
transform 1 0 193719 0 1 7965
box 0 0 540 900
use font_49  font_49_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598765816
transform 1 0 194956 0 1 7973
box 0 0 540 1260
use font_43  font_43_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598763351
transform 1 0 195675 0 1 7969
box 0 0 540 1260
use font_73  font_73_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598777283
transform 1 0 196393 0 1 7963
box 0 0 540 900
use font_22  font_22_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598785768
transform 1 0 186753 0 1 8245
box 0 540 540 1260
use font_22  font_22_1
timestamp 1598785768
transform 1 0 197105 0 1 8265
box 0 540 540 1260
<< end >>
