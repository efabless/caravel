magic
tech sky130A
magscale 1 2
timestamp 1637274817
<< locali >>
rect 4537 5695 4571 5797
rect 15853 5695 15887 5865
rect 10149 3927 10183 4029
rect 18981 2975 19015 3893
rect 12541 2431 12575 2601
<< viali >>
rect 1317 9537 1351 9571
rect 8033 9537 8067 9571
rect 8677 9537 8711 9571
rect 9229 9537 9263 9571
rect 9505 9537 9539 9571
rect 9597 9537 9631 9571
rect 9781 9537 9815 9571
rect 10057 9537 10091 9571
rect 10425 9537 10459 9571
rect 10793 9537 10827 9571
rect 13277 9537 13311 9571
rect 15577 9537 15611 9571
rect 17923 9537 17957 9571
rect 18153 9537 18187 9571
rect 18337 9537 18371 9571
rect 2329 9469 2363 9503
rect 5825 9469 5859 9503
rect 6101 9469 6135 9503
rect 8769 9469 8803 9503
rect 11069 9469 11103 9503
rect 11345 9469 11379 9503
rect 13553 9469 13587 9503
rect 13921 9469 13955 9503
rect 16129 9469 16163 9503
rect 16497 9469 16531 9503
rect 18245 9469 18279 9503
rect 7849 9401 7883 9435
rect 9413 9401 9447 9435
rect 9505 9401 9539 9435
rect 13093 9401 13127 9435
rect 7573 9333 7607 9367
rect 9965 9333 9999 9367
rect 10609 9333 10643 9367
rect 10885 9333 10919 9367
rect 12817 9333 12851 9367
rect 15347 9333 15381 9367
rect 16911 9129 16945 9163
rect 18337 9129 18371 9163
rect 10287 9061 10321 9095
rect 10701 9061 10735 9095
rect 14933 9061 14967 9095
rect 7021 8993 7055 9027
rect 8125 8993 8159 9027
rect 8401 8993 8435 9027
rect 8493 8993 8527 9027
rect 13001 8993 13035 9027
rect 15117 8993 15151 9027
rect 15485 8993 15519 9027
rect 673 8925 707 8959
rect 2697 8925 2731 8959
rect 8033 8925 8067 8959
rect 8861 8925 8895 8959
rect 10517 8925 10551 8959
rect 10701 8925 10735 8959
rect 10977 8925 11011 8959
rect 12817 8925 12851 8959
rect 15025 8925 15059 8959
rect 17969 8925 18003 8959
rect 18521 8925 18555 8959
rect 2973 8857 3007 8891
rect 6745 8857 6779 8891
rect 12541 8857 12575 8891
rect 13277 8857 13311 8891
rect 581 8789 615 8823
rect 4445 8789 4479 8823
rect 5273 8789 5307 8823
rect 11069 8789 11103 8823
rect 14749 8789 14783 8823
rect 17785 8789 17819 8823
rect 2973 8585 3007 8619
rect 5733 8585 5767 8619
rect 5825 8585 5859 8619
rect 6469 8585 6503 8619
rect 6929 8585 6963 8619
rect 8125 8585 8159 8619
rect 8493 8585 8527 8619
rect 9321 8585 9355 8619
rect 14565 8585 14599 8619
rect 5457 8517 5491 8551
rect 5641 8517 5675 8551
rect 9045 8517 9079 8551
rect 10762 8517 10796 8551
rect 14289 8517 14323 8551
rect 16773 8517 16807 8551
rect 397 8449 431 8483
rect 2191 8449 2225 8483
rect 2513 8449 2547 8483
rect 3709 8449 3743 8483
rect 3893 8449 3927 8483
rect 4169 8449 4203 8483
rect 5733 8449 5767 8483
rect 7021 8449 7055 8483
rect 8953 8449 8987 8483
rect 9137 8449 9171 8483
rect 9597 8449 9631 8483
rect 10241 8449 10275 8483
rect 10517 8449 10551 8483
rect 12081 8449 12115 8483
rect 12173 8449 12207 8483
rect 12265 8449 12299 8483
rect 12541 8449 12575 8483
rect 14933 8449 14967 8483
rect 15577 8449 15611 8483
rect 765 8381 799 8415
rect 3157 8381 3191 8415
rect 3249 8381 3283 8415
rect 3617 8381 3651 8415
rect 6193 8381 6227 8415
rect 6285 8381 6319 8415
rect 7205 8381 7239 8415
rect 8585 8381 8619 8415
rect 8769 8381 8803 8415
rect 9505 8381 9539 8415
rect 9965 8381 9999 8415
rect 15025 8381 15059 8415
rect 15117 8381 15151 8415
rect 16497 8381 16531 8415
rect 18521 8381 18555 8415
rect 4077 8313 4111 8347
rect 6561 8313 6595 8347
rect 12449 8313 12483 8347
rect 15761 8313 15795 8347
rect 2421 8245 2455 8279
rect 3893 8245 3927 8279
rect 10149 8245 10183 8279
rect 11897 8245 11931 8279
rect 2237 8041 2271 8075
rect 3341 8041 3375 8075
rect 3893 8041 3927 8075
rect 5089 8041 5123 8075
rect 6009 8041 6043 8075
rect 6561 8041 6595 8075
rect 7021 8041 7055 8075
rect 11437 8041 11471 8075
rect 13001 8041 13035 8075
rect 16484 8041 16518 8075
rect 2145 7973 2179 8007
rect 3157 7973 3191 8007
rect 2329 7905 2363 7939
rect 4905 7905 4939 7939
rect 5733 7905 5767 7939
rect 6377 7905 6411 7939
rect 7205 7905 7239 7939
rect 9137 7905 9171 7939
rect 11989 7905 12023 7939
rect 13461 7905 13495 7939
rect 13645 7905 13679 7939
rect 14289 7905 14323 7939
rect 16221 7905 16255 7939
rect 1777 7837 1811 7871
rect 1961 7837 1995 7871
rect 2072 7837 2106 7871
rect 2697 7837 2731 7871
rect 2789 7837 2823 7871
rect 3249 7837 3283 7871
rect 3617 7837 3651 7871
rect 3801 7837 3835 7871
rect 4077 7837 4111 7871
rect 4169 7815 4203 7849
rect 4261 7837 4295 7871
rect 4813 7837 4847 7871
rect 4997 7837 5031 7871
rect 5457 7837 5491 7871
rect 5917 7837 5951 7871
rect 6101 7837 6135 7871
rect 6653 7837 6687 7871
rect 7297 7837 7331 7871
rect 7849 7837 7883 7871
rect 8125 7837 8159 7871
rect 11253 7837 11287 7871
rect 11713 7837 11747 7871
rect 12173 7837 12207 7871
rect 13369 7837 13403 7871
rect 13829 7837 13863 7871
rect 14105 7837 14139 7871
rect 14657 7837 14691 7871
rect 18521 7837 18555 7871
rect 7941 7769 7975 7803
rect 11897 7769 11931 7803
rect 13921 7769 13955 7803
rect 1961 7701 1995 7735
rect 2973 7701 3007 7735
rect 3525 7701 3559 7735
rect 5549 7701 5583 7735
rect 6377 7701 6411 7735
rect 7665 7701 7699 7735
rect 7849 7701 7883 7735
rect 8493 7701 8527 7735
rect 8861 7701 8895 7735
rect 8953 7701 8987 7735
rect 9965 7701 9999 7735
rect 12817 7701 12851 7735
rect 13829 7701 13863 7735
rect 16083 7701 16117 7735
rect 17969 7701 18003 7735
rect 18337 7701 18371 7735
rect 2605 7497 2639 7531
rect 3525 7497 3559 7531
rect 4721 7497 4755 7531
rect 7205 7497 7239 7531
rect 3985 7429 4019 7463
rect 6101 7429 6135 7463
rect 6469 7429 6503 7463
rect 6745 7429 6779 7463
rect 8309 7429 8343 7463
rect 8769 7429 8803 7463
rect 9137 7429 9171 7463
rect 14473 7429 14507 7463
rect 15209 7429 15243 7463
rect 18153 7429 18187 7463
rect 581 7361 615 7395
rect 2697 7361 2731 7395
rect 2789 7361 2823 7395
rect 2973 7361 3007 7395
rect 4813 7361 4847 7395
rect 4905 7361 4939 7395
rect 5089 7361 5123 7395
rect 5549 7361 5583 7395
rect 5641 7361 5675 7395
rect 5917 7361 5951 7395
rect 6285 7361 6319 7395
rect 6929 7361 6963 7395
rect 7021 7361 7055 7395
rect 7297 7361 7331 7395
rect 8953 7361 8987 7395
rect 9321 7361 9355 7395
rect 9413 7361 9447 7395
rect 9873 7361 9907 7395
rect 9965 7361 9999 7395
rect 10793 7361 10827 7395
rect 11621 7361 11655 7395
rect 14105 7361 14139 7395
rect 14749 7361 14783 7395
rect 15945 7361 15979 7395
rect 857 7293 891 7327
rect 2329 7293 2363 7327
rect 2881 7293 2915 7327
rect 6653 7293 6687 7327
rect 8401 7293 8435 7327
rect 8585 7293 8619 7327
rect 10149 7293 10183 7327
rect 10885 7293 10919 7327
rect 10977 7293 11011 7327
rect 11529 7293 11563 7327
rect 11989 7293 12023 7327
rect 12357 7293 12391 7327
rect 14013 7293 14047 7327
rect 14657 7293 14691 7327
rect 16037 7293 16071 7327
rect 16405 7293 16439 7327
rect 18429 7293 18463 7327
rect 3709 7225 3743 7259
rect 5733 7225 5767 7259
rect 7941 7225 7975 7259
rect 9505 7225 9539 7259
rect 10425 7225 10459 7259
rect 11253 7225 11287 7259
rect 15025 7225 15059 7259
rect 15577 7225 15611 7259
rect 4997 7157 5031 7191
rect 5825 7157 5859 7191
rect 7021 7157 7055 7191
rect 9413 7157 9447 7191
rect 13783 7157 13817 7191
rect 7205 6953 7239 6987
rect 13737 6953 13771 6987
rect 13829 6953 13863 6987
rect 15209 6953 15243 6987
rect 3801 6885 3835 6919
rect 6009 6885 6043 6919
rect 3157 6817 3191 6851
rect 3341 6817 3375 6851
rect 3985 6817 4019 6851
rect 5457 6817 5491 6851
rect 7021 6817 7055 6851
rect 8217 6817 8251 6851
rect 9643 6817 9677 6851
rect 11989 6817 12023 6851
rect 12449 6817 12483 6851
rect 12541 6817 12575 6851
rect 13093 6817 13127 6851
rect 13277 6817 13311 6851
rect 14427 6817 14461 6851
rect 16589 6817 16623 6851
rect 16957 6817 16991 6851
rect 17601 6817 17635 6851
rect 3065 6749 3099 6783
rect 3249 6749 3283 6783
rect 3525 6749 3559 6783
rect 3617 6749 3651 6783
rect 3893 6749 3927 6783
rect 4261 6749 4295 6783
rect 5273 6749 5307 6783
rect 5825 6749 5859 6783
rect 6009 6749 6043 6783
rect 6285 6749 6319 6783
rect 7205 6749 7239 6783
rect 7849 6749 7883 6783
rect 9873 6749 9907 6783
rect 11897 6749 11931 6783
rect 12081 6749 12115 6783
rect 12265 6749 12299 6783
rect 12725 6749 12759 6783
rect 12817 6749 12851 6783
rect 13369 6749 13403 6783
rect 14841 6749 14875 6783
rect 14933 6749 14967 6783
rect 17509 6749 17543 6783
rect 18153 6749 18187 6783
rect 3341 6681 3375 6715
rect 7297 6681 7331 6715
rect 7481 6681 7515 6715
rect 11621 6681 11655 6715
rect 14657 6681 14691 6715
rect 4905 6613 4939 6647
rect 5365 6613 5399 6647
rect 6377 6613 6411 6647
rect 6745 6613 6779 6647
rect 6837 6613 6871 6647
rect 12541 6613 12575 6647
rect 14197 6613 14231 6647
rect 14289 6613 14323 6647
rect 14749 6613 14783 6647
rect 17049 6613 17083 6647
rect 17417 6613 17451 6647
rect 18337 6613 18371 6647
rect 3893 6409 3927 6443
rect 4261 6409 4295 6443
rect 4353 6409 4387 6443
rect 6009 6409 6043 6443
rect 6469 6409 6503 6443
rect 8033 6409 8067 6443
rect 8401 6409 8435 6443
rect 11437 6409 11471 6443
rect 15025 6409 15059 6443
rect 17509 6409 17543 6443
rect 17969 6409 18003 6443
rect 1685 6341 1719 6375
rect 3525 6341 3559 6375
rect 3709 6341 3743 6375
rect 4813 6341 4847 6375
rect 6101 6341 6135 6375
rect 6929 6341 6963 6375
rect 8852 6341 8886 6375
rect 12081 6341 12115 6375
rect 14197 6341 14231 6375
rect 14381 6341 14415 6375
rect 17877 6341 17911 6375
rect 1409 6273 1443 6307
rect 3249 6273 3283 6307
rect 3433 6273 3467 6307
rect 3801 6273 3835 6307
rect 4905 6273 4939 6307
rect 5273 6273 5307 6307
rect 5457 6273 5491 6307
rect 6837 6273 6871 6307
rect 8125 6273 8159 6307
rect 8493 6273 8527 6307
rect 10057 6273 10091 6307
rect 10241 6273 10275 6307
rect 10885 6273 10919 6307
rect 11253 6273 11287 6307
rect 11713 6273 11747 6307
rect 11897 6273 11931 6307
rect 15117 6273 15151 6307
rect 15577 6273 15611 6307
rect 17371 6273 17405 6307
rect 18337 6273 18371 6307
rect 4445 6205 4479 6239
rect 6285 6205 6319 6239
rect 7021 6205 7055 6239
rect 8585 6205 8619 6239
rect 10977 6205 11011 6239
rect 11069 6205 11103 6239
rect 12173 6205 12207 6239
rect 12541 6205 12575 6239
rect 15209 6205 15243 6239
rect 15945 6205 15979 6239
rect 18153 6205 18187 6239
rect 18429 6205 18463 6239
rect 3157 6137 3191 6171
rect 5365 6137 5399 6171
rect 5641 6137 5675 6171
rect 9965 6137 9999 6171
rect 10241 6137 10275 6171
rect 14657 6137 14691 6171
rect 3341 6069 3375 6103
rect 3801 6069 3835 6103
rect 10425 6069 10459 6103
rect 10609 6069 10643 6103
rect 13967 6069 14001 6103
rect 6653 5865 6687 5899
rect 9505 5865 9539 5899
rect 12817 5865 12851 5899
rect 15761 5865 15795 5899
rect 15853 5865 15887 5899
rect 17233 5865 17267 5899
rect 18337 5865 18371 5899
rect 3249 5797 3283 5831
rect 4353 5797 4387 5831
rect 4537 5797 4571 5831
rect 765 5729 799 5763
rect 1041 5729 1075 5763
rect 3157 5729 3191 5763
rect 3893 5729 3927 5763
rect 5917 5729 5951 5763
rect 7205 5729 7239 5763
rect 8125 5729 8159 5763
rect 10977 5729 11011 5763
rect 14013 5729 14047 5763
rect 16129 5797 16163 5831
rect 17877 5729 17911 5763
rect 3341 5661 3375 5695
rect 3433 5661 3467 5695
rect 3617 5661 3651 5695
rect 3709 5661 3743 5695
rect 4169 5661 4203 5695
rect 4445 5661 4479 5695
rect 4537 5661 4571 5695
rect 4629 5661 4663 5695
rect 4997 5661 5031 5695
rect 5365 5661 5399 5695
rect 5549 5661 5583 5695
rect 5733 5661 5767 5695
rect 6009 5661 6043 5695
rect 7849 5661 7883 5695
rect 8033 5661 8067 5695
rect 8392 5661 8426 5695
rect 11069 5661 11103 5695
rect 13277 5661 13311 5695
rect 13553 5661 13587 5695
rect 13737 5661 13771 5695
rect 15853 5661 15887 5695
rect 15945 5661 15979 5695
rect 16221 5661 16255 5695
rect 16313 5661 16347 5695
rect 16681 5661 16715 5695
rect 17141 5661 17175 5695
rect 17601 5661 17635 5695
rect 18521 5661 18555 5695
rect 3893 5593 3927 5627
rect 4077 5593 4111 5627
rect 7113 5593 7147 5627
rect 10721 5593 10755 5627
rect 11345 5593 11379 5627
rect 14289 5593 14323 5627
rect 2513 5525 2547 5559
rect 5365 5525 5399 5559
rect 5641 5525 5675 5559
rect 6377 5525 6411 5559
rect 7021 5525 7055 5559
rect 7941 5525 7975 5559
rect 9597 5525 9631 5559
rect 13093 5525 13127 5559
rect 13461 5525 13495 5559
rect 13921 5525 13955 5559
rect 16221 5525 16255 5559
rect 16865 5525 16899 5559
rect 17693 5525 17727 5559
rect 4951 5321 4985 5355
rect 8033 5321 8067 5355
rect 10241 5321 10275 5355
rect 13185 5321 13219 5355
rect 16681 5321 16715 5355
rect 18521 5321 18555 5355
rect 9965 5253 9999 5287
rect 10149 5253 10183 5287
rect 3157 5185 3191 5219
rect 5917 5185 5951 5219
rect 7573 5185 7607 5219
rect 10241 5185 10275 5219
rect 10885 5185 10919 5219
rect 11161 5185 11195 5219
rect 13093 5185 13127 5219
rect 13553 5185 13587 5219
rect 16313 5185 16347 5219
rect 16773 5185 16807 5219
rect 3525 5117 3559 5151
rect 5825 5117 5859 5151
rect 6285 5117 6319 5151
rect 7665 5117 7699 5151
rect 7941 5117 7975 5151
rect 9505 5117 9539 5151
rect 9781 5117 9815 5151
rect 10425 5117 10459 5151
rect 11529 5117 11563 5151
rect 13829 5117 13863 5151
rect 16405 5117 16439 5151
rect 17049 5117 17083 5151
rect 12955 5049 12989 5083
rect 10793 4981 10827 5015
rect 15301 4981 15335 5015
rect 7941 4777 7975 4811
rect 11713 4777 11747 4811
rect 12725 4777 12759 4811
rect 14197 4777 14231 4811
rect 14473 4777 14507 4811
rect 14933 4777 14967 4811
rect 15761 4777 15795 4811
rect 7573 4709 7607 4743
rect 8033 4709 8067 4743
rect 10241 4709 10275 4743
rect 18337 4709 18371 4743
rect 8585 4641 8619 4675
rect 9597 4641 9631 4675
rect 11897 4641 11931 4675
rect 13645 4641 13679 4675
rect 13921 4641 13955 4675
rect 15485 4641 15519 4675
rect 5825 4573 5859 4607
rect 8125 4573 8159 4607
rect 8493 4573 8527 4607
rect 11989 4573 12023 4607
rect 12357 4573 12391 4607
rect 12633 4573 12667 4607
rect 12817 4573 12851 4607
rect 13369 4573 13403 4607
rect 13829 4573 13863 4607
rect 14007 4573 14041 4607
rect 14097 4575 14131 4609
rect 14381 4573 14415 4607
rect 14933 4573 14967 4607
rect 15117 4573 15151 4607
rect 15393 4573 15427 4607
rect 17601 4573 17635 4607
rect 17969 4573 18003 4607
rect 18521 4573 18555 4607
rect 6101 4505 6135 4539
rect 7849 4505 7883 4539
rect 9413 4505 9447 4539
rect 11529 4505 11563 4539
rect 12541 4505 12575 4539
rect 8861 4437 8895 4471
rect 8953 4437 8987 4471
rect 9321 4437 9355 4471
rect 13001 4437 13035 4471
rect 13461 4437 13495 4471
rect 14841 4437 14875 4471
rect 15853 4437 15887 4471
rect 6377 4233 6411 4267
rect 7389 4233 7423 4267
rect 8401 4233 8435 4267
rect 9321 4233 9355 4267
rect 13921 4233 13955 4267
rect 7297 4165 7331 4199
rect 9045 4165 9079 4199
rect 10885 4165 10919 4199
rect 11897 4165 11931 4199
rect 15577 4165 15611 4199
rect 6561 4097 6595 4131
rect 7757 4097 7791 4131
rect 8493 4097 8527 4131
rect 9689 4097 9723 4131
rect 10481 4097 10515 4131
rect 10609 4119 10643 4153
rect 10701 4087 10735 4121
rect 11069 4097 11103 4131
rect 11437 4097 11471 4131
rect 11621 4097 11655 4131
rect 12541 4097 12575 4131
rect 12808 4097 12842 4131
rect 14280 4097 14314 4131
rect 18521 4097 18555 4131
rect 7573 4029 7607 4063
rect 8677 4029 8711 4063
rect 9781 4029 9815 4063
rect 9965 4029 9999 4063
rect 10149 4029 10183 4063
rect 14013 4029 14047 4063
rect 17325 4029 17359 4063
rect 17601 4029 17635 4063
rect 6929 3961 6963 3995
rect 8033 3961 8067 3995
rect 11069 3961 11103 3995
rect 12265 3961 12299 3995
rect 7941 3893 7975 3927
rect 8953 3893 8987 3927
rect 10149 3893 10183 3927
rect 11529 3893 11563 3927
rect 12357 3893 12391 3927
rect 15393 3893 15427 3927
rect 18337 3893 18371 3927
rect 18981 3893 19015 3927
rect 9597 3689 9631 3723
rect 14657 3689 14691 3723
rect 5273 3621 5307 3655
rect 11713 3621 11747 3655
rect 13461 3621 13495 3655
rect 5089 3553 5123 3587
rect 5457 3553 5491 3587
rect 7849 3553 7883 3587
rect 12173 3553 12207 3587
rect 12357 3553 12391 3587
rect 12541 3553 12575 3587
rect 15945 3553 15979 3587
rect 3525 3485 3559 3519
rect 5365 3485 5399 3519
rect 8217 3485 8251 3519
rect 9965 3485 9999 3519
rect 10333 3485 10367 3519
rect 10600 3485 10634 3519
rect 11805 3485 11839 3519
rect 11989 3485 12023 3519
rect 12265 3485 12299 3519
rect 12633 3485 12667 3519
rect 12817 3485 12851 3519
rect 13001 3485 13035 3519
rect 13369 3485 13403 3519
rect 13645 3485 13679 3519
rect 14381 3485 14415 3519
rect 14933 3485 14967 3519
rect 15025 3485 15059 3519
rect 15209 3485 15243 3519
rect 5733 3417 5767 3451
rect 12725 3417 12759 3451
rect 16221 3417 16255 3451
rect 17969 3417 18003 3451
rect 3433 3349 3467 3383
rect 5089 3349 5123 3383
rect 7205 3349 7239 3383
rect 9873 3349 9907 3383
rect 12541 3349 12575 3383
rect 14841 3349 14875 3383
rect 14933 3349 14967 3383
rect 5825 3145 5859 3179
rect 6009 3145 6043 3179
rect 12449 3145 12483 3179
rect 12909 3145 12943 3179
rect 15393 3145 15427 3179
rect 15669 3145 15703 3179
rect 16451 3145 16485 3179
rect 6285 3077 6319 3111
rect 15117 3077 15151 3111
rect 3249 3009 3283 3043
rect 3617 3009 3651 3043
rect 5043 3009 5077 3043
rect 5457 3009 5491 3043
rect 5549 3009 5583 3043
rect 5733 3009 5767 3043
rect 6101 3009 6135 3043
rect 6193 3009 6227 3043
rect 6469 3009 6503 3043
rect 6653 3009 6687 3043
rect 6837 3009 6871 3043
rect 7021 3009 7055 3043
rect 7941 3009 7975 3043
rect 8125 3009 8159 3043
rect 8401 3009 8435 3043
rect 10609 3009 10643 3043
rect 12081 3009 12115 3043
rect 13093 3009 13127 3043
rect 13737 3009 13771 3043
rect 13921 3009 13955 3043
rect 14381 3009 14415 3043
rect 14565 3009 14599 3043
rect 14657 3009 14691 3043
rect 14841 3009 14875 3043
rect 15301 3009 15335 3043
rect 15393 3009 15427 3043
rect 18245 3009 18279 3043
rect 18521 3009 18555 3043
rect 6561 2941 6595 2975
rect 6929 2941 6963 2975
rect 8769 2941 8803 2975
rect 10195 2941 10229 2975
rect 11989 2941 12023 2975
rect 13369 2941 13403 2975
rect 16037 2941 16071 2975
rect 16129 2941 16163 2975
rect 16313 2941 16347 2975
rect 17877 2941 17911 2975
rect 18981 2941 19015 2975
rect 5365 2873 5399 2907
rect 10517 2873 10551 2907
rect 7941 2805 7975 2839
rect 13277 2805 13311 2839
rect 13461 2805 13495 2839
rect 13737 2805 13771 2839
rect 14197 2805 14231 2839
rect 14933 2805 14967 2839
rect 18337 2805 18371 2839
rect 5733 2601 5767 2635
rect 6469 2601 6503 2635
rect 9413 2601 9447 2635
rect 12403 2601 12437 2635
rect 12541 2601 12575 2635
rect 7849 2533 7883 2567
rect 4813 2465 4847 2499
rect 5273 2465 5307 2499
rect 8401 2465 8435 2499
rect 9137 2465 9171 2499
rect 9229 2465 9263 2499
rect 10609 2465 10643 2499
rect 12725 2533 12759 2567
rect 18153 2533 18187 2567
rect 14013 2465 14047 2499
rect 16129 2465 16163 2499
rect 16405 2465 16439 2499
rect 4905 2397 4939 2431
rect 5457 2397 5491 2431
rect 5733 2397 5767 2431
rect 5917 2397 5951 2431
rect 6101 2397 6135 2431
rect 6193 2397 6227 2431
rect 6285 2397 6319 2431
rect 6745 2397 6779 2431
rect 6837 2397 6871 2431
rect 7481 2397 7515 2431
rect 7665 2397 7699 2431
rect 9505 2397 9539 2431
rect 9597 2397 9631 2431
rect 9781 2397 9815 2431
rect 10057 2397 10091 2431
rect 10977 2397 11011 2431
rect 12541 2397 12575 2431
rect 12633 2397 12667 2431
rect 13093 2397 13127 2431
rect 13185 2397 13219 2431
rect 13277 2397 13311 2431
rect 13461 2397 13495 2431
rect 13553 2397 13587 2431
rect 13829 2397 13863 2431
rect 18153 2397 18187 2431
rect 8769 2329 8803 2363
rect 9045 2329 9079 2363
rect 13645 2329 13679 2363
rect 14289 2329 14323 2363
rect 16037 2329 16071 2363
rect 4629 2261 4663 2295
rect 7665 2261 7699 2295
rect 8217 2261 8251 2295
rect 8309 2261 8343 2295
rect 8861 2261 8895 2295
rect 9873 2261 9907 2295
rect 13553 2261 13587 2295
rect 17877 2261 17911 2295
rect 5089 2057 5123 2091
rect 5273 2057 5307 2091
rect 5917 2057 5951 2091
rect 6837 2057 6871 2091
rect 7297 2057 7331 2091
rect 7757 2057 7791 2091
rect 8769 2057 8803 2091
rect 8953 2057 8987 2091
rect 12541 2057 12575 2091
rect 12633 2057 12667 2091
rect 13829 2057 13863 2091
rect 14565 2057 14599 2091
rect 16773 2057 16807 2091
rect 3617 1989 3651 2023
rect 6193 1989 6227 2023
rect 6929 1989 6963 2023
rect 9045 1989 9079 2023
rect 9229 1989 9263 2023
rect 10609 1989 10643 2023
rect 12449 1989 12483 2023
rect 15853 1989 15887 2023
rect 18245 1989 18279 2023
rect 3341 1921 3375 1955
rect 5733 1921 5767 1955
rect 5825 1921 5859 1955
rect 6009 1921 6043 1955
rect 6285 1921 6319 1955
rect 7665 1921 7699 1955
rect 8217 1921 8251 1955
rect 8401 1921 8435 1955
rect 8585 1921 8619 1955
rect 8677 1921 8711 1955
rect 8861 1921 8895 1955
rect 8953 1921 8987 1955
rect 9321 1921 9355 1955
rect 9505 1921 9539 1955
rect 9597 1921 9631 1955
rect 9781 1921 9815 1955
rect 10701 1921 10735 1955
rect 10977 1921 11011 1955
rect 11437 1921 11471 1955
rect 12265 1921 12299 1955
rect 12541 1921 12575 1955
rect 13921 1921 13955 1955
rect 14289 1921 14323 1955
rect 14933 1921 14967 1955
rect 15577 1921 15611 1955
rect 15669 1921 15703 1955
rect 16313 1921 16347 1955
rect 18521 1921 18555 1955
rect 7113 1853 7147 1887
rect 7941 1853 7975 1887
rect 11161 1853 11195 1887
rect 13001 1853 13035 1887
rect 13093 1853 13127 1887
rect 14013 1853 14047 1887
rect 15025 1853 15059 1887
rect 15117 1853 15151 1887
rect 16405 1853 16439 1887
rect 16589 1853 16623 1887
rect 5457 1785 5491 1819
rect 13461 1785 13495 1819
rect 6469 1717 6503 1751
rect 8401 1717 8435 1751
rect 9413 1717 9447 1751
rect 9689 1717 9723 1751
rect 11529 1717 11563 1751
rect 13277 1717 13311 1751
rect 14381 1717 14415 1751
rect 15577 1717 15611 1751
rect 15945 1717 15979 1751
rect 14749 1513 14783 1547
rect 15025 1513 15059 1547
rect 17233 1513 17267 1547
rect 7389 1445 7423 1479
rect 5733 1377 5767 1411
rect 7297 1377 7331 1411
rect 7481 1377 7515 1411
rect 8125 1377 8159 1411
rect 9505 1377 9539 1411
rect 9597 1377 9631 1411
rect 10517 1377 10551 1411
rect 11161 1377 11195 1411
rect 11253 1377 11287 1411
rect 12081 1377 12115 1411
rect 14473 1377 14507 1411
rect 15669 1377 15703 1411
rect 16037 1377 16071 1411
rect 16129 1377 16163 1411
rect 16957 1377 16991 1411
rect 17693 1377 17727 1411
rect 17785 1377 17819 1411
rect 5457 1309 5491 1343
rect 7573 1309 7607 1343
rect 7849 1309 7883 1343
rect 8769 1309 8803 1343
rect 11989 1309 12023 1343
rect 14381 1309 14415 1343
rect 14841 1309 14875 1343
rect 14933 1309 14967 1343
rect 15301 1309 15335 1343
rect 15393 1309 15427 1343
rect 10241 1241 10275 1275
rect 15117 1241 15151 1275
rect 16865 1241 16899 1275
rect 7205 1173 7239 1207
rect 8861 1173 8895 1207
rect 9045 1173 9079 1207
rect 9413 1173 9447 1207
rect 9873 1173 9907 1207
rect 10333 1173 10367 1207
rect 10701 1173 10735 1207
rect 11069 1173 11103 1207
rect 11529 1173 11563 1207
rect 11897 1173 11931 1207
rect 16313 1173 16347 1207
rect 16405 1173 16439 1207
rect 16773 1173 16807 1207
rect 17601 1173 17635 1207
rect 6469 969 6503 1003
rect 8631 969 8665 1003
rect 9137 969 9171 1003
rect 10517 969 10551 1003
rect 11345 969 11379 1003
rect 12081 969 12115 1003
rect 15117 969 15151 1003
rect 17509 969 17543 1003
rect 17877 969 17911 1003
rect 17969 969 18003 1003
rect 18429 969 18463 1003
rect 8861 901 8895 935
rect 9045 901 9079 935
rect 9873 901 9907 935
rect 13553 901 13587 935
rect 6285 833 6319 867
rect 6469 833 6503 867
rect 6561 833 6595 867
rect 7205 833 7239 867
rect 9137 833 9171 867
rect 9505 833 9539 867
rect 9597 833 9631 867
rect 10057 833 10091 867
rect 10149 833 10183 867
rect 10425 833 10459 867
rect 10701 833 10735 867
rect 11253 833 11287 867
rect 11713 833 11747 867
rect 13829 833 13863 867
rect 15025 833 15059 867
rect 15209 833 15243 867
rect 15945 833 15979 867
rect 18337 833 18371 867
rect 6653 765 6687 799
rect 6837 765 6871 799
rect 9229 765 9263 799
rect 9873 765 9907 799
rect 11621 765 11655 799
rect 15577 765 15611 799
rect 18061 765 18095 799
rect 9413 697 9447 731
rect 9689 697 9723 731
rect 9321 629 9355 663
rect 17371 629 17405 663
rect 7389 425 7423 459
rect 10977 425 11011 459
rect 17417 425 17451 459
rect 18337 425 18371 459
rect 11069 357 11103 391
rect 8401 289 8435 323
rect 8677 289 8711 323
rect 10149 289 10183 323
rect 10701 289 10735 323
rect 17049 289 17083 323
rect 7481 221 7515 255
rect 10609 221 10643 255
rect 11069 221 11103 255
rect 11253 221 11287 255
rect 17141 221 17175 255
rect 18521 221 18555 255
<< metal1 >>
rect 0 9818 18860 9840
rect 0 9766 6144 9818
rect 6196 9766 6208 9818
rect 6260 9766 6272 9818
rect 6324 9766 6336 9818
rect 6388 9766 6400 9818
rect 6452 9766 12443 9818
rect 12495 9766 12507 9818
rect 12559 9766 12571 9818
rect 12623 9766 12635 9818
rect 12687 9766 12699 9818
rect 12751 9766 18860 9818
rect 0 9744 18860 9766
rect 11330 9664 11336 9716
rect 11388 9704 11394 9716
rect 11388 9676 12664 9704
rect 11388 9664 11394 9676
rect 5626 9596 5632 9648
rect 5684 9636 5690 9648
rect 11422 9636 11428 9648
rect 5684 9608 6578 9636
rect 8036 9608 11428 9636
rect 5684 9596 5690 9608
rect 1302 9568 1308 9580
rect 1263 9540 1308 9568
rect 1302 9528 1308 9540
rect 1360 9528 1366 9580
rect 8036 9577 8064 9608
rect 11422 9596 11428 9608
rect 11480 9596 11486 9648
rect 11606 9596 11612 9648
rect 11664 9636 11670 9648
rect 12636 9636 12664 9676
rect 13648 9676 15056 9704
rect 13078 9636 13084 9648
rect 11664 9608 11822 9636
rect 12636 9608 13084 9636
rect 11664 9596 11670 9608
rect 13078 9596 13084 9608
rect 13136 9596 13142 9648
rect 8021 9571 8079 9577
rect 8021 9537 8033 9571
rect 8067 9537 8079 9571
rect 8021 9531 8079 9537
rect 8294 9528 8300 9580
rect 8352 9568 8358 9580
rect 8665 9571 8723 9577
rect 8665 9568 8677 9571
rect 8352 9540 8677 9568
rect 8352 9528 8358 9540
rect 8665 9537 8677 9540
rect 8711 9537 8723 9571
rect 9214 9568 9220 9580
rect 9175 9540 9220 9568
rect 8665 9531 8723 9537
rect 9214 9528 9220 9540
rect 9272 9528 9278 9580
rect 9493 9571 9551 9577
rect 9493 9568 9505 9571
rect 9324 9540 9505 9568
rect 2314 9500 2320 9512
rect 2275 9472 2320 9500
rect 2314 9460 2320 9472
rect 2372 9460 2378 9512
rect 2682 9460 2688 9512
rect 2740 9500 2746 9512
rect 5718 9500 5724 9512
rect 2740 9472 5724 9500
rect 2740 9460 2746 9472
rect 5718 9460 5724 9472
rect 5776 9500 5782 9512
rect 5813 9503 5871 9509
rect 5813 9500 5825 9503
rect 5776 9472 5825 9500
rect 5776 9460 5782 9472
rect 5813 9469 5825 9472
rect 5859 9469 5871 9503
rect 5813 9463 5871 9469
rect 6089 9503 6147 9509
rect 6089 9469 6101 9503
rect 6135 9500 6147 9503
rect 7282 9500 7288 9512
rect 6135 9472 7288 9500
rect 6135 9469 6147 9472
rect 6089 9463 6147 9469
rect 7282 9460 7288 9472
rect 7340 9460 7346 9512
rect 8757 9503 8815 9509
rect 8757 9469 8769 9503
rect 8803 9500 8815 9503
rect 9324 9500 9352 9540
rect 9493 9537 9505 9540
rect 9539 9537 9551 9571
rect 9493 9531 9551 9537
rect 9585 9571 9643 9577
rect 9585 9537 9597 9571
rect 9631 9568 9643 9571
rect 9674 9568 9680 9580
rect 9631 9540 9680 9568
rect 9631 9537 9643 9540
rect 9585 9531 9643 9537
rect 9674 9528 9680 9540
rect 9732 9528 9738 9580
rect 9766 9528 9772 9580
rect 9824 9568 9830 9580
rect 10042 9568 10048 9580
rect 9824 9540 9869 9568
rect 10003 9540 10048 9568
rect 9824 9528 9830 9540
rect 10042 9528 10048 9540
rect 10100 9528 10106 9580
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9537 10471 9571
rect 10413 9531 10471 9537
rect 10781 9571 10839 9577
rect 10781 9537 10793 9571
rect 10827 9568 10839 9571
rect 10962 9568 10968 9580
rect 10827 9540 10968 9568
rect 10827 9537 10839 9540
rect 10781 9531 10839 9537
rect 9950 9500 9956 9512
rect 8803 9472 9352 9500
rect 9416 9472 9956 9500
rect 8803 9469 8815 9472
rect 8757 9463 8815 9469
rect 7098 9392 7104 9444
rect 7156 9432 7162 9444
rect 9416 9441 9444 9472
rect 9950 9460 9956 9472
rect 10008 9460 10014 9512
rect 10428 9500 10456 9531
rect 10962 9528 10968 9540
rect 11020 9528 11026 9580
rect 13265 9571 13323 9577
rect 13265 9537 13277 9571
rect 13311 9568 13323 9571
rect 13648 9568 13676 9676
rect 14274 9596 14280 9648
rect 14332 9596 14338 9648
rect 15028 9636 15056 9676
rect 15028 9608 15700 9636
rect 15565 9571 15623 9577
rect 15565 9568 15577 9571
rect 13311 9540 13676 9568
rect 14660 9540 15577 9568
rect 13311 9537 13323 9540
rect 13265 9531 13323 9537
rect 10870 9500 10876 9512
rect 10428 9472 10876 9500
rect 10870 9460 10876 9472
rect 10928 9460 10934 9512
rect 11057 9503 11115 9509
rect 11057 9469 11069 9503
rect 11103 9469 11115 9503
rect 11330 9500 11336 9512
rect 11291 9472 11336 9500
rect 11057 9463 11115 9469
rect 7837 9435 7895 9441
rect 7837 9432 7849 9435
rect 7156 9404 7849 9432
rect 7156 9392 7162 9404
rect 7837 9401 7849 9404
rect 7883 9401 7895 9435
rect 7837 9395 7895 9401
rect 9401 9435 9459 9441
rect 9401 9401 9413 9435
rect 9447 9401 9459 9435
rect 9401 9395 9459 9401
rect 9493 9435 9551 9441
rect 9493 9401 9505 9435
rect 9539 9432 9551 9435
rect 10686 9432 10692 9444
rect 9539 9404 10692 9432
rect 9539 9401 9551 9404
rect 9493 9395 9551 9401
rect 10686 9392 10692 9404
rect 10744 9392 10750 9444
rect 10778 9392 10784 9444
rect 10836 9432 10842 9444
rect 11072 9432 11100 9463
rect 11330 9460 11336 9472
rect 11388 9460 11394 9512
rect 11422 9460 11428 9512
rect 11480 9500 11486 9512
rect 13541 9503 13599 9509
rect 13541 9500 13553 9503
rect 11480 9472 13553 9500
rect 11480 9460 11486 9472
rect 13541 9469 13553 9472
rect 13587 9469 13599 9503
rect 13541 9463 13599 9469
rect 13909 9503 13967 9509
rect 13909 9469 13921 9503
rect 13955 9500 13967 9503
rect 14660 9500 14688 9540
rect 15565 9537 15577 9540
rect 15611 9537 15623 9571
rect 15672 9568 15700 9608
rect 16850 9596 16856 9648
rect 16908 9596 16914 9648
rect 17911 9571 17969 9577
rect 15672 9540 16620 9568
rect 15565 9531 15623 9537
rect 16117 9503 16175 9509
rect 16117 9500 16129 9503
rect 13955 9472 14688 9500
rect 14752 9472 16129 9500
rect 13955 9469 13967 9472
rect 13909 9463 13967 9469
rect 10836 9404 11100 9432
rect 10836 9392 10842 9404
rect 12894 9392 12900 9444
rect 12952 9432 12958 9444
rect 13081 9435 13139 9441
rect 13081 9432 13093 9435
rect 12952 9404 13093 9432
rect 12952 9392 12958 9404
rect 13081 9401 13093 9404
rect 13127 9401 13139 9435
rect 13081 9395 13139 9401
rect 7561 9367 7619 9373
rect 7561 9333 7573 9367
rect 7607 9364 7619 9367
rect 8110 9364 8116 9376
rect 7607 9336 8116 9364
rect 7607 9333 7619 9336
rect 7561 9327 7619 9333
rect 8110 9324 8116 9336
rect 8168 9324 8174 9376
rect 9674 9324 9680 9376
rect 9732 9364 9738 9376
rect 9953 9367 10011 9373
rect 9953 9364 9965 9367
rect 9732 9336 9965 9364
rect 9732 9324 9738 9336
rect 9953 9333 9965 9336
rect 9999 9333 10011 9367
rect 10594 9364 10600 9376
rect 10555 9336 10600 9364
rect 9953 9327 10011 9333
rect 10594 9324 10600 9336
rect 10652 9324 10658 9376
rect 10873 9367 10931 9373
rect 10873 9333 10885 9367
rect 10919 9364 10931 9367
rect 11790 9364 11796 9376
rect 10919 9336 11796 9364
rect 10919 9333 10931 9336
rect 10873 9327 10931 9333
rect 11790 9324 11796 9336
rect 11848 9324 11854 9376
rect 12805 9367 12863 9373
rect 12805 9333 12817 9367
rect 12851 9364 12863 9367
rect 13170 9364 13176 9376
rect 12851 9336 13176 9364
rect 12851 9333 12863 9336
rect 12805 9327 12863 9333
rect 13170 9324 13176 9336
rect 13228 9324 13234 9376
rect 13556 9364 13584 9463
rect 14458 9364 14464 9376
rect 13556 9336 14464 9364
rect 14458 9324 14464 9336
rect 14516 9364 14522 9376
rect 14752 9364 14780 9472
rect 16117 9469 16129 9472
rect 16163 9469 16175 9503
rect 16482 9500 16488 9512
rect 16443 9472 16488 9500
rect 16117 9463 16175 9469
rect 16482 9460 16488 9472
rect 16540 9460 16546 9512
rect 16592 9500 16620 9540
rect 17911 9537 17923 9571
rect 17957 9568 17969 9571
rect 18141 9571 18199 9577
rect 18141 9568 18153 9571
rect 17957 9540 18153 9568
rect 17957 9537 17969 9540
rect 17911 9531 17969 9537
rect 18141 9537 18153 9540
rect 18187 9537 18199 9571
rect 18322 9568 18328 9580
rect 18283 9540 18328 9568
rect 18141 9531 18199 9537
rect 18322 9528 18328 9540
rect 18380 9528 18386 9580
rect 18233 9503 18291 9509
rect 18233 9500 18245 9503
rect 16592 9472 18245 9500
rect 18233 9469 18245 9472
rect 18279 9469 18291 9503
rect 18233 9463 18291 9469
rect 14516 9336 14780 9364
rect 15335 9367 15393 9373
rect 14516 9324 14522 9336
rect 15335 9333 15347 9367
rect 15381 9364 15393 9367
rect 15470 9364 15476 9376
rect 15381 9336 15476 9364
rect 15381 9333 15393 9336
rect 15335 9327 15393 9333
rect 15470 9324 15476 9336
rect 15528 9324 15534 9376
rect 16022 9324 16028 9376
rect 16080 9364 16086 9376
rect 16850 9364 16856 9376
rect 16080 9336 16856 9364
rect 16080 9324 16086 9336
rect 16850 9324 16856 9336
rect 16908 9324 16914 9376
rect 0 9274 18860 9296
rect 0 9222 2995 9274
rect 3047 9222 3059 9274
rect 3111 9222 3123 9274
rect 3175 9222 3187 9274
rect 3239 9222 3251 9274
rect 3303 9222 9294 9274
rect 9346 9222 9358 9274
rect 9410 9222 9422 9274
rect 9474 9222 9486 9274
rect 9538 9222 9550 9274
rect 9602 9222 15592 9274
rect 15644 9222 15656 9274
rect 15708 9222 15720 9274
rect 15772 9222 15784 9274
rect 15836 9222 15848 9274
rect 15900 9222 18860 9274
rect 0 9200 18860 9222
rect 2314 9120 2320 9172
rect 2372 9160 2378 9172
rect 2372 9132 4108 9160
rect 2372 9120 2378 9132
rect 566 8916 572 8968
rect 624 8956 630 8968
rect 661 8959 719 8965
rect 661 8956 673 8959
rect 624 8928 673 8956
rect 624 8916 630 8928
rect 661 8925 673 8928
rect 707 8956 719 8959
rect 2682 8956 2688 8968
rect 707 8928 2688 8956
rect 707 8925 719 8928
rect 661 8919 719 8925
rect 2682 8916 2688 8928
rect 2740 8916 2746 8968
rect 4080 8956 4108 9132
rect 5626 9120 5632 9172
rect 5684 9160 5690 9172
rect 9122 9160 9128 9172
rect 5684 9132 9128 9160
rect 5684 9120 5690 9132
rect 9122 9120 9128 9132
rect 9180 9120 9186 9172
rect 9214 9120 9220 9172
rect 9272 9160 9278 9172
rect 12986 9160 12992 9172
rect 9272 9132 12992 9160
rect 9272 9120 9278 9132
rect 12986 9120 12992 9132
rect 13044 9120 13050 9172
rect 15286 9160 15292 9172
rect 13096 9132 15292 9160
rect 7208 9064 8524 9092
rect 7208 9036 7236 9064
rect 5718 8984 5724 9036
rect 5776 9024 5782 9036
rect 7009 9027 7067 9033
rect 7009 9024 7021 9027
rect 5776 8996 7021 9024
rect 5776 8984 5782 8996
rect 7009 8993 7021 8996
rect 7055 9024 7067 9027
rect 7190 9024 7196 9036
rect 7055 8996 7196 9024
rect 7055 8993 7067 8996
rect 7009 8987 7067 8993
rect 7190 8984 7196 8996
rect 7248 8984 7254 9036
rect 8113 9027 8171 9033
rect 8113 8993 8125 9027
rect 8159 9024 8171 9027
rect 8202 9024 8208 9036
rect 8159 8996 8208 9024
rect 8159 8993 8171 8996
rect 8113 8987 8171 8993
rect 8202 8984 8208 8996
rect 8260 8984 8266 9036
rect 8386 9024 8392 9036
rect 8347 8996 8392 9024
rect 8386 8984 8392 8996
rect 8444 8984 8450 9036
rect 8496 9033 8524 9064
rect 9674 9052 9680 9104
rect 9732 9092 9738 9104
rect 10042 9092 10048 9104
rect 9732 9064 10048 9092
rect 9732 9052 9738 9064
rect 10042 9052 10048 9064
rect 10100 9092 10106 9104
rect 10275 9095 10333 9101
rect 10275 9092 10287 9095
rect 10100 9064 10287 9092
rect 10100 9052 10106 9064
rect 10275 9061 10287 9064
rect 10321 9061 10333 9095
rect 10275 9055 10333 9061
rect 10689 9095 10747 9101
rect 10689 9061 10701 9095
rect 10735 9092 10747 9095
rect 11514 9092 11520 9104
rect 10735 9064 11520 9092
rect 10735 9061 10747 9064
rect 10689 9055 10747 9061
rect 11514 9052 11520 9064
rect 11572 9052 11578 9104
rect 12802 9052 12808 9104
rect 12860 9092 12866 9104
rect 13096 9092 13124 9132
rect 15286 9120 15292 9132
rect 15344 9120 15350 9172
rect 16482 9120 16488 9172
rect 16540 9160 16546 9172
rect 16899 9163 16957 9169
rect 16899 9160 16911 9163
rect 16540 9132 16911 9160
rect 16540 9120 16546 9132
rect 16899 9129 16911 9132
rect 16945 9129 16957 9163
rect 18322 9160 18328 9172
rect 18283 9132 18328 9160
rect 16899 9123 16957 9129
rect 18322 9120 18328 9132
rect 18380 9120 18386 9172
rect 14921 9095 14979 9101
rect 14921 9092 14933 9095
rect 12860 9064 13124 9092
rect 14292 9064 14933 9092
rect 12860 9052 12866 9064
rect 8481 9027 8539 9033
rect 8481 8993 8493 9027
rect 8527 8993 8539 9027
rect 9766 9024 9772 9036
rect 8481 8987 8539 8993
rect 8956 8996 9772 9024
rect 8956 8968 8984 8996
rect 9766 8984 9772 8996
rect 9824 8984 9830 9036
rect 10778 8984 10784 9036
rect 10836 9024 10842 9036
rect 11146 9024 11152 9036
rect 10836 8996 11152 9024
rect 10836 8984 10842 8996
rect 11146 8984 11152 8996
rect 11204 9024 11210 9036
rect 12989 9027 13047 9033
rect 12989 9024 13001 9027
rect 11204 8996 13001 9024
rect 11204 8984 11210 8996
rect 12989 8993 13001 8996
rect 13035 8993 13047 9027
rect 12989 8987 13047 8993
rect 13262 8984 13268 9036
rect 13320 9024 13326 9036
rect 14292 9024 14320 9064
rect 14921 9061 14933 9064
rect 14967 9061 14979 9095
rect 14921 9055 14979 9061
rect 13320 8996 14320 9024
rect 13320 8984 13326 8996
rect 14458 8984 14464 9036
rect 14516 9024 14522 9036
rect 15105 9027 15163 9033
rect 15105 9024 15117 9027
rect 14516 8996 15117 9024
rect 14516 8984 14522 8996
rect 15105 8993 15117 8996
rect 15151 8993 15163 9027
rect 15470 9024 15476 9036
rect 15431 8996 15476 9024
rect 15105 8987 15163 8993
rect 15470 8984 15476 8996
rect 15528 8984 15534 9036
rect 17862 8984 17868 9036
rect 17920 9024 17926 9036
rect 17920 8996 18552 9024
rect 17920 8984 17926 8996
rect 5626 8956 5632 8968
rect 4080 8942 5632 8956
rect 4094 8928 5632 8942
rect 5626 8916 5632 8928
rect 5684 8916 5690 8968
rect 8021 8959 8079 8965
rect 8021 8925 8033 8959
rect 8067 8956 8079 8959
rect 8294 8956 8300 8968
rect 8067 8928 8300 8956
rect 8067 8925 8079 8928
rect 8021 8919 8079 8925
rect 2958 8888 2964 8900
rect 2919 8860 2964 8888
rect 2958 8848 2964 8860
rect 3016 8848 3022 8900
rect 6730 8888 6736 8900
rect 6691 8860 6736 8888
rect 6730 8848 6736 8860
rect 6788 8848 6794 8900
rect 382 8780 388 8832
rect 440 8820 446 8832
rect 569 8823 627 8829
rect 569 8820 581 8823
rect 440 8792 581 8820
rect 440 8780 446 8792
rect 569 8789 581 8792
rect 615 8789 627 8823
rect 569 8783 627 8789
rect 3878 8780 3884 8832
rect 3936 8820 3942 8832
rect 4338 8820 4344 8832
rect 3936 8792 4344 8820
rect 3936 8780 3942 8792
rect 4338 8780 4344 8792
rect 4396 8820 4402 8832
rect 4433 8823 4491 8829
rect 4433 8820 4445 8823
rect 4396 8792 4445 8820
rect 4396 8780 4402 8792
rect 4433 8789 4445 8792
rect 4479 8789 4491 8823
rect 4433 8783 4491 8789
rect 5261 8823 5319 8829
rect 5261 8789 5273 8823
rect 5307 8820 5319 8823
rect 5442 8820 5448 8832
rect 5307 8792 5448 8820
rect 5307 8789 5319 8792
rect 5261 8783 5319 8789
rect 5442 8780 5448 8792
rect 5500 8820 5506 8832
rect 8036 8820 8064 8919
rect 8294 8916 8300 8928
rect 8352 8916 8358 8968
rect 8846 8956 8852 8968
rect 8807 8928 8852 8956
rect 8846 8916 8852 8928
rect 8904 8916 8910 8968
rect 8938 8916 8944 8968
rect 8996 8916 9002 8968
rect 10502 8956 10508 8968
rect 10463 8928 10508 8956
rect 10502 8916 10508 8928
rect 10560 8916 10566 8968
rect 10686 8956 10692 8968
rect 10647 8928 10692 8956
rect 10686 8916 10692 8928
rect 10744 8916 10750 8968
rect 10965 8959 11023 8965
rect 10965 8925 10977 8959
rect 11011 8956 11023 8959
rect 11238 8956 11244 8968
rect 11011 8928 11244 8956
rect 11011 8925 11023 8928
rect 10965 8919 11023 8925
rect 11238 8916 11244 8928
rect 11296 8916 11302 8968
rect 12802 8916 12808 8968
rect 12860 8956 12866 8968
rect 12860 8928 12905 8956
rect 12860 8916 12866 8928
rect 14918 8916 14924 8968
rect 14976 8956 14982 8968
rect 15013 8959 15071 8965
rect 15013 8956 15025 8959
rect 14976 8928 15025 8956
rect 14976 8916 14982 8928
rect 15013 8925 15025 8928
rect 15059 8925 15071 8959
rect 15013 8919 15071 8925
rect 17770 8916 17776 8968
rect 17828 8956 17834 8968
rect 18524 8965 18552 8996
rect 17957 8959 18015 8965
rect 17957 8956 17969 8959
rect 17828 8928 17969 8956
rect 17828 8916 17834 8928
rect 17957 8925 17969 8928
rect 18003 8925 18015 8959
rect 17957 8919 18015 8925
rect 18509 8959 18567 8965
rect 18509 8925 18521 8959
rect 18555 8925 18567 8959
rect 18509 8919 18567 8925
rect 9214 8848 9220 8900
rect 9272 8848 9278 8900
rect 10410 8848 10416 8900
rect 10468 8888 10474 8900
rect 10704 8888 10732 8916
rect 11514 8892 11520 8900
rect 11348 8888 11520 8892
rect 10468 8860 10732 8888
rect 10980 8864 11520 8888
rect 10980 8860 11362 8864
rect 10468 8848 10474 8860
rect 5500 8792 8064 8820
rect 9232 8820 9260 8848
rect 10042 8820 10048 8832
rect 9232 8792 10048 8820
rect 5500 8780 5506 8792
rect 10042 8780 10048 8792
rect 10100 8820 10106 8832
rect 10980 8820 11008 8860
rect 11514 8848 11520 8864
rect 11572 8848 11578 8900
rect 12434 8888 12440 8900
rect 12406 8848 12440 8888
rect 12492 8848 12498 8900
rect 12529 8891 12587 8897
rect 12529 8857 12541 8891
rect 12575 8857 12587 8891
rect 12529 8851 12587 8857
rect 10100 8792 11008 8820
rect 11057 8823 11115 8829
rect 10100 8780 10106 8792
rect 11057 8789 11069 8823
rect 11103 8820 11115 8823
rect 12406 8820 12434 8848
rect 11103 8792 12434 8820
rect 12544 8820 12572 8851
rect 12894 8848 12900 8900
rect 12952 8888 12958 8900
rect 13265 8891 13323 8897
rect 13265 8888 13277 8891
rect 12952 8860 13277 8888
rect 12952 8848 12958 8860
rect 13265 8857 13277 8860
rect 13311 8857 13323 8891
rect 13265 8851 13323 8857
rect 13722 8848 13728 8900
rect 13780 8848 13786 8900
rect 14568 8860 15148 8888
rect 14568 8820 14596 8860
rect 14734 8820 14740 8832
rect 12544 8792 14596 8820
rect 14695 8792 14740 8820
rect 11103 8789 11115 8792
rect 11057 8783 11115 8789
rect 14734 8780 14740 8792
rect 14792 8780 14798 8832
rect 15120 8820 15148 8860
rect 16022 8848 16028 8900
rect 16080 8848 16086 8900
rect 17773 8823 17831 8829
rect 17773 8820 17785 8823
rect 15120 8792 17785 8820
rect 17773 8789 17785 8792
rect 17819 8789 17831 8823
rect 17773 8783 17831 8789
rect 0 8730 18860 8752
rect 0 8678 6144 8730
rect 6196 8678 6208 8730
rect 6260 8678 6272 8730
rect 6324 8678 6336 8730
rect 6388 8678 6400 8730
rect 6452 8678 12443 8730
rect 12495 8678 12507 8730
rect 12559 8678 12571 8730
rect 12623 8678 12635 8730
rect 12687 8678 12699 8730
rect 12751 8678 18860 8730
rect 0 8656 18860 8678
rect 2958 8616 2964 8628
rect 2919 8588 2964 8616
rect 2958 8576 2964 8588
rect 3016 8576 3022 8628
rect 5721 8619 5779 8625
rect 5721 8585 5733 8619
rect 5767 8616 5779 8619
rect 5813 8619 5871 8625
rect 5813 8616 5825 8619
rect 5767 8588 5825 8616
rect 5767 8585 5779 8588
rect 5721 8579 5779 8585
rect 5813 8585 5825 8588
rect 5859 8585 5871 8619
rect 5813 8579 5871 8585
rect 6457 8619 6515 8625
rect 6457 8585 6469 8619
rect 6503 8616 6515 8619
rect 6730 8616 6736 8628
rect 6503 8588 6736 8616
rect 6503 8585 6515 8588
rect 6457 8579 6515 8585
rect 6730 8576 6736 8588
rect 6788 8576 6794 8628
rect 6917 8619 6975 8625
rect 6917 8585 6929 8619
rect 6963 8616 6975 8619
rect 8113 8619 8171 8625
rect 8113 8616 8125 8619
rect 6963 8588 8125 8616
rect 6963 8585 6975 8588
rect 6917 8579 6975 8585
rect 8113 8585 8125 8588
rect 8159 8585 8171 8619
rect 8113 8579 8171 8585
rect 8386 8576 8392 8628
rect 8444 8616 8450 8628
rect 8481 8619 8539 8625
rect 8481 8616 8493 8619
rect 8444 8588 8493 8616
rect 8444 8576 8450 8588
rect 8481 8585 8493 8588
rect 8527 8585 8539 8619
rect 8481 8579 8539 8585
rect 8846 8576 8852 8628
rect 8904 8616 8910 8628
rect 9309 8619 9367 8625
rect 9309 8616 9321 8619
rect 8904 8588 9321 8616
rect 8904 8576 8910 8588
rect 9309 8585 9321 8588
rect 9355 8585 9367 8619
rect 9309 8579 9367 8585
rect 9582 8576 9588 8628
rect 9640 8576 9646 8628
rect 10410 8576 10416 8628
rect 10468 8616 10474 8628
rect 10468 8588 10916 8616
rect 10468 8576 10474 8588
rect 1946 8548 1952 8560
rect 1794 8520 1952 8548
rect 1946 8508 1952 8520
rect 2004 8548 2010 8560
rect 2314 8548 2320 8560
rect 2004 8520 2320 8548
rect 2004 8508 2010 8520
rect 2314 8508 2320 8520
rect 2372 8508 2378 8560
rect 5442 8548 5448 8560
rect 3068 8520 3924 8548
rect 5403 8520 5448 8548
rect 382 8480 388 8492
rect 343 8452 388 8480
rect 382 8440 388 8452
rect 440 8440 446 8492
rect 2179 8483 2237 8489
rect 2179 8449 2191 8483
rect 2225 8480 2237 8483
rect 2501 8483 2559 8489
rect 2501 8480 2513 8483
rect 2225 8452 2513 8480
rect 2225 8449 2237 8452
rect 2179 8443 2237 8449
rect 2501 8449 2513 8452
rect 2547 8480 2559 8483
rect 2958 8480 2964 8492
rect 2547 8452 2964 8480
rect 2547 8449 2559 8452
rect 2501 8443 2559 8449
rect 2958 8440 2964 8452
rect 3016 8440 3022 8492
rect 750 8412 756 8424
rect 711 8384 756 8412
rect 750 8372 756 8384
rect 808 8372 814 8424
rect 3068 8412 3096 8520
rect 3896 8492 3924 8520
rect 5442 8508 5448 8520
rect 5500 8508 5506 8560
rect 5629 8551 5687 8557
rect 5629 8517 5641 8551
rect 5675 8548 5687 8551
rect 5675 8520 6776 8548
rect 5675 8517 5687 8520
rect 5629 8511 5687 8517
rect 6748 8492 6776 8520
rect 8202 8508 8208 8560
rect 8260 8548 8266 8560
rect 9033 8551 9091 8557
rect 9033 8548 9045 8551
rect 8260 8520 9045 8548
rect 8260 8508 8266 8520
rect 9033 8517 9045 8520
rect 9079 8517 9091 8551
rect 9600 8548 9628 8576
rect 9033 8511 9091 8517
rect 9140 8520 9628 8548
rect 9140 8492 9168 8520
rect 10594 8508 10600 8560
rect 10652 8548 10658 8560
rect 10750 8551 10808 8557
rect 10750 8548 10762 8551
rect 10652 8520 10762 8548
rect 10652 8508 10658 8520
rect 10750 8517 10762 8520
rect 10796 8517 10808 8551
rect 10888 8548 10916 8588
rect 10962 8576 10968 8628
rect 11020 8616 11026 8628
rect 11020 8588 14320 8616
rect 11020 8576 11026 8588
rect 12434 8548 12440 8560
rect 10888 8520 12112 8548
rect 10750 8511 10808 8517
rect 3326 8440 3332 8492
rect 3384 8480 3390 8492
rect 3697 8483 3755 8489
rect 3697 8480 3709 8483
rect 3384 8452 3709 8480
rect 3384 8440 3390 8452
rect 3697 8449 3709 8452
rect 3743 8449 3755 8483
rect 3878 8480 3884 8492
rect 3839 8452 3884 8480
rect 3697 8443 3755 8449
rect 3878 8440 3884 8452
rect 3936 8440 3942 8492
rect 4154 8480 4160 8492
rect 4115 8452 4160 8480
rect 4154 8440 4160 8452
rect 4212 8440 4218 8492
rect 5721 8483 5779 8489
rect 5721 8449 5733 8483
rect 5767 8480 5779 8483
rect 6638 8480 6644 8492
rect 5767 8452 6644 8480
rect 5767 8449 5779 8452
rect 5721 8443 5779 8449
rect 6638 8440 6644 8452
rect 6696 8440 6702 8492
rect 6730 8440 6736 8492
rect 6788 8440 6794 8492
rect 7009 8483 7067 8489
rect 7009 8449 7021 8483
rect 7055 8480 7067 8483
rect 8938 8480 8944 8492
rect 7055 8452 8616 8480
rect 8899 8452 8944 8480
rect 7055 8449 7067 8452
rect 7009 8443 7067 8449
rect 3145 8415 3203 8421
rect 3145 8412 3157 8415
rect 3068 8384 3157 8412
rect 3145 8381 3157 8384
rect 3191 8381 3203 8415
rect 3145 8375 3203 8381
rect 3237 8415 3295 8421
rect 3237 8381 3249 8415
rect 3283 8381 3295 8415
rect 3237 8375 3295 8381
rect 3605 8415 3663 8421
rect 3605 8381 3617 8415
rect 3651 8412 3663 8415
rect 3786 8412 3792 8424
rect 3651 8384 3792 8412
rect 3651 8381 3663 8384
rect 3605 8375 3663 8381
rect 3252 8344 3280 8375
rect 3786 8372 3792 8384
rect 3844 8372 3850 8424
rect 6181 8415 6239 8421
rect 6181 8381 6193 8415
rect 6227 8381 6239 8415
rect 6181 8375 6239 8381
rect 6273 8415 6331 8421
rect 6273 8381 6285 8415
rect 6319 8412 6331 8415
rect 6454 8412 6460 8424
rect 6319 8384 6460 8412
rect 6319 8381 6331 8384
rect 6273 8375 6331 8381
rect 3326 8344 3332 8356
rect 3239 8316 3332 8344
rect 3326 8304 3332 8316
rect 3384 8344 3390 8356
rect 4065 8347 4123 8353
rect 4065 8344 4077 8347
rect 3384 8316 4077 8344
rect 3384 8304 3390 8316
rect 4065 8313 4077 8316
rect 4111 8313 4123 8347
rect 6196 8344 6224 8375
rect 6454 8372 6460 8384
rect 6512 8372 6518 8424
rect 6549 8347 6607 8353
rect 6549 8344 6561 8347
rect 6196 8316 6561 8344
rect 4065 8307 4123 8313
rect 6549 8313 6561 8316
rect 6595 8313 6607 8347
rect 7024 8344 7052 8443
rect 8588 8421 8616 8452
rect 8938 8440 8944 8452
rect 8996 8440 9002 8492
rect 9122 8480 9128 8492
rect 9083 8452 9128 8480
rect 9122 8440 9128 8452
rect 9180 8440 9186 8492
rect 9214 8440 9220 8492
rect 9272 8480 9278 8492
rect 9585 8483 9643 8489
rect 9585 8480 9597 8483
rect 9272 8452 9597 8480
rect 9272 8440 9278 8452
rect 9585 8449 9597 8452
rect 9631 8449 9643 8483
rect 9585 8443 9643 8449
rect 10229 8483 10287 8489
rect 10229 8449 10241 8483
rect 10275 8480 10287 8483
rect 10410 8480 10416 8492
rect 10275 8452 10416 8480
rect 10275 8449 10287 8452
rect 10229 8443 10287 8449
rect 10410 8440 10416 8452
rect 10468 8440 10474 8492
rect 10505 8483 10563 8489
rect 10505 8449 10517 8483
rect 10551 8480 10563 8483
rect 11146 8480 11152 8492
rect 10551 8452 11152 8480
rect 10551 8449 10563 8452
rect 10505 8443 10563 8449
rect 11146 8440 11152 8452
rect 11204 8440 11210 8492
rect 11238 8440 11244 8492
rect 11296 8480 11302 8492
rect 12084 8489 12112 8520
rect 12176 8520 12440 8548
rect 12176 8489 12204 8520
rect 12434 8508 12440 8520
rect 12492 8508 12498 8560
rect 12710 8508 12716 8560
rect 12768 8548 12774 8560
rect 13722 8548 13728 8560
rect 12768 8520 13728 8548
rect 12768 8508 12774 8520
rect 13722 8508 13728 8520
rect 13780 8548 13786 8560
rect 14182 8548 14188 8560
rect 13780 8520 14188 8548
rect 13780 8508 13786 8520
rect 14182 8508 14188 8520
rect 14240 8508 14246 8560
rect 14292 8557 14320 8588
rect 14458 8576 14464 8628
rect 14516 8616 14522 8628
rect 14553 8619 14611 8625
rect 14553 8616 14565 8619
rect 14516 8588 14565 8616
rect 14516 8576 14522 8588
rect 14553 8585 14565 8588
rect 14599 8585 14611 8619
rect 14553 8579 14611 8585
rect 14277 8551 14335 8557
rect 14277 8517 14289 8551
rect 14323 8548 14335 8551
rect 15194 8548 15200 8560
rect 14323 8520 15200 8548
rect 14323 8517 14335 8520
rect 14277 8511 14335 8517
rect 15194 8508 15200 8520
rect 15252 8508 15258 8560
rect 15286 8508 15292 8560
rect 15344 8548 15350 8560
rect 16761 8551 16819 8557
rect 16761 8548 16773 8551
rect 15344 8520 16773 8548
rect 15344 8508 15350 8520
rect 16761 8517 16773 8520
rect 16807 8517 16819 8551
rect 16761 8511 16819 8517
rect 16850 8508 16856 8560
rect 16908 8548 16914 8560
rect 16908 8520 17250 8548
rect 16908 8508 16914 8520
rect 12069 8483 12127 8489
rect 11296 8452 12020 8480
rect 11296 8440 11302 8452
rect 7193 8415 7251 8421
rect 7193 8381 7205 8415
rect 7239 8381 7251 8415
rect 7193 8375 7251 8381
rect 8573 8415 8631 8421
rect 8573 8381 8585 8415
rect 8619 8412 8631 8415
rect 8662 8412 8668 8424
rect 8619 8384 8668 8412
rect 8619 8381 8631 8384
rect 8573 8375 8631 8381
rect 6549 8307 6607 8313
rect 6840 8316 7052 8344
rect 6840 8288 6868 8316
rect 2406 8276 2412 8288
rect 2367 8248 2412 8276
rect 2406 8236 2412 8248
rect 2464 8236 2470 8288
rect 3602 8236 3608 8288
rect 3660 8276 3666 8288
rect 3881 8279 3939 8285
rect 3881 8276 3893 8279
rect 3660 8248 3893 8276
rect 3660 8236 3666 8248
rect 3881 8245 3893 8248
rect 3927 8245 3939 8279
rect 3881 8239 3939 8245
rect 6822 8236 6828 8288
rect 6880 8236 6886 8288
rect 7208 8276 7236 8375
rect 8662 8372 8668 8384
rect 8720 8372 8726 8424
rect 8757 8415 8815 8421
rect 8757 8381 8769 8415
rect 8803 8381 8815 8415
rect 8757 8375 8815 8381
rect 8772 8344 8800 8375
rect 9030 8372 9036 8424
rect 9088 8412 9094 8424
rect 9493 8415 9551 8421
rect 9493 8412 9505 8415
rect 9088 8384 9505 8412
rect 9088 8372 9094 8384
rect 9493 8381 9505 8384
rect 9539 8381 9551 8415
rect 9493 8375 9551 8381
rect 9674 8372 9680 8424
rect 9732 8412 9738 8424
rect 9953 8415 10011 8421
rect 9953 8412 9965 8415
rect 9732 8384 9965 8412
rect 9732 8372 9738 8384
rect 9953 8381 9965 8384
rect 9999 8381 10011 8415
rect 11992 8412 12020 8452
rect 12069 8449 12081 8483
rect 12115 8449 12127 8483
rect 12069 8443 12127 8449
rect 12161 8483 12219 8489
rect 12161 8449 12173 8483
rect 12207 8449 12219 8483
rect 12161 8443 12219 8449
rect 12253 8483 12311 8489
rect 12253 8449 12265 8483
rect 12299 8449 12311 8483
rect 12526 8480 12532 8492
rect 12487 8452 12532 8480
rect 12253 8443 12311 8449
rect 12268 8412 12296 8443
rect 12526 8440 12532 8452
rect 12584 8440 12590 8492
rect 13354 8440 13360 8492
rect 13412 8480 13418 8492
rect 14921 8483 14979 8489
rect 14921 8480 14933 8483
rect 13412 8452 14933 8480
rect 13412 8440 13418 8452
rect 14921 8449 14933 8452
rect 14967 8449 14979 8483
rect 14921 8443 14979 8449
rect 15565 8483 15623 8489
rect 15565 8449 15577 8483
rect 15611 8449 15623 8483
rect 15565 8443 15623 8449
rect 13262 8412 13268 8424
rect 11992 8384 13268 8412
rect 9953 8375 10011 8381
rect 13262 8372 13268 8384
rect 13320 8372 13326 8424
rect 13538 8372 13544 8424
rect 13596 8412 13602 8424
rect 15013 8415 15071 8421
rect 15013 8412 15025 8415
rect 13596 8384 15025 8412
rect 13596 8372 13602 8384
rect 15013 8381 15025 8384
rect 15059 8381 15071 8415
rect 15013 8375 15071 8381
rect 15105 8415 15163 8421
rect 15105 8381 15117 8415
rect 15151 8381 15163 8415
rect 15580 8412 15608 8443
rect 16482 8412 16488 8424
rect 15580 8384 16344 8412
rect 16443 8384 16488 8412
rect 15105 8375 15163 8381
rect 8772 8316 10180 8344
rect 10152 8288 10180 8316
rect 11606 8304 11612 8356
rect 11664 8344 11670 8356
rect 11974 8344 11980 8356
rect 11664 8316 11980 8344
rect 11664 8304 11670 8316
rect 11974 8304 11980 8316
rect 12032 8304 12038 8356
rect 12437 8347 12495 8353
rect 12437 8313 12449 8347
rect 12483 8344 12495 8347
rect 13814 8344 13820 8356
rect 12483 8316 13820 8344
rect 12483 8313 12495 8316
rect 12437 8307 12495 8313
rect 13814 8304 13820 8316
rect 13872 8304 13878 8356
rect 14182 8304 14188 8356
rect 14240 8344 14246 8356
rect 14734 8344 14740 8356
rect 14240 8316 14740 8344
rect 14240 8304 14246 8316
rect 14734 8304 14740 8316
rect 14792 8344 14798 8356
rect 15120 8344 15148 8375
rect 14792 8316 15148 8344
rect 15749 8347 15807 8353
rect 14792 8304 14798 8316
rect 15749 8313 15761 8347
rect 15795 8344 15807 8347
rect 15930 8344 15936 8356
rect 15795 8316 15936 8344
rect 15795 8313 15807 8316
rect 15749 8307 15807 8313
rect 15930 8304 15936 8316
rect 15988 8304 15994 8356
rect 16316 8344 16344 8384
rect 16482 8372 16488 8384
rect 16540 8372 16546 8424
rect 16850 8412 16856 8424
rect 16592 8384 16856 8412
rect 16592 8344 16620 8384
rect 16850 8372 16856 8384
rect 16908 8372 16914 8424
rect 17770 8372 17776 8424
rect 17828 8412 17834 8424
rect 18509 8415 18567 8421
rect 18509 8412 18521 8415
rect 17828 8384 18521 8412
rect 17828 8372 17834 8384
rect 18509 8381 18521 8384
rect 18555 8381 18567 8415
rect 18509 8375 18567 8381
rect 16316 8316 16620 8344
rect 8570 8276 8576 8288
rect 7208 8248 8576 8276
rect 8570 8236 8576 8248
rect 8628 8236 8634 8288
rect 10134 8276 10140 8288
rect 10047 8248 10140 8276
rect 10134 8236 10140 8248
rect 10192 8276 10198 8288
rect 10870 8276 10876 8288
rect 10192 8248 10876 8276
rect 10192 8236 10198 8248
rect 10870 8236 10876 8248
rect 10928 8236 10934 8288
rect 11698 8236 11704 8288
rect 11756 8276 11762 8288
rect 11885 8279 11943 8285
rect 11885 8276 11897 8279
rect 11756 8248 11897 8276
rect 11756 8236 11762 8248
rect 11885 8245 11897 8248
rect 11931 8276 11943 8279
rect 12158 8276 12164 8288
rect 11931 8248 12164 8276
rect 11931 8245 11943 8248
rect 11885 8239 11943 8245
rect 12158 8236 12164 8248
rect 12216 8236 12222 8288
rect 13262 8236 13268 8288
rect 13320 8276 13326 8288
rect 18506 8276 18512 8288
rect 13320 8248 18512 8276
rect 13320 8236 13326 8248
rect 18506 8236 18512 8248
rect 18564 8236 18570 8288
rect 0 8186 18860 8208
rect 0 8134 2995 8186
rect 3047 8134 3059 8186
rect 3111 8134 3123 8186
rect 3175 8134 3187 8186
rect 3239 8134 3251 8186
rect 3303 8134 9294 8186
rect 9346 8134 9358 8186
rect 9410 8134 9422 8186
rect 9474 8134 9486 8186
rect 9538 8134 9550 8186
rect 9602 8134 15592 8186
rect 15644 8134 15656 8186
rect 15708 8134 15720 8186
rect 15772 8134 15784 8186
rect 15836 8134 15848 8186
rect 15900 8134 18860 8186
rect 0 8112 18860 8134
rect 750 8032 756 8084
rect 808 8072 814 8084
rect 2225 8075 2283 8081
rect 2225 8072 2237 8075
rect 808 8044 2237 8072
rect 808 8032 814 8044
rect 2225 8041 2237 8044
rect 2271 8041 2283 8075
rect 2225 8035 2283 8041
rect 2314 8032 2320 8084
rect 2372 8072 2378 8084
rect 3326 8072 3332 8084
rect 2372 8044 3188 8072
rect 3287 8044 3332 8072
rect 2372 8032 2378 8044
rect 2133 8007 2191 8013
rect 2133 7973 2145 8007
rect 2179 8004 2191 8007
rect 3050 8004 3056 8016
rect 2179 7976 3056 8004
rect 2179 7973 2191 7976
rect 2133 7967 2191 7973
rect 3050 7964 3056 7976
rect 3108 7964 3114 8016
rect 3160 8013 3188 8044
rect 3326 8032 3332 8044
rect 3384 8032 3390 8084
rect 3786 8032 3792 8084
rect 3844 8072 3850 8084
rect 3881 8075 3939 8081
rect 3881 8072 3893 8075
rect 3844 8044 3893 8072
rect 3844 8032 3850 8044
rect 3881 8041 3893 8044
rect 3927 8041 3939 8075
rect 3881 8035 3939 8041
rect 4154 8032 4160 8084
rect 4212 8072 4218 8084
rect 5077 8075 5135 8081
rect 5077 8072 5089 8075
rect 4212 8044 5089 8072
rect 4212 8032 4218 8044
rect 5077 8041 5089 8044
rect 5123 8041 5135 8075
rect 5077 8035 5135 8041
rect 5534 8032 5540 8084
rect 5592 8072 5598 8084
rect 5997 8075 6055 8081
rect 5997 8072 6009 8075
rect 5592 8044 6009 8072
rect 5592 8032 5598 8044
rect 5997 8041 6009 8044
rect 6043 8072 6055 8075
rect 6454 8072 6460 8084
rect 6043 8044 6460 8072
rect 6043 8041 6055 8044
rect 5997 8035 6055 8041
rect 6454 8032 6460 8044
rect 6512 8032 6518 8084
rect 6549 8075 6607 8081
rect 6549 8041 6561 8075
rect 6595 8072 6607 8075
rect 6822 8072 6828 8084
rect 6595 8044 6828 8072
rect 6595 8041 6607 8044
rect 6549 8035 6607 8041
rect 6822 8032 6828 8044
rect 6880 8032 6886 8084
rect 7009 8075 7067 8081
rect 7009 8041 7021 8075
rect 7055 8072 7067 8075
rect 7282 8072 7288 8084
rect 7055 8044 7288 8072
rect 7055 8041 7067 8044
rect 7009 8035 7067 8041
rect 7282 8032 7288 8044
rect 7340 8032 7346 8084
rect 7834 8032 7840 8084
rect 7892 8072 7898 8084
rect 9766 8072 9772 8084
rect 7892 8044 9772 8072
rect 7892 8032 7898 8044
rect 9766 8032 9772 8044
rect 9824 8032 9830 8084
rect 11054 8032 11060 8084
rect 11112 8072 11118 8084
rect 11425 8075 11483 8081
rect 11425 8072 11437 8075
rect 11112 8044 11437 8072
rect 11112 8032 11118 8044
rect 11425 8041 11437 8044
rect 11471 8041 11483 8075
rect 12526 8072 12532 8084
rect 11425 8035 11483 8041
rect 11532 8044 12532 8072
rect 3145 8007 3203 8013
rect 3145 7973 3157 8007
rect 3191 8004 3203 8007
rect 3191 7976 3924 8004
rect 3191 7973 3203 7976
rect 3145 7967 3203 7973
rect 2317 7939 2375 7945
rect 2317 7905 2329 7939
rect 2363 7936 2375 7939
rect 3694 7936 3700 7948
rect 2363 7908 2820 7936
rect 2363 7905 2375 7908
rect 2317 7899 2375 7905
rect 1765 7871 1823 7877
rect 1765 7837 1777 7871
rect 1811 7837 1823 7871
rect 1765 7831 1823 7837
rect 1780 7800 1808 7831
rect 1854 7828 1860 7880
rect 1912 7868 1918 7880
rect 1949 7871 2007 7877
rect 1949 7868 1961 7871
rect 1912 7840 1961 7868
rect 1912 7828 1918 7840
rect 1949 7837 1961 7840
rect 1995 7837 2007 7871
rect 1949 7831 2007 7837
rect 2060 7871 2118 7877
rect 2060 7837 2072 7871
rect 2106 7868 2118 7871
rect 2406 7868 2412 7880
rect 2106 7840 2412 7868
rect 2106 7837 2118 7840
rect 2060 7831 2118 7837
rect 2148 7800 2176 7840
rect 2406 7828 2412 7840
rect 2464 7828 2470 7880
rect 2682 7868 2688 7880
rect 2643 7840 2688 7868
rect 2682 7828 2688 7840
rect 2740 7828 2746 7880
rect 2792 7877 2820 7908
rect 3252 7908 3700 7936
rect 3252 7877 3280 7908
rect 3694 7896 3700 7908
rect 3752 7896 3758 7948
rect 3896 7936 3924 7976
rect 4246 7964 4252 8016
rect 4304 8004 4310 8016
rect 11532 8004 11560 8044
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 12986 8072 12992 8084
rect 12947 8044 12992 8072
rect 12986 8032 12992 8044
rect 13044 8032 13050 8084
rect 14182 8072 14188 8084
rect 13648 8044 14188 8072
rect 13262 8004 13268 8016
rect 4304 7976 11560 8004
rect 11900 7976 13268 8004
rect 4304 7964 4310 7976
rect 4893 7939 4951 7945
rect 3896 7908 4844 7936
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7868 2835 7871
rect 3237 7871 3295 7877
rect 2823 7840 3096 7868
rect 2823 7837 2835 7840
rect 2777 7831 2835 7837
rect 3068 7800 3096 7840
rect 3237 7837 3249 7871
rect 3283 7837 3295 7871
rect 3602 7868 3608 7880
rect 3563 7840 3608 7868
rect 3237 7831 3295 7837
rect 3602 7828 3608 7840
rect 3660 7828 3666 7880
rect 3789 7871 3847 7877
rect 3789 7837 3801 7871
rect 3835 7837 3847 7871
rect 4062 7868 4068 7880
rect 4023 7840 4068 7868
rect 3789 7831 3847 7837
rect 1780 7772 2176 7800
rect 2746 7772 3004 7800
rect 3068 7772 3556 7800
rect 1949 7735 2007 7741
rect 1949 7701 1961 7735
rect 1995 7732 2007 7735
rect 2314 7732 2320 7744
rect 1995 7704 2320 7732
rect 1995 7701 2007 7704
rect 1949 7695 2007 7701
rect 2314 7692 2320 7704
rect 2372 7692 2378 7744
rect 2498 7692 2504 7744
rect 2556 7732 2562 7744
rect 2746 7732 2774 7772
rect 2976 7741 3004 7772
rect 3528 7741 3556 7772
rect 2556 7704 2774 7732
rect 2961 7735 3019 7741
rect 2556 7692 2562 7704
rect 2961 7701 2973 7735
rect 3007 7701 3019 7735
rect 2961 7695 3019 7701
rect 3513 7735 3571 7741
rect 3513 7701 3525 7735
rect 3559 7701 3571 7735
rect 3804 7732 3832 7831
rect 4062 7828 4068 7840
rect 4120 7828 4126 7880
rect 4249 7871 4307 7877
rect 4157 7849 4215 7855
rect 4157 7815 4169 7849
rect 4203 7815 4215 7849
rect 4249 7837 4261 7871
rect 4295 7868 4307 7871
rect 4338 7868 4344 7880
rect 4295 7840 4344 7868
rect 4295 7837 4307 7840
rect 4249 7831 4307 7837
rect 4338 7828 4344 7840
rect 4396 7828 4402 7880
rect 4816 7877 4844 7908
rect 4893 7905 4905 7939
rect 4939 7936 4951 7939
rect 5721 7939 5779 7945
rect 5721 7936 5733 7939
rect 4939 7908 5733 7936
rect 4939 7905 4951 7908
rect 4893 7899 4951 7905
rect 5721 7905 5733 7908
rect 5767 7936 5779 7939
rect 6362 7936 6368 7948
rect 5767 7908 6224 7936
rect 6323 7908 6368 7936
rect 5767 7905 5779 7908
rect 5721 7899 5779 7905
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7837 4859 7871
rect 4801 7831 4859 7837
rect 4985 7871 5043 7877
rect 4985 7837 4997 7871
rect 5031 7837 5043 7871
rect 4985 7831 5043 7837
rect 5445 7871 5503 7877
rect 5445 7837 5457 7871
rect 5491 7868 5503 7871
rect 5534 7868 5540 7880
rect 5491 7840 5540 7868
rect 5491 7837 5503 7840
rect 5445 7831 5503 7837
rect 4157 7812 4215 7815
rect 4154 7760 4160 7812
rect 4212 7760 4218 7812
rect 5000 7800 5028 7831
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 5902 7868 5908 7880
rect 5863 7840 5908 7868
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 6089 7871 6147 7877
rect 6089 7837 6101 7871
rect 6135 7837 6147 7871
rect 6196 7868 6224 7908
rect 6362 7896 6368 7908
rect 6420 7896 6426 7948
rect 6454 7896 6460 7948
rect 6512 7936 6518 7948
rect 7193 7939 7251 7945
rect 7193 7936 7205 7939
rect 6512 7908 7205 7936
rect 6512 7896 6518 7908
rect 7193 7905 7205 7908
rect 7239 7936 7251 7939
rect 9030 7936 9036 7948
rect 7239 7908 9036 7936
rect 7239 7905 7251 7908
rect 7193 7899 7251 7905
rect 9030 7896 9036 7908
rect 9088 7896 9094 7948
rect 9125 7939 9183 7945
rect 9125 7905 9137 7939
rect 9171 7936 9183 7939
rect 10134 7936 10140 7948
rect 9171 7908 10140 7936
rect 9171 7905 9183 7908
rect 9125 7899 9183 7905
rect 10134 7896 10140 7908
rect 10192 7896 10198 7948
rect 11900 7936 11928 7976
rect 13262 7964 13268 7976
rect 13320 7964 13326 8016
rect 11256 7908 11928 7936
rect 6641 7871 6699 7877
rect 6196 7840 6408 7868
rect 6089 7831 6147 7837
rect 6104 7800 6132 7831
rect 5000 7772 6132 7800
rect 6380 7800 6408 7840
rect 6641 7837 6653 7871
rect 6687 7868 6699 7871
rect 6822 7868 6828 7880
rect 6687 7840 6828 7868
rect 6687 7837 6699 7840
rect 6641 7831 6699 7837
rect 6822 7828 6828 7840
rect 6880 7828 6886 7880
rect 7282 7828 7288 7880
rect 7340 7868 7346 7880
rect 7834 7868 7840 7880
rect 7340 7840 7385 7868
rect 7795 7840 7840 7868
rect 7340 7828 7346 7840
rect 7834 7828 7840 7840
rect 7892 7828 7898 7880
rect 8110 7868 8116 7880
rect 8071 7840 8116 7868
rect 8110 7828 8116 7840
rect 8168 7868 8174 7880
rect 8938 7868 8944 7880
rect 8168 7840 8944 7868
rect 8168 7828 8174 7840
rect 8938 7828 8944 7840
rect 8996 7868 9002 7880
rect 9582 7868 9588 7880
rect 8996 7840 9588 7868
rect 8996 7828 9002 7840
rect 9582 7828 9588 7840
rect 9640 7828 9646 7880
rect 11256 7877 11284 7908
rect 11974 7896 11980 7948
rect 12032 7936 12038 7948
rect 12710 7936 12716 7948
rect 12032 7908 12716 7936
rect 12032 7896 12038 7908
rect 12710 7896 12716 7908
rect 12768 7896 12774 7948
rect 12802 7896 12808 7948
rect 12860 7936 12866 7948
rect 13648 7945 13676 8044
rect 14182 8032 14188 8044
rect 14240 8032 14246 8084
rect 16472 8075 16530 8081
rect 16472 8041 16484 8075
rect 16518 8072 16530 8075
rect 18322 8072 18328 8084
rect 16518 8044 18328 8072
rect 16518 8041 16530 8044
rect 16472 8035 16530 8041
rect 18322 8032 18328 8044
rect 18380 8032 18386 8084
rect 13449 7939 13507 7945
rect 13449 7936 13461 7939
rect 12860 7908 13461 7936
rect 12860 7896 12866 7908
rect 13449 7905 13461 7908
rect 13495 7905 13507 7939
rect 13449 7899 13507 7905
rect 13633 7939 13691 7945
rect 13633 7905 13645 7939
rect 13679 7905 13691 7939
rect 14277 7939 14335 7945
rect 14277 7936 14289 7939
rect 13633 7899 13691 7905
rect 13740 7908 14289 7936
rect 11241 7871 11299 7877
rect 11241 7837 11253 7871
rect 11287 7837 11299 7871
rect 11698 7868 11704 7880
rect 11659 7840 11704 7868
rect 11241 7831 11299 7837
rect 11698 7828 11704 7840
rect 11756 7828 11762 7880
rect 12158 7868 12164 7880
rect 12119 7840 12164 7868
rect 12158 7828 12164 7840
rect 12216 7828 12222 7880
rect 13354 7868 13360 7880
rect 13315 7840 13360 7868
rect 13354 7828 13360 7840
rect 13412 7828 13418 7880
rect 13464 7868 13492 7899
rect 13740 7880 13768 7908
rect 14277 7905 14289 7908
rect 14323 7936 14335 7939
rect 16209 7939 16267 7945
rect 16209 7936 16221 7939
rect 14323 7908 16221 7936
rect 14323 7905 14335 7908
rect 14277 7899 14335 7905
rect 16209 7905 16221 7908
rect 16255 7936 16267 7939
rect 16482 7936 16488 7948
rect 16255 7908 16488 7936
rect 16255 7905 16267 7908
rect 16209 7899 16267 7905
rect 16482 7896 16488 7908
rect 16540 7936 16546 7948
rect 16942 7936 16948 7948
rect 16540 7908 16948 7936
rect 16540 7896 16546 7908
rect 16942 7896 16948 7908
rect 17000 7896 17006 7948
rect 13722 7868 13728 7880
rect 13464 7840 13728 7868
rect 13722 7828 13728 7840
rect 13780 7828 13786 7880
rect 13814 7828 13820 7880
rect 13872 7868 13878 7880
rect 13872 7840 13917 7868
rect 13872 7828 13878 7840
rect 13998 7828 14004 7880
rect 14056 7868 14062 7880
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 14056 7840 14105 7868
rect 14056 7828 14062 7840
rect 14093 7837 14105 7840
rect 14139 7837 14151 7871
rect 14642 7868 14648 7880
rect 14603 7840 14648 7868
rect 14093 7831 14151 7837
rect 14642 7828 14648 7840
rect 14700 7828 14706 7880
rect 16022 7868 16028 7880
rect 15764 7840 16028 7868
rect 7098 7800 7104 7812
rect 6380 7772 7104 7800
rect 4338 7732 4344 7744
rect 3804 7704 4344 7732
rect 3513 7695 3571 7701
rect 4338 7692 4344 7704
rect 4396 7732 4402 7744
rect 4798 7732 4804 7744
rect 4396 7704 4804 7732
rect 4396 7692 4402 7704
rect 4798 7692 4804 7704
rect 4856 7732 4862 7744
rect 5442 7732 5448 7744
rect 4856 7704 5448 7732
rect 4856 7692 4862 7704
rect 5442 7692 5448 7704
rect 5500 7732 5506 7744
rect 5537 7735 5595 7741
rect 5537 7732 5549 7735
rect 5500 7704 5549 7732
rect 5500 7692 5506 7704
rect 5537 7701 5549 7704
rect 5583 7701 5595 7735
rect 6104 7732 6132 7772
rect 7098 7760 7104 7772
rect 7156 7760 7162 7812
rect 7929 7803 7987 7809
rect 7929 7800 7941 7803
rect 7208 7772 7941 7800
rect 6365 7735 6423 7741
rect 6365 7732 6377 7735
rect 6104 7704 6377 7732
rect 5537 7695 5595 7701
rect 6365 7701 6377 7704
rect 6411 7732 6423 7735
rect 6546 7732 6552 7744
rect 6411 7704 6552 7732
rect 6411 7701 6423 7704
rect 6365 7695 6423 7701
rect 6546 7692 6552 7704
rect 6604 7692 6610 7744
rect 6730 7692 6736 7744
rect 6788 7732 6794 7744
rect 7208 7732 7236 7772
rect 7929 7769 7941 7772
rect 7975 7800 7987 7803
rect 9306 7800 9312 7812
rect 7975 7772 9312 7800
rect 7975 7769 7987 7772
rect 7929 7763 7987 7769
rect 9306 7760 9312 7772
rect 9364 7800 9370 7812
rect 9364 7772 11744 7800
rect 9364 7760 9370 7772
rect 6788 7704 7236 7732
rect 7653 7735 7711 7741
rect 6788 7692 6794 7704
rect 7653 7701 7665 7735
rect 7699 7732 7711 7735
rect 7837 7735 7895 7741
rect 7837 7732 7849 7735
rect 7699 7704 7849 7732
rect 7699 7701 7711 7704
rect 7653 7695 7711 7701
rect 7837 7701 7849 7704
rect 7883 7701 7895 7735
rect 7837 7695 7895 7701
rect 8294 7692 8300 7744
rect 8352 7732 8358 7744
rect 8481 7735 8539 7741
rect 8481 7732 8493 7735
rect 8352 7704 8493 7732
rect 8352 7692 8358 7704
rect 8481 7701 8493 7704
rect 8527 7701 8539 7735
rect 8481 7695 8539 7701
rect 8754 7692 8760 7744
rect 8812 7732 8818 7744
rect 8849 7735 8907 7741
rect 8849 7732 8861 7735
rect 8812 7704 8861 7732
rect 8812 7692 8818 7704
rect 8849 7701 8861 7704
rect 8895 7701 8907 7735
rect 8849 7695 8907 7701
rect 8941 7735 8999 7741
rect 8941 7701 8953 7735
rect 8987 7732 8999 7735
rect 9398 7732 9404 7744
rect 8987 7704 9404 7732
rect 8987 7701 8999 7704
rect 8941 7695 8999 7701
rect 9398 7692 9404 7704
rect 9456 7692 9462 7744
rect 9950 7732 9956 7744
rect 9911 7704 9956 7732
rect 9950 7692 9956 7704
rect 10008 7692 10014 7744
rect 11716 7732 11744 7772
rect 11790 7760 11796 7812
rect 11848 7800 11854 7812
rect 11885 7803 11943 7809
rect 11885 7800 11897 7803
rect 11848 7772 11897 7800
rect 11848 7760 11854 7772
rect 11885 7769 11897 7772
rect 11931 7769 11943 7803
rect 13909 7803 13967 7809
rect 13909 7800 13921 7803
rect 11885 7763 11943 7769
rect 12728 7772 13921 7800
rect 12728 7732 12756 7772
rect 13909 7769 13921 7772
rect 13955 7769 13967 7803
rect 13909 7763 13967 7769
rect 11716 7704 12756 7732
rect 12805 7735 12863 7741
rect 12805 7701 12817 7735
rect 12851 7732 12863 7735
rect 13078 7732 13084 7744
rect 12851 7704 13084 7732
rect 12851 7701 12863 7704
rect 12805 7695 12863 7701
rect 13078 7692 13084 7704
rect 13136 7692 13142 7744
rect 13814 7732 13820 7744
rect 13775 7704 13820 7732
rect 13814 7692 13820 7704
rect 13872 7692 13878 7744
rect 14274 7692 14280 7744
rect 14332 7732 14338 7744
rect 15028 7732 15056 7786
rect 15286 7732 15292 7744
rect 14332 7704 15292 7732
rect 14332 7692 14338 7704
rect 15286 7692 15292 7704
rect 15344 7732 15350 7744
rect 15764 7732 15792 7840
rect 16022 7828 16028 7840
rect 16080 7828 16086 7880
rect 18509 7871 18567 7877
rect 18509 7837 18521 7871
rect 18555 7868 18567 7871
rect 18598 7868 18604 7880
rect 18555 7840 18604 7868
rect 18555 7837 18567 7840
rect 18509 7831 18567 7837
rect 18598 7828 18604 7840
rect 18656 7828 18662 7880
rect 16040 7800 16068 7828
rect 16454 7800 16620 7810
rect 16758 7800 16764 7812
rect 16040 7782 16764 7800
rect 16040 7772 16482 7782
rect 16592 7772 16764 7782
rect 16758 7760 16764 7772
rect 16816 7800 16822 7812
rect 16816 7772 16974 7800
rect 16816 7760 16822 7772
rect 15344 7704 15792 7732
rect 16071 7735 16129 7741
rect 15344 7692 15350 7704
rect 16071 7701 16083 7735
rect 16117 7732 16129 7735
rect 16390 7732 16396 7744
rect 16117 7704 16396 7732
rect 16117 7701 16129 7704
rect 16071 7695 16129 7701
rect 16390 7692 16396 7704
rect 16448 7692 16454 7744
rect 17957 7735 18015 7741
rect 17957 7701 17969 7735
rect 18003 7732 18015 7735
rect 18138 7732 18144 7744
rect 18003 7704 18144 7732
rect 18003 7701 18015 7704
rect 17957 7695 18015 7701
rect 18138 7692 18144 7704
rect 18196 7692 18202 7744
rect 18230 7692 18236 7744
rect 18288 7732 18294 7744
rect 18325 7735 18383 7741
rect 18325 7732 18337 7735
rect 18288 7704 18337 7732
rect 18288 7692 18294 7704
rect 18325 7701 18337 7704
rect 18371 7701 18383 7735
rect 18325 7695 18383 7701
rect 0 7642 18860 7664
rect 0 7590 6144 7642
rect 6196 7590 6208 7642
rect 6260 7590 6272 7642
rect 6324 7590 6336 7642
rect 6388 7590 6400 7642
rect 6452 7590 12443 7642
rect 12495 7590 12507 7642
rect 12559 7590 12571 7642
rect 12623 7590 12635 7642
rect 12687 7590 12699 7642
rect 12751 7590 18860 7642
rect 0 7568 18860 7590
rect 1854 7488 1860 7540
rect 1912 7528 1918 7540
rect 2593 7531 2651 7537
rect 2593 7528 2605 7531
rect 1912 7500 2605 7528
rect 1912 7488 1918 7500
rect 2593 7497 2605 7500
rect 2639 7497 2651 7531
rect 2593 7491 2651 7497
rect 3050 7488 3056 7540
rect 3108 7528 3114 7540
rect 3513 7531 3571 7537
rect 3513 7528 3525 7531
rect 3108 7500 3525 7528
rect 3108 7488 3114 7500
rect 3513 7497 3525 7500
rect 3559 7497 3571 7531
rect 3513 7491 3571 7497
rect 4062 7488 4068 7540
rect 4120 7528 4126 7540
rect 4709 7531 4767 7537
rect 4709 7528 4721 7531
rect 4120 7500 4721 7528
rect 4120 7488 4126 7500
rect 4709 7497 4721 7500
rect 4755 7528 4767 7531
rect 5902 7528 5908 7540
rect 4755 7500 5908 7528
rect 4755 7497 4767 7500
rect 4709 7491 4767 7497
rect 2498 7460 2504 7472
rect 2148 7432 2504 7460
rect 566 7392 572 7404
rect 527 7364 572 7392
rect 566 7352 572 7364
rect 624 7352 630 7404
rect 1946 7352 1952 7404
rect 2004 7352 2010 7404
rect 845 7327 903 7333
rect 845 7293 857 7327
rect 891 7324 903 7327
rect 2148 7324 2176 7432
rect 2498 7420 2504 7432
rect 2556 7420 2562 7472
rect 2866 7420 2872 7472
rect 2924 7420 2930 7472
rect 3973 7463 4031 7469
rect 3973 7429 3985 7463
rect 4019 7460 4031 7463
rect 4246 7460 4252 7472
rect 4019 7432 4252 7460
rect 4019 7429 4031 7432
rect 3973 7423 4031 7429
rect 4246 7420 4252 7432
rect 4304 7420 4310 7472
rect 2682 7392 2688 7404
rect 2332 7364 2688 7392
rect 2332 7333 2360 7364
rect 2682 7352 2688 7364
rect 2740 7392 2746 7404
rect 2777 7395 2835 7401
rect 2777 7392 2789 7395
rect 2740 7364 2789 7392
rect 2740 7352 2746 7364
rect 2777 7361 2789 7364
rect 2823 7361 2835 7395
rect 2884 7392 2912 7420
rect 2961 7395 3019 7401
rect 2961 7392 2973 7395
rect 2884 7364 2973 7392
rect 2777 7355 2835 7361
rect 2961 7361 2973 7364
rect 3007 7361 3019 7395
rect 4798 7392 4804 7404
rect 4759 7364 4804 7392
rect 2961 7355 3019 7361
rect 4798 7352 4804 7364
rect 4856 7352 4862 7404
rect 4908 7401 4936 7500
rect 5902 7488 5908 7500
rect 5960 7528 5966 7540
rect 6822 7528 6828 7540
rect 5960 7500 6132 7528
rect 5960 7488 5966 7500
rect 6104 7469 6132 7500
rect 6196 7500 6828 7528
rect 6089 7463 6147 7469
rect 5000 7432 5580 7460
rect 4893 7395 4951 7401
rect 4893 7361 4905 7395
rect 4939 7361 4951 7395
rect 4893 7355 4951 7361
rect 891 7296 2176 7324
rect 2317 7327 2375 7333
rect 891 7293 903 7296
rect 845 7287 903 7293
rect 2317 7293 2329 7327
rect 2363 7293 2375 7327
rect 2317 7287 2375 7293
rect 2869 7327 2927 7333
rect 2869 7293 2881 7327
rect 2915 7324 2927 7327
rect 5000 7324 5028 7432
rect 5552 7401 5580 7432
rect 6089 7429 6101 7463
rect 6135 7429 6147 7463
rect 6089 7423 6147 7429
rect 5077 7395 5135 7401
rect 5077 7361 5089 7395
rect 5123 7361 5135 7395
rect 5077 7355 5135 7361
rect 5537 7395 5595 7401
rect 5537 7361 5549 7395
rect 5583 7361 5595 7395
rect 5537 7355 5595 7361
rect 2915 7296 5028 7324
rect 2915 7293 2927 7296
rect 2869 7287 2927 7293
rect 1946 7216 1952 7268
rect 2004 7256 2010 7268
rect 2590 7256 2596 7268
rect 2004 7228 2596 7256
rect 2004 7216 2010 7228
rect 2590 7216 2596 7228
rect 2648 7216 2654 7268
rect 3697 7259 3755 7265
rect 3697 7225 3709 7259
rect 3743 7256 3755 7259
rect 4154 7256 4160 7268
rect 3743 7228 4160 7256
rect 3743 7225 3755 7228
rect 3697 7219 3755 7225
rect 4154 7216 4160 7228
rect 4212 7216 4218 7268
rect 5092 7256 5120 7355
rect 5626 7352 5632 7404
rect 5684 7392 5690 7404
rect 5905 7395 5963 7401
rect 5684 7364 5729 7392
rect 5684 7352 5690 7364
rect 5905 7361 5917 7395
rect 5951 7392 5963 7395
rect 6196 7392 6224 7500
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 7190 7528 7196 7540
rect 7151 7500 7196 7528
rect 7190 7488 7196 7500
rect 7248 7488 7254 7540
rect 9950 7528 9956 7540
rect 8588 7500 9956 7528
rect 6457 7463 6515 7469
rect 6457 7429 6469 7463
rect 6503 7460 6515 7463
rect 6546 7460 6552 7472
rect 6503 7432 6552 7460
rect 6503 7429 6515 7432
rect 6457 7423 6515 7429
rect 6546 7420 6552 7432
rect 6604 7420 6610 7472
rect 6730 7460 6736 7472
rect 6691 7432 6736 7460
rect 6730 7420 6736 7432
rect 6788 7420 6794 7472
rect 8294 7460 8300 7472
rect 8255 7432 8300 7460
rect 8294 7420 8300 7432
rect 8352 7420 8358 7472
rect 5951 7364 6224 7392
rect 6273 7395 6331 7401
rect 5951 7361 5963 7364
rect 5905 7355 5963 7361
rect 6273 7361 6285 7395
rect 6319 7392 6331 7395
rect 6748 7392 6776 7420
rect 6319 7364 6776 7392
rect 6917 7395 6975 7401
rect 6319 7361 6331 7364
rect 6273 7355 6331 7361
rect 6917 7361 6929 7395
rect 6963 7361 6975 7395
rect 6917 7355 6975 7361
rect 6638 7324 6644 7336
rect 6599 7296 6644 7324
rect 6638 7284 6644 7296
rect 6696 7284 6702 7336
rect 5721 7259 5779 7265
rect 5721 7256 5733 7259
rect 5092 7228 5733 7256
rect 5721 7225 5733 7228
rect 5767 7256 5779 7259
rect 5994 7256 6000 7268
rect 5767 7228 6000 7256
rect 5767 7225 5779 7228
rect 5721 7219 5779 7225
rect 5994 7216 6000 7228
rect 6052 7216 6058 7268
rect 4982 7188 4988 7200
rect 4943 7160 4988 7188
rect 4982 7148 4988 7160
rect 5040 7148 5046 7200
rect 5813 7191 5871 7197
rect 5813 7157 5825 7191
rect 5859 7188 5871 7191
rect 5902 7188 5908 7200
rect 5859 7160 5908 7188
rect 5859 7157 5871 7160
rect 5813 7151 5871 7157
rect 5902 7148 5908 7160
rect 5960 7148 5966 7200
rect 6086 7148 6092 7200
rect 6144 7188 6150 7200
rect 6932 7188 6960 7355
rect 7006 7352 7012 7404
rect 7064 7392 7070 7404
rect 7285 7395 7343 7401
rect 7064 7364 7109 7392
rect 7064 7352 7070 7364
rect 7285 7361 7297 7395
rect 7331 7392 7343 7395
rect 8588 7392 8616 7500
rect 9950 7488 9956 7500
rect 10008 7528 10014 7540
rect 14182 7528 14188 7540
rect 10008 7500 14188 7528
rect 10008 7488 10014 7500
rect 14182 7488 14188 7500
rect 14240 7488 14246 7540
rect 8754 7460 8760 7472
rect 8715 7432 8760 7460
rect 8754 7420 8760 7432
rect 8812 7420 8818 7472
rect 9122 7460 9128 7472
rect 9035 7432 9128 7460
rect 9122 7420 9128 7432
rect 9180 7460 9186 7472
rect 9180 7432 11652 7460
rect 9180 7420 9186 7432
rect 8938 7392 8944 7404
rect 7331 7364 8616 7392
rect 8899 7364 8944 7392
rect 7331 7361 7343 7364
rect 7285 7355 7343 7361
rect 8938 7352 8944 7364
rect 8996 7352 9002 7404
rect 9306 7392 9312 7404
rect 9267 7364 9312 7392
rect 9306 7352 9312 7364
rect 9364 7352 9370 7404
rect 9401 7395 9459 7401
rect 9401 7361 9413 7395
rect 9447 7392 9459 7395
rect 9766 7392 9772 7404
rect 9447 7364 9772 7392
rect 9447 7361 9459 7364
rect 9401 7355 9459 7361
rect 9766 7352 9772 7364
rect 9824 7352 9830 7404
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7361 9919 7395
rect 9861 7355 9919 7361
rect 8386 7324 8392 7336
rect 8347 7296 8392 7324
rect 8386 7284 8392 7296
rect 8444 7284 8450 7336
rect 8570 7324 8576 7336
rect 8531 7296 8576 7324
rect 8570 7284 8576 7296
rect 8628 7284 8634 7336
rect 9214 7284 9220 7336
rect 9272 7284 9278 7336
rect 9582 7284 9588 7336
rect 9640 7324 9646 7336
rect 9640 7296 9812 7324
rect 9640 7284 9646 7296
rect 7282 7216 7288 7268
rect 7340 7256 7346 7268
rect 7929 7259 7987 7265
rect 7929 7256 7941 7259
rect 7340 7228 7941 7256
rect 7340 7216 7346 7228
rect 7929 7225 7941 7228
rect 7975 7225 7987 7259
rect 9232 7256 9260 7284
rect 9493 7259 9551 7265
rect 9493 7256 9505 7259
rect 9232 7228 9505 7256
rect 7929 7219 7987 7225
rect 9493 7225 9505 7228
rect 9539 7225 9551 7259
rect 9674 7256 9680 7268
rect 9493 7219 9551 7225
rect 9646 7216 9680 7256
rect 9732 7216 9738 7268
rect 6144 7160 6960 7188
rect 7009 7191 7067 7197
rect 6144 7148 6150 7160
rect 7009 7157 7021 7191
rect 7055 7188 7067 7191
rect 8202 7188 8208 7200
rect 7055 7160 8208 7188
rect 7055 7157 7067 7160
rect 7009 7151 7067 7157
rect 8202 7148 8208 7160
rect 8260 7148 8266 7200
rect 9401 7191 9459 7197
rect 9401 7157 9413 7191
rect 9447 7188 9459 7191
rect 9646 7188 9674 7216
rect 9447 7160 9674 7188
rect 9784 7188 9812 7296
rect 9876 7256 9904 7355
rect 9950 7352 9956 7404
rect 10008 7392 10014 7404
rect 11624 7401 11652 7432
rect 12710 7420 12716 7472
rect 12768 7420 12774 7472
rect 13722 7420 13728 7472
rect 13780 7460 13786 7472
rect 14461 7463 14519 7469
rect 14461 7460 14473 7463
rect 13780 7432 14473 7460
rect 13780 7420 13786 7432
rect 14461 7429 14473 7432
rect 14507 7429 14519 7463
rect 15194 7460 15200 7472
rect 15155 7432 15200 7460
rect 14461 7423 14519 7429
rect 15194 7420 15200 7432
rect 15252 7420 15258 7472
rect 16758 7420 16764 7472
rect 16816 7460 16822 7472
rect 18138 7460 18144 7472
rect 16816 7432 16974 7460
rect 18099 7432 18144 7460
rect 16816 7420 16822 7432
rect 18138 7420 18144 7432
rect 18196 7420 18202 7472
rect 10781 7395 10839 7401
rect 10008 7364 10272 7392
rect 10008 7352 10014 7364
rect 10134 7324 10140 7336
rect 10095 7296 10140 7324
rect 10134 7284 10140 7296
rect 10192 7284 10198 7336
rect 10244 7324 10272 7364
rect 10781 7361 10793 7395
rect 10827 7392 10839 7395
rect 11609 7395 11667 7401
rect 10827 7364 11284 7392
rect 10827 7361 10839 7364
rect 10781 7355 10839 7361
rect 10873 7327 10931 7333
rect 10873 7324 10885 7327
rect 10244 7296 10885 7324
rect 10873 7293 10885 7296
rect 10919 7293 10931 7327
rect 10873 7287 10931 7293
rect 10962 7284 10968 7336
rect 11020 7324 11026 7336
rect 11020 7296 11065 7324
rect 11020 7284 11026 7296
rect 11256 7265 11284 7364
rect 11609 7361 11621 7395
rect 11655 7361 11667 7395
rect 14090 7392 14096 7404
rect 14051 7364 14096 7392
rect 11609 7355 11667 7361
rect 14090 7352 14096 7364
rect 14148 7352 14154 7404
rect 14737 7395 14795 7401
rect 14737 7361 14749 7395
rect 14783 7392 14795 7395
rect 15933 7395 15991 7401
rect 15933 7392 15945 7395
rect 14783 7364 15608 7392
rect 14783 7361 14795 7364
rect 14737 7355 14795 7361
rect 11517 7327 11575 7333
rect 11517 7293 11529 7327
rect 11563 7293 11575 7327
rect 11517 7287 11575 7293
rect 10413 7259 10471 7265
rect 10413 7256 10425 7259
rect 9876 7228 10425 7256
rect 10413 7225 10425 7228
rect 10459 7225 10471 7259
rect 10413 7219 10471 7225
rect 11241 7259 11299 7265
rect 11241 7225 11253 7259
rect 11287 7225 11299 7259
rect 11241 7219 11299 7225
rect 11532 7188 11560 7287
rect 11882 7284 11888 7336
rect 11940 7324 11946 7336
rect 11977 7327 12035 7333
rect 11977 7324 11989 7327
rect 11940 7296 11989 7324
rect 11940 7284 11946 7296
rect 11977 7293 11989 7296
rect 12023 7293 12035 7327
rect 11977 7287 12035 7293
rect 12345 7327 12403 7333
rect 12345 7293 12357 7327
rect 12391 7324 12403 7327
rect 13814 7324 13820 7336
rect 12391 7296 13820 7324
rect 12391 7293 12403 7296
rect 12345 7287 12403 7293
rect 13814 7284 13820 7296
rect 13872 7284 13878 7336
rect 13998 7324 14004 7336
rect 13959 7296 14004 7324
rect 13998 7284 14004 7296
rect 14056 7284 14062 7336
rect 14645 7327 14703 7333
rect 14645 7324 14657 7327
rect 14108 7296 14657 7324
rect 14108 7256 14136 7296
rect 14645 7293 14657 7296
rect 14691 7293 14703 7327
rect 14645 7287 14703 7293
rect 13096 7228 14136 7256
rect 9784 7160 11560 7188
rect 9447 7157 9459 7160
rect 9401 7151 9459 7157
rect 12526 7148 12532 7200
rect 12584 7188 12590 7200
rect 13096 7188 13124 7228
rect 14274 7216 14280 7268
rect 14332 7256 14338 7268
rect 15580 7265 15608 7364
rect 15672 7364 15945 7392
rect 15013 7259 15071 7265
rect 15013 7256 15025 7259
rect 14332 7228 15025 7256
rect 14332 7216 14338 7228
rect 15013 7225 15025 7228
rect 15059 7225 15071 7259
rect 15013 7219 15071 7225
rect 15565 7259 15623 7265
rect 15565 7225 15577 7259
rect 15611 7225 15623 7259
rect 15565 7219 15623 7225
rect 12584 7160 13124 7188
rect 13771 7191 13829 7197
rect 12584 7148 12590 7160
rect 13771 7157 13783 7191
rect 13817 7188 13829 7191
rect 14918 7188 14924 7200
rect 13817 7160 14924 7188
rect 13817 7157 13829 7160
rect 13771 7151 13829 7157
rect 14918 7148 14924 7160
rect 14976 7188 14982 7200
rect 15672 7188 15700 7364
rect 15933 7361 15945 7364
rect 15979 7361 15991 7395
rect 15933 7355 15991 7361
rect 16022 7324 16028 7336
rect 15983 7296 16028 7324
rect 16022 7284 16028 7296
rect 16080 7284 16086 7336
rect 16393 7327 16451 7333
rect 16393 7293 16405 7327
rect 16439 7324 16451 7327
rect 16666 7324 16672 7336
rect 16439 7296 16672 7324
rect 16439 7293 16451 7296
rect 16393 7287 16451 7293
rect 16666 7284 16672 7296
rect 16724 7284 16730 7336
rect 18417 7327 18475 7333
rect 18417 7324 18429 7327
rect 18340 7296 18429 7324
rect 14976 7160 15700 7188
rect 14976 7148 14982 7160
rect 16942 7148 16948 7200
rect 17000 7188 17006 7200
rect 18340 7188 18368 7296
rect 18417 7293 18429 7296
rect 18463 7293 18475 7327
rect 18417 7287 18475 7293
rect 17000 7160 18368 7188
rect 17000 7148 17006 7160
rect 0 7098 18860 7120
rect 0 7046 2995 7098
rect 3047 7046 3059 7098
rect 3111 7046 3123 7098
rect 3175 7046 3187 7098
rect 3239 7046 3251 7098
rect 3303 7046 9294 7098
rect 9346 7046 9358 7098
rect 9410 7046 9422 7098
rect 9474 7046 9486 7098
rect 9538 7046 9550 7098
rect 9602 7046 15592 7098
rect 15644 7046 15656 7098
rect 15708 7046 15720 7098
rect 15772 7046 15784 7098
rect 15836 7046 15848 7098
rect 15900 7046 18860 7098
rect 0 7024 18860 7046
rect 5442 6944 5448 6996
rect 5500 6984 5506 6996
rect 5500 6956 6592 6984
rect 5500 6944 5506 6956
rect 6564 6928 6592 6956
rect 7006 6944 7012 6996
rect 7064 6984 7070 6996
rect 7193 6987 7251 6993
rect 7193 6984 7205 6987
rect 7064 6956 7205 6984
rect 7064 6944 7070 6956
rect 7193 6953 7205 6956
rect 7239 6953 7251 6987
rect 8570 6984 8576 6996
rect 7193 6947 7251 6953
rect 7300 6956 8576 6984
rect 3602 6876 3608 6928
rect 3660 6916 3666 6928
rect 3789 6919 3847 6925
rect 3789 6916 3801 6919
rect 3660 6888 3801 6916
rect 3660 6876 3666 6888
rect 3789 6885 3801 6888
rect 3835 6916 3847 6919
rect 5997 6919 6055 6925
rect 3835 6888 5304 6916
rect 3835 6885 3847 6888
rect 3789 6879 3847 6885
rect 3145 6851 3203 6857
rect 3145 6817 3157 6851
rect 3191 6848 3203 6851
rect 3329 6851 3387 6857
rect 3329 6848 3341 6851
rect 3191 6820 3341 6848
rect 3191 6817 3203 6820
rect 3145 6811 3203 6817
rect 3329 6817 3341 6820
rect 3375 6817 3387 6851
rect 3973 6851 4031 6857
rect 3973 6848 3985 6851
rect 3329 6811 3387 6817
rect 3436 6820 3985 6848
rect 3050 6780 3056 6792
rect 3011 6752 3056 6780
rect 3050 6740 3056 6752
rect 3108 6740 3114 6792
rect 3237 6783 3295 6789
rect 3237 6749 3249 6783
rect 3283 6780 3295 6783
rect 3436 6780 3464 6820
rect 3973 6817 3985 6820
rect 4019 6848 4031 6851
rect 4982 6848 4988 6860
rect 4019 6820 4988 6848
rect 4019 6817 4031 6820
rect 3973 6811 4031 6817
rect 4982 6808 4988 6820
rect 5040 6808 5046 6860
rect 3283 6752 3464 6780
rect 3513 6783 3571 6789
rect 3283 6749 3295 6752
rect 3237 6743 3295 6749
rect 3513 6749 3525 6783
rect 3559 6749 3571 6783
rect 3513 6743 3571 6749
rect 3329 6715 3387 6721
rect 3329 6712 3341 6715
rect 2746 6684 3341 6712
rect 1670 6604 1676 6656
rect 1728 6644 1734 6656
rect 2746 6644 2774 6684
rect 3329 6681 3341 6684
rect 3375 6681 3387 6715
rect 3329 6675 3387 6681
rect 1728 6616 2774 6644
rect 1728 6604 1734 6616
rect 3234 6604 3240 6656
rect 3292 6644 3298 6656
rect 3528 6644 3556 6743
rect 3602 6740 3608 6792
rect 3660 6780 3666 6792
rect 3878 6780 3884 6792
rect 3660 6752 3705 6780
rect 3839 6752 3884 6780
rect 3660 6740 3666 6752
rect 3878 6740 3884 6752
rect 3936 6740 3942 6792
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6780 4307 6783
rect 5074 6780 5080 6792
rect 4295 6752 5080 6780
rect 4295 6749 4307 6752
rect 4249 6743 4307 6749
rect 4264 6712 4292 6743
rect 5074 6740 5080 6752
rect 5132 6740 5138 6792
rect 5276 6789 5304 6888
rect 5997 6885 6009 6919
rect 6043 6916 6055 6919
rect 6086 6916 6092 6928
rect 6043 6888 6092 6916
rect 6043 6885 6055 6888
rect 5997 6879 6055 6885
rect 6086 6876 6092 6888
rect 6144 6876 6150 6928
rect 6546 6876 6552 6928
rect 6604 6916 6610 6928
rect 7300 6916 7328 6956
rect 8570 6944 8576 6956
rect 8628 6984 8634 6996
rect 8628 6956 8984 6984
rect 8628 6944 8634 6956
rect 6604 6888 7328 6916
rect 8956 6916 8984 6956
rect 9766 6944 9772 6996
rect 9824 6984 9830 6996
rect 10502 6984 10508 6996
rect 9824 6956 10508 6984
rect 9824 6944 9830 6956
rect 10502 6944 10508 6956
rect 10560 6984 10566 6996
rect 12342 6984 12348 6996
rect 10560 6956 12348 6984
rect 10560 6944 10566 6956
rect 12342 6944 12348 6956
rect 12400 6944 12406 6996
rect 13354 6944 13360 6996
rect 13412 6984 13418 6996
rect 13725 6987 13783 6993
rect 13725 6984 13737 6987
rect 13412 6956 13737 6984
rect 13412 6944 13418 6956
rect 13725 6953 13737 6956
rect 13771 6953 13783 6987
rect 13725 6947 13783 6953
rect 13817 6987 13875 6993
rect 13817 6953 13829 6987
rect 13863 6984 13875 6987
rect 14090 6984 14096 6996
rect 13863 6956 14096 6984
rect 13863 6953 13875 6956
rect 13817 6947 13875 6953
rect 14090 6944 14096 6956
rect 14148 6944 14154 6996
rect 15102 6984 15108 6996
rect 14200 6956 15108 6984
rect 10134 6916 10140 6928
rect 8956 6888 10140 6916
rect 6604 6876 6610 6888
rect 5350 6808 5356 6860
rect 5408 6848 5414 6860
rect 7024 6857 7052 6888
rect 10134 6876 10140 6888
rect 10192 6876 10198 6928
rect 12360 6888 13400 6916
rect 5445 6851 5503 6857
rect 5445 6848 5457 6851
rect 5408 6820 5457 6848
rect 5408 6808 5414 6820
rect 5445 6817 5457 6820
rect 5491 6817 5503 6851
rect 5445 6811 5503 6817
rect 7009 6851 7067 6857
rect 7009 6817 7021 6851
rect 7055 6817 7067 6851
rect 7009 6811 7067 6817
rect 7098 6808 7104 6860
rect 7156 6848 7162 6860
rect 8202 6848 8208 6860
rect 7156 6820 7236 6848
rect 8163 6820 8208 6848
rect 7156 6808 7162 6820
rect 5261 6783 5319 6789
rect 5261 6749 5273 6783
rect 5307 6749 5319 6783
rect 5810 6780 5816 6792
rect 5771 6752 5816 6780
rect 5261 6743 5319 6749
rect 5810 6740 5816 6752
rect 5868 6740 5874 6792
rect 5994 6780 6000 6792
rect 5955 6752 6000 6780
rect 5994 6740 6000 6752
rect 6052 6740 6058 6792
rect 7208 6789 7236 6820
rect 8202 6808 8208 6820
rect 8260 6808 8266 6860
rect 8478 6808 8484 6860
rect 8536 6848 8542 6860
rect 9631 6851 9689 6857
rect 9631 6848 9643 6851
rect 8536 6820 9643 6848
rect 8536 6808 8542 6820
rect 9631 6817 9643 6820
rect 9677 6848 9689 6851
rect 11606 6848 11612 6860
rect 9677 6820 11612 6848
rect 9677 6817 9689 6820
rect 9631 6811 9689 6817
rect 11606 6808 11612 6820
rect 11664 6808 11670 6860
rect 11974 6848 11980 6860
rect 11935 6820 11980 6848
rect 11974 6808 11980 6820
rect 12032 6848 12038 6860
rect 12360 6848 12388 6888
rect 12032 6820 12388 6848
rect 12032 6808 12038 6820
rect 12434 6808 12440 6860
rect 12492 6848 12498 6860
rect 12529 6851 12587 6857
rect 12529 6848 12541 6851
rect 12492 6820 12541 6848
rect 12492 6808 12498 6820
rect 12529 6817 12541 6820
rect 12575 6817 12587 6851
rect 12529 6811 12587 6817
rect 12986 6808 12992 6860
rect 13044 6848 13050 6860
rect 13081 6851 13139 6857
rect 13081 6848 13093 6851
rect 13044 6820 13093 6848
rect 13044 6808 13050 6820
rect 13081 6817 13093 6820
rect 13127 6817 13139 6851
rect 13081 6811 13139 6817
rect 13170 6808 13176 6860
rect 13228 6848 13234 6860
rect 13265 6851 13323 6857
rect 13265 6848 13277 6851
rect 13228 6820 13277 6848
rect 13228 6808 13234 6820
rect 13265 6817 13277 6820
rect 13311 6817 13323 6851
rect 13372 6848 13400 6888
rect 14200 6848 14228 6956
rect 15102 6944 15108 6956
rect 15160 6984 15166 6996
rect 15197 6987 15255 6993
rect 15197 6984 15209 6987
rect 15160 6956 15209 6984
rect 15160 6944 15166 6956
rect 15197 6953 15209 6956
rect 15243 6953 15255 6987
rect 15197 6947 15255 6953
rect 14458 6857 14464 6860
rect 13372 6820 14228 6848
rect 14415 6851 14464 6857
rect 13265 6811 13323 6817
rect 14415 6817 14427 6851
rect 14461 6817 14464 6851
rect 14415 6811 14464 6817
rect 14458 6808 14464 6811
rect 14516 6808 14522 6860
rect 16022 6848 16028 6860
rect 14660 6837 16028 6848
rect 14568 6820 16028 6837
rect 14568 6809 14688 6820
rect 6273 6783 6331 6789
rect 6273 6749 6285 6783
rect 6319 6780 6331 6783
rect 7193 6783 7251 6789
rect 6319 6752 7144 6780
rect 6319 6749 6331 6752
rect 6273 6743 6331 6749
rect 4080 6684 4292 6712
rect 4080 6644 4108 6684
rect 5442 6672 5448 6724
rect 5500 6712 5506 6724
rect 7116 6712 7144 6752
rect 7193 6749 7205 6783
rect 7239 6749 7251 6783
rect 7834 6780 7840 6792
rect 7795 6752 7840 6780
rect 7193 6743 7251 6749
rect 7834 6740 7840 6752
rect 7892 6740 7898 6792
rect 9861 6783 9919 6789
rect 9861 6749 9873 6783
rect 9907 6780 9919 6783
rect 10134 6780 10140 6792
rect 9907 6752 10140 6780
rect 9907 6749 9919 6752
rect 9861 6743 9919 6749
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 11882 6740 11888 6792
rect 11940 6780 11946 6792
rect 12069 6783 12127 6789
rect 11940 6752 11985 6780
rect 11940 6740 11946 6752
rect 12069 6749 12081 6783
rect 12115 6749 12127 6783
rect 12069 6743 12127 6749
rect 7285 6715 7343 6721
rect 7285 6712 7297 6715
rect 5500 6684 6408 6712
rect 7116 6684 7297 6712
rect 5500 6672 5506 6684
rect 3292 6616 4108 6644
rect 3292 6604 3298 6616
rect 4246 6604 4252 6656
rect 4304 6644 4310 6656
rect 4893 6647 4951 6653
rect 4893 6644 4905 6647
rect 4304 6616 4905 6644
rect 4304 6604 4310 6616
rect 4893 6613 4905 6616
rect 4939 6613 4951 6647
rect 4893 6607 4951 6613
rect 5353 6647 5411 6653
rect 5353 6613 5365 6647
rect 5399 6644 5411 6647
rect 5626 6644 5632 6656
rect 5399 6616 5632 6644
rect 5399 6613 5411 6616
rect 5353 6607 5411 6613
rect 5626 6604 5632 6616
rect 5684 6604 5690 6656
rect 6380 6653 6408 6684
rect 7285 6681 7297 6684
rect 7331 6681 7343 6715
rect 7285 6675 7343 6681
rect 6365 6647 6423 6653
rect 6365 6613 6377 6647
rect 6411 6613 6423 6647
rect 6365 6607 6423 6613
rect 6638 6604 6644 6656
rect 6696 6644 6702 6656
rect 6733 6647 6791 6653
rect 6733 6644 6745 6647
rect 6696 6616 6745 6644
rect 6696 6604 6702 6616
rect 6733 6613 6745 6616
rect 6779 6613 6791 6647
rect 6733 6607 6791 6613
rect 6822 6604 6828 6656
rect 6880 6644 6886 6656
rect 7098 6644 7104 6656
rect 6880 6616 7104 6644
rect 6880 6604 6886 6616
rect 7098 6604 7104 6616
rect 7156 6604 7162 6656
rect 7300 6644 7328 6675
rect 7374 6672 7380 6724
rect 7432 6712 7438 6724
rect 7469 6715 7527 6721
rect 7469 6712 7481 6715
rect 7432 6684 7481 6712
rect 7432 6672 7438 6684
rect 7469 6681 7481 6684
rect 7515 6681 7527 6715
rect 7469 6675 7527 6681
rect 9214 6672 9220 6724
rect 9272 6712 9278 6724
rect 10042 6712 10048 6724
rect 9272 6684 10048 6712
rect 9272 6672 9278 6684
rect 10042 6672 10048 6684
rect 10100 6672 10106 6724
rect 11606 6712 11612 6724
rect 11178 6684 11468 6712
rect 11567 6684 11612 6712
rect 8110 6644 8116 6656
rect 7300 6616 8116 6644
rect 8110 6604 8116 6616
rect 8168 6604 8174 6656
rect 9030 6604 9036 6656
rect 9088 6644 9094 6656
rect 11238 6644 11244 6656
rect 9088 6616 11244 6644
rect 9088 6604 9094 6616
rect 11238 6604 11244 6616
rect 11296 6604 11302 6656
rect 11440 6644 11468 6684
rect 11606 6672 11612 6684
rect 11664 6672 11670 6724
rect 12084 6712 12112 6743
rect 12158 6740 12164 6792
rect 12216 6780 12222 6792
rect 12253 6783 12311 6789
rect 12253 6780 12265 6783
rect 12216 6752 12265 6780
rect 12216 6740 12222 6752
rect 12253 6749 12265 6752
rect 12299 6749 12311 6783
rect 12713 6783 12771 6789
rect 12713 6780 12725 6783
rect 12253 6743 12311 6749
rect 12406 6752 12725 6780
rect 12406 6712 12434 6752
rect 12713 6749 12725 6752
rect 12759 6749 12771 6783
rect 12713 6743 12771 6749
rect 12805 6783 12863 6789
rect 12805 6749 12817 6783
rect 12851 6780 12863 6783
rect 12894 6780 12900 6792
rect 12851 6752 12900 6780
rect 12851 6749 12863 6752
rect 12805 6743 12863 6749
rect 12894 6740 12900 6752
rect 12952 6740 12958 6792
rect 13357 6783 13415 6789
rect 13357 6749 13369 6783
rect 13403 6780 13415 6783
rect 14274 6780 14280 6792
rect 13403 6752 14280 6780
rect 13403 6749 13415 6752
rect 13357 6743 13415 6749
rect 14274 6740 14280 6752
rect 14332 6740 14338 6792
rect 14568 6780 14596 6809
rect 16022 6808 16028 6820
rect 16080 6808 16086 6860
rect 16574 6848 16580 6860
rect 16535 6820 16580 6848
rect 16574 6808 16580 6820
rect 16632 6808 16638 6860
rect 16942 6848 16948 6860
rect 16903 6820 16948 6848
rect 16942 6808 16948 6820
rect 17000 6808 17006 6860
rect 17589 6851 17647 6857
rect 17589 6848 17601 6851
rect 17052 6820 17601 6848
rect 14476 6774 14596 6780
rect 14384 6752 14596 6774
rect 14384 6746 14504 6752
rect 11808 6684 12112 6712
rect 12176 6684 12434 6712
rect 11808 6656 11836 6684
rect 11514 6644 11520 6656
rect 11440 6616 11520 6644
rect 11514 6604 11520 6616
rect 11572 6604 11578 6656
rect 11790 6604 11796 6656
rect 11848 6604 11854 6656
rect 12066 6604 12072 6656
rect 12124 6644 12130 6656
rect 12176 6644 12204 6684
rect 12618 6672 12624 6724
rect 12676 6712 12682 6724
rect 14384 6712 14412 6746
rect 14734 6740 14740 6792
rect 14792 6780 14798 6792
rect 14829 6783 14887 6789
rect 14829 6780 14841 6783
rect 14792 6752 14841 6780
rect 14792 6740 14798 6752
rect 14829 6749 14841 6752
rect 14875 6749 14887 6783
rect 14829 6743 14887 6749
rect 14918 6740 14924 6792
rect 14976 6780 14982 6792
rect 14976 6752 15021 6780
rect 14976 6740 14982 6752
rect 16666 6740 16672 6792
rect 16724 6780 16730 6792
rect 17052 6780 17080 6820
rect 17589 6817 17601 6820
rect 17635 6817 17647 6851
rect 17589 6811 17647 6817
rect 17494 6780 17500 6792
rect 16724 6752 17080 6780
rect 17407 6752 17500 6780
rect 16724 6740 16730 6752
rect 17494 6740 17500 6752
rect 17552 6780 17558 6792
rect 18141 6783 18199 6789
rect 18141 6780 18153 6783
rect 17552 6752 18153 6780
rect 17552 6740 17558 6752
rect 18141 6749 18153 6752
rect 18187 6749 18199 6783
rect 18141 6743 18199 6749
rect 14642 6712 14648 6724
rect 12676 6684 14412 6712
rect 14603 6684 14648 6712
rect 12676 6672 12682 6684
rect 14642 6672 14648 6684
rect 14700 6672 14706 6724
rect 15286 6672 15292 6724
rect 15344 6712 15350 6724
rect 15344 6706 15594 6712
rect 15344 6684 15700 6706
rect 15344 6672 15350 6684
rect 15580 6678 15700 6684
rect 12124 6616 12204 6644
rect 12124 6604 12130 6616
rect 12250 6604 12256 6656
rect 12308 6644 12314 6656
rect 12529 6647 12587 6653
rect 12529 6644 12541 6647
rect 12308 6616 12541 6644
rect 12308 6604 12314 6616
rect 12529 6613 12541 6616
rect 12575 6613 12587 6647
rect 12529 6607 12587 6613
rect 12802 6604 12808 6656
rect 12860 6644 12866 6656
rect 13078 6644 13084 6656
rect 12860 6616 13084 6644
rect 12860 6604 12866 6616
rect 13078 6604 13084 6616
rect 13136 6604 13142 6656
rect 14090 6604 14096 6656
rect 14148 6644 14154 6656
rect 14185 6647 14243 6653
rect 14185 6644 14197 6647
rect 14148 6616 14197 6644
rect 14148 6604 14154 6616
rect 14185 6613 14197 6616
rect 14231 6613 14243 6647
rect 14185 6607 14243 6613
rect 14277 6647 14335 6653
rect 14277 6613 14289 6647
rect 14323 6644 14335 6647
rect 14366 6644 14372 6656
rect 14323 6616 14372 6644
rect 14323 6613 14335 6616
rect 14277 6607 14335 6613
rect 14366 6604 14372 6616
rect 14424 6604 14430 6656
rect 14734 6644 14740 6656
rect 14695 6616 14740 6644
rect 14734 6604 14740 6616
rect 14792 6604 14798 6656
rect 15672 6644 15700 6678
rect 16298 6644 16304 6656
rect 15672 6616 16304 6644
rect 16298 6604 16304 6616
rect 16356 6604 16362 6656
rect 16850 6604 16856 6656
rect 16908 6644 16914 6656
rect 17037 6647 17095 6653
rect 17037 6644 17049 6647
rect 16908 6616 17049 6644
rect 16908 6604 16914 6616
rect 17037 6613 17049 6616
rect 17083 6613 17095 6647
rect 17402 6644 17408 6656
rect 17363 6616 17408 6644
rect 17037 6607 17095 6613
rect 17402 6604 17408 6616
rect 17460 6604 17466 6656
rect 17954 6604 17960 6656
rect 18012 6644 18018 6656
rect 18325 6647 18383 6653
rect 18325 6644 18337 6647
rect 18012 6616 18337 6644
rect 18012 6604 18018 6616
rect 18325 6613 18337 6616
rect 18371 6613 18383 6647
rect 18325 6607 18383 6613
rect 0 6554 18860 6576
rect 0 6502 6144 6554
rect 6196 6502 6208 6554
rect 6260 6502 6272 6554
rect 6324 6502 6336 6554
rect 6388 6502 6400 6554
rect 6452 6502 12443 6554
rect 12495 6502 12507 6554
rect 12559 6502 12571 6554
rect 12623 6502 12635 6554
rect 12687 6502 12699 6554
rect 12751 6502 18860 6554
rect 0 6480 18860 6502
rect 2590 6400 2596 6452
rect 2648 6400 2654 6452
rect 3050 6400 3056 6452
rect 3108 6440 3114 6452
rect 3881 6443 3939 6449
rect 3881 6440 3893 6443
rect 3108 6412 3893 6440
rect 3108 6400 3114 6412
rect 3881 6409 3893 6412
rect 3927 6409 3939 6443
rect 4246 6440 4252 6452
rect 4207 6412 4252 6440
rect 3881 6403 3939 6409
rect 4246 6400 4252 6412
rect 4304 6400 4310 6452
rect 4341 6443 4399 6449
rect 4341 6409 4353 6443
rect 4387 6440 4399 6443
rect 5626 6440 5632 6452
rect 4387 6412 5632 6440
rect 4387 6409 4399 6412
rect 4341 6403 4399 6409
rect 5626 6400 5632 6412
rect 5684 6400 5690 6452
rect 5997 6443 6055 6449
rect 5997 6409 6009 6443
rect 6043 6440 6055 6443
rect 6457 6443 6515 6449
rect 6457 6440 6469 6443
rect 6043 6412 6469 6440
rect 6043 6409 6055 6412
rect 5997 6403 6055 6409
rect 6457 6409 6469 6412
rect 6503 6409 6515 6443
rect 6457 6403 6515 6409
rect 7834 6400 7840 6452
rect 7892 6440 7898 6452
rect 8021 6443 8079 6449
rect 8021 6440 8033 6443
rect 7892 6412 8033 6440
rect 7892 6400 7898 6412
rect 8021 6409 8033 6412
rect 8067 6409 8079 6443
rect 8021 6403 8079 6409
rect 8110 6400 8116 6452
rect 8168 6440 8174 6452
rect 8389 6443 8447 6449
rect 8389 6440 8401 6443
rect 8168 6412 8401 6440
rect 8168 6400 8174 6412
rect 8389 6409 8401 6412
rect 8435 6409 8447 6443
rect 10226 6440 10232 6452
rect 8389 6403 8447 6409
rect 9646 6412 10232 6440
rect 1670 6372 1676 6384
rect 1631 6344 1676 6372
rect 1670 6332 1676 6344
rect 1728 6332 1734 6384
rect 2608 6358 2636 6400
rect 3513 6375 3571 6381
rect 3513 6372 3525 6375
rect 3344 6344 3525 6372
rect 566 6264 572 6316
rect 624 6304 630 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 624 6276 1409 6304
rect 624 6264 630 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 3234 6304 3240 6316
rect 3195 6276 3240 6304
rect 1397 6267 1455 6273
rect 3234 6264 3240 6276
rect 3292 6264 3298 6316
rect 3145 6171 3203 6177
rect 3145 6137 3157 6171
rect 3191 6168 3203 6171
rect 3344 6168 3372 6344
rect 3513 6341 3525 6344
rect 3559 6341 3571 6375
rect 3513 6335 3571 6341
rect 3602 6332 3608 6384
rect 3660 6372 3666 6384
rect 3697 6375 3755 6381
rect 3697 6372 3709 6375
rect 3660 6344 3709 6372
rect 3660 6332 3666 6344
rect 3697 6341 3709 6344
rect 3743 6372 3755 6375
rect 4801 6375 4859 6381
rect 4801 6372 4813 6375
rect 3743 6344 4813 6372
rect 3743 6341 3755 6344
rect 3697 6335 3755 6341
rect 4801 6341 4813 6344
rect 4847 6341 4859 6375
rect 4801 6335 4859 6341
rect 5350 6332 5356 6384
rect 5408 6372 5414 6384
rect 5408 6344 5856 6372
rect 5408 6332 5414 6344
rect 3421 6307 3479 6313
rect 3421 6273 3433 6307
rect 3467 6273 3479 6307
rect 3786 6304 3792 6316
rect 3747 6276 3792 6304
rect 3421 6267 3479 6273
rect 3436 6236 3464 6267
rect 3786 6264 3792 6276
rect 3844 6264 3850 6316
rect 4890 6304 4896 6316
rect 3896 6276 4660 6304
rect 4851 6276 4896 6304
rect 3896 6236 3924 6276
rect 4246 6236 4252 6248
rect 3436 6208 3924 6236
rect 3988 6208 4252 6236
rect 3878 6168 3884 6180
rect 3191 6140 3884 6168
rect 3191 6137 3203 6140
rect 3145 6131 3203 6137
rect 3878 6128 3884 6140
rect 3936 6168 3942 6180
rect 3988 6168 4016 6208
rect 4246 6196 4252 6208
rect 4304 6196 4310 6248
rect 4338 6196 4344 6248
rect 4396 6236 4402 6248
rect 4433 6239 4491 6245
rect 4433 6236 4445 6239
rect 4396 6208 4445 6236
rect 4396 6196 4402 6208
rect 4433 6205 4445 6208
rect 4479 6205 4491 6239
rect 4632 6236 4660 6276
rect 4890 6264 4896 6276
rect 4948 6264 4954 6316
rect 5074 6264 5080 6316
rect 5132 6304 5138 6316
rect 5261 6307 5319 6313
rect 5261 6304 5273 6307
rect 5132 6276 5273 6304
rect 5132 6264 5138 6276
rect 5261 6273 5273 6276
rect 5307 6273 5319 6307
rect 5442 6304 5448 6316
rect 5403 6276 5448 6304
rect 5261 6267 5319 6273
rect 5442 6264 5448 6276
rect 5500 6264 5506 6316
rect 4632 6208 5672 6236
rect 4433 6199 4491 6205
rect 3936 6140 4016 6168
rect 3936 6128 3942 6140
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 5644 6177 5672 6208
rect 5353 6171 5411 6177
rect 5353 6168 5365 6171
rect 4120 6140 5365 6168
rect 4120 6128 4126 6140
rect 5353 6137 5365 6140
rect 5399 6137 5411 6171
rect 5353 6131 5411 6137
rect 5629 6171 5687 6177
rect 5629 6137 5641 6171
rect 5675 6137 5687 6171
rect 5828 6168 5856 6344
rect 5902 6332 5908 6384
rect 5960 6372 5966 6384
rect 6089 6375 6147 6381
rect 6089 6372 6101 6375
rect 5960 6344 6101 6372
rect 5960 6332 5966 6344
rect 6089 6341 6101 6344
rect 6135 6372 6147 6375
rect 6917 6375 6975 6381
rect 6917 6372 6929 6375
rect 6135 6344 6929 6372
rect 6135 6341 6147 6344
rect 6089 6335 6147 6341
rect 6917 6341 6929 6344
rect 6963 6372 6975 6375
rect 8662 6372 8668 6384
rect 6963 6344 8668 6372
rect 6963 6341 6975 6344
rect 6917 6335 6975 6341
rect 8662 6332 8668 6344
rect 8720 6372 8726 6384
rect 8840 6375 8898 6381
rect 8840 6372 8852 6375
rect 8720 6344 8852 6372
rect 8720 6332 8726 6344
rect 8840 6341 8852 6344
rect 8886 6372 8898 6375
rect 9646 6372 9674 6412
rect 10226 6400 10232 6412
rect 10284 6400 10290 6452
rect 11425 6443 11483 6449
rect 11425 6409 11437 6443
rect 11471 6440 11483 6443
rect 11606 6440 11612 6452
rect 11471 6412 11612 6440
rect 11471 6409 11483 6412
rect 11425 6403 11483 6409
rect 11606 6400 11612 6412
rect 11664 6400 11670 6452
rect 11698 6400 11704 6452
rect 11756 6440 11762 6452
rect 11882 6440 11888 6452
rect 11756 6412 11888 6440
rect 11756 6400 11762 6412
rect 11882 6400 11888 6412
rect 11940 6440 11946 6452
rect 15010 6440 15016 6452
rect 11940 6412 14412 6440
rect 14971 6412 15016 6440
rect 11940 6400 11946 6412
rect 12066 6372 12072 6384
rect 8886 6344 9674 6372
rect 10603 6344 11744 6372
rect 12027 6344 12072 6372
rect 8886 6341 8898 6344
rect 8840 6335 8898 6341
rect 6822 6304 6828 6316
rect 6783 6276 6828 6304
rect 6822 6264 6828 6276
rect 6880 6264 6886 6316
rect 7190 6264 7196 6316
rect 7248 6304 7254 6316
rect 8110 6304 8116 6316
rect 7248 6276 8116 6304
rect 7248 6264 7254 6276
rect 8110 6264 8116 6276
rect 8168 6264 8174 6316
rect 8478 6304 8484 6316
rect 8439 6276 8484 6304
rect 8478 6264 8484 6276
rect 8536 6264 8542 6316
rect 10045 6307 10103 6313
rect 10045 6273 10057 6307
rect 10091 6273 10103 6307
rect 10045 6267 10103 6273
rect 6273 6239 6331 6245
rect 6273 6205 6285 6239
rect 6319 6236 6331 6239
rect 6546 6236 6552 6248
rect 6319 6208 6552 6236
rect 6319 6205 6331 6208
rect 6273 6199 6331 6205
rect 6546 6196 6552 6208
rect 6604 6196 6610 6248
rect 7009 6239 7067 6245
rect 7009 6205 7021 6239
rect 7055 6205 7067 6239
rect 8128 6236 8156 6264
rect 8573 6239 8631 6245
rect 8573 6236 8585 6239
rect 8128 6208 8585 6236
rect 7009 6199 7067 6205
rect 8573 6205 8585 6208
rect 8619 6205 8631 6239
rect 10060 6236 10088 6267
rect 10226 6264 10232 6316
rect 10284 6304 10290 6316
rect 10284 6276 10329 6304
rect 10284 6264 10290 6276
rect 10603 6236 10631 6344
rect 10778 6264 10784 6316
rect 10836 6304 10842 6316
rect 10873 6307 10931 6313
rect 10873 6304 10885 6307
rect 10836 6276 10885 6304
rect 10836 6264 10842 6276
rect 10873 6273 10885 6276
rect 10919 6273 10931 6307
rect 11238 6304 11244 6316
rect 11199 6276 11244 6304
rect 10873 6267 10931 6273
rect 11238 6264 11244 6276
rect 11296 6264 11302 6316
rect 11716 6313 11744 6344
rect 12066 6332 12072 6344
rect 12124 6332 12130 6384
rect 11701 6307 11759 6313
rect 11701 6273 11713 6307
rect 11747 6273 11759 6307
rect 11882 6304 11888 6316
rect 11843 6276 11888 6304
rect 11701 6267 11759 6273
rect 11882 6264 11888 6276
rect 11940 6264 11946 6316
rect 10962 6236 10968 6248
rect 8573 6199 8631 6205
rect 9968 6208 10631 6236
rect 10923 6208 10968 6236
rect 7024 6168 7052 6199
rect 7190 6168 7196 6180
rect 5828 6140 7196 6168
rect 5629 6131 5687 6137
rect 7190 6128 7196 6140
rect 7248 6128 7254 6180
rect 9968 6177 9996 6208
rect 10962 6196 10968 6208
rect 11020 6196 11026 6248
rect 11057 6239 11115 6245
rect 11057 6205 11069 6239
rect 11103 6236 11115 6239
rect 11606 6236 11612 6248
rect 11103 6208 11612 6236
rect 11103 6205 11115 6208
rect 11057 6199 11115 6205
rect 11606 6196 11612 6208
rect 11664 6196 11670 6248
rect 12161 6239 12219 6245
rect 12161 6205 12173 6239
rect 12207 6236 12219 6239
rect 12268 6236 12296 6412
rect 14384 6384 14412 6412
rect 15010 6400 15016 6412
rect 15068 6400 15074 6452
rect 15102 6400 15108 6452
rect 15160 6440 15166 6452
rect 15160 6412 17080 6440
rect 15160 6400 15166 6412
rect 13078 6332 13084 6384
rect 13136 6332 13142 6384
rect 14182 6372 14188 6384
rect 14143 6344 14188 6372
rect 14182 6332 14188 6344
rect 14240 6332 14246 6384
rect 14366 6332 14372 6384
rect 14424 6372 14430 6384
rect 14424 6344 15608 6372
rect 14424 6332 14430 6344
rect 13354 6264 13360 6316
rect 13412 6304 13418 6316
rect 15105 6307 15163 6313
rect 13412 6276 15056 6304
rect 13412 6264 13418 6276
rect 12207 6208 12296 6236
rect 12529 6239 12587 6245
rect 12207 6205 12219 6208
rect 12161 6199 12219 6205
rect 12529 6205 12541 6239
rect 12575 6236 12587 6239
rect 12802 6236 12808 6248
rect 12575 6208 12808 6236
rect 12575 6205 12587 6208
rect 12529 6199 12587 6205
rect 12802 6196 12808 6208
rect 12860 6196 12866 6248
rect 13630 6196 13636 6248
rect 13688 6236 13694 6248
rect 14918 6236 14924 6248
rect 13688 6208 14924 6236
rect 13688 6196 13694 6208
rect 14918 6196 14924 6208
rect 14976 6196 14982 6248
rect 15028 6236 15056 6276
rect 15105 6273 15117 6307
rect 15151 6304 15163 6307
rect 15470 6304 15476 6316
rect 15151 6276 15476 6304
rect 15151 6273 15163 6276
rect 15105 6267 15163 6273
rect 15470 6264 15476 6276
rect 15528 6264 15534 6316
rect 15580 6313 15608 6344
rect 16298 6332 16304 6384
rect 16356 6332 16362 6384
rect 17052 6372 17080 6412
rect 17402 6400 17408 6452
rect 17460 6440 17466 6452
rect 17497 6443 17555 6449
rect 17497 6440 17509 6443
rect 17460 6412 17509 6440
rect 17460 6400 17466 6412
rect 17497 6409 17509 6412
rect 17543 6409 17555 6443
rect 17954 6440 17960 6452
rect 17915 6412 17960 6440
rect 17497 6403 17555 6409
rect 17954 6400 17960 6412
rect 18012 6400 18018 6452
rect 17865 6375 17923 6381
rect 17865 6372 17877 6375
rect 17052 6344 17877 6372
rect 17865 6341 17877 6344
rect 17911 6341 17923 6375
rect 17865 6335 17923 6341
rect 15565 6307 15623 6313
rect 15565 6273 15577 6307
rect 15611 6304 15623 6307
rect 16022 6304 16028 6316
rect 15611 6276 16028 6304
rect 15611 6273 15623 6276
rect 15565 6267 15623 6273
rect 16022 6264 16028 6276
rect 16080 6264 16086 6316
rect 17359 6307 17417 6313
rect 17359 6273 17371 6307
rect 17405 6304 17417 6307
rect 17494 6304 17500 6316
rect 17405 6276 17500 6304
rect 17405 6273 17417 6276
rect 17359 6267 17417 6273
rect 17494 6264 17500 6276
rect 17552 6264 17558 6316
rect 17586 6264 17592 6316
rect 17644 6304 17650 6316
rect 18325 6307 18383 6313
rect 18325 6304 18337 6307
rect 17644 6276 18337 6304
rect 17644 6264 17650 6276
rect 18325 6273 18337 6276
rect 18371 6273 18383 6307
rect 18325 6267 18383 6273
rect 15197 6239 15255 6245
rect 15197 6236 15209 6239
rect 15028 6208 15209 6236
rect 15197 6205 15209 6208
rect 15243 6236 15255 6239
rect 15286 6236 15292 6248
rect 15243 6208 15292 6236
rect 15243 6205 15255 6208
rect 15197 6199 15255 6205
rect 15286 6196 15292 6208
rect 15344 6196 15350 6248
rect 15930 6236 15936 6248
rect 15891 6208 15936 6236
rect 15930 6196 15936 6208
rect 15988 6196 15994 6248
rect 18138 6236 18144 6248
rect 18051 6208 18144 6236
rect 18138 6196 18144 6208
rect 18196 6236 18202 6248
rect 18417 6239 18475 6245
rect 18417 6236 18429 6239
rect 18196 6208 18429 6236
rect 18196 6196 18202 6208
rect 18417 6205 18429 6208
rect 18463 6205 18475 6239
rect 18417 6199 18475 6205
rect 9953 6171 10011 6177
rect 9953 6137 9965 6171
rect 9999 6137 10011 6171
rect 9953 6131 10011 6137
rect 10229 6171 10287 6177
rect 10229 6137 10241 6171
rect 10275 6168 10287 6171
rect 10275 6140 12204 6168
rect 10275 6137 10287 6140
rect 10229 6131 10287 6137
rect 3326 6100 3332 6112
rect 3287 6072 3332 6100
rect 3326 6060 3332 6072
rect 3384 6060 3390 6112
rect 3789 6103 3847 6109
rect 3789 6069 3801 6103
rect 3835 6100 3847 6103
rect 5810 6100 5816 6112
rect 3835 6072 5816 6100
rect 3835 6069 3847 6072
rect 3789 6063 3847 6069
rect 5810 6060 5816 6072
rect 5868 6060 5874 6112
rect 8386 6060 8392 6112
rect 8444 6100 8450 6112
rect 10134 6100 10140 6112
rect 8444 6072 10140 6100
rect 8444 6060 8450 6072
rect 10134 6060 10140 6072
rect 10192 6060 10198 6112
rect 10410 6100 10416 6112
rect 10371 6072 10416 6100
rect 10410 6060 10416 6072
rect 10468 6060 10474 6112
rect 10502 6060 10508 6112
rect 10560 6100 10566 6112
rect 10597 6103 10655 6109
rect 10597 6100 10609 6103
rect 10560 6072 10609 6100
rect 10560 6060 10566 6072
rect 10597 6069 10609 6072
rect 10643 6100 10655 6103
rect 11974 6100 11980 6112
rect 10643 6072 11980 6100
rect 10643 6069 10655 6072
rect 10597 6063 10655 6069
rect 11974 6060 11980 6072
rect 12032 6060 12038 6112
rect 12176 6100 12204 6140
rect 13722 6128 13728 6180
rect 13780 6168 13786 6180
rect 14645 6171 14703 6177
rect 14645 6168 14657 6171
rect 13780 6140 14657 6168
rect 13780 6128 13786 6140
rect 14645 6137 14657 6140
rect 14691 6137 14703 6171
rect 14645 6131 14703 6137
rect 12894 6100 12900 6112
rect 12176 6072 12900 6100
rect 12894 6060 12900 6072
rect 12952 6060 12958 6112
rect 13955 6103 14013 6109
rect 13955 6069 13967 6103
rect 14001 6100 14013 6103
rect 14182 6100 14188 6112
rect 14001 6072 14188 6100
rect 14001 6069 14013 6072
rect 13955 6063 14013 6069
rect 14182 6060 14188 6072
rect 14240 6060 14246 6112
rect 15010 6060 15016 6112
rect 15068 6100 15074 6112
rect 17218 6100 17224 6112
rect 15068 6072 17224 6100
rect 15068 6060 15074 6072
rect 17218 6060 17224 6072
rect 17276 6060 17282 6112
rect 0 6010 18860 6032
rect 0 5958 2995 6010
rect 3047 5958 3059 6010
rect 3111 5958 3123 6010
rect 3175 5958 3187 6010
rect 3239 5958 3251 6010
rect 3303 5958 9294 6010
rect 9346 5958 9358 6010
rect 9410 5958 9422 6010
rect 9474 5958 9486 6010
rect 9538 5958 9550 6010
rect 9602 5958 15592 6010
rect 15644 5958 15656 6010
rect 15708 5958 15720 6010
rect 15772 5958 15784 6010
rect 15836 5958 15848 6010
rect 15900 5958 18860 6010
rect 0 5936 18860 5958
rect 4154 5896 4160 5908
rect 768 5868 4160 5896
rect 566 5720 572 5772
rect 624 5760 630 5772
rect 768 5769 796 5868
rect 4154 5856 4160 5868
rect 4212 5856 4218 5908
rect 4246 5856 4252 5908
rect 4304 5896 4310 5908
rect 6638 5896 6644 5908
rect 4304 5868 4568 5896
rect 6599 5868 6644 5896
rect 4304 5856 4310 5868
rect 3237 5831 3295 5837
rect 3237 5828 3249 5831
rect 2056 5800 3249 5828
rect 753 5763 811 5769
rect 753 5760 765 5763
rect 624 5732 765 5760
rect 624 5720 630 5732
rect 753 5729 765 5732
rect 799 5729 811 5763
rect 753 5723 811 5729
rect 1029 5763 1087 5769
rect 1029 5729 1041 5763
rect 1075 5760 1087 5763
rect 2056 5760 2084 5800
rect 3237 5797 3249 5800
rect 3283 5797 3295 5831
rect 3237 5791 3295 5797
rect 3326 5788 3332 5840
rect 3384 5788 3390 5840
rect 3786 5828 3792 5840
rect 3528 5800 3792 5828
rect 1075 5732 2084 5760
rect 3145 5763 3203 5769
rect 1075 5729 1087 5732
rect 1029 5723 1087 5729
rect 3145 5729 3157 5763
rect 3191 5760 3203 5763
rect 3344 5760 3372 5788
rect 3528 5760 3556 5800
rect 3786 5788 3792 5800
rect 3844 5828 3850 5840
rect 4540 5837 4568 5868
rect 6638 5856 6644 5868
rect 6696 5856 6702 5908
rect 9493 5899 9551 5905
rect 9493 5865 9505 5899
rect 9539 5896 9551 5899
rect 10778 5896 10784 5908
rect 9539 5868 10784 5896
rect 9539 5865 9551 5868
rect 9493 5859 9551 5865
rect 10778 5856 10784 5868
rect 10836 5856 10842 5908
rect 12805 5899 12863 5905
rect 12805 5865 12817 5899
rect 12851 5896 12863 5899
rect 12986 5896 12992 5908
rect 12851 5868 12992 5896
rect 12851 5865 12863 5868
rect 12805 5859 12863 5865
rect 12986 5856 12992 5868
rect 13044 5856 13050 5908
rect 13262 5856 13268 5908
rect 13320 5896 13326 5908
rect 14274 5896 14280 5908
rect 13320 5868 14280 5896
rect 13320 5856 13326 5868
rect 14274 5856 14280 5868
rect 14332 5896 14338 5908
rect 14642 5896 14648 5908
rect 14332 5868 14648 5896
rect 14332 5856 14338 5868
rect 14642 5856 14648 5868
rect 14700 5856 14706 5908
rect 15470 5856 15476 5908
rect 15528 5896 15534 5908
rect 15749 5899 15807 5905
rect 15749 5896 15761 5899
rect 15528 5868 15761 5896
rect 15528 5856 15534 5868
rect 15749 5865 15761 5868
rect 15795 5896 15807 5899
rect 15841 5899 15899 5905
rect 15841 5896 15853 5899
rect 15795 5868 15853 5896
rect 15795 5865 15807 5868
rect 15749 5859 15807 5865
rect 15841 5865 15853 5868
rect 15887 5865 15899 5899
rect 15841 5859 15899 5865
rect 16298 5856 16304 5908
rect 16356 5896 16362 5908
rect 16942 5896 16948 5908
rect 16356 5868 16948 5896
rect 16356 5856 16362 5868
rect 16942 5856 16948 5868
rect 17000 5856 17006 5908
rect 17218 5896 17224 5908
rect 17179 5868 17224 5896
rect 17218 5856 17224 5868
rect 17276 5856 17282 5908
rect 18322 5896 18328 5908
rect 18283 5868 18328 5896
rect 18322 5856 18328 5868
rect 18380 5856 18386 5908
rect 4341 5831 4399 5837
rect 4341 5828 4353 5831
rect 3844 5800 4353 5828
rect 3844 5788 3850 5800
rect 4341 5797 4353 5800
rect 4387 5797 4399 5831
rect 4341 5791 4399 5797
rect 4525 5831 4583 5837
rect 4525 5797 4537 5831
rect 4571 5828 4583 5831
rect 4571 5800 5948 5828
rect 4571 5797 4583 5800
rect 4525 5791 4583 5797
rect 3191 5732 3372 5760
rect 3436 5732 3556 5760
rect 3881 5763 3939 5769
rect 3191 5729 3203 5732
rect 3145 5723 3203 5729
rect 3326 5692 3332 5704
rect 3287 5664 3332 5692
rect 3326 5652 3332 5664
rect 3384 5652 3390 5704
rect 3436 5701 3464 5732
rect 3881 5729 3893 5763
rect 3927 5760 3939 5763
rect 3970 5760 3976 5772
rect 3927 5732 3976 5760
rect 3927 5729 3939 5732
rect 3881 5723 3939 5729
rect 3970 5720 3976 5732
rect 4028 5720 4034 5772
rect 5626 5760 5632 5772
rect 4448 5732 5632 5760
rect 3421 5695 3479 5701
rect 3421 5661 3433 5695
rect 3467 5661 3479 5695
rect 3602 5692 3608 5704
rect 3563 5664 3608 5692
rect 3421 5655 3479 5661
rect 3602 5652 3608 5664
rect 3660 5652 3666 5704
rect 3697 5695 3755 5701
rect 3697 5661 3709 5695
rect 3743 5661 3755 5695
rect 3697 5655 3755 5661
rect 2590 5624 2596 5636
rect 2254 5596 2596 5624
rect 2590 5584 2596 5596
rect 2648 5584 2654 5636
rect 3344 5624 3372 5652
rect 3712 5624 3740 5655
rect 3786 5652 3792 5704
rect 3844 5692 3850 5704
rect 4154 5692 4160 5704
rect 3844 5664 3924 5692
rect 4115 5664 4160 5692
rect 3844 5652 3850 5664
rect 3896 5633 3924 5664
rect 4154 5652 4160 5664
rect 4212 5652 4218 5704
rect 4448 5701 4476 5732
rect 4433 5695 4491 5701
rect 4433 5661 4445 5695
rect 4479 5661 4491 5695
rect 4433 5655 4491 5661
rect 4525 5695 4583 5701
rect 4525 5661 4537 5695
rect 4571 5692 4583 5695
rect 4617 5695 4675 5701
rect 4617 5692 4629 5695
rect 4571 5664 4629 5692
rect 4571 5661 4583 5664
rect 4525 5655 4583 5661
rect 4617 5661 4629 5664
rect 4663 5661 4675 5695
rect 4617 5655 4675 5661
rect 3344 5596 3740 5624
rect 3881 5627 3939 5633
rect 3881 5593 3893 5627
rect 3927 5593 3939 5627
rect 4062 5624 4068 5636
rect 4023 5596 4068 5624
rect 3881 5587 3939 5593
rect 4062 5584 4068 5596
rect 4120 5584 4126 5636
rect 2501 5559 2559 5565
rect 2501 5525 2513 5559
rect 2547 5556 2559 5559
rect 4448 5556 4476 5655
rect 4890 5652 4896 5704
rect 4948 5692 4954 5704
rect 5368 5701 5396 5732
rect 5626 5720 5632 5732
rect 5684 5720 5690 5772
rect 5920 5769 5948 5800
rect 15286 5788 15292 5840
rect 15344 5828 15350 5840
rect 16117 5831 16175 5837
rect 16117 5828 16129 5831
rect 15344 5800 16129 5828
rect 15344 5788 15350 5800
rect 16117 5797 16129 5800
rect 16163 5828 16175 5831
rect 16574 5828 16580 5840
rect 16163 5800 16580 5828
rect 16163 5797 16175 5800
rect 16117 5791 16175 5797
rect 16574 5788 16580 5800
rect 16632 5788 16638 5840
rect 5905 5763 5963 5769
rect 5905 5729 5917 5763
rect 5951 5729 5963 5763
rect 7190 5760 7196 5772
rect 7151 5732 7196 5760
rect 5905 5723 5963 5729
rect 4985 5695 5043 5701
rect 4985 5692 4997 5695
rect 4948 5664 4997 5692
rect 4948 5652 4954 5664
rect 4985 5661 4997 5664
rect 5031 5661 5043 5695
rect 4985 5655 5043 5661
rect 5353 5695 5411 5701
rect 5353 5661 5365 5695
rect 5399 5661 5411 5695
rect 5353 5655 5411 5661
rect 5537 5695 5595 5701
rect 5537 5661 5549 5695
rect 5583 5661 5595 5695
rect 5537 5655 5595 5661
rect 5721 5695 5779 5701
rect 5721 5661 5733 5695
rect 5767 5692 5779 5695
rect 5920 5692 5948 5723
rect 7190 5720 7196 5732
rect 7248 5720 7254 5772
rect 8110 5760 8116 5772
rect 8071 5732 8116 5760
rect 8110 5720 8116 5732
rect 8168 5720 8174 5772
rect 10965 5763 11023 5769
rect 10965 5729 10977 5763
rect 11011 5760 11023 5763
rect 11698 5760 11704 5772
rect 11011 5732 11704 5760
rect 11011 5729 11023 5732
rect 10965 5723 11023 5729
rect 11698 5720 11704 5732
rect 11756 5720 11762 5772
rect 13906 5760 13912 5772
rect 13556 5732 13912 5760
rect 5767 5664 5948 5692
rect 5997 5695 6055 5701
rect 5767 5661 5779 5664
rect 5721 5655 5779 5661
rect 5997 5661 6009 5695
rect 6043 5661 6055 5695
rect 7834 5692 7840 5704
rect 7795 5664 7840 5692
rect 5997 5655 6055 5661
rect 5000 5624 5028 5655
rect 5552 5624 5580 5655
rect 6012 5624 6040 5655
rect 7834 5652 7840 5664
rect 7892 5652 7898 5704
rect 8018 5692 8024 5704
rect 7979 5664 8024 5692
rect 8018 5652 8024 5664
rect 8076 5652 8082 5704
rect 8380 5695 8438 5701
rect 8380 5692 8392 5695
rect 8128 5664 8392 5692
rect 7098 5624 7104 5636
rect 5000 5596 6040 5624
rect 7011 5596 7104 5624
rect 7098 5584 7104 5596
rect 7156 5624 7162 5636
rect 8128 5624 8156 5664
rect 8380 5661 8392 5664
rect 8426 5692 8438 5695
rect 9950 5692 9956 5704
rect 8426 5664 9956 5692
rect 8426 5661 8438 5664
rect 8380 5655 8438 5661
rect 9950 5652 9956 5664
rect 10008 5652 10014 5704
rect 10134 5652 10140 5704
rect 10192 5692 10198 5704
rect 11054 5692 11060 5704
rect 10192 5664 10640 5692
rect 11015 5664 11060 5692
rect 10192 5652 10198 5664
rect 10502 5624 10508 5636
rect 7156 5596 8156 5624
rect 9508 5596 10508 5624
rect 7156 5584 7162 5596
rect 5350 5556 5356 5568
rect 2547 5528 4476 5556
rect 5311 5528 5356 5556
rect 2547 5525 2559 5528
rect 2501 5519 2559 5525
rect 5350 5516 5356 5528
rect 5408 5516 5414 5568
rect 5629 5559 5687 5565
rect 5629 5525 5641 5559
rect 5675 5556 5687 5559
rect 5810 5556 5816 5568
rect 5675 5528 5816 5556
rect 5675 5525 5687 5528
rect 5629 5519 5687 5525
rect 5810 5516 5816 5528
rect 5868 5516 5874 5568
rect 6365 5559 6423 5565
rect 6365 5525 6377 5559
rect 6411 5556 6423 5559
rect 7009 5559 7067 5565
rect 7009 5556 7021 5559
rect 6411 5528 7021 5556
rect 6411 5525 6423 5528
rect 6365 5519 6423 5525
rect 7009 5525 7021 5528
rect 7055 5525 7067 5559
rect 7009 5519 7067 5525
rect 7929 5559 7987 5565
rect 7929 5525 7941 5559
rect 7975 5556 7987 5559
rect 9508 5556 9536 5596
rect 10502 5584 10508 5596
rect 10560 5584 10566 5636
rect 10612 5624 10640 5664
rect 11054 5652 11060 5664
rect 11112 5652 11118 5704
rect 12342 5652 12348 5704
rect 12400 5692 12406 5704
rect 13078 5692 13084 5704
rect 12400 5664 13084 5692
rect 12400 5652 12406 5664
rect 13078 5652 13084 5664
rect 13136 5652 13142 5704
rect 13262 5692 13268 5704
rect 13223 5664 13268 5692
rect 13262 5652 13268 5664
rect 13320 5652 13326 5704
rect 13446 5652 13452 5704
rect 13504 5692 13510 5704
rect 13556 5701 13584 5732
rect 13906 5720 13912 5732
rect 13964 5720 13970 5772
rect 14001 5763 14059 5769
rect 14001 5729 14013 5763
rect 14047 5760 14059 5763
rect 14366 5760 14372 5772
rect 14047 5732 14372 5760
rect 14047 5729 14059 5732
rect 14001 5723 14059 5729
rect 14366 5720 14372 5732
rect 14424 5720 14430 5772
rect 16390 5760 16396 5772
rect 16224 5732 16396 5760
rect 13541 5695 13599 5701
rect 13541 5692 13553 5695
rect 13504 5664 13553 5692
rect 13504 5652 13510 5664
rect 13541 5661 13553 5664
rect 13587 5661 13599 5695
rect 13722 5692 13728 5704
rect 13683 5664 13728 5692
rect 13541 5655 13599 5661
rect 13722 5652 13728 5664
rect 13780 5652 13786 5704
rect 16224 5701 16252 5732
rect 16390 5720 16396 5732
rect 16448 5760 16454 5772
rect 17865 5763 17923 5769
rect 16448 5732 17172 5760
rect 16448 5720 16454 5732
rect 15841 5695 15899 5701
rect 15841 5661 15853 5695
rect 15887 5692 15899 5695
rect 15933 5695 15991 5701
rect 15933 5692 15945 5695
rect 15887 5664 15945 5692
rect 15887 5661 15899 5664
rect 15841 5655 15899 5661
rect 15933 5661 15945 5664
rect 15979 5661 15991 5695
rect 15933 5655 15991 5661
rect 16209 5695 16267 5701
rect 16209 5661 16221 5695
rect 16255 5661 16267 5695
rect 16209 5655 16267 5661
rect 10709 5627 10767 5633
rect 10709 5624 10721 5627
rect 10612 5596 10721 5624
rect 10709 5593 10721 5596
rect 10755 5624 10767 5627
rect 11330 5624 11336 5636
rect 10755 5596 10824 5624
rect 11291 5596 11336 5624
rect 10755 5593 10767 5596
rect 10709 5587 10767 5593
rect 7975 5528 9536 5556
rect 9585 5559 9643 5565
rect 7975 5525 7987 5528
rect 7929 5519 7987 5525
rect 9585 5525 9597 5559
rect 9631 5556 9643 5559
rect 9950 5556 9956 5568
rect 9631 5528 9956 5556
rect 9631 5525 9643 5528
rect 9585 5519 9643 5525
rect 9950 5516 9956 5528
rect 10008 5516 10014 5568
rect 10796 5556 10824 5596
rect 11330 5584 11336 5596
rect 11388 5584 11394 5636
rect 14277 5627 14335 5633
rect 14277 5624 14289 5627
rect 14272 5593 14289 5624
rect 14323 5593 14335 5627
rect 14272 5587 14335 5593
rect 12158 5556 12164 5568
rect 10796 5528 12164 5556
rect 12158 5516 12164 5528
rect 12216 5516 12222 5568
rect 13078 5556 13084 5568
rect 13039 5528 13084 5556
rect 13078 5516 13084 5528
rect 13136 5516 13142 5568
rect 13449 5559 13507 5565
rect 13449 5525 13461 5559
rect 13495 5556 13507 5559
rect 13630 5556 13636 5568
rect 13495 5528 13636 5556
rect 13495 5525 13507 5528
rect 13449 5519 13507 5525
rect 13630 5516 13636 5528
rect 13688 5516 13694 5568
rect 13909 5559 13967 5565
rect 13909 5525 13921 5559
rect 13955 5556 13967 5559
rect 14272 5556 14300 5587
rect 14366 5584 14372 5636
rect 14424 5624 14430 5636
rect 15948 5624 15976 5655
rect 16298 5652 16304 5704
rect 16356 5692 16362 5704
rect 16666 5692 16672 5704
rect 16356 5664 16449 5692
rect 16627 5664 16672 5692
rect 16356 5652 16362 5664
rect 16408 5624 16436 5664
rect 16666 5652 16672 5664
rect 16724 5652 16730 5704
rect 17144 5701 17172 5732
rect 17865 5729 17877 5763
rect 17911 5760 17923 5763
rect 18138 5760 18144 5772
rect 17911 5732 18144 5760
rect 17911 5729 17923 5732
rect 17865 5723 17923 5729
rect 18138 5720 18144 5732
rect 18196 5720 18202 5772
rect 17129 5695 17187 5701
rect 17129 5661 17141 5695
rect 17175 5692 17187 5695
rect 17494 5692 17500 5704
rect 17175 5664 17500 5692
rect 17175 5661 17187 5664
rect 17129 5655 17187 5661
rect 17494 5652 17500 5664
rect 17552 5652 17558 5704
rect 17589 5695 17647 5701
rect 17589 5661 17601 5695
rect 17635 5692 17647 5695
rect 17770 5692 17776 5704
rect 17635 5664 17776 5692
rect 17635 5661 17647 5664
rect 17589 5655 17647 5661
rect 17770 5652 17776 5664
rect 17828 5652 17834 5704
rect 18506 5692 18512 5704
rect 18467 5664 18512 5692
rect 18506 5652 18512 5664
rect 18564 5652 18570 5704
rect 14424 5596 14766 5624
rect 15948 5596 16436 5624
rect 16684 5624 16712 5652
rect 17862 5624 17868 5636
rect 16684 5596 17868 5624
rect 14424 5584 14430 5596
rect 17862 5584 17868 5596
rect 17920 5584 17926 5636
rect 16206 5556 16212 5568
rect 13955 5528 14300 5556
rect 16167 5528 16212 5556
rect 13955 5525 13967 5528
rect 13909 5519 13967 5525
rect 16206 5516 16212 5528
rect 16264 5516 16270 5568
rect 16853 5559 16911 5565
rect 16853 5525 16865 5559
rect 16899 5556 16911 5559
rect 17586 5556 17592 5568
rect 16899 5528 17592 5556
rect 16899 5525 16911 5528
rect 16853 5519 16911 5525
rect 17586 5516 17592 5528
rect 17644 5516 17650 5568
rect 17678 5516 17684 5568
rect 17736 5556 17742 5568
rect 17736 5528 17781 5556
rect 17736 5516 17742 5528
rect 0 5466 18860 5488
rect 0 5414 6144 5466
rect 6196 5414 6208 5466
rect 6260 5414 6272 5466
rect 6324 5414 6336 5466
rect 6388 5414 6400 5466
rect 6452 5414 12443 5466
rect 12495 5414 12507 5466
rect 12559 5414 12571 5466
rect 12623 5414 12635 5466
rect 12687 5414 12699 5466
rect 12751 5414 18860 5466
rect 0 5392 18860 5414
rect 4062 5352 4068 5364
rect 3160 5324 4068 5352
rect 3160 5225 3188 5324
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 4890 5312 4896 5364
rect 4948 5361 4954 5364
rect 4948 5355 4997 5361
rect 4948 5321 4951 5355
rect 4985 5321 4997 5355
rect 4948 5315 4997 5321
rect 8021 5355 8079 5361
rect 8021 5321 8033 5355
rect 8067 5321 8079 5355
rect 8021 5315 8079 5321
rect 10229 5355 10287 5361
rect 10229 5321 10241 5355
rect 10275 5352 10287 5355
rect 10962 5352 10968 5364
rect 10275 5324 10968 5352
rect 10275 5321 10287 5324
rect 10229 5315 10287 5321
rect 4948 5312 4954 5315
rect 4338 5244 4344 5296
rect 4396 5244 4402 5296
rect 3145 5219 3203 5225
rect 3145 5185 3157 5219
rect 3191 5185 3203 5219
rect 3145 5179 3203 5185
rect 5626 5176 5632 5228
rect 5684 5216 5690 5228
rect 5905 5219 5963 5225
rect 5905 5216 5917 5219
rect 5684 5188 5917 5216
rect 5684 5176 5690 5188
rect 5905 5185 5917 5188
rect 5951 5185 5963 5219
rect 5905 5179 5963 5185
rect 7561 5219 7619 5225
rect 7561 5185 7573 5219
rect 7607 5216 7619 5219
rect 7834 5216 7840 5228
rect 7607 5188 7840 5216
rect 7607 5185 7619 5188
rect 7561 5179 7619 5185
rect 7834 5176 7840 5188
rect 7892 5216 7898 5228
rect 8036 5216 8064 5315
rect 10962 5312 10968 5324
rect 11020 5312 11026 5364
rect 11790 5312 11796 5364
rect 11848 5352 11854 5364
rect 12342 5352 12348 5364
rect 11848 5324 12348 5352
rect 11848 5312 11854 5324
rect 12342 5312 12348 5324
rect 12400 5352 12406 5364
rect 13173 5355 13231 5361
rect 12400 5324 13124 5352
rect 12400 5312 12406 5324
rect 9214 5284 9220 5296
rect 9062 5256 9220 5284
rect 9214 5244 9220 5256
rect 9272 5244 9278 5296
rect 9950 5284 9956 5296
rect 9911 5256 9956 5284
rect 9950 5244 9956 5256
rect 10008 5244 10014 5296
rect 10137 5287 10195 5293
rect 10137 5253 10149 5287
rect 10183 5284 10195 5287
rect 10410 5284 10416 5296
rect 10183 5256 10416 5284
rect 10183 5253 10195 5256
rect 10137 5247 10195 5253
rect 10410 5244 10416 5256
rect 10468 5244 10474 5296
rect 12360 5270 12388 5312
rect 13096 5284 13124 5324
rect 13173 5321 13185 5355
rect 13219 5352 13231 5355
rect 13446 5352 13452 5364
rect 13219 5324 13452 5352
rect 13219 5321 13231 5324
rect 13173 5315 13231 5321
rect 13446 5312 13452 5324
rect 13504 5312 13510 5364
rect 13814 5312 13820 5364
rect 13872 5352 13878 5364
rect 14734 5352 14740 5364
rect 13872 5324 14740 5352
rect 13872 5312 13878 5324
rect 14734 5312 14740 5324
rect 14792 5312 14798 5364
rect 16669 5355 16727 5361
rect 16669 5321 16681 5355
rect 16715 5352 16727 5355
rect 17678 5352 17684 5364
rect 16715 5324 17684 5352
rect 16715 5321 16727 5324
rect 16669 5315 16727 5321
rect 17678 5312 17684 5324
rect 17736 5312 17742 5364
rect 17862 5312 17868 5364
rect 17920 5352 17926 5364
rect 18509 5355 18567 5361
rect 18509 5352 18521 5355
rect 17920 5324 18521 5352
rect 17920 5312 17926 5324
rect 18509 5321 18521 5324
rect 18555 5321 18567 5355
rect 18509 5315 18567 5321
rect 14366 5290 14372 5296
rect 14292 5284 14372 5290
rect 13096 5262 14372 5284
rect 13096 5256 14306 5262
rect 14366 5244 14372 5262
rect 14424 5244 14430 5296
rect 16022 5244 16028 5296
rect 16080 5284 16086 5296
rect 16080 5256 16804 5284
rect 16080 5244 16086 5256
rect 7892 5188 8064 5216
rect 10229 5219 10287 5225
rect 7892 5176 7898 5188
rect 10229 5185 10241 5219
rect 10275 5216 10287 5219
rect 10275 5188 10456 5216
rect 10275 5185 10287 5188
rect 10229 5179 10287 5185
rect 3513 5151 3571 5157
rect 3513 5117 3525 5151
rect 3559 5148 3571 5151
rect 3694 5148 3700 5160
rect 3559 5120 3700 5148
rect 3559 5117 3571 5120
rect 3513 5111 3571 5117
rect 3694 5108 3700 5120
rect 3752 5108 3758 5160
rect 5810 5148 5816 5160
rect 5771 5120 5816 5148
rect 5810 5108 5816 5120
rect 5868 5108 5874 5160
rect 6273 5151 6331 5157
rect 6273 5117 6285 5151
rect 6319 5148 6331 5151
rect 6822 5148 6828 5160
rect 6319 5120 6828 5148
rect 6319 5117 6331 5120
rect 6273 5111 6331 5117
rect 6822 5108 6828 5120
rect 6880 5108 6886 5160
rect 7650 5148 7656 5160
rect 7611 5120 7656 5148
rect 7650 5108 7656 5120
rect 7708 5108 7714 5160
rect 7929 5151 7987 5157
rect 7929 5117 7941 5151
rect 7975 5148 7987 5151
rect 9493 5151 9551 5157
rect 9493 5148 9505 5151
rect 7975 5120 9505 5148
rect 7975 5117 7987 5120
rect 7929 5111 7987 5117
rect 9493 5117 9505 5120
rect 9539 5117 9551 5151
rect 9766 5148 9772 5160
rect 9727 5120 9772 5148
rect 9493 5111 9551 5117
rect 9766 5108 9772 5120
rect 9824 5108 9830 5160
rect 10428 5157 10456 5188
rect 10594 5176 10600 5228
rect 10652 5216 10658 5228
rect 10873 5219 10931 5225
rect 10873 5216 10885 5219
rect 10652 5188 10885 5216
rect 10652 5176 10658 5188
rect 10873 5185 10885 5188
rect 10919 5185 10931 5219
rect 10873 5179 10931 5185
rect 11054 5176 11060 5228
rect 11112 5216 11118 5228
rect 11149 5219 11207 5225
rect 11149 5216 11161 5219
rect 11112 5188 11161 5216
rect 11112 5176 11118 5188
rect 11149 5185 11161 5188
rect 11195 5216 11207 5219
rect 13081 5219 13139 5225
rect 13081 5216 13093 5219
rect 11195 5188 11652 5216
rect 11195 5185 11207 5188
rect 11149 5179 11207 5185
rect 10413 5151 10471 5157
rect 10413 5117 10425 5151
rect 10459 5117 10471 5151
rect 11514 5148 11520 5160
rect 11475 5120 11520 5148
rect 10413 5111 10471 5117
rect 11514 5108 11520 5120
rect 11572 5108 11578 5160
rect 11624 5148 11652 5188
rect 12452 5188 13093 5216
rect 12452 5160 12480 5188
rect 13081 5185 13093 5188
rect 13127 5216 13139 5219
rect 13354 5216 13360 5228
rect 13127 5188 13360 5216
rect 13127 5185 13139 5188
rect 13081 5179 13139 5185
rect 13354 5176 13360 5188
rect 13412 5176 13418 5228
rect 13538 5216 13544 5228
rect 13499 5188 13544 5216
rect 13538 5176 13544 5188
rect 13596 5176 13602 5228
rect 16298 5216 16304 5228
rect 16259 5188 16304 5216
rect 16298 5176 16304 5188
rect 16356 5176 16362 5228
rect 16776 5225 16804 5256
rect 16942 5244 16948 5296
rect 17000 5284 17006 5296
rect 17000 5256 17526 5284
rect 17000 5244 17006 5256
rect 16761 5219 16819 5225
rect 16761 5185 16773 5219
rect 16807 5185 16819 5219
rect 16761 5179 16819 5185
rect 12342 5148 12348 5160
rect 11624 5120 12348 5148
rect 12342 5108 12348 5120
rect 12400 5108 12406 5160
rect 12434 5108 12440 5160
rect 12492 5108 12498 5160
rect 13817 5151 13875 5157
rect 13817 5117 13829 5151
rect 13863 5148 13875 5151
rect 16390 5148 16396 5160
rect 13863 5120 16160 5148
rect 16351 5120 16396 5148
rect 13863 5117 13875 5120
rect 13817 5111 13875 5117
rect 12943 5083 13001 5089
rect 12943 5080 12955 5083
rect 12406 5052 12955 5080
rect 10778 5012 10784 5024
rect 10739 4984 10784 5012
rect 10778 4972 10784 4984
rect 10836 4972 10842 5024
rect 11974 4972 11980 5024
rect 12032 5012 12038 5024
rect 12406 5012 12434 5052
rect 12943 5049 12955 5052
rect 12989 5080 13001 5083
rect 13354 5080 13360 5092
rect 12989 5052 13360 5080
rect 12989 5049 13001 5052
rect 12943 5043 13001 5049
rect 13354 5040 13360 5052
rect 13412 5040 13418 5092
rect 16132 5080 16160 5120
rect 16390 5108 16396 5120
rect 16448 5108 16454 5160
rect 17034 5148 17040 5160
rect 16995 5120 17040 5148
rect 17034 5108 17040 5120
rect 17092 5108 17098 5160
rect 16758 5080 16764 5092
rect 16132 5052 16764 5080
rect 16758 5040 16764 5052
rect 16816 5040 16822 5092
rect 12032 4984 12434 5012
rect 15289 5015 15347 5021
rect 12032 4972 12038 4984
rect 15289 4981 15301 5015
rect 15335 5012 15347 5015
rect 17218 5012 17224 5024
rect 15335 4984 17224 5012
rect 15335 4981 15347 4984
rect 15289 4975 15347 4981
rect 17218 4972 17224 4984
rect 17276 4972 17282 5024
rect 0 4922 18860 4944
rect 0 4870 2995 4922
rect 3047 4870 3059 4922
rect 3111 4870 3123 4922
rect 3175 4870 3187 4922
rect 3239 4870 3251 4922
rect 3303 4870 9294 4922
rect 9346 4870 9358 4922
rect 9410 4870 9422 4922
rect 9474 4870 9486 4922
rect 9538 4870 9550 4922
rect 9602 4870 15592 4922
rect 15644 4870 15656 4922
rect 15708 4870 15720 4922
rect 15772 4870 15784 4922
rect 15836 4870 15848 4922
rect 15900 4870 18860 4922
rect 0 4848 18860 4870
rect 7650 4768 7656 4820
rect 7708 4808 7714 4820
rect 7929 4811 7987 4817
rect 7929 4808 7941 4811
rect 7708 4780 7941 4808
rect 7708 4768 7714 4780
rect 7929 4777 7941 4780
rect 7975 4777 7987 4811
rect 7929 4771 7987 4777
rect 11514 4768 11520 4820
rect 11572 4808 11578 4820
rect 11701 4811 11759 4817
rect 11701 4808 11713 4811
rect 11572 4780 11713 4808
rect 11572 4768 11578 4780
rect 11701 4777 11713 4780
rect 11747 4777 11759 4811
rect 11701 4771 11759 4777
rect 12342 4768 12348 4820
rect 12400 4808 12406 4820
rect 12526 4808 12532 4820
rect 12400 4780 12532 4808
rect 12400 4768 12406 4780
rect 12526 4768 12532 4780
rect 12584 4768 12590 4820
rect 12713 4811 12771 4817
rect 12713 4777 12725 4811
rect 12759 4808 12771 4811
rect 12802 4808 12808 4820
rect 12759 4780 12808 4808
rect 12759 4777 12771 4780
rect 12713 4771 12771 4777
rect 12802 4768 12808 4780
rect 12860 4768 12866 4820
rect 14185 4811 14243 4817
rect 14185 4777 14197 4811
rect 14231 4808 14243 4811
rect 14274 4808 14280 4820
rect 14231 4780 14280 4808
rect 14231 4777 14243 4780
rect 14185 4771 14243 4777
rect 14274 4768 14280 4780
rect 14332 4768 14338 4820
rect 14458 4808 14464 4820
rect 14419 4780 14464 4808
rect 14458 4768 14464 4780
rect 14516 4768 14522 4820
rect 14550 4768 14556 4820
rect 14608 4808 14614 4820
rect 14921 4811 14979 4817
rect 14921 4808 14933 4811
rect 14608 4780 14933 4808
rect 14608 4768 14614 4780
rect 14921 4777 14933 4780
rect 14967 4777 14979 4811
rect 14921 4771 14979 4777
rect 15749 4811 15807 4817
rect 15749 4777 15761 4811
rect 15795 4808 15807 4811
rect 17034 4808 17040 4820
rect 15795 4780 17040 4808
rect 15795 4777 15807 4780
rect 15749 4771 15807 4777
rect 17034 4768 17040 4780
rect 17092 4768 17098 4820
rect 7374 4700 7380 4752
rect 7432 4740 7438 4752
rect 7561 4743 7619 4749
rect 7561 4740 7573 4743
rect 7432 4712 7573 4740
rect 7432 4700 7438 4712
rect 7561 4709 7573 4712
rect 7607 4740 7619 4743
rect 8018 4740 8024 4752
rect 7607 4712 8024 4740
rect 7607 4709 7619 4712
rect 7561 4703 7619 4709
rect 8018 4700 8024 4712
rect 8076 4740 8082 4752
rect 8076 4712 8524 4740
rect 8076 4700 8082 4712
rect 5534 4564 5540 4616
rect 5592 4604 5598 4616
rect 5813 4607 5871 4613
rect 5813 4604 5825 4607
rect 5592 4576 5825 4604
rect 5592 4564 5598 4576
rect 5813 4573 5825 4576
rect 5859 4573 5871 4607
rect 5813 4567 5871 4573
rect 8113 4607 8171 4613
rect 8113 4573 8125 4607
rect 8159 4604 8171 4607
rect 8294 4604 8300 4616
rect 8159 4576 8300 4604
rect 8159 4573 8171 4576
rect 8113 4567 8171 4573
rect 8294 4564 8300 4576
rect 8352 4564 8358 4616
rect 8496 4613 8524 4712
rect 9030 4700 9036 4752
rect 9088 4740 9094 4752
rect 10229 4743 10287 4749
rect 10229 4740 10241 4743
rect 9088 4712 10241 4740
rect 9088 4700 9094 4712
rect 10229 4709 10241 4712
rect 10275 4740 10287 4743
rect 15378 4740 15384 4752
rect 10275 4712 12388 4740
rect 10275 4709 10287 4712
rect 10229 4703 10287 4709
rect 8570 4632 8576 4684
rect 8628 4672 8634 4684
rect 9585 4675 9643 4681
rect 8628 4644 8673 4672
rect 8628 4632 8634 4644
rect 9585 4641 9597 4675
rect 9631 4672 9643 4675
rect 9950 4672 9956 4684
rect 9631 4644 9956 4672
rect 9631 4641 9643 4644
rect 9585 4635 9643 4641
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 10870 4632 10876 4684
rect 10928 4672 10934 4684
rect 11885 4675 11943 4681
rect 11885 4672 11897 4675
rect 10928 4644 11897 4672
rect 10928 4632 10934 4644
rect 11885 4641 11897 4644
rect 11931 4641 11943 4675
rect 11885 4635 11943 4641
rect 8481 4607 8539 4613
rect 8481 4573 8493 4607
rect 8527 4573 8539 4607
rect 9214 4604 9220 4616
rect 8481 4567 8539 4573
rect 8588 4576 9220 4604
rect 5994 4496 6000 4548
rect 6052 4536 6058 4548
rect 6089 4539 6147 4545
rect 6089 4536 6101 4539
rect 6052 4508 6101 4536
rect 6052 4496 6058 4508
rect 6089 4505 6101 4508
rect 6135 4505 6147 4539
rect 6089 4499 6147 4505
rect 7300 4468 7328 4522
rect 7558 4496 7564 4548
rect 7616 4536 7622 4548
rect 7837 4539 7895 4545
rect 7837 4536 7849 4539
rect 7616 4508 7849 4536
rect 7616 4496 7622 4508
rect 7837 4505 7849 4508
rect 7883 4536 7895 4539
rect 8202 4536 8208 4548
rect 7883 4508 8208 4536
rect 7883 4505 7895 4508
rect 7837 4499 7895 4505
rect 8202 4496 8208 4508
rect 8260 4496 8266 4548
rect 8294 4468 8300 4480
rect 7300 4440 8300 4468
rect 8294 4428 8300 4440
rect 8352 4468 8358 4480
rect 8588 4468 8616 4576
rect 9214 4564 9220 4576
rect 9272 4564 9278 4616
rect 11974 4604 11980 4616
rect 11935 4576 11980 4604
rect 11974 4564 11980 4576
rect 12032 4564 12038 4616
rect 12360 4613 12388 4712
rect 12452 4712 15384 4740
rect 12345 4607 12403 4613
rect 12345 4573 12357 4607
rect 12391 4573 12403 4607
rect 12345 4567 12403 4573
rect 9401 4539 9459 4545
rect 9401 4536 9413 4539
rect 8864 4508 9413 4536
rect 8864 4477 8892 4508
rect 9401 4505 9413 4508
rect 9447 4505 9459 4539
rect 9401 4499 9459 4505
rect 11517 4539 11575 4545
rect 11517 4505 11529 4539
rect 11563 4536 11575 4539
rect 12452 4536 12480 4712
rect 15378 4700 15384 4712
rect 15436 4700 15442 4752
rect 18325 4743 18383 4749
rect 18325 4709 18337 4743
rect 18371 4709 18383 4743
rect 18325 4703 18383 4709
rect 13078 4672 13084 4684
rect 12636 4644 13084 4672
rect 12636 4613 12664 4644
rect 13078 4632 13084 4644
rect 13136 4632 13142 4684
rect 13633 4675 13691 4681
rect 13188 4644 13492 4672
rect 12621 4607 12679 4613
rect 12621 4573 12633 4607
rect 12667 4573 12679 4607
rect 12621 4567 12679 4573
rect 12805 4607 12863 4613
rect 12805 4573 12817 4607
rect 12851 4604 12863 4607
rect 13188 4604 13216 4644
rect 13354 4604 13360 4616
rect 12851 4576 13216 4604
rect 13315 4576 13360 4604
rect 12851 4573 12863 4576
rect 12805 4567 12863 4573
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 13464 4604 13492 4644
rect 13633 4641 13645 4675
rect 13679 4672 13691 4675
rect 13909 4675 13967 4681
rect 13909 4672 13921 4675
rect 13679 4644 13921 4672
rect 13679 4641 13691 4644
rect 13633 4635 13691 4641
rect 13909 4641 13921 4644
rect 13955 4641 13967 4675
rect 15194 4672 15200 4684
rect 13909 4635 13967 4641
rect 14016 4644 15200 4672
rect 13722 4604 13728 4616
rect 13464 4576 13728 4604
rect 13722 4564 13728 4576
rect 13780 4564 13786 4616
rect 14016 4613 14044 4644
rect 15194 4632 15200 4644
rect 15252 4632 15258 4684
rect 15473 4675 15531 4681
rect 15473 4641 15485 4675
rect 15519 4672 15531 4675
rect 16206 4672 16212 4684
rect 15519 4644 16212 4672
rect 15519 4641 15531 4644
rect 15473 4635 15531 4641
rect 16206 4632 16212 4644
rect 16264 4632 16270 4684
rect 16758 4632 16764 4684
rect 16816 4672 16822 4684
rect 18340 4672 18368 4703
rect 16816 4644 18368 4672
rect 16816 4632 16822 4644
rect 13817 4607 13875 4613
rect 13817 4573 13829 4607
rect 13863 4604 13875 4607
rect 13995 4607 14053 4613
rect 13863 4576 13952 4604
rect 13863 4573 13875 4576
rect 13817 4567 13875 4573
rect 11563 4508 12480 4536
rect 11563 4505 11575 4508
rect 11517 4499 11575 4505
rect 12526 4496 12532 4548
rect 12584 4536 12590 4548
rect 13924 4536 13952 4576
rect 13995 4573 14007 4607
rect 14041 4573 14053 4607
rect 13995 4567 14053 4573
rect 14085 4609 14143 4615
rect 14085 4575 14097 4609
rect 14131 4604 14143 4609
rect 14182 4604 14188 4616
rect 14131 4576 14188 4604
rect 14131 4575 14143 4576
rect 14085 4569 14143 4575
rect 14182 4564 14188 4576
rect 14240 4564 14246 4616
rect 14369 4607 14427 4613
rect 14369 4573 14381 4607
rect 14415 4573 14427 4607
rect 14918 4604 14924 4616
rect 14879 4576 14924 4604
rect 14369 4567 14427 4573
rect 14384 4536 14412 4567
rect 14918 4564 14924 4576
rect 14976 4564 14982 4616
rect 15102 4604 15108 4616
rect 15063 4576 15108 4604
rect 15102 4564 15108 4576
rect 15160 4564 15166 4616
rect 15381 4607 15439 4613
rect 15381 4573 15393 4607
rect 15427 4604 15439 4607
rect 16666 4604 16672 4616
rect 15427 4576 16672 4604
rect 15427 4573 15439 4576
rect 15381 4567 15439 4573
rect 16666 4564 16672 4576
rect 16724 4564 16730 4616
rect 17586 4604 17592 4616
rect 17547 4576 17592 4604
rect 17586 4564 17592 4576
rect 17644 4564 17650 4616
rect 17954 4604 17960 4616
rect 17915 4576 17960 4604
rect 17954 4564 17960 4576
rect 18012 4564 18018 4616
rect 18506 4604 18512 4616
rect 18467 4576 18512 4604
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 12584 4508 13492 4536
rect 13924 4508 15148 4536
rect 12584 4496 12590 4508
rect 8352 4440 8616 4468
rect 8849 4471 8907 4477
rect 8352 4428 8358 4440
rect 8849 4437 8861 4471
rect 8895 4437 8907 4471
rect 8849 4431 8907 4437
rect 8938 4428 8944 4480
rect 8996 4468 9002 4480
rect 8996 4440 9041 4468
rect 8996 4428 9002 4440
rect 9122 4428 9128 4480
rect 9180 4468 9186 4480
rect 9309 4471 9367 4477
rect 9309 4468 9321 4471
rect 9180 4440 9321 4468
rect 9180 4428 9186 4440
rect 9309 4437 9321 4440
rect 9355 4437 9367 4471
rect 12986 4468 12992 4480
rect 12947 4440 12992 4468
rect 9309 4431 9367 4437
rect 12986 4428 12992 4440
rect 13044 4428 13050 4480
rect 13464 4477 13492 4508
rect 15120 4480 15148 4508
rect 16960 4480 16988 4522
rect 13449 4471 13507 4477
rect 13449 4437 13461 4471
rect 13495 4468 13507 4471
rect 13998 4468 14004 4480
rect 13495 4440 14004 4468
rect 13495 4437 13507 4440
rect 13449 4431 13507 4437
rect 13998 4428 14004 4440
rect 14056 4428 14062 4480
rect 14829 4471 14887 4477
rect 14829 4437 14841 4471
rect 14875 4468 14887 4471
rect 14918 4468 14924 4480
rect 14875 4440 14924 4468
rect 14875 4437 14887 4440
rect 14829 4431 14887 4437
rect 14918 4428 14924 4440
rect 14976 4428 14982 4480
rect 15102 4428 15108 4480
rect 15160 4468 15166 4480
rect 15841 4471 15899 4477
rect 15841 4468 15853 4471
rect 15160 4440 15853 4468
rect 15160 4428 15166 4440
rect 15841 4437 15853 4440
rect 15887 4468 15899 4471
rect 16298 4468 16304 4480
rect 15887 4440 16304 4468
rect 15887 4437 15899 4440
rect 15841 4431 15899 4437
rect 16298 4428 16304 4440
rect 16356 4428 16362 4480
rect 16942 4428 16948 4480
rect 17000 4428 17006 4480
rect 0 4378 18860 4400
rect 0 4326 6144 4378
rect 6196 4326 6208 4378
rect 6260 4326 6272 4378
rect 6324 4326 6336 4378
rect 6388 4326 6400 4378
rect 6452 4326 12443 4378
rect 12495 4326 12507 4378
rect 12559 4326 12571 4378
rect 12623 4326 12635 4378
rect 12687 4326 12699 4378
rect 12751 4326 18860 4378
rect 0 4304 18860 4326
rect 5994 4224 6000 4276
rect 6052 4264 6058 4276
rect 6365 4267 6423 4273
rect 6365 4264 6377 4267
rect 6052 4236 6377 4264
rect 6052 4224 6058 4236
rect 6365 4233 6377 4236
rect 6411 4233 6423 4267
rect 7374 4264 7380 4276
rect 7335 4236 7380 4264
rect 6365 4227 6423 4233
rect 7374 4224 7380 4236
rect 7432 4224 7438 4276
rect 8389 4267 8447 4273
rect 8389 4233 8401 4267
rect 8435 4264 8447 4267
rect 9309 4267 9367 4273
rect 9309 4264 9321 4267
rect 8435 4236 9321 4264
rect 8435 4233 8447 4236
rect 8389 4227 8447 4233
rect 9309 4233 9321 4236
rect 9355 4233 9367 4267
rect 9309 4227 9367 4233
rect 10686 4224 10692 4276
rect 10744 4264 10750 4276
rect 13909 4267 13967 4273
rect 10744 4236 11468 4264
rect 10744 4224 10750 4236
rect 7285 4199 7343 4205
rect 7285 4165 7297 4199
rect 7331 4196 7343 4199
rect 8846 4196 8852 4208
rect 7331 4168 8852 4196
rect 7331 4165 7343 4168
rect 7285 4159 7343 4165
rect 8846 4156 8852 4168
rect 8904 4156 8910 4208
rect 9030 4196 9036 4208
rect 8991 4168 9036 4196
rect 9030 4156 9036 4168
rect 9088 4156 9094 4208
rect 10594 4156 10600 4208
rect 10652 4156 10658 4208
rect 10870 4156 10876 4208
rect 10928 4196 10934 4208
rect 10928 4168 10973 4196
rect 10928 4156 10934 4168
rect 10597 4153 10655 4156
rect 6549 4131 6607 4137
rect 6549 4097 6561 4131
rect 6595 4128 6607 4131
rect 7745 4131 7803 4137
rect 6595 4100 6960 4128
rect 6595 4097 6607 4100
rect 6549 4091 6607 4097
rect 6932 4001 6960 4100
rect 7745 4097 7757 4131
rect 7791 4128 7803 4131
rect 8478 4128 8484 4140
rect 7791 4100 8064 4128
rect 8439 4100 8484 4128
rect 7791 4097 7803 4100
rect 7745 4091 7803 4097
rect 7558 4060 7564 4072
rect 7519 4032 7564 4060
rect 7558 4020 7564 4032
rect 7616 4020 7622 4072
rect 8036 4001 8064 4100
rect 8478 4088 8484 4100
rect 8536 4088 8542 4140
rect 9674 4128 9680 4140
rect 9635 4100 9680 4128
rect 9674 4088 9680 4100
rect 9732 4088 9738 4140
rect 10410 4088 10416 4140
rect 10468 4137 10474 4140
rect 10468 4131 10527 4137
rect 10468 4097 10481 4131
rect 10515 4097 10527 4131
rect 10597 4119 10609 4153
rect 10643 4119 10655 4153
rect 10597 4113 10655 4119
rect 10468 4091 10527 4097
rect 10468 4088 10474 4091
rect 10686 4078 10692 4130
rect 10744 4118 10750 4130
rect 11054 4128 11060 4140
rect 10744 4090 10789 4118
rect 11015 4100 11060 4128
rect 10744 4078 10750 4090
rect 11054 4088 11060 4100
rect 11112 4088 11118 4140
rect 11440 4137 11468 4236
rect 11900 4236 13124 4264
rect 11514 4156 11520 4208
rect 11572 4196 11578 4208
rect 11900 4205 11928 4236
rect 11885 4199 11943 4205
rect 11885 4196 11897 4199
rect 11572 4168 11897 4196
rect 11572 4156 11578 4168
rect 11885 4165 11897 4168
rect 11931 4165 11943 4199
rect 12986 4196 12992 4208
rect 11885 4159 11943 4165
rect 12636 4168 12992 4196
rect 11425 4131 11483 4137
rect 11425 4097 11437 4131
rect 11471 4097 11483 4131
rect 11425 4091 11483 4097
rect 11609 4131 11667 4137
rect 11609 4097 11621 4131
rect 11655 4097 11667 4131
rect 11609 4091 11667 4097
rect 8202 4020 8208 4072
rect 8260 4060 8266 4072
rect 8665 4063 8723 4069
rect 8665 4060 8677 4063
rect 8260 4032 8677 4060
rect 8260 4020 8266 4032
rect 8665 4029 8677 4032
rect 8711 4060 8723 4063
rect 9214 4060 9220 4072
rect 8711 4032 9220 4060
rect 8711 4029 8723 4032
rect 8665 4023 8723 4029
rect 9214 4020 9220 4032
rect 9272 4020 9278 4072
rect 9769 4063 9827 4069
rect 9769 4029 9781 4063
rect 9815 4029 9827 4063
rect 9769 4023 9827 4029
rect 6917 3995 6975 4001
rect 6917 3961 6929 3995
rect 6963 3961 6975 3995
rect 6917 3955 6975 3961
rect 8021 3995 8079 4001
rect 8021 3961 8033 3995
rect 8067 3961 8079 3995
rect 9784 3992 9812 4023
rect 9950 4020 9956 4072
rect 10008 4060 10014 4072
rect 10137 4063 10195 4069
rect 10137 4060 10149 4063
rect 10008 4032 10149 4060
rect 10008 4020 10014 4032
rect 10137 4029 10149 4032
rect 10183 4029 10195 4063
rect 11072 4060 11100 4088
rect 11624 4060 11652 4091
rect 12434 4088 12440 4140
rect 12492 4128 12498 4140
rect 12529 4131 12587 4137
rect 12529 4128 12541 4131
rect 12492 4100 12541 4128
rect 12492 4088 12498 4100
rect 12529 4097 12541 4100
rect 12575 4097 12587 4131
rect 12529 4091 12587 4097
rect 12636 4060 12664 4168
rect 12986 4156 12992 4168
rect 13044 4156 13050 4208
rect 13096 4140 13124 4236
rect 13909 4233 13921 4267
rect 13955 4264 13967 4267
rect 14458 4264 14464 4276
rect 13955 4236 14464 4264
rect 13955 4233 13967 4236
rect 13909 4227 13967 4233
rect 14458 4224 14464 4236
rect 14516 4224 14522 4276
rect 16942 4224 16948 4276
rect 17000 4224 17006 4276
rect 13446 4156 13452 4208
rect 13504 4196 13510 4208
rect 15194 4196 15200 4208
rect 13504 4168 15200 4196
rect 13504 4156 13510 4168
rect 15194 4156 15200 4168
rect 15252 4196 15258 4208
rect 15565 4199 15623 4205
rect 15565 4196 15577 4199
rect 15252 4168 15577 4196
rect 15252 4156 15258 4168
rect 15565 4165 15577 4168
rect 15611 4165 15623 4199
rect 16960 4196 16988 4224
rect 16882 4168 16988 4196
rect 15565 4159 15623 4165
rect 12802 4137 12808 4140
rect 12796 4128 12808 4137
rect 12763 4100 12808 4128
rect 12796 4091 12808 4100
rect 12802 4088 12808 4091
rect 12860 4088 12866 4140
rect 13078 4088 13084 4140
rect 13136 4128 13142 4140
rect 14268 4131 14326 4137
rect 14268 4128 14280 4131
rect 13136 4100 14280 4128
rect 13136 4088 13142 4100
rect 14268 4097 14280 4100
rect 14314 4128 14326 4131
rect 18506 4128 18512 4140
rect 14314 4100 15516 4128
rect 18467 4100 18512 4128
rect 14314 4097 14326 4100
rect 14268 4091 14326 4097
rect 13998 4060 14004 4072
rect 11072 4032 11652 4060
rect 12268 4032 12664 4060
rect 13959 4032 14004 4060
rect 10137 4023 10195 4029
rect 12268 4001 12296 4032
rect 13998 4020 14004 4032
rect 14056 4020 14062 4072
rect 11057 3995 11115 4001
rect 11057 3992 11069 3995
rect 9784 3964 11069 3992
rect 8021 3955 8079 3961
rect 11057 3961 11069 3964
rect 11103 3961 11115 3995
rect 11057 3955 11115 3961
rect 12253 3995 12311 4001
rect 12253 3961 12265 3995
rect 12299 3961 12311 3995
rect 12253 3955 12311 3961
rect 7929 3927 7987 3933
rect 7929 3893 7941 3927
rect 7975 3924 7987 3927
rect 8202 3924 8208 3936
rect 7975 3896 8208 3924
rect 7975 3893 7987 3896
rect 7929 3887 7987 3893
rect 8202 3884 8208 3896
rect 8260 3884 8266 3936
rect 8938 3924 8944 3936
rect 8899 3896 8944 3924
rect 8938 3884 8944 3896
rect 8996 3884 9002 3936
rect 10137 3927 10195 3933
rect 10137 3893 10149 3927
rect 10183 3924 10195 3927
rect 11517 3927 11575 3933
rect 11517 3924 11529 3927
rect 10183 3896 11529 3924
rect 10183 3893 10195 3896
rect 10137 3887 10195 3893
rect 11517 3893 11529 3896
rect 11563 3893 11575 3927
rect 11517 3887 11575 3893
rect 12345 3927 12403 3933
rect 12345 3893 12357 3927
rect 12391 3924 12403 3927
rect 12894 3924 12900 3936
rect 12391 3896 12900 3924
rect 12391 3893 12403 3896
rect 12345 3887 12403 3893
rect 12894 3884 12900 3896
rect 12952 3884 12958 3936
rect 15194 3884 15200 3936
rect 15252 3924 15258 3936
rect 15381 3927 15439 3933
rect 15381 3924 15393 3927
rect 15252 3896 15393 3924
rect 15252 3884 15258 3896
rect 15381 3893 15393 3896
rect 15427 3893 15439 3927
rect 15488 3924 15516 4100
rect 18506 4088 18512 4100
rect 18564 4088 18570 4140
rect 17218 4020 17224 4072
rect 17276 4060 17282 4072
rect 17313 4063 17371 4069
rect 17313 4060 17325 4063
rect 17276 4032 17325 4060
rect 17276 4020 17282 4032
rect 17313 4029 17325 4032
rect 17359 4029 17371 4063
rect 17313 4023 17371 4029
rect 17589 4063 17647 4069
rect 17589 4029 17601 4063
rect 17635 4060 17647 4063
rect 17954 4060 17960 4072
rect 17635 4032 17960 4060
rect 17635 4029 17647 4032
rect 17589 4023 17647 4029
rect 17954 4020 17960 4032
rect 18012 4020 18018 4072
rect 18046 3924 18052 3936
rect 15488 3896 18052 3924
rect 15381 3887 15439 3893
rect 18046 3884 18052 3896
rect 18104 3884 18110 3936
rect 18325 3927 18383 3933
rect 18325 3893 18337 3927
rect 18371 3924 18383 3927
rect 18969 3927 19027 3933
rect 18969 3924 18981 3927
rect 18371 3896 18981 3924
rect 18371 3893 18383 3896
rect 18325 3887 18383 3893
rect 18969 3893 18981 3896
rect 19015 3893 19027 3927
rect 18969 3887 19027 3893
rect 0 3834 18860 3856
rect 0 3782 2995 3834
rect 3047 3782 3059 3834
rect 3111 3782 3123 3834
rect 3175 3782 3187 3834
rect 3239 3782 3251 3834
rect 3303 3782 9294 3834
rect 9346 3782 9358 3834
rect 9410 3782 9422 3834
rect 9474 3782 9486 3834
rect 9538 3782 9550 3834
rect 9602 3782 15592 3834
rect 15644 3782 15656 3834
rect 15708 3782 15720 3834
rect 15772 3782 15784 3834
rect 15836 3782 15848 3834
rect 15900 3782 18860 3834
rect 0 3760 18860 3782
rect 5902 3720 5908 3732
rect 5092 3692 5908 3720
rect 5092 3593 5120 3692
rect 5902 3680 5908 3692
rect 5960 3680 5966 3732
rect 8478 3680 8484 3732
rect 8536 3720 8542 3732
rect 9585 3723 9643 3729
rect 9585 3720 9597 3723
rect 8536 3692 9597 3720
rect 8536 3680 8542 3692
rect 9585 3689 9597 3692
rect 9631 3720 9643 3723
rect 10594 3720 10600 3732
rect 9631 3692 10600 3720
rect 9631 3689 9643 3692
rect 9585 3683 9643 3689
rect 10594 3680 10600 3692
rect 10652 3720 10658 3732
rect 11054 3720 11060 3732
rect 10652 3692 11060 3720
rect 10652 3680 10658 3692
rect 11054 3680 11060 3692
rect 11112 3680 11118 3732
rect 11624 3692 12848 3720
rect 5258 3652 5264 3664
rect 5219 3624 5264 3652
rect 5258 3612 5264 3624
rect 5316 3612 5322 3664
rect 5077 3587 5135 3593
rect 5077 3553 5089 3587
rect 5123 3553 5135 3587
rect 5445 3587 5503 3593
rect 5445 3584 5457 3587
rect 5077 3547 5135 3553
rect 5184 3556 5457 3584
rect 3326 3476 3332 3528
rect 3384 3516 3390 3528
rect 3513 3519 3571 3525
rect 3513 3516 3525 3519
rect 3384 3488 3525 3516
rect 3384 3476 3390 3488
rect 3513 3485 3525 3488
rect 3559 3516 3571 3519
rect 5184 3516 5212 3556
rect 5445 3553 5457 3556
rect 5491 3584 5503 3587
rect 7837 3587 7895 3593
rect 7837 3584 7849 3587
rect 5491 3556 7849 3584
rect 5491 3553 5503 3556
rect 5445 3547 5503 3553
rect 7837 3553 7849 3556
rect 7883 3584 7895 3587
rect 8938 3584 8944 3596
rect 7883 3556 8944 3584
rect 7883 3553 7895 3556
rect 7837 3547 7895 3553
rect 5350 3516 5356 3528
rect 3559 3488 5212 3516
rect 5311 3488 5356 3516
rect 3559 3485 3571 3488
rect 3513 3479 3571 3485
rect 5350 3476 5356 3488
rect 5408 3476 5414 3528
rect 5460 3448 5488 3547
rect 8938 3544 8944 3556
rect 8996 3544 9002 3596
rect 8202 3516 8208 3528
rect 8163 3488 8208 3516
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 8956 3516 8984 3544
rect 9766 3516 9772 3528
rect 8956 3488 9772 3516
rect 9766 3476 9772 3488
rect 9824 3516 9830 3528
rect 9953 3519 10011 3525
rect 9953 3516 9965 3519
rect 9824 3488 9965 3516
rect 9824 3476 9830 3488
rect 9953 3485 9965 3488
rect 9999 3516 10011 3519
rect 10321 3519 10379 3525
rect 10321 3516 10333 3519
rect 9999 3488 10333 3516
rect 9999 3485 10011 3488
rect 9953 3479 10011 3485
rect 10321 3485 10333 3488
rect 10367 3485 10379 3519
rect 10321 3479 10379 3485
rect 10588 3519 10646 3525
rect 10588 3485 10600 3519
rect 10634 3516 10646 3519
rect 11624 3516 11652 3692
rect 11701 3655 11759 3661
rect 11701 3621 11713 3655
rect 11747 3652 11759 3655
rect 11747 3624 12664 3652
rect 11747 3621 11759 3624
rect 11701 3615 11759 3621
rect 11793 3519 11851 3525
rect 11793 3516 11805 3519
rect 10634 3488 11805 3516
rect 10634 3485 10646 3488
rect 10588 3479 10646 3485
rect 11793 3485 11805 3488
rect 11839 3516 11851 3519
rect 11882 3516 11888 3528
rect 11839 3488 11888 3516
rect 11839 3485 11851 3488
rect 11793 3479 11851 3485
rect 11882 3476 11888 3488
rect 11940 3476 11946 3528
rect 11992 3525 12020 3624
rect 12161 3587 12219 3593
rect 12161 3553 12173 3587
rect 12207 3584 12219 3587
rect 12345 3587 12403 3593
rect 12345 3584 12357 3587
rect 12207 3556 12357 3584
rect 12207 3553 12219 3556
rect 12161 3547 12219 3553
rect 12345 3553 12357 3556
rect 12391 3553 12403 3587
rect 12526 3584 12532 3596
rect 12487 3556 12532 3584
rect 12345 3547 12403 3553
rect 12526 3544 12532 3556
rect 12584 3544 12590 3596
rect 12636 3525 12664 3624
rect 12820 3525 12848 3692
rect 12986 3680 12992 3732
rect 13044 3720 13050 3732
rect 13262 3720 13268 3732
rect 13044 3692 13268 3720
rect 13044 3680 13050 3692
rect 13262 3680 13268 3692
rect 13320 3720 13326 3732
rect 14645 3723 14703 3729
rect 14645 3720 14657 3723
rect 13320 3692 14657 3720
rect 13320 3680 13326 3692
rect 14645 3689 14657 3692
rect 14691 3720 14703 3723
rect 15102 3720 15108 3732
rect 14691 3692 15108 3720
rect 14691 3689 14703 3692
rect 14645 3683 14703 3689
rect 15102 3680 15108 3692
rect 15160 3680 15166 3732
rect 13449 3655 13507 3661
rect 13449 3621 13461 3655
rect 13495 3652 13507 3655
rect 13538 3652 13544 3664
rect 13495 3624 13544 3652
rect 13495 3621 13507 3624
rect 13449 3615 13507 3621
rect 13538 3612 13544 3624
rect 13596 3612 13602 3664
rect 13630 3612 13636 3664
rect 13688 3652 13694 3664
rect 15378 3652 15384 3664
rect 13688 3624 15384 3652
rect 13688 3612 13694 3624
rect 15378 3612 15384 3624
rect 15436 3612 15442 3664
rect 13556 3584 13584 3612
rect 15933 3587 15991 3593
rect 15933 3584 15945 3587
rect 13556 3556 15945 3584
rect 15933 3553 15945 3556
rect 15979 3584 15991 3587
rect 17954 3584 17960 3596
rect 15979 3556 17960 3584
rect 15979 3553 15991 3556
rect 15933 3547 15991 3553
rect 17954 3544 17960 3556
rect 18012 3544 18018 3596
rect 11977 3519 12035 3525
rect 11977 3485 11989 3519
rect 12023 3485 12035 3519
rect 11977 3479 12035 3485
rect 12253 3519 12311 3525
rect 12253 3485 12265 3519
rect 12299 3485 12311 3519
rect 12253 3479 12311 3485
rect 12621 3519 12679 3525
rect 12621 3485 12633 3519
rect 12667 3485 12679 3519
rect 12621 3479 12679 3485
rect 12805 3519 12863 3525
rect 12805 3485 12817 3519
rect 12851 3485 12863 3519
rect 12805 3479 12863 3485
rect 5534 3448 5540 3460
rect 5460 3420 5540 3448
rect 5534 3408 5540 3420
rect 5592 3408 5598 3460
rect 5721 3451 5779 3457
rect 5721 3417 5733 3451
rect 5767 3448 5779 3451
rect 5810 3448 5816 3460
rect 5767 3420 5816 3448
rect 5767 3417 5779 3420
rect 5721 3411 5779 3417
rect 5810 3408 5816 3420
rect 5868 3408 5874 3460
rect 8570 3448 8576 3460
rect 6946 3420 7972 3448
rect 3234 3340 3240 3392
rect 3292 3380 3298 3392
rect 3421 3383 3479 3389
rect 3421 3380 3433 3383
rect 3292 3352 3433 3380
rect 3292 3340 3298 3352
rect 3421 3349 3433 3352
rect 3467 3349 3479 3383
rect 3421 3343 3479 3349
rect 3602 3340 3608 3392
rect 3660 3380 3666 3392
rect 5077 3383 5135 3389
rect 5077 3380 5089 3383
rect 3660 3352 5089 3380
rect 3660 3340 3666 3352
rect 5077 3349 5089 3352
rect 5123 3349 5135 3383
rect 5077 3343 5135 3349
rect 7006 3340 7012 3392
rect 7064 3380 7070 3392
rect 7193 3383 7251 3389
rect 7193 3380 7205 3383
rect 7064 3352 7205 3380
rect 7064 3340 7070 3352
rect 7193 3349 7205 3352
rect 7239 3349 7251 3383
rect 7944 3380 7972 3420
rect 8496 3420 8576 3448
rect 8294 3380 8300 3392
rect 7944 3352 8300 3380
rect 7193 3343 7251 3349
rect 8294 3340 8300 3352
rect 8352 3380 8358 3392
rect 8496 3380 8524 3420
rect 8570 3408 8576 3420
rect 8628 3408 8634 3460
rect 12268 3448 12296 3479
rect 12713 3451 12771 3457
rect 12713 3448 12725 3451
rect 12268 3420 12725 3448
rect 12713 3417 12725 3420
rect 12759 3417 12771 3451
rect 12820 3448 12848 3479
rect 12894 3476 12900 3528
rect 12952 3516 12958 3528
rect 12989 3519 13047 3525
rect 12989 3516 13001 3519
rect 12952 3488 13001 3516
rect 12952 3476 12958 3488
rect 12989 3485 13001 3488
rect 13035 3485 13047 3519
rect 13354 3516 13360 3528
rect 13315 3488 13360 3516
rect 12989 3479 13047 3485
rect 13354 3476 13360 3488
rect 13412 3476 13418 3528
rect 13630 3516 13636 3528
rect 13591 3488 13636 3516
rect 13630 3476 13636 3488
rect 13688 3476 13694 3528
rect 14369 3519 14427 3525
rect 14369 3485 14381 3519
rect 14415 3516 14427 3519
rect 14458 3516 14464 3528
rect 14415 3488 14464 3516
rect 14415 3485 14427 3488
rect 14369 3479 14427 3485
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 14921 3519 14979 3525
rect 14921 3516 14933 3519
rect 14844 3488 14933 3516
rect 13446 3448 13452 3460
rect 12820 3420 13452 3448
rect 12713 3411 12771 3417
rect 13446 3408 13452 3420
rect 13504 3408 13510 3460
rect 8352 3352 8524 3380
rect 8352 3340 8358 3352
rect 8846 3340 8852 3392
rect 8904 3380 8910 3392
rect 9861 3383 9919 3389
rect 9861 3380 9873 3383
rect 8904 3352 9873 3380
rect 8904 3340 8910 3352
rect 9861 3349 9873 3352
rect 9907 3349 9919 3383
rect 9861 3343 9919 3349
rect 12529 3383 12587 3389
rect 12529 3349 12541 3383
rect 12575 3380 12587 3383
rect 14550 3380 14556 3392
rect 12575 3352 14556 3380
rect 12575 3349 12587 3352
rect 12529 3343 12587 3349
rect 14550 3340 14556 3352
rect 14608 3340 14614 3392
rect 14844 3389 14872 3488
rect 14921 3485 14933 3488
rect 14967 3485 14979 3519
rect 14921 3479 14979 3485
rect 15010 3476 15016 3528
rect 15068 3516 15074 3528
rect 15194 3516 15200 3528
rect 15068 3488 15113 3516
rect 15155 3488 15200 3516
rect 15068 3476 15074 3488
rect 15194 3476 15200 3488
rect 15252 3476 15258 3528
rect 16209 3451 16267 3457
rect 16209 3417 16221 3451
rect 16255 3448 16267 3451
rect 16255 3420 16620 3448
rect 16255 3417 16267 3420
rect 16209 3411 16267 3417
rect 16592 3392 16620 3420
rect 16942 3408 16948 3460
rect 17000 3408 17006 3460
rect 17957 3451 18015 3457
rect 17957 3417 17969 3451
rect 18003 3448 18015 3451
rect 18046 3448 18052 3460
rect 18003 3420 18052 3448
rect 18003 3417 18015 3420
rect 17957 3411 18015 3417
rect 18046 3408 18052 3420
rect 18104 3408 18110 3460
rect 14829 3383 14887 3389
rect 14829 3349 14841 3383
rect 14875 3349 14887 3383
rect 14829 3343 14887 3349
rect 14918 3340 14924 3392
rect 14976 3380 14982 3392
rect 14976 3352 15021 3380
rect 14976 3340 14982 3352
rect 16574 3340 16580 3392
rect 16632 3340 16638 3392
rect 0 3290 18860 3312
rect 0 3238 6144 3290
rect 6196 3238 6208 3290
rect 6260 3238 6272 3290
rect 6324 3238 6336 3290
rect 6388 3238 6400 3290
rect 6452 3238 12443 3290
rect 12495 3238 12507 3290
rect 12559 3238 12571 3290
rect 12623 3238 12635 3290
rect 12687 3238 12699 3290
rect 12751 3238 18860 3290
rect 0 3216 18860 3238
rect 5810 3176 5816 3188
rect 5771 3148 5816 3176
rect 5810 3136 5816 3148
rect 5868 3136 5874 3188
rect 5902 3136 5908 3188
rect 5960 3176 5966 3188
rect 5997 3179 6055 3185
rect 5997 3176 6009 3179
rect 5960 3148 6009 3176
rect 5960 3136 5966 3148
rect 5997 3145 6009 3148
rect 6043 3145 6055 3179
rect 7006 3176 7012 3188
rect 5997 3139 6055 3145
rect 6196 3148 7012 3176
rect 4338 3068 4344 3120
rect 4396 3068 4402 3120
rect 5460 3080 5948 3108
rect 3234 3040 3240 3052
rect 3195 3012 3240 3040
rect 3234 3000 3240 3012
rect 3292 3000 3298 3052
rect 3602 3040 3608 3052
rect 3563 3012 3608 3040
rect 3602 3000 3608 3012
rect 3660 3000 3666 3052
rect 4356 3040 4384 3068
rect 4890 3040 4896 3052
rect 4356 3012 4896 3040
rect 4890 3000 4896 3012
rect 4948 3000 4954 3052
rect 5460 3049 5488 3080
rect 5920 3052 5948 3080
rect 5031 3043 5089 3049
rect 5031 3009 5043 3043
rect 5077 3040 5089 3043
rect 5445 3043 5503 3049
rect 5445 3040 5457 3043
rect 5077 3012 5457 3040
rect 5077 3009 5089 3012
rect 5031 3003 5089 3009
rect 5445 3009 5457 3012
rect 5491 3009 5503 3043
rect 5445 3003 5503 3009
rect 5537 3043 5595 3049
rect 5537 3009 5549 3043
rect 5583 3040 5595 3043
rect 5626 3040 5632 3052
rect 5583 3012 5632 3040
rect 5583 3009 5595 3012
rect 5537 3003 5595 3009
rect 5626 3000 5632 3012
rect 5684 3000 5690 3052
rect 5721 3043 5779 3049
rect 5721 3009 5733 3043
rect 5767 3009 5779 3043
rect 5721 3003 5779 3009
rect 5736 2972 5764 3003
rect 5902 3000 5908 3052
rect 5960 3000 5966 3052
rect 6196 3049 6224 3148
rect 7006 3136 7012 3148
rect 7064 3136 7070 3188
rect 8294 3136 8300 3188
rect 8352 3176 8358 3188
rect 8352 3148 9168 3176
rect 8352 3136 8358 3148
rect 6273 3111 6331 3117
rect 6273 3077 6285 3111
rect 6319 3108 6331 3111
rect 6319 3080 6684 3108
rect 6319 3077 6331 3080
rect 6273 3071 6331 3077
rect 6089 3043 6147 3049
rect 6089 3009 6101 3043
rect 6135 3040 6147 3043
rect 6181 3043 6239 3049
rect 6181 3040 6193 3043
rect 6135 3012 6193 3040
rect 6135 3009 6147 3012
rect 6089 3003 6147 3009
rect 6181 3009 6193 3012
rect 6227 3009 6239 3043
rect 6454 3040 6460 3052
rect 6415 3012 6460 3040
rect 6181 3003 6239 3009
rect 6454 3000 6460 3012
rect 6512 3000 6518 3052
rect 6656 3049 6684 3080
rect 6748 3080 7972 3108
rect 9140 3094 9168 3148
rect 9214 3136 9220 3188
rect 9272 3176 9278 3188
rect 10410 3176 10416 3188
rect 9272 3148 10416 3176
rect 9272 3136 9278 3148
rect 10410 3136 10416 3148
rect 10468 3176 10474 3188
rect 11514 3176 11520 3188
rect 10468 3148 11520 3176
rect 10468 3136 10474 3148
rect 11514 3136 11520 3148
rect 11572 3136 11578 3188
rect 12437 3179 12495 3185
rect 12437 3145 12449 3179
rect 12483 3145 12495 3179
rect 12437 3139 12495 3145
rect 12452 3108 12480 3139
rect 12802 3136 12808 3188
rect 12860 3176 12866 3188
rect 12897 3179 12955 3185
rect 12897 3176 12909 3179
rect 12860 3148 12909 3176
rect 12860 3136 12866 3148
rect 12897 3145 12909 3148
rect 12943 3145 12955 3179
rect 12897 3139 12955 3145
rect 13906 3136 13912 3188
rect 13964 3176 13970 3188
rect 14826 3176 14832 3188
rect 13964 3148 14832 3176
rect 13964 3136 13970 3148
rect 14826 3136 14832 3148
rect 14884 3176 14890 3188
rect 15381 3179 15439 3185
rect 14884 3148 15148 3176
rect 14884 3136 14890 3148
rect 13354 3108 13360 3120
rect 12452 3080 13360 3108
rect 6641 3043 6699 3049
rect 6641 3009 6653 3043
rect 6687 3009 6699 3043
rect 6641 3003 6699 3009
rect 6362 2972 6368 2984
rect 5736 2944 6368 2972
rect 6362 2932 6368 2944
rect 6420 2932 6426 2984
rect 6546 2932 6552 2984
rect 6604 2972 6610 2984
rect 6748 2972 6776 3080
rect 6825 3043 6883 3049
rect 6825 3009 6837 3043
rect 6871 3009 6883 3043
rect 7006 3040 7012 3052
rect 6967 3012 7012 3040
rect 6825 3003 6883 3009
rect 6604 2944 6776 2972
rect 6604 2932 6610 2944
rect 5350 2904 5356 2916
rect 5263 2876 5356 2904
rect 5350 2864 5356 2876
rect 5408 2904 5414 2916
rect 6454 2904 6460 2916
rect 5408 2876 6460 2904
rect 5408 2864 5414 2876
rect 6454 2864 6460 2876
rect 6512 2864 6518 2916
rect 5902 2796 5908 2848
rect 5960 2836 5966 2848
rect 6840 2836 6868 3003
rect 7006 3000 7012 3012
rect 7064 3000 7070 3052
rect 7944 3049 7972 3080
rect 13354 3068 13360 3080
rect 13412 3068 13418 3120
rect 13630 3108 13636 3120
rect 13543 3080 13636 3108
rect 13630 3068 13636 3080
rect 13688 3108 13694 3120
rect 14918 3108 14924 3120
rect 13688 3080 13952 3108
rect 13688 3068 13694 3080
rect 7929 3043 7987 3049
rect 7929 3009 7941 3043
rect 7975 3009 7987 3043
rect 8110 3040 8116 3052
rect 8071 3012 8116 3040
rect 7929 3003 7987 3009
rect 8110 3000 8116 3012
rect 8168 3000 8174 3052
rect 8389 3043 8447 3049
rect 8389 3009 8401 3043
rect 8435 3040 8447 3043
rect 8846 3040 8852 3052
rect 8435 3012 8852 3040
rect 8435 3009 8447 3012
rect 8389 3003 8447 3009
rect 8846 3000 8852 3012
rect 8904 3000 8910 3052
rect 10597 3043 10655 3049
rect 10597 3009 10609 3043
rect 10643 3009 10655 3043
rect 12066 3040 12072 3052
rect 12027 3012 12072 3040
rect 10597 3003 10655 3009
rect 6917 2975 6975 2981
rect 6917 2941 6929 2975
rect 6963 2972 6975 2975
rect 8662 2972 8668 2984
rect 6963 2944 8668 2972
rect 6963 2941 6975 2944
rect 6917 2935 6975 2941
rect 8662 2932 8668 2944
rect 8720 2932 8726 2984
rect 8757 2975 8815 2981
rect 8757 2941 8769 2975
rect 8803 2972 8815 2975
rect 8938 2972 8944 2984
rect 8803 2944 8944 2972
rect 8803 2941 8815 2944
rect 8757 2935 8815 2941
rect 8938 2932 8944 2944
rect 8996 2932 9002 2984
rect 10183 2975 10241 2981
rect 10183 2941 10195 2975
rect 10229 2972 10241 2975
rect 10612 2972 10640 3003
rect 12066 3000 12072 3012
rect 12124 3000 12130 3052
rect 13078 3040 13084 3052
rect 13039 3012 13084 3040
rect 13078 3000 13084 3012
rect 13136 3000 13142 3052
rect 13648 3040 13676 3068
rect 13924 3049 13952 3080
rect 14660 3080 14924 3108
rect 13280 3012 13676 3040
rect 13725 3043 13783 3049
rect 11977 2975 12035 2981
rect 11977 2972 11989 2975
rect 10229 2944 11989 2972
rect 10229 2941 10241 2944
rect 10183 2935 10241 2941
rect 11977 2941 11989 2944
rect 12023 2941 12035 2975
rect 11977 2935 12035 2941
rect 12802 2932 12808 2984
rect 12860 2972 12866 2984
rect 13280 2972 13308 3012
rect 13725 3009 13737 3043
rect 13771 3009 13783 3043
rect 13725 3003 13783 3009
rect 13909 3043 13967 3049
rect 13909 3009 13921 3043
rect 13955 3009 13967 3043
rect 14366 3040 14372 3052
rect 14327 3012 14372 3040
rect 13909 3003 13967 3009
rect 12860 2944 13308 2972
rect 13357 2975 13415 2981
rect 12860 2932 12866 2944
rect 13357 2941 13369 2975
rect 13403 2972 13415 2975
rect 13446 2972 13452 2984
rect 13403 2944 13452 2972
rect 13403 2941 13415 2944
rect 13357 2935 13415 2941
rect 13446 2932 13452 2944
rect 13504 2932 13510 2984
rect 10042 2864 10048 2916
rect 10100 2904 10106 2916
rect 10505 2907 10563 2913
rect 10505 2904 10517 2907
rect 10100 2876 10517 2904
rect 10100 2864 10106 2876
rect 10505 2873 10517 2876
rect 10551 2873 10563 2907
rect 10505 2867 10563 2873
rect 13078 2864 13084 2916
rect 13136 2904 13142 2916
rect 13740 2904 13768 3003
rect 14366 3000 14372 3012
rect 14424 3000 14430 3052
rect 14550 3040 14556 3052
rect 14511 3012 14556 3040
rect 14550 3000 14556 3012
rect 14608 3000 14614 3052
rect 14660 3049 14688 3080
rect 14918 3068 14924 3080
rect 14976 3068 14982 3120
rect 15120 3117 15148 3148
rect 15381 3145 15393 3179
rect 15427 3176 15439 3179
rect 15657 3179 15715 3185
rect 15657 3176 15669 3179
rect 15427 3148 15669 3176
rect 15427 3145 15439 3148
rect 15381 3139 15439 3145
rect 15657 3145 15669 3148
rect 15703 3145 15715 3179
rect 15657 3139 15715 3145
rect 16439 3179 16497 3185
rect 16439 3145 16451 3179
rect 16485 3176 16497 3179
rect 17586 3176 17592 3188
rect 16485 3148 17592 3176
rect 16485 3145 16497 3148
rect 16439 3139 16497 3145
rect 17586 3136 17592 3148
rect 17644 3136 17650 3188
rect 15105 3111 15163 3117
rect 15105 3077 15117 3111
rect 15151 3077 15163 3111
rect 15105 3071 15163 3077
rect 16942 3068 16948 3120
rect 17000 3068 17006 3120
rect 14645 3043 14703 3049
rect 14645 3009 14657 3043
rect 14691 3009 14703 3043
rect 14645 3003 14703 3009
rect 14829 3043 14887 3049
rect 14829 3009 14841 3043
rect 14875 3040 14887 3043
rect 15010 3040 15016 3052
rect 14875 3012 15016 3040
rect 14875 3009 14887 3012
rect 14829 3003 14887 3009
rect 15010 3000 15016 3012
rect 15068 3000 15074 3052
rect 15289 3043 15347 3049
rect 15289 3009 15301 3043
rect 15335 3009 15347 3043
rect 15289 3003 15347 3009
rect 14734 2932 14740 2984
rect 14792 2972 14798 2984
rect 15304 2972 15332 3003
rect 15378 3000 15384 3052
rect 15436 3040 15442 3052
rect 15436 3012 15481 3040
rect 15436 3000 15442 3012
rect 17954 3000 17960 3052
rect 18012 3040 18018 3052
rect 18233 3043 18291 3049
rect 18233 3040 18245 3043
rect 18012 3012 18245 3040
rect 18012 3000 18018 3012
rect 18233 3009 18245 3012
rect 18279 3040 18291 3043
rect 18414 3040 18420 3052
rect 18279 3012 18420 3040
rect 18279 3009 18291 3012
rect 18233 3003 18291 3009
rect 18414 3000 18420 3012
rect 18472 3000 18478 3052
rect 18509 3043 18567 3049
rect 18509 3009 18521 3043
rect 18555 3040 18567 3043
rect 18598 3040 18604 3052
rect 18555 3012 18604 3040
rect 18555 3009 18567 3012
rect 18509 3003 18567 3009
rect 18598 3000 18604 3012
rect 18656 3000 18662 3052
rect 16022 2972 16028 2984
rect 14792 2944 15332 2972
rect 15983 2944 16028 2972
rect 14792 2932 14798 2944
rect 16022 2932 16028 2944
rect 16080 2932 16086 2984
rect 16114 2932 16120 2984
rect 16172 2972 16178 2984
rect 16301 2975 16359 2981
rect 16172 2944 16217 2972
rect 16172 2932 16178 2944
rect 16301 2941 16313 2975
rect 16347 2972 16359 2975
rect 16390 2972 16396 2984
rect 16347 2944 16396 2972
rect 16347 2941 16359 2944
rect 16301 2935 16359 2941
rect 16390 2932 16396 2944
rect 16448 2932 16454 2984
rect 17865 2975 17923 2981
rect 17865 2941 17877 2975
rect 17911 2972 17923 2975
rect 18969 2975 19027 2981
rect 18969 2972 18981 2975
rect 17911 2944 18981 2972
rect 17911 2941 17923 2944
rect 17865 2935 17923 2941
rect 18969 2941 18981 2944
rect 19015 2941 19027 2975
rect 18969 2935 19027 2941
rect 15010 2904 15016 2916
rect 13136 2876 15016 2904
rect 13136 2864 13142 2876
rect 15010 2864 15016 2876
rect 15068 2864 15074 2916
rect 7926 2836 7932 2848
rect 5960 2808 6868 2836
rect 7887 2808 7932 2836
rect 5960 2796 5966 2808
rect 7926 2796 7932 2808
rect 7984 2796 7990 2848
rect 9674 2796 9680 2848
rect 9732 2836 9738 2848
rect 10962 2836 10968 2848
rect 9732 2808 10968 2836
rect 9732 2796 9738 2808
rect 10962 2796 10968 2808
rect 11020 2836 11026 2848
rect 13262 2836 13268 2848
rect 11020 2808 13268 2836
rect 11020 2796 11026 2808
rect 13262 2796 13268 2808
rect 13320 2796 13326 2848
rect 13354 2796 13360 2848
rect 13412 2836 13418 2848
rect 13449 2839 13507 2845
rect 13449 2836 13461 2839
rect 13412 2808 13461 2836
rect 13412 2796 13418 2808
rect 13449 2805 13461 2808
rect 13495 2805 13507 2839
rect 13449 2799 13507 2805
rect 13725 2839 13783 2845
rect 13725 2805 13737 2839
rect 13771 2836 13783 2839
rect 13814 2836 13820 2848
rect 13771 2808 13820 2836
rect 13771 2805 13783 2808
rect 13725 2799 13783 2805
rect 13814 2796 13820 2808
rect 13872 2796 13878 2848
rect 14185 2839 14243 2845
rect 14185 2805 14197 2839
rect 14231 2836 14243 2839
rect 14274 2836 14280 2848
rect 14231 2808 14280 2836
rect 14231 2805 14243 2808
rect 14185 2799 14243 2805
rect 14274 2796 14280 2808
rect 14332 2796 14338 2848
rect 14921 2839 14979 2845
rect 14921 2805 14933 2839
rect 14967 2836 14979 2839
rect 15102 2836 15108 2848
rect 14967 2808 15108 2836
rect 14967 2805 14979 2808
rect 14921 2799 14979 2805
rect 15102 2796 15108 2808
rect 15160 2796 15166 2848
rect 18322 2836 18328 2848
rect 18283 2808 18328 2836
rect 18322 2796 18328 2808
rect 18380 2796 18386 2848
rect 0 2746 18860 2768
rect 0 2694 2995 2746
rect 3047 2694 3059 2746
rect 3111 2694 3123 2746
rect 3175 2694 3187 2746
rect 3239 2694 3251 2746
rect 3303 2694 9294 2746
rect 9346 2694 9358 2746
rect 9410 2694 9422 2746
rect 9474 2694 9486 2746
rect 9538 2694 9550 2746
rect 9602 2694 15592 2746
rect 15644 2694 15656 2746
rect 15708 2694 15720 2746
rect 15772 2694 15784 2746
rect 15836 2694 15848 2746
rect 15900 2694 18860 2746
rect 0 2672 18860 2694
rect 5721 2635 5779 2641
rect 5721 2601 5733 2635
rect 5767 2632 5779 2635
rect 5994 2632 6000 2644
rect 5767 2604 6000 2632
rect 5767 2601 5779 2604
rect 5721 2595 5779 2601
rect 5994 2592 6000 2604
rect 6052 2592 6058 2644
rect 6457 2635 6515 2641
rect 6457 2632 6469 2635
rect 6104 2604 6469 2632
rect 4801 2499 4859 2505
rect 4801 2465 4813 2499
rect 4847 2496 4859 2499
rect 5074 2496 5080 2508
rect 4847 2468 5080 2496
rect 4847 2465 4859 2468
rect 4801 2459 4859 2465
rect 5074 2456 5080 2468
rect 5132 2456 5138 2508
rect 5261 2499 5319 2505
rect 5261 2465 5273 2499
rect 5307 2496 5319 2499
rect 5626 2496 5632 2508
rect 5307 2468 5632 2496
rect 5307 2465 5319 2468
rect 5261 2459 5319 2465
rect 5626 2456 5632 2468
rect 5684 2496 5690 2508
rect 6104 2496 6132 2604
rect 6457 2601 6469 2604
rect 6503 2601 6515 2635
rect 6457 2595 6515 2601
rect 9401 2635 9459 2641
rect 9401 2601 9413 2635
rect 9447 2632 9459 2635
rect 9674 2632 9680 2644
rect 9447 2604 9680 2632
rect 9447 2601 9459 2604
rect 9401 2595 9459 2601
rect 9674 2592 9680 2604
rect 9732 2592 9738 2644
rect 11882 2632 11888 2644
rect 9784 2604 11888 2632
rect 6546 2564 6552 2576
rect 5684 2468 6132 2496
rect 6196 2536 6552 2564
rect 5684 2456 5690 2468
rect 4893 2431 4951 2437
rect 4893 2397 4905 2431
rect 4939 2428 4951 2431
rect 5442 2428 5448 2440
rect 4939 2400 5448 2428
rect 4939 2397 4951 2400
rect 4893 2391 4951 2397
rect 5442 2388 5448 2400
rect 5500 2388 5506 2440
rect 5718 2428 5724 2440
rect 5679 2400 5724 2428
rect 5718 2388 5724 2400
rect 5776 2388 5782 2440
rect 5905 2431 5963 2437
rect 5905 2397 5917 2431
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 5920 2360 5948 2391
rect 5994 2388 6000 2440
rect 6052 2428 6058 2440
rect 6196 2437 6224 2536
rect 6546 2524 6552 2536
rect 6604 2564 6610 2576
rect 7837 2567 7895 2573
rect 7837 2564 7849 2567
rect 6604 2536 7849 2564
rect 6604 2524 6610 2536
rect 7837 2533 7849 2536
rect 7883 2533 7895 2567
rect 7837 2527 7895 2533
rect 8018 2524 8024 2576
rect 8076 2564 8082 2576
rect 8076 2536 9260 2564
rect 8076 2524 8082 2536
rect 9232 2508 9260 2536
rect 6748 2468 7512 2496
rect 6748 2437 6776 2468
rect 6089 2431 6147 2437
rect 6089 2428 6101 2431
rect 6052 2400 6101 2428
rect 6052 2388 6058 2400
rect 6089 2397 6101 2400
rect 6135 2397 6147 2431
rect 6089 2391 6147 2397
rect 6181 2431 6239 2437
rect 6181 2397 6193 2431
rect 6227 2397 6239 2431
rect 6181 2391 6239 2397
rect 6273 2431 6331 2437
rect 6273 2397 6285 2431
rect 6319 2428 6331 2431
rect 6733 2431 6791 2437
rect 6733 2428 6745 2431
rect 6319 2400 6745 2428
rect 6319 2397 6331 2400
rect 6273 2391 6331 2397
rect 6733 2397 6745 2400
rect 6779 2397 6791 2431
rect 6733 2391 6791 2397
rect 6822 2388 6828 2440
rect 6880 2428 6886 2440
rect 7484 2437 7512 2468
rect 7926 2456 7932 2508
rect 7984 2496 7990 2508
rect 8389 2499 8447 2505
rect 8389 2496 8401 2499
rect 7984 2468 8401 2496
rect 7984 2456 7990 2468
rect 8389 2465 8401 2468
rect 8435 2465 8447 2499
rect 8389 2459 8447 2465
rect 8662 2456 8668 2508
rect 8720 2496 8726 2508
rect 9125 2499 9183 2505
rect 9125 2496 9137 2499
rect 8720 2468 9137 2496
rect 8720 2456 8726 2468
rect 9125 2465 9137 2468
rect 9171 2465 9183 2499
rect 9125 2459 9183 2465
rect 9214 2456 9220 2508
rect 9272 2496 9278 2508
rect 9784 2496 9812 2604
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 12066 2592 12072 2644
rect 12124 2632 12130 2644
rect 12391 2635 12449 2641
rect 12391 2632 12403 2635
rect 12124 2604 12403 2632
rect 12124 2592 12130 2604
rect 12391 2601 12403 2604
rect 12437 2632 12449 2635
rect 12529 2635 12587 2641
rect 12529 2632 12541 2635
rect 12437 2604 12541 2632
rect 12437 2601 12449 2604
rect 12391 2595 12449 2601
rect 12529 2601 12541 2604
rect 12575 2601 12587 2635
rect 12529 2595 12587 2601
rect 13170 2592 13176 2644
rect 13228 2632 13234 2644
rect 14366 2632 14372 2644
rect 13228 2604 14372 2632
rect 13228 2592 13234 2604
rect 14366 2592 14372 2604
rect 14424 2632 14430 2644
rect 16114 2632 16120 2644
rect 14424 2604 16120 2632
rect 14424 2592 14430 2604
rect 16114 2592 16120 2604
rect 16172 2592 16178 2644
rect 12713 2567 12771 2573
rect 12713 2533 12725 2567
rect 12759 2564 12771 2567
rect 13354 2564 13360 2576
rect 12759 2536 13360 2564
rect 12759 2533 12771 2536
rect 12713 2527 12771 2533
rect 13354 2524 13360 2536
rect 13412 2524 13418 2576
rect 17862 2524 17868 2576
rect 17920 2564 17926 2576
rect 18141 2567 18199 2573
rect 18141 2564 18153 2567
rect 17920 2536 18153 2564
rect 17920 2524 17926 2536
rect 18141 2533 18153 2536
rect 18187 2533 18199 2567
rect 18141 2527 18199 2533
rect 9272 2468 9317 2496
rect 9508 2468 9812 2496
rect 10597 2499 10655 2505
rect 9272 2456 9278 2468
rect 7469 2431 7527 2437
rect 6880 2400 6925 2428
rect 6880 2388 6886 2400
rect 7469 2397 7481 2431
rect 7515 2397 7527 2431
rect 7469 2391 7527 2397
rect 7653 2431 7711 2437
rect 7653 2397 7665 2431
rect 7699 2428 7711 2431
rect 7699 2400 9076 2428
rect 7699 2397 7711 2400
rect 7653 2391 7711 2397
rect 6840 2360 6868 2388
rect 5920 2332 6868 2360
rect 7484 2360 7512 2391
rect 8386 2360 8392 2372
rect 7484 2332 8392 2360
rect 8386 2320 8392 2332
rect 8444 2360 8450 2372
rect 9048 2369 9076 2400
rect 9306 2388 9312 2440
rect 9364 2428 9370 2440
rect 9508 2437 9536 2468
rect 10597 2465 10609 2499
rect 10643 2496 10655 2499
rect 13998 2496 14004 2508
rect 10643 2468 14004 2496
rect 10643 2465 10655 2468
rect 10597 2459 10655 2465
rect 13998 2456 14004 2468
rect 14056 2496 14062 2508
rect 16117 2499 16175 2505
rect 16117 2496 16129 2499
rect 14056 2468 16129 2496
rect 14056 2456 14062 2468
rect 16117 2465 16129 2468
rect 16163 2465 16175 2499
rect 16390 2496 16396 2508
rect 16351 2468 16396 2496
rect 16117 2459 16175 2465
rect 16390 2456 16396 2468
rect 16448 2456 16454 2508
rect 9493 2431 9551 2437
rect 9493 2428 9505 2431
rect 9364 2400 9505 2428
rect 9364 2388 9370 2400
rect 9493 2397 9505 2400
rect 9539 2397 9551 2431
rect 9493 2391 9551 2397
rect 9582 2388 9588 2440
rect 9640 2428 9646 2440
rect 9769 2431 9827 2437
rect 9640 2400 9685 2428
rect 9640 2388 9646 2400
rect 9769 2397 9781 2431
rect 9815 2397 9827 2431
rect 10042 2428 10048 2440
rect 10003 2400 10048 2428
rect 9769 2391 9827 2397
rect 8757 2363 8815 2369
rect 8757 2360 8769 2363
rect 8444 2332 8769 2360
rect 8444 2320 8450 2332
rect 8757 2329 8769 2332
rect 8803 2329 8815 2363
rect 8757 2323 8815 2329
rect 9033 2363 9091 2369
rect 9033 2329 9045 2363
rect 9079 2360 9091 2363
rect 9784 2360 9812 2391
rect 10042 2388 10048 2400
rect 10100 2388 10106 2440
rect 10965 2431 11023 2437
rect 10965 2428 10977 2431
rect 10704 2400 10977 2428
rect 9079 2332 9812 2360
rect 9079 2329 9091 2332
rect 9033 2323 9091 2329
rect 3602 2252 3608 2304
rect 3660 2292 3666 2304
rect 4617 2295 4675 2301
rect 4617 2292 4629 2295
rect 3660 2264 4629 2292
rect 3660 2252 3666 2264
rect 4617 2261 4629 2264
rect 4663 2261 4675 2295
rect 4617 2255 4675 2261
rect 7653 2295 7711 2301
rect 7653 2261 7665 2295
rect 7699 2292 7711 2295
rect 7742 2292 7748 2304
rect 7699 2264 7748 2292
rect 7699 2261 7711 2264
rect 7653 2255 7711 2261
rect 7742 2252 7748 2264
rect 7800 2252 7806 2304
rect 8202 2292 8208 2304
rect 8163 2264 8208 2292
rect 8202 2252 8208 2264
rect 8260 2252 8266 2304
rect 8297 2295 8355 2301
rect 8297 2261 8309 2295
rect 8343 2292 8355 2295
rect 8478 2292 8484 2304
rect 8343 2264 8484 2292
rect 8343 2261 8355 2264
rect 8297 2255 8355 2261
rect 8478 2252 8484 2264
rect 8536 2252 8542 2304
rect 8849 2295 8907 2301
rect 8849 2261 8861 2295
rect 8895 2292 8907 2295
rect 9122 2292 9128 2304
rect 8895 2264 9128 2292
rect 8895 2261 8907 2264
rect 8849 2255 8907 2261
rect 9122 2252 9128 2264
rect 9180 2292 9186 2304
rect 9490 2292 9496 2304
rect 9180 2264 9496 2292
rect 9180 2252 9186 2264
rect 9490 2252 9496 2264
rect 9548 2252 9554 2304
rect 9858 2292 9864 2304
rect 9819 2264 9864 2292
rect 9858 2252 9864 2264
rect 9916 2252 9922 2304
rect 10704 2292 10732 2400
rect 10965 2397 10977 2400
rect 11011 2397 11023 2431
rect 10965 2391 11023 2397
rect 12529 2431 12587 2437
rect 12529 2397 12541 2431
rect 12575 2428 12587 2431
rect 12621 2431 12679 2437
rect 12621 2428 12633 2431
rect 12575 2400 12633 2428
rect 12575 2397 12587 2400
rect 12529 2391 12587 2397
rect 12621 2397 12633 2400
rect 12667 2397 12679 2431
rect 13078 2428 13084 2440
rect 13039 2400 13084 2428
rect 12621 2391 12679 2397
rect 13078 2388 13084 2400
rect 13136 2388 13142 2440
rect 13173 2431 13231 2437
rect 13173 2397 13185 2431
rect 13219 2397 13231 2431
rect 13173 2391 13231 2397
rect 13265 2431 13323 2437
rect 13265 2397 13277 2431
rect 13311 2428 13323 2431
rect 13354 2428 13360 2440
rect 13311 2400 13360 2428
rect 13311 2397 13323 2400
rect 13265 2391 13323 2397
rect 11790 2320 11796 2372
rect 11848 2320 11854 2372
rect 12636 2332 12848 2360
rect 12636 2292 12664 2332
rect 10704 2264 12664 2292
rect 12820 2292 12848 2332
rect 12894 2320 12900 2372
rect 12952 2360 12958 2372
rect 13188 2360 13216 2391
rect 13354 2388 13360 2400
rect 13412 2388 13418 2440
rect 13449 2431 13507 2437
rect 13449 2397 13461 2431
rect 13495 2428 13507 2431
rect 13541 2431 13599 2437
rect 13541 2428 13553 2431
rect 13495 2400 13553 2428
rect 13495 2397 13507 2400
rect 13449 2391 13507 2397
rect 13541 2397 13553 2400
rect 13587 2397 13599 2431
rect 13814 2428 13820 2440
rect 13775 2400 13820 2428
rect 13541 2391 13599 2397
rect 13814 2388 13820 2400
rect 13872 2388 13878 2440
rect 18141 2431 18199 2437
rect 18141 2397 18153 2431
rect 18187 2397 18199 2431
rect 18141 2391 18199 2397
rect 12952 2332 13216 2360
rect 13633 2363 13691 2369
rect 12952 2320 12958 2332
rect 13633 2329 13645 2363
rect 13679 2329 13691 2363
rect 14274 2360 14280 2372
rect 14235 2332 14280 2360
rect 13633 2323 13691 2329
rect 13541 2295 13599 2301
rect 13541 2292 13553 2295
rect 12820 2264 13553 2292
rect 13541 2261 13553 2264
rect 13587 2261 13599 2295
rect 13648 2292 13676 2323
rect 14274 2320 14280 2332
rect 14332 2320 14338 2372
rect 15562 2360 15568 2372
rect 15502 2332 15568 2360
rect 15562 2320 15568 2332
rect 15620 2320 15626 2372
rect 16025 2363 16083 2369
rect 16025 2329 16037 2363
rect 16071 2360 16083 2363
rect 16482 2360 16488 2372
rect 16071 2332 16488 2360
rect 16071 2329 16083 2332
rect 16025 2323 16083 2329
rect 16482 2320 16488 2332
rect 16540 2320 16546 2372
rect 16942 2320 16948 2372
rect 17000 2320 17006 2372
rect 17678 2320 17684 2372
rect 17736 2360 17742 2372
rect 18156 2360 18184 2391
rect 17736 2332 18184 2360
rect 17736 2320 17742 2332
rect 13814 2292 13820 2304
rect 13648 2264 13820 2292
rect 13541 2255 13599 2261
rect 13814 2252 13820 2264
rect 13872 2252 13878 2304
rect 15102 2252 15108 2304
rect 15160 2292 15166 2304
rect 17770 2292 17776 2304
rect 15160 2264 17776 2292
rect 15160 2252 15166 2264
rect 17770 2252 17776 2264
rect 17828 2252 17834 2304
rect 17880 2301 17908 2332
rect 17865 2295 17923 2301
rect 17865 2261 17877 2295
rect 17911 2261 17923 2295
rect 17865 2255 17923 2261
rect 0 2202 18860 2224
rect 0 2150 6144 2202
rect 6196 2150 6208 2202
rect 6260 2150 6272 2202
rect 6324 2150 6336 2202
rect 6388 2150 6400 2202
rect 6452 2150 12443 2202
rect 12495 2150 12507 2202
rect 12559 2150 12571 2202
rect 12623 2150 12635 2202
rect 12687 2150 12699 2202
rect 12751 2150 18860 2202
rect 0 2128 18860 2150
rect 5074 2088 5080 2100
rect 5035 2060 5080 2088
rect 5074 2048 5080 2060
rect 5132 2048 5138 2100
rect 5258 2088 5264 2100
rect 5219 2060 5264 2088
rect 5258 2048 5264 2060
rect 5316 2048 5322 2100
rect 5718 2048 5724 2100
rect 5776 2088 5782 2100
rect 5905 2091 5963 2097
rect 5905 2088 5917 2091
rect 5776 2060 5917 2088
rect 5776 2048 5782 2060
rect 5905 2057 5917 2060
rect 5951 2057 5963 2091
rect 5905 2051 5963 2057
rect 6825 2091 6883 2097
rect 6825 2057 6837 2091
rect 6871 2088 6883 2091
rect 7285 2091 7343 2097
rect 7285 2088 7297 2091
rect 6871 2060 7297 2088
rect 6871 2057 6883 2060
rect 6825 2051 6883 2057
rect 7285 2057 7297 2060
rect 7331 2057 7343 2091
rect 7285 2051 7343 2057
rect 7745 2091 7803 2097
rect 7745 2057 7757 2091
rect 7791 2088 7803 2091
rect 8018 2088 8024 2100
rect 7791 2060 8024 2088
rect 7791 2057 7803 2060
rect 7745 2051 7803 2057
rect 3602 2020 3608 2032
rect 3563 1992 3608 2020
rect 3602 1980 3608 1992
rect 3660 1980 3666 2032
rect 4890 2020 4896 2032
rect 4830 1992 4896 2020
rect 4890 1980 4896 1992
rect 4948 1980 4954 2032
rect 3326 1952 3332 1964
rect 3287 1924 3332 1952
rect 3326 1912 3332 1924
rect 3384 1912 3390 1964
rect 5092 1952 5120 2048
rect 5442 1980 5448 2032
rect 5500 2020 5506 2032
rect 6181 2023 6239 2029
rect 6181 2020 6193 2023
rect 5500 1992 6193 2020
rect 5500 1980 5506 1992
rect 6181 1989 6193 1992
rect 6227 1989 6239 2023
rect 6181 1983 6239 1989
rect 6917 2023 6975 2029
rect 6917 1989 6929 2023
rect 6963 2020 6975 2023
rect 7760 2020 7788 2051
rect 8018 2048 8024 2060
rect 8076 2048 8082 2100
rect 8757 2091 8815 2097
rect 8757 2057 8769 2091
rect 8803 2057 8815 2091
rect 8938 2088 8944 2100
rect 8899 2060 8944 2088
rect 8757 2051 8815 2057
rect 6963 1992 7788 2020
rect 6963 1989 6975 1992
rect 6917 1983 6975 1989
rect 7926 1980 7932 2032
rect 7984 2020 7990 2032
rect 8772 2020 8800 2051
rect 8938 2048 8944 2060
rect 8996 2048 9002 2100
rect 9048 2060 9444 2088
rect 9048 2029 9076 2060
rect 9033 2023 9091 2029
rect 7984 1992 8616 2020
rect 8772 1992 8984 2020
rect 7984 1980 7990 1992
rect 5721 1955 5779 1961
rect 5721 1952 5733 1955
rect 5092 1924 5733 1952
rect 5721 1921 5733 1924
rect 5767 1952 5779 1955
rect 5810 1952 5816 1964
rect 5767 1924 5816 1952
rect 5767 1921 5779 1924
rect 5721 1915 5779 1921
rect 5810 1912 5816 1924
rect 5868 1912 5874 1964
rect 5902 1912 5908 1964
rect 5960 1952 5966 1964
rect 5997 1955 6055 1961
rect 5997 1952 6009 1955
rect 5960 1924 6009 1952
rect 5960 1912 5966 1924
rect 5997 1921 6009 1924
rect 6043 1921 6055 1955
rect 5997 1915 6055 1921
rect 6273 1955 6331 1961
rect 6273 1921 6285 1955
rect 6319 1952 6331 1955
rect 6546 1952 6552 1964
rect 6319 1924 6552 1952
rect 6319 1921 6331 1924
rect 6273 1915 6331 1921
rect 5445 1819 5503 1825
rect 5445 1785 5457 1819
rect 5491 1816 5503 1819
rect 6288 1816 6316 1915
rect 6546 1912 6552 1924
rect 6604 1912 6610 1964
rect 7558 1912 7564 1964
rect 7616 1952 7622 1964
rect 7653 1955 7711 1961
rect 7653 1952 7665 1955
rect 7616 1924 7665 1952
rect 7616 1912 7622 1924
rect 7653 1921 7665 1924
rect 7699 1921 7711 1955
rect 7653 1915 7711 1921
rect 8110 1912 8116 1964
rect 8168 1952 8174 1964
rect 8205 1955 8263 1961
rect 8205 1952 8217 1955
rect 8168 1924 8217 1952
rect 8168 1912 8174 1924
rect 8205 1921 8217 1924
rect 8251 1921 8263 1955
rect 8386 1952 8392 1964
rect 8347 1924 8392 1952
rect 8205 1915 8263 1921
rect 8386 1912 8392 1924
rect 8444 1912 8450 1964
rect 8588 1961 8616 1992
rect 8573 1955 8631 1961
rect 8573 1921 8585 1955
rect 8619 1921 8631 1955
rect 8573 1915 8631 1921
rect 8662 1912 8668 1964
rect 8720 1952 8726 1964
rect 8956 1961 8984 1992
rect 9033 1989 9045 2023
rect 9079 1989 9091 2023
rect 9033 1983 9091 1989
rect 9122 1980 9128 2032
rect 9180 2020 9186 2032
rect 9217 2023 9275 2029
rect 9217 2020 9229 2023
rect 9180 1992 9229 2020
rect 9180 1980 9186 1992
rect 9217 1989 9229 1992
rect 9263 1989 9275 2023
rect 9416 2020 9444 2060
rect 9490 2048 9496 2100
rect 9548 2088 9554 2100
rect 12529 2091 12587 2097
rect 9548 2060 12020 2088
rect 9548 2048 9554 2060
rect 9858 2020 9864 2032
rect 9416 1992 9864 2020
rect 9217 1983 9275 1989
rect 9858 1980 9864 1992
rect 9916 1980 9922 2032
rect 10597 2023 10655 2029
rect 10597 1989 10609 2023
rect 10643 2020 10655 2023
rect 11514 2020 11520 2032
rect 10643 1992 11520 2020
rect 10643 1989 10655 1992
rect 10597 1983 10655 1989
rect 11514 1980 11520 1992
rect 11572 1980 11578 2032
rect 8849 1955 8907 1961
rect 8720 1924 8765 1952
rect 8720 1912 8726 1924
rect 8849 1921 8861 1955
rect 8895 1921 8907 1955
rect 8849 1915 8907 1921
rect 8941 1955 8999 1961
rect 8941 1921 8953 1955
rect 8987 1921 8999 1955
rect 8941 1915 8999 1921
rect 6822 1844 6828 1896
rect 6880 1884 6886 1896
rect 7101 1887 7159 1893
rect 7101 1884 7113 1887
rect 6880 1856 7113 1884
rect 6880 1844 6886 1856
rect 7101 1853 7113 1856
rect 7147 1853 7159 1887
rect 7101 1847 7159 1853
rect 7929 1887 7987 1893
rect 7929 1853 7941 1887
rect 7975 1884 7987 1887
rect 8864 1884 8892 1915
rect 9306 1912 9312 1964
rect 9364 1952 9370 1964
rect 9364 1924 9409 1952
rect 9364 1912 9370 1924
rect 9490 1912 9496 1964
rect 9548 1952 9554 1964
rect 9585 1955 9643 1961
rect 9585 1952 9597 1955
rect 9548 1924 9597 1952
rect 9548 1912 9554 1924
rect 9585 1921 9597 1924
rect 9631 1921 9643 1955
rect 9766 1952 9772 1964
rect 9727 1924 9772 1952
rect 9585 1915 9643 1921
rect 9766 1912 9772 1924
rect 9824 1912 9830 1964
rect 9950 1912 9956 1964
rect 10008 1952 10014 1964
rect 10689 1955 10747 1961
rect 10689 1952 10701 1955
rect 10008 1924 10701 1952
rect 10008 1912 10014 1924
rect 10689 1921 10701 1924
rect 10735 1921 10747 1955
rect 10962 1952 10968 1964
rect 10923 1924 10968 1952
rect 10689 1915 10747 1921
rect 10502 1884 10508 1896
rect 7975 1856 10508 1884
rect 7975 1853 7987 1856
rect 7929 1847 7987 1853
rect 5491 1788 6316 1816
rect 7116 1816 7144 1847
rect 10502 1844 10508 1856
rect 10560 1844 10566 1896
rect 10704 1884 10732 1915
rect 10962 1912 10968 1924
rect 11020 1912 11026 1964
rect 11425 1955 11483 1961
rect 11425 1952 11437 1955
rect 11072 1924 11437 1952
rect 11072 1884 11100 1924
rect 11425 1921 11437 1924
rect 11471 1921 11483 1955
rect 11992 1952 12020 2060
rect 12529 2057 12541 2091
rect 12575 2088 12587 2091
rect 12621 2091 12679 2097
rect 12621 2088 12633 2091
rect 12575 2060 12633 2088
rect 12575 2057 12587 2060
rect 12529 2051 12587 2057
rect 12621 2057 12633 2060
rect 12667 2057 12679 2091
rect 12621 2051 12679 2057
rect 13817 2091 13875 2097
rect 13817 2057 13829 2091
rect 13863 2088 13875 2091
rect 14553 2091 14611 2097
rect 14553 2088 14565 2091
rect 13863 2060 14565 2088
rect 13863 2057 13875 2060
rect 13817 2051 13875 2057
rect 14553 2057 14565 2060
rect 14599 2057 14611 2091
rect 14553 2051 14611 2057
rect 16574 2048 16580 2100
rect 16632 2088 16638 2100
rect 16761 2091 16819 2097
rect 16761 2088 16773 2091
rect 16632 2060 16773 2088
rect 16632 2048 16638 2060
rect 16761 2057 16773 2060
rect 16807 2057 16819 2091
rect 16761 2051 16819 2057
rect 16942 2048 16948 2100
rect 17000 2088 17006 2100
rect 17000 2060 17172 2088
rect 17000 2048 17006 2060
rect 12066 1980 12072 2032
rect 12124 2020 12130 2032
rect 12437 2023 12495 2029
rect 12437 2020 12449 2023
rect 12124 1992 12449 2020
rect 12124 1980 12130 1992
rect 12437 1989 12449 1992
rect 12483 2020 12495 2023
rect 12483 1992 14320 2020
rect 12483 1989 12495 1992
rect 12437 1983 12495 1989
rect 14292 1964 14320 1992
rect 14826 1980 14832 2032
rect 14884 2020 14890 2032
rect 15841 2023 15899 2029
rect 15841 2020 15853 2023
rect 14884 1992 15853 2020
rect 14884 1980 14890 1992
rect 15841 1989 15853 1992
rect 15887 1989 15899 2023
rect 17144 2006 17172 2060
rect 18233 2023 18291 2029
rect 15841 1983 15899 1989
rect 18233 1989 18245 2023
rect 18279 2020 18291 2023
rect 18322 2020 18328 2032
rect 18279 1992 18328 2020
rect 18279 1989 18291 1992
rect 18233 1983 18291 1989
rect 18322 1980 18328 1992
rect 18380 1980 18386 2032
rect 12253 1955 12311 1961
rect 12253 1952 12265 1955
rect 11992 1924 12265 1952
rect 11425 1915 11483 1921
rect 12253 1921 12265 1924
rect 12299 1952 12311 1955
rect 12529 1955 12587 1961
rect 12299 1924 12434 1952
rect 12299 1921 12311 1924
rect 12253 1915 12311 1921
rect 10704 1856 11100 1884
rect 11149 1887 11207 1893
rect 11149 1853 11161 1887
rect 11195 1884 11207 1887
rect 11882 1884 11888 1896
rect 11195 1856 11888 1884
rect 11195 1853 11207 1856
rect 11149 1847 11207 1853
rect 11882 1844 11888 1856
rect 11940 1844 11946 1896
rect 8478 1816 8484 1828
rect 7116 1788 8484 1816
rect 5491 1785 5503 1788
rect 5445 1779 5503 1785
rect 8478 1776 8484 1788
rect 8536 1776 8542 1828
rect 10042 1816 10048 1828
rect 9140 1788 10048 1816
rect 6457 1751 6515 1757
rect 6457 1717 6469 1751
rect 6503 1748 6515 1751
rect 6638 1748 6644 1760
rect 6503 1720 6644 1748
rect 6503 1717 6515 1720
rect 6457 1711 6515 1717
rect 6638 1708 6644 1720
rect 6696 1708 6702 1760
rect 8294 1708 8300 1760
rect 8352 1748 8358 1760
rect 8389 1751 8447 1757
rect 8389 1748 8401 1751
rect 8352 1720 8401 1748
rect 8352 1708 8358 1720
rect 8389 1717 8401 1720
rect 8435 1717 8447 1751
rect 8389 1711 8447 1717
rect 8662 1708 8668 1760
rect 8720 1748 8726 1760
rect 9140 1748 9168 1788
rect 10042 1776 10048 1788
rect 10100 1776 10106 1828
rect 12406 1816 12434 1924
rect 12529 1921 12541 1955
rect 12575 1952 12587 1955
rect 12802 1952 12808 1964
rect 12575 1924 12808 1952
rect 12575 1921 12587 1924
rect 12529 1915 12587 1921
rect 12802 1912 12808 1924
rect 12860 1912 12866 1964
rect 12912 1924 13492 1952
rect 12912 1816 12940 1924
rect 12989 1887 13047 1893
rect 12989 1853 13001 1887
rect 13035 1853 13047 1887
rect 12989 1847 13047 1853
rect 12406 1788 12940 1816
rect 13004 1816 13032 1847
rect 13078 1844 13084 1896
rect 13136 1884 13142 1896
rect 13464 1884 13492 1924
rect 13538 1912 13544 1964
rect 13596 1952 13602 1964
rect 13909 1955 13967 1961
rect 13909 1952 13921 1955
rect 13596 1924 13921 1952
rect 13596 1912 13602 1924
rect 13909 1921 13921 1924
rect 13955 1952 13967 1955
rect 14274 1952 14280 1964
rect 13955 1924 14136 1952
rect 14235 1924 14280 1952
rect 13955 1921 13967 1924
rect 13909 1915 13967 1921
rect 13814 1884 13820 1896
rect 13136 1856 13181 1884
rect 13464 1856 13820 1884
rect 13136 1844 13142 1856
rect 13814 1844 13820 1856
rect 13872 1844 13878 1896
rect 14001 1887 14059 1893
rect 14001 1853 14013 1887
rect 14047 1853 14059 1887
rect 14108 1884 14136 1924
rect 14274 1912 14280 1924
rect 14332 1912 14338 1964
rect 14918 1952 14924 1964
rect 14879 1924 14924 1952
rect 14918 1912 14924 1924
rect 14976 1912 14982 1964
rect 15378 1912 15384 1964
rect 15436 1952 15442 1964
rect 15565 1955 15623 1961
rect 15565 1952 15577 1955
rect 15436 1924 15577 1952
rect 15436 1912 15442 1924
rect 15565 1921 15577 1924
rect 15611 1921 15623 1955
rect 15565 1915 15623 1921
rect 15657 1955 15715 1961
rect 15657 1921 15669 1955
rect 15703 1921 15715 1955
rect 15657 1915 15715 1921
rect 16301 1955 16359 1961
rect 16301 1921 16313 1955
rect 16347 1952 16359 1955
rect 16942 1952 16948 1964
rect 16347 1924 16948 1952
rect 16347 1921 16359 1924
rect 16301 1915 16359 1921
rect 15013 1887 15071 1893
rect 15013 1884 15025 1887
rect 14108 1856 15025 1884
rect 14001 1847 14059 1853
rect 15013 1853 15025 1856
rect 15059 1853 15071 1887
rect 15013 1847 15071 1853
rect 13449 1819 13507 1825
rect 13449 1816 13461 1819
rect 13004 1788 13461 1816
rect 13449 1785 13461 1788
rect 13495 1785 13507 1819
rect 14016 1816 14044 1847
rect 15102 1844 15108 1896
rect 15160 1884 15166 1896
rect 15672 1884 15700 1915
rect 16942 1912 16948 1924
rect 17000 1912 17006 1964
rect 18506 1912 18512 1964
rect 18564 1952 18570 1964
rect 18564 1924 18609 1952
rect 18564 1912 18570 1924
rect 15160 1856 15205 1884
rect 15396 1856 15700 1884
rect 16393 1887 16451 1893
rect 15160 1844 15166 1856
rect 15396 1828 15424 1856
rect 16393 1853 16405 1887
rect 16439 1853 16451 1887
rect 16574 1884 16580 1896
rect 16535 1856 16580 1884
rect 16393 1847 16451 1853
rect 14182 1816 14188 1828
rect 14016 1788 14188 1816
rect 13449 1779 13507 1785
rect 14182 1776 14188 1788
rect 14240 1776 14246 1828
rect 15378 1776 15384 1828
rect 15436 1776 15442 1828
rect 16298 1776 16304 1828
rect 16356 1816 16362 1828
rect 16408 1816 16436 1847
rect 16574 1844 16580 1856
rect 16632 1844 16638 1896
rect 17034 1816 17040 1828
rect 16356 1788 17040 1816
rect 16356 1776 16362 1788
rect 17034 1776 17040 1788
rect 17092 1776 17098 1828
rect 8720 1720 9168 1748
rect 8720 1708 8726 1720
rect 9214 1708 9220 1760
rect 9272 1748 9278 1760
rect 9401 1751 9459 1757
rect 9401 1748 9413 1751
rect 9272 1720 9413 1748
rect 9272 1708 9278 1720
rect 9401 1717 9413 1720
rect 9447 1717 9459 1751
rect 9401 1711 9459 1717
rect 9677 1751 9735 1757
rect 9677 1717 9689 1751
rect 9723 1748 9735 1751
rect 9858 1748 9864 1760
rect 9723 1720 9864 1748
rect 9723 1717 9735 1720
rect 9677 1711 9735 1717
rect 9858 1708 9864 1720
rect 9916 1708 9922 1760
rect 11517 1751 11575 1757
rect 11517 1717 11529 1751
rect 11563 1748 11575 1751
rect 12802 1748 12808 1760
rect 11563 1720 12808 1748
rect 11563 1717 11575 1720
rect 11517 1711 11575 1717
rect 12802 1708 12808 1720
rect 12860 1708 12866 1760
rect 13262 1748 13268 1760
rect 13223 1720 13268 1748
rect 13262 1708 13268 1720
rect 13320 1708 13326 1760
rect 14369 1751 14427 1757
rect 14369 1717 14381 1751
rect 14415 1748 14427 1751
rect 14826 1748 14832 1760
rect 14415 1720 14832 1748
rect 14415 1717 14427 1720
rect 14369 1711 14427 1717
rect 14826 1708 14832 1720
rect 14884 1708 14890 1760
rect 15470 1708 15476 1760
rect 15528 1748 15534 1760
rect 15565 1751 15623 1757
rect 15565 1748 15577 1751
rect 15528 1720 15577 1748
rect 15528 1708 15534 1720
rect 15565 1717 15577 1720
rect 15611 1717 15623 1751
rect 15930 1748 15936 1760
rect 15891 1720 15936 1748
rect 15565 1711 15623 1717
rect 15930 1708 15936 1720
rect 15988 1708 15994 1760
rect 0 1658 18860 1680
rect 0 1606 2995 1658
rect 3047 1606 3059 1658
rect 3111 1606 3123 1658
rect 3175 1606 3187 1658
rect 3239 1606 3251 1658
rect 3303 1606 9294 1658
rect 9346 1606 9358 1658
rect 9410 1606 9422 1658
rect 9474 1606 9486 1658
rect 9538 1606 9550 1658
rect 9602 1606 15592 1658
rect 15644 1606 15656 1658
rect 15708 1606 15720 1658
rect 15772 1606 15784 1658
rect 15836 1606 15848 1658
rect 15900 1606 18860 1658
rect 0 1584 18860 1606
rect 14737 1547 14795 1553
rect 10336 1516 14228 1544
rect 7377 1479 7435 1485
rect 7377 1476 7389 1479
rect 6748 1448 7389 1476
rect 5721 1411 5779 1417
rect 5721 1377 5733 1411
rect 5767 1408 5779 1411
rect 6748 1408 6776 1448
rect 7377 1445 7389 1448
rect 7423 1445 7435 1479
rect 7377 1439 7435 1445
rect 8478 1436 8484 1488
rect 8536 1476 8542 1488
rect 10336 1476 10364 1516
rect 14200 1488 14228 1516
rect 14737 1513 14749 1547
rect 14783 1544 14795 1547
rect 14918 1544 14924 1556
rect 14783 1516 14924 1544
rect 14783 1513 14795 1516
rect 14737 1507 14795 1513
rect 14918 1504 14924 1516
rect 14976 1504 14982 1556
rect 15010 1504 15016 1556
rect 15068 1544 15074 1556
rect 15068 1516 15113 1544
rect 15068 1504 15074 1516
rect 16942 1504 16948 1556
rect 17000 1544 17006 1556
rect 17221 1547 17279 1553
rect 17221 1544 17233 1547
rect 17000 1516 17233 1544
rect 17000 1504 17006 1516
rect 17221 1513 17233 1516
rect 17267 1513 17279 1547
rect 17221 1507 17279 1513
rect 8536 1448 10364 1476
rect 8536 1436 8542 1448
rect 5767 1380 6776 1408
rect 5767 1377 5779 1380
rect 5721 1371 5779 1377
rect 6914 1368 6920 1420
rect 6972 1408 6978 1420
rect 7285 1411 7343 1417
rect 7285 1408 7297 1411
rect 6972 1380 7297 1408
rect 6972 1368 6978 1380
rect 7285 1377 7297 1380
rect 7331 1377 7343 1411
rect 7285 1371 7343 1377
rect 7469 1411 7527 1417
rect 7469 1377 7481 1411
rect 7515 1408 7527 1411
rect 8018 1408 8024 1420
rect 7515 1380 8024 1408
rect 7515 1377 7527 1380
rect 7469 1371 7527 1377
rect 8018 1368 8024 1380
rect 8076 1408 8082 1420
rect 9600 1417 9628 1448
rect 8113 1411 8171 1417
rect 8113 1408 8125 1411
rect 8076 1380 8125 1408
rect 8076 1368 8082 1380
rect 8113 1377 8125 1380
rect 8159 1377 8171 1411
rect 9493 1411 9551 1417
rect 9493 1408 9505 1411
rect 8113 1371 8171 1377
rect 9324 1380 9505 1408
rect 5445 1343 5503 1349
rect 5445 1309 5457 1343
rect 5491 1309 5503 1343
rect 5445 1303 5503 1309
rect 5460 1204 5488 1303
rect 7558 1300 7564 1352
rect 7616 1340 7622 1352
rect 7616 1312 7661 1340
rect 7616 1300 7622 1312
rect 7742 1300 7748 1352
rect 7800 1340 7806 1352
rect 7837 1343 7895 1349
rect 7837 1340 7849 1343
rect 7800 1312 7849 1340
rect 7800 1300 7806 1312
rect 7837 1309 7849 1312
rect 7883 1309 7895 1343
rect 8754 1340 8760 1352
rect 8715 1312 8760 1340
rect 7837 1303 7895 1309
rect 8754 1300 8760 1312
rect 8812 1300 8818 1352
rect 9030 1300 9036 1352
rect 9088 1340 9094 1352
rect 9324 1340 9352 1380
rect 9493 1377 9505 1380
rect 9539 1377 9551 1411
rect 9493 1371 9551 1377
rect 9585 1411 9643 1417
rect 9585 1377 9597 1411
rect 9631 1377 9643 1411
rect 10336 1408 10364 1448
rect 10410 1436 10416 1488
rect 10468 1476 10474 1488
rect 10468 1448 11284 1476
rect 10468 1436 10474 1448
rect 10505 1411 10563 1417
rect 10505 1408 10517 1411
rect 10336 1380 10517 1408
rect 9585 1371 9643 1377
rect 10505 1377 10517 1380
rect 10551 1377 10563 1411
rect 10505 1371 10563 1377
rect 10686 1368 10692 1420
rect 10744 1408 10750 1420
rect 10962 1408 10968 1420
rect 10744 1380 10968 1408
rect 10744 1368 10750 1380
rect 10962 1368 10968 1380
rect 11020 1408 11026 1420
rect 11256 1417 11284 1448
rect 14182 1436 14188 1488
rect 14240 1476 14246 1488
rect 14240 1448 16620 1476
rect 14240 1436 14246 1448
rect 16592 1420 16620 1448
rect 11149 1411 11207 1417
rect 11149 1408 11161 1411
rect 11020 1380 11161 1408
rect 11020 1368 11026 1380
rect 11149 1377 11161 1380
rect 11195 1377 11207 1411
rect 11149 1371 11207 1377
rect 11241 1411 11299 1417
rect 11241 1377 11253 1411
rect 11287 1408 11299 1411
rect 12069 1411 12127 1417
rect 12069 1408 12081 1411
rect 11287 1380 12081 1408
rect 11287 1377 11299 1380
rect 11241 1371 11299 1377
rect 12069 1377 12081 1380
rect 12115 1377 12127 1411
rect 14458 1408 14464 1420
rect 14419 1380 14464 1408
rect 12069 1371 12127 1377
rect 14458 1368 14464 1380
rect 14516 1368 14522 1420
rect 15470 1368 15476 1420
rect 15528 1408 15534 1420
rect 15657 1411 15715 1417
rect 15657 1408 15669 1411
rect 15528 1380 15669 1408
rect 15528 1368 15534 1380
rect 15657 1377 15669 1380
rect 15703 1377 15715 1411
rect 15657 1371 15715 1377
rect 15930 1368 15936 1420
rect 15988 1408 15994 1420
rect 16025 1411 16083 1417
rect 16025 1408 16037 1411
rect 15988 1380 16037 1408
rect 15988 1368 15994 1380
rect 16025 1377 16037 1380
rect 16071 1377 16083 1411
rect 16025 1371 16083 1377
rect 16114 1368 16120 1420
rect 16172 1408 16178 1420
rect 16172 1380 16217 1408
rect 16172 1368 16178 1380
rect 16574 1368 16580 1420
rect 16632 1408 16638 1420
rect 16945 1411 17003 1417
rect 16945 1408 16957 1411
rect 16632 1380 16957 1408
rect 16632 1368 16638 1380
rect 16945 1377 16957 1380
rect 16991 1377 17003 1411
rect 16945 1371 17003 1377
rect 17034 1368 17040 1420
rect 17092 1408 17098 1420
rect 17681 1411 17739 1417
rect 17681 1408 17693 1411
rect 17092 1380 17693 1408
rect 17092 1368 17098 1380
rect 17681 1377 17693 1380
rect 17727 1377 17739 1411
rect 17681 1371 17739 1377
rect 17770 1368 17776 1420
rect 17828 1408 17834 1420
rect 17828 1380 17873 1408
rect 17828 1368 17834 1380
rect 9088 1312 9352 1340
rect 9692 1312 11560 1340
rect 9088 1300 9094 1312
rect 7006 1272 7012 1284
rect 6946 1244 7012 1272
rect 7006 1232 7012 1244
rect 7064 1232 7070 1284
rect 5534 1204 5540 1216
rect 5447 1176 5540 1204
rect 5534 1164 5540 1176
rect 5592 1204 5598 1216
rect 6546 1204 6552 1216
rect 5592 1176 6552 1204
rect 5592 1164 5598 1176
rect 6546 1164 6552 1176
rect 6604 1164 6610 1216
rect 7193 1207 7251 1213
rect 7193 1173 7205 1207
rect 7239 1204 7251 1207
rect 7466 1204 7472 1216
rect 7239 1176 7472 1204
rect 7239 1173 7251 1176
rect 7193 1167 7251 1173
rect 7466 1164 7472 1176
rect 7524 1164 7530 1216
rect 8849 1207 8907 1213
rect 8849 1173 8861 1207
rect 8895 1204 8907 1207
rect 8938 1204 8944 1216
rect 8895 1176 8944 1204
rect 8895 1173 8907 1176
rect 8849 1167 8907 1173
rect 8938 1164 8944 1176
rect 8996 1164 9002 1216
rect 9033 1207 9091 1213
rect 9033 1173 9045 1207
rect 9079 1204 9091 1207
rect 9122 1204 9128 1216
rect 9079 1176 9128 1204
rect 9079 1173 9091 1176
rect 9033 1167 9091 1173
rect 9122 1164 9128 1176
rect 9180 1164 9186 1216
rect 9401 1207 9459 1213
rect 9401 1173 9413 1207
rect 9447 1204 9459 1207
rect 9692 1204 9720 1312
rect 10229 1275 10287 1281
rect 10229 1241 10241 1275
rect 10275 1272 10287 1275
rect 10275 1244 10732 1272
rect 10275 1241 10287 1244
rect 10229 1235 10287 1241
rect 9447 1176 9720 1204
rect 9447 1173 9459 1176
rect 9401 1167 9459 1173
rect 9766 1164 9772 1216
rect 9824 1204 9830 1216
rect 9861 1207 9919 1213
rect 9861 1204 9873 1207
rect 9824 1176 9873 1204
rect 9824 1164 9830 1176
rect 9861 1173 9873 1176
rect 9907 1173 9919 1207
rect 9861 1167 9919 1173
rect 10321 1207 10379 1213
rect 10321 1173 10333 1207
rect 10367 1204 10379 1207
rect 10594 1204 10600 1216
rect 10367 1176 10600 1204
rect 10367 1173 10379 1176
rect 10321 1167 10379 1173
rect 10594 1164 10600 1176
rect 10652 1164 10658 1216
rect 10704 1213 10732 1244
rect 10689 1207 10747 1213
rect 10689 1173 10701 1207
rect 10735 1173 10747 1207
rect 11054 1204 11060 1216
rect 11015 1176 11060 1204
rect 10689 1167 10747 1173
rect 11054 1164 11060 1176
rect 11112 1164 11118 1216
rect 11532 1213 11560 1312
rect 11882 1300 11888 1352
rect 11940 1340 11946 1352
rect 11977 1343 12035 1349
rect 11977 1340 11989 1343
rect 11940 1312 11989 1340
rect 11940 1300 11946 1312
rect 11977 1309 11989 1312
rect 12023 1309 12035 1343
rect 11977 1303 12035 1309
rect 14274 1300 14280 1352
rect 14332 1340 14338 1352
rect 14369 1343 14427 1349
rect 14369 1340 14381 1343
rect 14332 1312 14381 1340
rect 14332 1300 14338 1312
rect 14369 1309 14381 1312
rect 14415 1309 14427 1343
rect 14826 1340 14832 1352
rect 14787 1312 14832 1340
rect 14369 1303 14427 1309
rect 14826 1300 14832 1312
rect 14884 1300 14890 1352
rect 14921 1343 14979 1349
rect 14921 1309 14933 1343
rect 14967 1340 14979 1343
rect 15289 1343 15347 1349
rect 15289 1340 15301 1343
rect 14967 1312 15301 1340
rect 14967 1309 14979 1312
rect 14921 1303 14979 1309
rect 15289 1309 15301 1312
rect 15335 1309 15347 1343
rect 15289 1303 15347 1309
rect 15378 1300 15384 1352
rect 15436 1340 15442 1352
rect 15436 1312 15481 1340
rect 15436 1300 15442 1312
rect 14734 1232 14740 1284
rect 14792 1272 14798 1284
rect 15105 1275 15163 1281
rect 15105 1272 15117 1275
rect 14792 1244 15117 1272
rect 14792 1232 14798 1244
rect 15105 1241 15117 1244
rect 15151 1241 15163 1275
rect 15105 1235 15163 1241
rect 16022 1232 16028 1284
rect 16080 1272 16086 1284
rect 16853 1275 16911 1281
rect 16080 1244 16436 1272
rect 16080 1232 16086 1244
rect 11517 1207 11575 1213
rect 11517 1173 11529 1207
rect 11563 1173 11575 1207
rect 11882 1204 11888 1216
rect 11843 1176 11888 1204
rect 11517 1167 11575 1173
rect 11882 1164 11888 1176
rect 11940 1164 11946 1216
rect 15930 1164 15936 1216
rect 15988 1204 15994 1216
rect 16408 1213 16436 1244
rect 16853 1241 16865 1275
rect 16899 1272 16911 1275
rect 17954 1272 17960 1284
rect 16899 1244 17960 1272
rect 16899 1241 16911 1244
rect 16853 1235 16911 1241
rect 17954 1232 17960 1244
rect 18012 1232 18018 1284
rect 16301 1207 16359 1213
rect 16301 1204 16313 1207
rect 15988 1176 16313 1204
rect 15988 1164 15994 1176
rect 16301 1173 16313 1176
rect 16347 1173 16359 1207
rect 16301 1167 16359 1173
rect 16393 1207 16451 1213
rect 16393 1173 16405 1207
rect 16439 1173 16451 1207
rect 16758 1204 16764 1216
rect 16719 1176 16764 1204
rect 16393 1167 16451 1173
rect 16758 1164 16764 1176
rect 16816 1164 16822 1216
rect 17402 1164 17408 1216
rect 17460 1204 17466 1216
rect 17589 1207 17647 1213
rect 17589 1204 17601 1207
rect 17460 1176 17601 1204
rect 17460 1164 17466 1176
rect 17589 1173 17601 1176
rect 17635 1173 17647 1207
rect 17589 1167 17647 1173
rect 0 1114 18860 1136
rect 0 1062 6144 1114
rect 6196 1062 6208 1114
rect 6260 1062 6272 1114
rect 6324 1062 6336 1114
rect 6388 1062 6400 1114
rect 6452 1062 12443 1114
rect 12495 1062 12507 1114
rect 12559 1062 12571 1114
rect 12623 1062 12635 1114
rect 12687 1062 12699 1114
rect 12751 1062 18860 1114
rect 0 1040 18860 1062
rect 6457 1003 6515 1009
rect 6457 969 6469 1003
rect 6503 1000 6515 1003
rect 6822 1000 6828 1012
rect 6503 972 6828 1000
rect 6503 969 6515 972
rect 6457 963 6515 969
rect 6822 960 6828 972
rect 6880 960 6886 1012
rect 7466 960 7472 1012
rect 7524 1000 7530 1012
rect 8619 1003 8677 1009
rect 7524 972 8524 1000
rect 7524 960 7530 972
rect 6638 932 6644 944
rect 6288 904 6644 932
rect 6288 873 6316 904
rect 6638 892 6644 904
rect 6696 892 6702 944
rect 8202 892 8208 944
rect 8260 892 8266 944
rect 8496 932 8524 972
rect 8619 969 8631 1003
rect 8665 1000 8677 1003
rect 8754 1000 8760 1012
rect 8665 972 8760 1000
rect 8665 969 8677 972
rect 8619 963 8677 969
rect 8754 960 8760 972
rect 8812 960 8818 1012
rect 9125 1003 9183 1009
rect 9125 969 9137 1003
rect 9171 1000 9183 1003
rect 9582 1000 9588 1012
rect 9171 972 9588 1000
rect 9171 969 9183 972
rect 9125 963 9183 969
rect 9582 960 9588 972
rect 9640 960 9646 1012
rect 10502 1000 10508 1012
rect 10463 972 10508 1000
rect 10502 960 10508 972
rect 10560 960 10566 1012
rect 11054 960 11060 1012
rect 11112 1000 11118 1012
rect 11333 1003 11391 1009
rect 11333 1000 11345 1003
rect 11112 972 11345 1000
rect 11112 960 11118 972
rect 11333 969 11345 972
rect 11379 969 11391 1003
rect 12066 1000 12072 1012
rect 12027 972 12072 1000
rect 11333 963 11391 969
rect 12066 960 12072 972
rect 12124 960 12130 1012
rect 14458 960 14464 1012
rect 14516 1000 14522 1012
rect 15105 1003 15163 1009
rect 15105 1000 15117 1003
rect 14516 972 15117 1000
rect 14516 960 14522 972
rect 15105 969 15117 972
rect 15151 969 15163 1003
rect 15105 963 15163 969
rect 16758 960 16764 1012
rect 16816 1000 16822 1012
rect 17497 1003 17555 1009
rect 17497 1000 17509 1003
rect 16816 972 17509 1000
rect 16816 960 16822 972
rect 17497 969 17509 972
rect 17543 969 17555 1003
rect 17862 1000 17868 1012
rect 17823 972 17868 1000
rect 17497 963 17555 969
rect 17862 960 17868 972
rect 17920 960 17926 1012
rect 17954 960 17960 1012
rect 18012 1000 18018 1012
rect 18414 1000 18420 1012
rect 18012 972 18057 1000
rect 18375 972 18420 1000
rect 18012 960 18018 972
rect 18414 960 18420 972
rect 18472 960 18478 1012
rect 8846 932 8852 944
rect 8496 904 8852 932
rect 8846 892 8852 904
rect 8904 892 8910 944
rect 8938 892 8944 944
rect 8996 932 9002 944
rect 9033 935 9091 941
rect 9033 932 9045 935
rect 8996 904 9045 932
rect 8996 892 9002 904
rect 9033 901 9045 904
rect 9079 932 9091 935
rect 9079 904 9628 932
rect 9079 901 9091 904
rect 9033 895 9091 901
rect 6273 867 6331 873
rect 6273 833 6285 867
rect 6319 833 6331 867
rect 6273 827 6331 833
rect 6457 867 6515 873
rect 6457 833 6469 867
rect 6503 833 6515 867
rect 6457 827 6515 833
rect 6472 660 6500 827
rect 6546 824 6552 876
rect 6604 864 6610 876
rect 7190 864 7196 876
rect 6604 836 6649 864
rect 7151 836 7196 864
rect 6604 824 6610 836
rect 7190 824 7196 836
rect 7248 824 7254 876
rect 9600 873 9628 904
rect 9674 892 9680 944
rect 9732 932 9738 944
rect 9861 935 9919 941
rect 9861 932 9873 935
rect 9732 904 9873 932
rect 9732 892 9738 904
rect 9861 901 9873 904
rect 9907 901 9919 935
rect 11146 932 11152 944
rect 9861 895 9919 901
rect 10704 904 11152 932
rect 10704 876 10732 904
rect 11146 892 11152 904
rect 11204 932 11210 944
rect 11204 904 11744 932
rect 11204 892 11210 904
rect 9125 867 9183 873
rect 9125 833 9137 867
rect 9171 864 9183 867
rect 9493 867 9551 873
rect 9493 864 9505 867
rect 9171 836 9505 864
rect 9171 833 9183 836
rect 9125 827 9183 833
rect 9493 833 9505 836
rect 9539 833 9551 867
rect 9493 827 9551 833
rect 9585 867 9643 873
rect 9585 833 9597 867
rect 9631 833 9643 867
rect 10045 867 10103 873
rect 10045 864 10057 867
rect 9585 827 9643 833
rect 9692 836 10057 864
rect 6641 799 6699 805
rect 6641 765 6653 799
rect 6687 796 6699 799
rect 6825 799 6883 805
rect 6825 796 6837 799
rect 6687 768 6837 796
rect 6687 765 6699 768
rect 6641 759 6699 765
rect 6825 765 6837 768
rect 6871 765 6883 799
rect 9214 796 9220 808
rect 9175 768 9220 796
rect 6825 759 6883 765
rect 9214 756 9220 768
rect 9272 756 9278 808
rect 9508 796 9536 827
rect 9692 796 9720 836
rect 10045 833 10057 836
rect 10091 833 10103 867
rect 10045 827 10103 833
rect 10134 824 10140 876
rect 10192 864 10198 876
rect 10413 867 10471 873
rect 10413 864 10425 867
rect 10192 836 10425 864
rect 10192 824 10198 836
rect 10413 833 10425 836
rect 10459 833 10471 867
rect 10686 864 10692 876
rect 10647 836 10692 864
rect 10413 827 10471 833
rect 10686 824 10692 836
rect 10744 824 10750 876
rect 11716 873 11744 904
rect 11790 892 11796 944
rect 11848 932 11854 944
rect 11848 904 12374 932
rect 11848 892 11854 904
rect 13262 892 13268 944
rect 13320 932 13326 944
rect 13541 935 13599 941
rect 13541 932 13553 935
rect 13320 904 13553 932
rect 13320 892 13326 904
rect 13541 901 13553 904
rect 13587 901 13599 935
rect 13541 895 13599 901
rect 16850 892 16856 944
rect 16908 892 16914 944
rect 11241 867 11299 873
rect 11241 833 11253 867
rect 11287 833 11299 867
rect 11241 827 11299 833
rect 11701 867 11759 873
rect 11701 833 11713 867
rect 11747 833 11759 867
rect 11701 827 11759 833
rect 13817 867 13875 873
rect 13817 833 13829 867
rect 13863 864 13875 867
rect 13998 864 14004 876
rect 13863 836 14004 864
rect 13863 833 13875 836
rect 13817 827 13875 833
rect 9858 796 9864 808
rect 9508 768 9720 796
rect 9819 768 9864 796
rect 9858 756 9864 768
rect 9916 756 9922 808
rect 11054 756 11060 808
rect 11112 796 11118 808
rect 11256 796 11284 827
rect 13998 824 14004 836
rect 14056 824 14062 876
rect 14734 824 14740 876
rect 14792 864 14798 876
rect 15013 867 15071 873
rect 15013 864 15025 867
rect 14792 836 15025 864
rect 14792 824 14798 836
rect 15013 833 15025 836
rect 15059 833 15071 867
rect 15013 827 15071 833
rect 15197 867 15255 873
rect 15197 833 15209 867
rect 15243 864 15255 867
rect 15378 864 15384 876
rect 15243 836 15384 864
rect 15243 833 15255 836
rect 15197 827 15255 833
rect 15378 824 15384 836
rect 15436 864 15442 876
rect 15930 864 15936 876
rect 15436 836 15792 864
rect 15891 836 15936 864
rect 15436 824 15442 836
rect 11609 799 11667 805
rect 11609 796 11621 799
rect 11112 768 11621 796
rect 11112 756 11118 768
rect 11609 765 11621 768
rect 11655 765 11667 799
rect 14016 796 14044 824
rect 15565 799 15623 805
rect 15565 796 15577 799
rect 14016 768 15577 796
rect 11609 759 11667 765
rect 15565 765 15577 768
rect 15611 765 15623 799
rect 15764 796 15792 836
rect 15930 824 15936 836
rect 15988 824 15994 876
rect 18322 864 18328 876
rect 18283 836 18328 864
rect 18322 824 18328 836
rect 18380 824 18386 876
rect 15764 768 17172 796
rect 15565 759 15623 765
rect 8018 688 8024 740
rect 8076 728 8082 740
rect 9401 731 9459 737
rect 9401 728 9413 731
rect 8076 700 9413 728
rect 8076 688 8082 700
rect 9401 697 9413 700
rect 9447 728 9459 731
rect 9677 731 9735 737
rect 9677 728 9689 731
rect 9447 700 9689 728
rect 9447 697 9459 700
rect 9401 691 9459 697
rect 9677 697 9689 700
rect 9723 697 9735 731
rect 9677 691 9735 697
rect 17144 672 17172 768
rect 17770 756 17776 808
rect 17828 796 17834 808
rect 18049 799 18107 805
rect 18049 796 18061 799
rect 17828 768 18061 796
rect 17828 756 17834 768
rect 18049 765 18061 768
rect 18095 765 18107 799
rect 18049 759 18107 765
rect 7742 660 7748 672
rect 6472 632 7748 660
rect 7742 620 7748 632
rect 7800 620 7806 672
rect 9030 620 9036 672
rect 9088 660 9094 672
rect 9309 663 9367 669
rect 9309 660 9321 663
rect 9088 632 9321 660
rect 9088 620 9094 632
rect 9309 629 9321 632
rect 9355 629 9367 663
rect 9309 623 9367 629
rect 17126 620 17132 672
rect 17184 660 17190 672
rect 17359 663 17417 669
rect 17359 660 17371 663
rect 17184 632 17371 660
rect 17184 620 17190 632
rect 17359 629 17371 632
rect 17405 629 17417 663
rect 17359 623 17417 629
rect 0 570 18860 592
rect 0 518 2995 570
rect 3047 518 3059 570
rect 3111 518 3123 570
rect 3175 518 3187 570
rect 3239 518 3251 570
rect 3303 518 9294 570
rect 9346 518 9358 570
rect 9410 518 9422 570
rect 9474 518 9486 570
rect 9538 518 9550 570
rect 9602 518 15592 570
rect 15644 518 15656 570
rect 15708 518 15720 570
rect 15772 518 15784 570
rect 15836 518 15848 570
rect 15900 518 18860 570
rect 0 496 18860 518
rect 7377 459 7435 465
rect 7377 425 7389 459
rect 7423 456 7435 459
rect 7558 456 7564 468
rect 7423 428 7564 456
rect 7423 425 7435 428
rect 7377 419 7435 425
rect 7558 416 7564 428
rect 7616 416 7622 468
rect 10965 459 11023 465
rect 10965 425 10977 459
rect 11011 456 11023 459
rect 11882 456 11888 468
rect 11011 428 11888 456
rect 11011 425 11023 428
rect 10965 419 11023 425
rect 11882 416 11888 428
rect 11940 416 11946 468
rect 17402 456 17408 468
rect 17363 428 17408 456
rect 17402 416 17408 428
rect 17460 416 17466 468
rect 18322 456 18328 468
rect 18283 428 18328 456
rect 18322 416 18328 428
rect 18380 416 18386 468
rect 11057 391 11115 397
rect 11057 388 11069 391
rect 10704 360 11069 388
rect 8386 320 8392 332
rect 8347 292 8392 320
rect 8386 280 8392 292
rect 8444 280 8450 332
rect 8665 323 8723 329
rect 8665 289 8677 323
rect 8711 320 8723 323
rect 9030 320 9036 332
rect 8711 292 9036 320
rect 8711 289 8723 292
rect 8665 283 8723 289
rect 9030 280 9036 292
rect 9088 280 9094 332
rect 10134 320 10140 332
rect 10047 292 10140 320
rect 10134 280 10140 292
rect 10192 320 10198 332
rect 10704 329 10732 360
rect 11057 357 11069 360
rect 11103 357 11115 391
rect 11057 351 11115 357
rect 10689 323 10747 329
rect 10192 292 10640 320
rect 10192 280 10198 292
rect 7466 252 7472 264
rect 7427 224 7472 252
rect 7466 212 7472 224
rect 7524 212 7530 264
rect 10612 261 10640 292
rect 10689 289 10701 323
rect 10735 289 10747 323
rect 10689 283 10747 289
rect 14734 280 14740 332
rect 14792 320 14798 332
rect 17037 323 17095 329
rect 17037 320 17049 323
rect 14792 292 17049 320
rect 14792 280 14798 292
rect 17037 289 17049 292
rect 17083 320 17095 323
rect 17678 320 17684 332
rect 17083 292 17684 320
rect 17083 289 17095 292
rect 17037 283 17095 289
rect 17678 280 17684 292
rect 17736 280 17742 332
rect 10597 255 10655 261
rect 10597 221 10609 255
rect 10643 221 10655 255
rect 11054 252 11060 264
rect 11015 224 11060 252
rect 10597 215 10655 221
rect 11054 212 11060 224
rect 11112 212 11118 264
rect 11146 212 11152 264
rect 11204 252 11210 264
rect 11241 255 11299 261
rect 11241 252 11253 255
rect 11204 224 11253 252
rect 11204 212 11210 224
rect 11241 221 11253 224
rect 11287 221 11299 255
rect 17126 252 17132 264
rect 17087 224 17132 252
rect 11241 215 11299 221
rect 17126 212 17132 224
rect 17184 212 17190 264
rect 18506 252 18512 264
rect 18467 224 18512 252
rect 18506 212 18512 224
rect 18564 212 18570 264
rect 8202 144 8208 196
rect 8260 184 8266 196
rect 8260 156 9154 184
rect 8260 144 8266 156
rect 0 26 18860 48
rect 0 -26 6144 26
rect 6196 -26 6208 26
rect 6260 -26 6272 26
rect 6324 -26 6336 26
rect 6388 -26 6400 26
rect 6452 -26 12443 26
rect 12495 -26 12507 26
rect 12559 -26 12571 26
rect 12623 -26 12635 26
rect 12687 -26 12699 26
rect 12751 -26 18860 26
rect 0 -48 18860 -26
<< via1 >>
rect 6144 9766 6196 9818
rect 6208 9766 6260 9818
rect 6272 9766 6324 9818
rect 6336 9766 6388 9818
rect 6400 9766 6452 9818
rect 12443 9766 12495 9818
rect 12507 9766 12559 9818
rect 12571 9766 12623 9818
rect 12635 9766 12687 9818
rect 12699 9766 12751 9818
rect 11336 9664 11388 9716
rect 5632 9596 5684 9648
rect 1308 9571 1360 9580
rect 1308 9537 1317 9571
rect 1317 9537 1351 9571
rect 1351 9537 1360 9571
rect 1308 9528 1360 9537
rect 11428 9596 11480 9648
rect 11612 9596 11664 9648
rect 13084 9596 13136 9648
rect 8300 9528 8352 9580
rect 9220 9571 9272 9580
rect 9220 9537 9229 9571
rect 9229 9537 9263 9571
rect 9263 9537 9272 9571
rect 9220 9528 9272 9537
rect 2320 9503 2372 9512
rect 2320 9469 2329 9503
rect 2329 9469 2363 9503
rect 2363 9469 2372 9503
rect 2320 9460 2372 9469
rect 2688 9460 2740 9512
rect 5724 9460 5776 9512
rect 7288 9460 7340 9512
rect 9680 9528 9732 9580
rect 9772 9571 9824 9580
rect 9772 9537 9781 9571
rect 9781 9537 9815 9571
rect 9815 9537 9824 9571
rect 10048 9571 10100 9580
rect 9772 9528 9824 9537
rect 10048 9537 10057 9571
rect 10057 9537 10091 9571
rect 10091 9537 10100 9571
rect 10048 9528 10100 9537
rect 7104 9392 7156 9444
rect 9956 9460 10008 9512
rect 10968 9528 11020 9580
rect 14280 9596 14332 9648
rect 10876 9460 10928 9512
rect 11336 9503 11388 9512
rect 10692 9392 10744 9444
rect 10784 9392 10836 9444
rect 11336 9469 11345 9503
rect 11345 9469 11379 9503
rect 11379 9469 11388 9503
rect 11336 9460 11388 9469
rect 11428 9460 11480 9512
rect 16856 9596 16908 9648
rect 12900 9392 12952 9444
rect 8116 9324 8168 9376
rect 9680 9324 9732 9376
rect 10600 9367 10652 9376
rect 10600 9333 10609 9367
rect 10609 9333 10643 9367
rect 10643 9333 10652 9367
rect 10600 9324 10652 9333
rect 11796 9324 11848 9376
rect 13176 9324 13228 9376
rect 14464 9324 14516 9376
rect 16488 9503 16540 9512
rect 16488 9469 16497 9503
rect 16497 9469 16531 9503
rect 16531 9469 16540 9503
rect 16488 9460 16540 9469
rect 18328 9571 18380 9580
rect 18328 9537 18337 9571
rect 18337 9537 18371 9571
rect 18371 9537 18380 9571
rect 18328 9528 18380 9537
rect 15476 9324 15528 9376
rect 16028 9324 16080 9376
rect 16856 9324 16908 9376
rect 2995 9222 3047 9274
rect 3059 9222 3111 9274
rect 3123 9222 3175 9274
rect 3187 9222 3239 9274
rect 3251 9222 3303 9274
rect 9294 9222 9346 9274
rect 9358 9222 9410 9274
rect 9422 9222 9474 9274
rect 9486 9222 9538 9274
rect 9550 9222 9602 9274
rect 15592 9222 15644 9274
rect 15656 9222 15708 9274
rect 15720 9222 15772 9274
rect 15784 9222 15836 9274
rect 15848 9222 15900 9274
rect 2320 9120 2372 9172
rect 572 8916 624 8968
rect 2688 8959 2740 8968
rect 2688 8925 2697 8959
rect 2697 8925 2731 8959
rect 2731 8925 2740 8959
rect 2688 8916 2740 8925
rect 5632 9120 5684 9172
rect 9128 9120 9180 9172
rect 9220 9120 9272 9172
rect 12992 9120 13044 9172
rect 5724 8984 5776 9036
rect 7196 8984 7248 9036
rect 8208 8984 8260 9036
rect 8392 9027 8444 9036
rect 8392 8993 8401 9027
rect 8401 8993 8435 9027
rect 8435 8993 8444 9027
rect 8392 8984 8444 8993
rect 9680 9052 9732 9104
rect 10048 9052 10100 9104
rect 11520 9052 11572 9104
rect 12808 9052 12860 9104
rect 15292 9120 15344 9172
rect 16488 9120 16540 9172
rect 18328 9163 18380 9172
rect 18328 9129 18337 9163
rect 18337 9129 18371 9163
rect 18371 9129 18380 9163
rect 18328 9120 18380 9129
rect 9772 8984 9824 9036
rect 10784 8984 10836 9036
rect 11152 8984 11204 9036
rect 13268 8984 13320 9036
rect 14464 8984 14516 9036
rect 15476 9027 15528 9036
rect 15476 8993 15485 9027
rect 15485 8993 15519 9027
rect 15519 8993 15528 9027
rect 15476 8984 15528 8993
rect 17868 8984 17920 9036
rect 5632 8916 5684 8968
rect 2964 8891 3016 8900
rect 2964 8857 2973 8891
rect 2973 8857 3007 8891
rect 3007 8857 3016 8891
rect 2964 8848 3016 8857
rect 6736 8891 6788 8900
rect 6736 8857 6745 8891
rect 6745 8857 6779 8891
rect 6779 8857 6788 8891
rect 6736 8848 6788 8857
rect 388 8780 440 8832
rect 3884 8780 3936 8832
rect 4344 8780 4396 8832
rect 5448 8780 5500 8832
rect 8300 8916 8352 8968
rect 8852 8959 8904 8968
rect 8852 8925 8861 8959
rect 8861 8925 8895 8959
rect 8895 8925 8904 8959
rect 8852 8916 8904 8925
rect 8944 8916 8996 8968
rect 10508 8959 10560 8968
rect 10508 8925 10517 8959
rect 10517 8925 10551 8959
rect 10551 8925 10560 8959
rect 10508 8916 10560 8925
rect 10692 8959 10744 8968
rect 10692 8925 10701 8959
rect 10701 8925 10735 8959
rect 10735 8925 10744 8959
rect 10692 8916 10744 8925
rect 11244 8916 11296 8968
rect 12808 8959 12860 8968
rect 12808 8925 12817 8959
rect 12817 8925 12851 8959
rect 12851 8925 12860 8959
rect 12808 8916 12860 8925
rect 14924 8916 14976 8968
rect 17776 8916 17828 8968
rect 9220 8848 9272 8900
rect 10416 8848 10468 8900
rect 10048 8780 10100 8832
rect 11520 8848 11572 8900
rect 12440 8848 12492 8900
rect 12900 8848 12952 8900
rect 13728 8848 13780 8900
rect 14740 8823 14792 8832
rect 14740 8789 14749 8823
rect 14749 8789 14783 8823
rect 14783 8789 14792 8823
rect 14740 8780 14792 8789
rect 16028 8848 16080 8900
rect 6144 8678 6196 8730
rect 6208 8678 6260 8730
rect 6272 8678 6324 8730
rect 6336 8678 6388 8730
rect 6400 8678 6452 8730
rect 12443 8678 12495 8730
rect 12507 8678 12559 8730
rect 12571 8678 12623 8730
rect 12635 8678 12687 8730
rect 12699 8678 12751 8730
rect 2964 8619 3016 8628
rect 2964 8585 2973 8619
rect 2973 8585 3007 8619
rect 3007 8585 3016 8619
rect 2964 8576 3016 8585
rect 6736 8576 6788 8628
rect 8392 8576 8444 8628
rect 8852 8576 8904 8628
rect 9588 8576 9640 8628
rect 10416 8576 10468 8628
rect 1952 8508 2004 8560
rect 2320 8508 2372 8560
rect 5448 8551 5500 8560
rect 388 8483 440 8492
rect 388 8449 397 8483
rect 397 8449 431 8483
rect 431 8449 440 8483
rect 388 8440 440 8449
rect 2964 8440 3016 8492
rect 756 8415 808 8424
rect 756 8381 765 8415
rect 765 8381 799 8415
rect 799 8381 808 8415
rect 756 8372 808 8381
rect 5448 8517 5457 8551
rect 5457 8517 5491 8551
rect 5491 8517 5500 8551
rect 5448 8508 5500 8517
rect 8208 8508 8260 8560
rect 10600 8508 10652 8560
rect 10968 8576 11020 8628
rect 3332 8440 3384 8492
rect 3884 8483 3936 8492
rect 3884 8449 3893 8483
rect 3893 8449 3927 8483
rect 3927 8449 3936 8483
rect 3884 8440 3936 8449
rect 4160 8483 4212 8492
rect 4160 8449 4169 8483
rect 4169 8449 4203 8483
rect 4203 8449 4212 8483
rect 4160 8440 4212 8449
rect 6644 8440 6696 8492
rect 6736 8440 6788 8492
rect 8944 8483 8996 8492
rect 3792 8372 3844 8424
rect 3332 8304 3384 8356
rect 6460 8372 6512 8424
rect 8944 8449 8953 8483
rect 8953 8449 8987 8483
rect 8987 8449 8996 8483
rect 8944 8440 8996 8449
rect 9128 8483 9180 8492
rect 9128 8449 9137 8483
rect 9137 8449 9171 8483
rect 9171 8449 9180 8483
rect 9128 8440 9180 8449
rect 9220 8440 9272 8492
rect 10416 8440 10468 8492
rect 11152 8440 11204 8492
rect 11244 8440 11296 8492
rect 12440 8508 12492 8560
rect 12716 8508 12768 8560
rect 13728 8508 13780 8560
rect 14188 8508 14240 8560
rect 14464 8576 14516 8628
rect 15200 8508 15252 8560
rect 15292 8508 15344 8560
rect 16856 8508 16908 8560
rect 2412 8279 2464 8288
rect 2412 8245 2421 8279
rect 2421 8245 2455 8279
rect 2455 8245 2464 8279
rect 2412 8236 2464 8245
rect 3608 8236 3660 8288
rect 6828 8236 6880 8288
rect 8668 8372 8720 8424
rect 9036 8372 9088 8424
rect 9680 8372 9732 8424
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 13360 8440 13412 8492
rect 13268 8372 13320 8424
rect 13544 8372 13596 8424
rect 16488 8415 16540 8424
rect 11612 8304 11664 8356
rect 11980 8304 12032 8356
rect 13820 8304 13872 8356
rect 14188 8304 14240 8356
rect 14740 8304 14792 8356
rect 15936 8304 15988 8356
rect 16488 8381 16497 8415
rect 16497 8381 16531 8415
rect 16531 8381 16540 8415
rect 16488 8372 16540 8381
rect 16856 8372 16908 8424
rect 17776 8372 17828 8424
rect 8576 8236 8628 8288
rect 10140 8279 10192 8288
rect 10140 8245 10149 8279
rect 10149 8245 10183 8279
rect 10183 8245 10192 8279
rect 10140 8236 10192 8245
rect 10876 8236 10928 8288
rect 11704 8236 11756 8288
rect 12164 8236 12216 8288
rect 13268 8236 13320 8288
rect 18512 8236 18564 8288
rect 2995 8134 3047 8186
rect 3059 8134 3111 8186
rect 3123 8134 3175 8186
rect 3187 8134 3239 8186
rect 3251 8134 3303 8186
rect 9294 8134 9346 8186
rect 9358 8134 9410 8186
rect 9422 8134 9474 8186
rect 9486 8134 9538 8186
rect 9550 8134 9602 8186
rect 15592 8134 15644 8186
rect 15656 8134 15708 8186
rect 15720 8134 15772 8186
rect 15784 8134 15836 8186
rect 15848 8134 15900 8186
rect 756 8032 808 8084
rect 2320 8032 2372 8084
rect 3332 8075 3384 8084
rect 3056 7964 3108 8016
rect 3332 8041 3341 8075
rect 3341 8041 3375 8075
rect 3375 8041 3384 8075
rect 3332 8032 3384 8041
rect 3792 8032 3844 8084
rect 4160 8032 4212 8084
rect 5540 8032 5592 8084
rect 6460 8032 6512 8084
rect 6828 8032 6880 8084
rect 7288 8032 7340 8084
rect 7840 8032 7892 8084
rect 9772 8032 9824 8084
rect 11060 8032 11112 8084
rect 1860 7828 1912 7880
rect 2412 7828 2464 7880
rect 2688 7871 2740 7880
rect 2688 7837 2697 7871
rect 2697 7837 2731 7871
rect 2731 7837 2740 7871
rect 2688 7828 2740 7837
rect 3700 7896 3752 7948
rect 4252 7964 4304 8016
rect 12532 8032 12584 8084
rect 12992 8075 13044 8084
rect 12992 8041 13001 8075
rect 13001 8041 13035 8075
rect 13035 8041 13044 8075
rect 12992 8032 13044 8041
rect 3608 7871 3660 7880
rect 3608 7837 3617 7871
rect 3617 7837 3651 7871
rect 3651 7837 3660 7871
rect 3608 7828 3660 7837
rect 4068 7871 4120 7880
rect 2320 7692 2372 7744
rect 2504 7692 2556 7744
rect 4068 7837 4077 7871
rect 4077 7837 4111 7871
rect 4111 7837 4120 7871
rect 4068 7828 4120 7837
rect 4344 7828 4396 7880
rect 6368 7939 6420 7948
rect 4160 7760 4212 7812
rect 5540 7828 5592 7880
rect 5908 7871 5960 7880
rect 5908 7837 5917 7871
rect 5917 7837 5951 7871
rect 5951 7837 5960 7871
rect 5908 7828 5960 7837
rect 6368 7905 6377 7939
rect 6377 7905 6411 7939
rect 6411 7905 6420 7939
rect 6368 7896 6420 7905
rect 6460 7896 6512 7948
rect 9036 7896 9088 7948
rect 10140 7896 10192 7948
rect 13268 7964 13320 8016
rect 6828 7828 6880 7880
rect 7288 7871 7340 7880
rect 7288 7837 7297 7871
rect 7297 7837 7331 7871
rect 7331 7837 7340 7871
rect 7840 7871 7892 7880
rect 7288 7828 7340 7837
rect 7840 7837 7849 7871
rect 7849 7837 7883 7871
rect 7883 7837 7892 7871
rect 7840 7828 7892 7837
rect 8116 7871 8168 7880
rect 8116 7837 8125 7871
rect 8125 7837 8159 7871
rect 8159 7837 8168 7871
rect 8116 7828 8168 7837
rect 8944 7828 8996 7880
rect 9588 7828 9640 7880
rect 11980 7939 12032 7948
rect 11980 7905 11989 7939
rect 11989 7905 12023 7939
rect 12023 7905 12032 7939
rect 11980 7896 12032 7905
rect 12716 7896 12768 7948
rect 12808 7896 12860 7948
rect 14188 8032 14240 8084
rect 18328 8032 18380 8084
rect 11704 7871 11756 7880
rect 11704 7837 11713 7871
rect 11713 7837 11747 7871
rect 11747 7837 11756 7871
rect 11704 7828 11756 7837
rect 12164 7871 12216 7880
rect 12164 7837 12173 7871
rect 12173 7837 12207 7871
rect 12207 7837 12216 7871
rect 12164 7828 12216 7837
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 16488 7896 16540 7948
rect 16948 7896 17000 7948
rect 13728 7828 13780 7880
rect 13820 7871 13872 7880
rect 13820 7837 13829 7871
rect 13829 7837 13863 7871
rect 13863 7837 13872 7871
rect 13820 7828 13872 7837
rect 14004 7828 14056 7880
rect 14648 7871 14700 7880
rect 14648 7837 14657 7871
rect 14657 7837 14691 7871
rect 14691 7837 14700 7871
rect 14648 7828 14700 7837
rect 4344 7692 4396 7744
rect 4804 7692 4856 7744
rect 5448 7692 5500 7744
rect 7104 7760 7156 7812
rect 6552 7692 6604 7744
rect 6736 7692 6788 7744
rect 9312 7760 9364 7812
rect 8300 7692 8352 7744
rect 8760 7692 8812 7744
rect 9404 7692 9456 7744
rect 9956 7735 10008 7744
rect 9956 7701 9965 7735
rect 9965 7701 9999 7735
rect 9999 7701 10008 7735
rect 9956 7692 10008 7701
rect 11796 7760 11848 7812
rect 13084 7692 13136 7744
rect 13820 7735 13872 7744
rect 13820 7701 13829 7735
rect 13829 7701 13863 7735
rect 13863 7701 13872 7735
rect 13820 7692 13872 7701
rect 14280 7692 14332 7744
rect 15292 7692 15344 7744
rect 16028 7828 16080 7880
rect 18604 7828 18656 7880
rect 16764 7760 16816 7812
rect 16396 7692 16448 7744
rect 18144 7692 18196 7744
rect 18236 7692 18288 7744
rect 6144 7590 6196 7642
rect 6208 7590 6260 7642
rect 6272 7590 6324 7642
rect 6336 7590 6388 7642
rect 6400 7590 6452 7642
rect 12443 7590 12495 7642
rect 12507 7590 12559 7642
rect 12571 7590 12623 7642
rect 12635 7590 12687 7642
rect 12699 7590 12751 7642
rect 1860 7488 1912 7540
rect 3056 7488 3108 7540
rect 4068 7488 4120 7540
rect 572 7395 624 7404
rect 572 7361 581 7395
rect 581 7361 615 7395
rect 615 7361 624 7395
rect 572 7352 624 7361
rect 1952 7352 2004 7404
rect 2504 7420 2556 7472
rect 2872 7420 2924 7472
rect 4252 7420 4304 7472
rect 2688 7395 2740 7404
rect 2688 7361 2697 7395
rect 2697 7361 2731 7395
rect 2731 7361 2740 7395
rect 2688 7352 2740 7361
rect 4804 7395 4856 7404
rect 4804 7361 4813 7395
rect 4813 7361 4847 7395
rect 4847 7361 4856 7395
rect 4804 7352 4856 7361
rect 5908 7488 5960 7540
rect 1952 7216 2004 7268
rect 2596 7216 2648 7268
rect 4160 7216 4212 7268
rect 5632 7395 5684 7404
rect 5632 7361 5641 7395
rect 5641 7361 5675 7395
rect 5675 7361 5684 7395
rect 5632 7352 5684 7361
rect 6828 7488 6880 7540
rect 7196 7531 7248 7540
rect 7196 7497 7205 7531
rect 7205 7497 7239 7531
rect 7239 7497 7248 7531
rect 7196 7488 7248 7497
rect 6552 7420 6604 7472
rect 6736 7463 6788 7472
rect 6736 7429 6745 7463
rect 6745 7429 6779 7463
rect 6779 7429 6788 7463
rect 6736 7420 6788 7429
rect 8300 7463 8352 7472
rect 8300 7429 8309 7463
rect 8309 7429 8343 7463
rect 8343 7429 8352 7463
rect 8300 7420 8352 7429
rect 6644 7327 6696 7336
rect 6644 7293 6653 7327
rect 6653 7293 6687 7327
rect 6687 7293 6696 7327
rect 6644 7284 6696 7293
rect 6000 7216 6052 7268
rect 4988 7191 5040 7200
rect 4988 7157 4997 7191
rect 4997 7157 5031 7191
rect 5031 7157 5040 7191
rect 4988 7148 5040 7157
rect 5908 7148 5960 7200
rect 6092 7148 6144 7200
rect 7012 7395 7064 7404
rect 7012 7361 7021 7395
rect 7021 7361 7055 7395
rect 7055 7361 7064 7395
rect 7012 7352 7064 7361
rect 9956 7488 10008 7540
rect 14188 7488 14240 7540
rect 8760 7463 8812 7472
rect 8760 7429 8769 7463
rect 8769 7429 8803 7463
rect 8803 7429 8812 7463
rect 8760 7420 8812 7429
rect 9128 7463 9180 7472
rect 9128 7429 9137 7463
rect 9137 7429 9171 7463
rect 9171 7429 9180 7463
rect 9128 7420 9180 7429
rect 8944 7395 8996 7404
rect 8944 7361 8953 7395
rect 8953 7361 8987 7395
rect 8987 7361 8996 7395
rect 8944 7352 8996 7361
rect 9312 7395 9364 7404
rect 9312 7361 9321 7395
rect 9321 7361 9355 7395
rect 9355 7361 9364 7395
rect 9312 7352 9364 7361
rect 9772 7352 9824 7404
rect 8392 7327 8444 7336
rect 8392 7293 8401 7327
rect 8401 7293 8435 7327
rect 8435 7293 8444 7327
rect 8392 7284 8444 7293
rect 8576 7327 8628 7336
rect 8576 7293 8585 7327
rect 8585 7293 8619 7327
rect 8619 7293 8628 7327
rect 8576 7284 8628 7293
rect 9220 7284 9272 7336
rect 9588 7284 9640 7336
rect 7288 7216 7340 7268
rect 9680 7216 9732 7268
rect 8208 7148 8260 7200
rect 9956 7395 10008 7404
rect 9956 7361 9965 7395
rect 9965 7361 9999 7395
rect 9999 7361 10008 7395
rect 12716 7420 12768 7472
rect 13728 7420 13780 7472
rect 15200 7463 15252 7472
rect 15200 7429 15209 7463
rect 15209 7429 15243 7463
rect 15243 7429 15252 7463
rect 15200 7420 15252 7429
rect 16764 7420 16816 7472
rect 18144 7463 18196 7472
rect 18144 7429 18153 7463
rect 18153 7429 18187 7463
rect 18187 7429 18196 7463
rect 18144 7420 18196 7429
rect 9956 7352 10008 7361
rect 10140 7327 10192 7336
rect 10140 7293 10149 7327
rect 10149 7293 10183 7327
rect 10183 7293 10192 7327
rect 10140 7284 10192 7293
rect 10968 7327 11020 7336
rect 10968 7293 10977 7327
rect 10977 7293 11011 7327
rect 11011 7293 11020 7327
rect 10968 7284 11020 7293
rect 14096 7395 14148 7404
rect 14096 7361 14105 7395
rect 14105 7361 14139 7395
rect 14139 7361 14148 7395
rect 14096 7352 14148 7361
rect 11888 7284 11940 7336
rect 13820 7284 13872 7336
rect 14004 7327 14056 7336
rect 14004 7293 14013 7327
rect 14013 7293 14047 7327
rect 14047 7293 14056 7327
rect 14004 7284 14056 7293
rect 12532 7148 12584 7200
rect 14280 7216 14332 7268
rect 14924 7148 14976 7200
rect 16028 7327 16080 7336
rect 16028 7293 16037 7327
rect 16037 7293 16071 7327
rect 16071 7293 16080 7327
rect 16028 7284 16080 7293
rect 16672 7284 16724 7336
rect 16948 7148 17000 7200
rect 2995 7046 3047 7098
rect 3059 7046 3111 7098
rect 3123 7046 3175 7098
rect 3187 7046 3239 7098
rect 3251 7046 3303 7098
rect 9294 7046 9346 7098
rect 9358 7046 9410 7098
rect 9422 7046 9474 7098
rect 9486 7046 9538 7098
rect 9550 7046 9602 7098
rect 15592 7046 15644 7098
rect 15656 7046 15708 7098
rect 15720 7046 15772 7098
rect 15784 7046 15836 7098
rect 15848 7046 15900 7098
rect 5448 6944 5500 6996
rect 7012 6944 7064 6996
rect 3608 6876 3660 6928
rect 3056 6783 3108 6792
rect 3056 6749 3065 6783
rect 3065 6749 3099 6783
rect 3099 6749 3108 6783
rect 3056 6740 3108 6749
rect 4988 6808 5040 6860
rect 1676 6604 1728 6656
rect 3240 6604 3292 6656
rect 3608 6783 3660 6792
rect 3608 6749 3617 6783
rect 3617 6749 3651 6783
rect 3651 6749 3660 6783
rect 3884 6783 3936 6792
rect 3608 6740 3660 6749
rect 3884 6749 3893 6783
rect 3893 6749 3927 6783
rect 3927 6749 3936 6783
rect 3884 6740 3936 6749
rect 5080 6740 5132 6792
rect 6092 6876 6144 6928
rect 6552 6876 6604 6928
rect 8576 6944 8628 6996
rect 9772 6944 9824 6996
rect 10508 6944 10560 6996
rect 12348 6944 12400 6996
rect 13360 6944 13412 6996
rect 14096 6944 14148 6996
rect 5356 6808 5408 6860
rect 10140 6876 10192 6928
rect 7104 6808 7156 6860
rect 8208 6851 8260 6860
rect 5816 6783 5868 6792
rect 5816 6749 5825 6783
rect 5825 6749 5859 6783
rect 5859 6749 5868 6783
rect 5816 6740 5868 6749
rect 6000 6783 6052 6792
rect 6000 6749 6009 6783
rect 6009 6749 6043 6783
rect 6043 6749 6052 6783
rect 6000 6740 6052 6749
rect 8208 6817 8217 6851
rect 8217 6817 8251 6851
rect 8251 6817 8260 6851
rect 8208 6808 8260 6817
rect 8484 6808 8536 6860
rect 11612 6808 11664 6860
rect 11980 6851 12032 6860
rect 11980 6817 11989 6851
rect 11989 6817 12023 6851
rect 12023 6817 12032 6851
rect 11980 6808 12032 6817
rect 12440 6851 12492 6860
rect 12440 6817 12449 6851
rect 12449 6817 12483 6851
rect 12483 6817 12492 6851
rect 12440 6808 12492 6817
rect 12992 6808 13044 6860
rect 13176 6808 13228 6860
rect 15108 6944 15160 6996
rect 14464 6808 14516 6860
rect 5448 6672 5500 6724
rect 7840 6783 7892 6792
rect 7840 6749 7849 6783
rect 7849 6749 7883 6783
rect 7883 6749 7892 6783
rect 7840 6740 7892 6749
rect 10140 6740 10192 6792
rect 11888 6783 11940 6792
rect 11888 6749 11897 6783
rect 11897 6749 11931 6783
rect 11931 6749 11940 6783
rect 11888 6740 11940 6749
rect 4252 6604 4304 6656
rect 5632 6604 5684 6656
rect 6644 6604 6696 6656
rect 6828 6647 6880 6656
rect 6828 6613 6837 6647
rect 6837 6613 6871 6647
rect 6871 6613 6880 6647
rect 6828 6604 6880 6613
rect 7104 6604 7156 6656
rect 7380 6672 7432 6724
rect 9220 6672 9272 6724
rect 10048 6672 10100 6724
rect 11612 6715 11664 6724
rect 8116 6604 8168 6656
rect 9036 6604 9088 6656
rect 11244 6604 11296 6656
rect 11612 6681 11621 6715
rect 11621 6681 11655 6715
rect 11655 6681 11664 6715
rect 11612 6672 11664 6681
rect 12164 6740 12216 6792
rect 12900 6740 12952 6792
rect 14280 6740 14332 6792
rect 16028 6808 16080 6860
rect 16580 6851 16632 6860
rect 16580 6817 16589 6851
rect 16589 6817 16623 6851
rect 16623 6817 16632 6851
rect 16580 6808 16632 6817
rect 16948 6851 17000 6860
rect 16948 6817 16957 6851
rect 16957 6817 16991 6851
rect 16991 6817 17000 6851
rect 16948 6808 17000 6817
rect 11520 6604 11572 6656
rect 11796 6604 11848 6656
rect 12072 6604 12124 6656
rect 12624 6672 12676 6724
rect 14740 6740 14792 6792
rect 14924 6783 14976 6792
rect 14924 6749 14933 6783
rect 14933 6749 14967 6783
rect 14967 6749 14976 6783
rect 14924 6740 14976 6749
rect 16672 6740 16724 6792
rect 17500 6783 17552 6792
rect 17500 6749 17509 6783
rect 17509 6749 17543 6783
rect 17543 6749 17552 6783
rect 17500 6740 17552 6749
rect 14648 6715 14700 6724
rect 14648 6681 14657 6715
rect 14657 6681 14691 6715
rect 14691 6681 14700 6715
rect 14648 6672 14700 6681
rect 15292 6672 15344 6724
rect 12256 6604 12308 6656
rect 12808 6604 12860 6656
rect 13084 6604 13136 6656
rect 14096 6604 14148 6656
rect 14372 6604 14424 6656
rect 14740 6647 14792 6656
rect 14740 6613 14749 6647
rect 14749 6613 14783 6647
rect 14783 6613 14792 6647
rect 14740 6604 14792 6613
rect 16304 6604 16356 6656
rect 16856 6604 16908 6656
rect 17408 6647 17460 6656
rect 17408 6613 17417 6647
rect 17417 6613 17451 6647
rect 17451 6613 17460 6647
rect 17408 6604 17460 6613
rect 17960 6604 18012 6656
rect 6144 6502 6196 6554
rect 6208 6502 6260 6554
rect 6272 6502 6324 6554
rect 6336 6502 6388 6554
rect 6400 6502 6452 6554
rect 12443 6502 12495 6554
rect 12507 6502 12559 6554
rect 12571 6502 12623 6554
rect 12635 6502 12687 6554
rect 12699 6502 12751 6554
rect 2596 6400 2648 6452
rect 3056 6400 3108 6452
rect 4252 6443 4304 6452
rect 4252 6409 4261 6443
rect 4261 6409 4295 6443
rect 4295 6409 4304 6443
rect 4252 6400 4304 6409
rect 5632 6400 5684 6452
rect 7840 6400 7892 6452
rect 8116 6400 8168 6452
rect 1676 6375 1728 6384
rect 1676 6341 1685 6375
rect 1685 6341 1719 6375
rect 1719 6341 1728 6375
rect 1676 6332 1728 6341
rect 572 6264 624 6316
rect 3240 6307 3292 6316
rect 3240 6273 3249 6307
rect 3249 6273 3283 6307
rect 3283 6273 3292 6307
rect 3240 6264 3292 6273
rect 3608 6332 3660 6384
rect 5356 6332 5408 6384
rect 3792 6307 3844 6316
rect 3792 6273 3801 6307
rect 3801 6273 3835 6307
rect 3835 6273 3844 6307
rect 3792 6264 3844 6273
rect 4896 6307 4948 6316
rect 3884 6128 3936 6180
rect 4252 6196 4304 6248
rect 4344 6196 4396 6248
rect 4896 6273 4905 6307
rect 4905 6273 4939 6307
rect 4939 6273 4948 6307
rect 4896 6264 4948 6273
rect 5080 6264 5132 6316
rect 5448 6307 5500 6316
rect 5448 6273 5457 6307
rect 5457 6273 5491 6307
rect 5491 6273 5500 6307
rect 5448 6264 5500 6273
rect 4068 6128 4120 6180
rect 5908 6332 5960 6384
rect 8668 6332 8720 6384
rect 10232 6400 10284 6452
rect 11612 6400 11664 6452
rect 11704 6400 11756 6452
rect 11888 6400 11940 6452
rect 15016 6443 15068 6452
rect 12072 6375 12124 6384
rect 6828 6307 6880 6316
rect 6828 6273 6837 6307
rect 6837 6273 6871 6307
rect 6871 6273 6880 6307
rect 6828 6264 6880 6273
rect 7196 6264 7248 6316
rect 8116 6307 8168 6316
rect 8116 6273 8125 6307
rect 8125 6273 8159 6307
rect 8159 6273 8168 6307
rect 8116 6264 8168 6273
rect 8484 6307 8536 6316
rect 8484 6273 8493 6307
rect 8493 6273 8527 6307
rect 8527 6273 8536 6307
rect 8484 6264 8536 6273
rect 6552 6196 6604 6248
rect 10232 6307 10284 6316
rect 10232 6273 10241 6307
rect 10241 6273 10275 6307
rect 10275 6273 10284 6307
rect 10232 6264 10284 6273
rect 10784 6264 10836 6316
rect 11244 6307 11296 6316
rect 11244 6273 11253 6307
rect 11253 6273 11287 6307
rect 11287 6273 11296 6307
rect 11244 6264 11296 6273
rect 12072 6341 12081 6375
rect 12081 6341 12115 6375
rect 12115 6341 12124 6375
rect 12072 6332 12124 6341
rect 11888 6307 11940 6316
rect 11888 6273 11897 6307
rect 11897 6273 11931 6307
rect 11931 6273 11940 6307
rect 11888 6264 11940 6273
rect 10968 6239 11020 6248
rect 7196 6128 7248 6180
rect 10968 6205 10977 6239
rect 10977 6205 11011 6239
rect 11011 6205 11020 6239
rect 10968 6196 11020 6205
rect 11612 6196 11664 6248
rect 15016 6409 15025 6443
rect 15025 6409 15059 6443
rect 15059 6409 15068 6443
rect 15016 6400 15068 6409
rect 15108 6400 15160 6452
rect 13084 6332 13136 6384
rect 14188 6375 14240 6384
rect 14188 6341 14197 6375
rect 14197 6341 14231 6375
rect 14231 6341 14240 6375
rect 14188 6332 14240 6341
rect 14372 6375 14424 6384
rect 14372 6341 14381 6375
rect 14381 6341 14415 6375
rect 14415 6341 14424 6375
rect 14372 6332 14424 6341
rect 13360 6264 13412 6316
rect 12808 6196 12860 6248
rect 13636 6196 13688 6248
rect 14924 6196 14976 6248
rect 15476 6264 15528 6316
rect 16304 6332 16356 6384
rect 17408 6400 17460 6452
rect 17960 6443 18012 6452
rect 17960 6409 17969 6443
rect 17969 6409 18003 6443
rect 18003 6409 18012 6443
rect 17960 6400 18012 6409
rect 16028 6264 16080 6316
rect 17500 6264 17552 6316
rect 17592 6264 17644 6316
rect 15292 6196 15344 6248
rect 15936 6239 15988 6248
rect 15936 6205 15945 6239
rect 15945 6205 15979 6239
rect 15979 6205 15988 6239
rect 15936 6196 15988 6205
rect 18144 6239 18196 6248
rect 18144 6205 18153 6239
rect 18153 6205 18187 6239
rect 18187 6205 18196 6239
rect 18144 6196 18196 6205
rect 3332 6103 3384 6112
rect 3332 6069 3341 6103
rect 3341 6069 3375 6103
rect 3375 6069 3384 6103
rect 3332 6060 3384 6069
rect 5816 6060 5868 6112
rect 8392 6060 8444 6112
rect 10140 6060 10192 6112
rect 10416 6103 10468 6112
rect 10416 6069 10425 6103
rect 10425 6069 10459 6103
rect 10459 6069 10468 6103
rect 10416 6060 10468 6069
rect 10508 6060 10560 6112
rect 11980 6060 12032 6112
rect 13728 6128 13780 6180
rect 12900 6060 12952 6112
rect 14188 6060 14240 6112
rect 15016 6060 15068 6112
rect 17224 6060 17276 6112
rect 2995 5958 3047 6010
rect 3059 5958 3111 6010
rect 3123 5958 3175 6010
rect 3187 5958 3239 6010
rect 3251 5958 3303 6010
rect 9294 5958 9346 6010
rect 9358 5958 9410 6010
rect 9422 5958 9474 6010
rect 9486 5958 9538 6010
rect 9550 5958 9602 6010
rect 15592 5958 15644 6010
rect 15656 5958 15708 6010
rect 15720 5958 15772 6010
rect 15784 5958 15836 6010
rect 15848 5958 15900 6010
rect 572 5720 624 5772
rect 4160 5856 4212 5908
rect 4252 5856 4304 5908
rect 6644 5899 6696 5908
rect 3332 5788 3384 5840
rect 3792 5788 3844 5840
rect 6644 5865 6653 5899
rect 6653 5865 6687 5899
rect 6687 5865 6696 5899
rect 6644 5856 6696 5865
rect 10784 5856 10836 5908
rect 12992 5856 13044 5908
rect 13268 5856 13320 5908
rect 14280 5856 14332 5908
rect 14648 5856 14700 5908
rect 15476 5856 15528 5908
rect 16304 5856 16356 5908
rect 16948 5856 17000 5908
rect 17224 5899 17276 5908
rect 17224 5865 17233 5899
rect 17233 5865 17267 5899
rect 17267 5865 17276 5899
rect 17224 5856 17276 5865
rect 18328 5899 18380 5908
rect 18328 5865 18337 5899
rect 18337 5865 18371 5899
rect 18371 5865 18380 5899
rect 18328 5856 18380 5865
rect 3332 5695 3384 5704
rect 3332 5661 3341 5695
rect 3341 5661 3375 5695
rect 3375 5661 3384 5695
rect 3332 5652 3384 5661
rect 3976 5720 4028 5772
rect 3608 5695 3660 5704
rect 3608 5661 3617 5695
rect 3617 5661 3651 5695
rect 3651 5661 3660 5695
rect 3608 5652 3660 5661
rect 2596 5584 2648 5636
rect 3792 5652 3844 5704
rect 4160 5695 4212 5704
rect 4160 5661 4169 5695
rect 4169 5661 4203 5695
rect 4203 5661 4212 5695
rect 4160 5652 4212 5661
rect 4068 5627 4120 5636
rect 4068 5593 4077 5627
rect 4077 5593 4111 5627
rect 4111 5593 4120 5627
rect 4068 5584 4120 5593
rect 4896 5652 4948 5704
rect 5632 5720 5684 5772
rect 15292 5788 15344 5840
rect 16580 5788 16632 5840
rect 7196 5763 7248 5772
rect 7196 5729 7205 5763
rect 7205 5729 7239 5763
rect 7239 5729 7248 5763
rect 7196 5720 7248 5729
rect 8116 5763 8168 5772
rect 8116 5729 8125 5763
rect 8125 5729 8159 5763
rect 8159 5729 8168 5763
rect 8116 5720 8168 5729
rect 11704 5720 11756 5772
rect 7840 5695 7892 5704
rect 7840 5661 7849 5695
rect 7849 5661 7883 5695
rect 7883 5661 7892 5695
rect 7840 5652 7892 5661
rect 8024 5695 8076 5704
rect 8024 5661 8033 5695
rect 8033 5661 8067 5695
rect 8067 5661 8076 5695
rect 8024 5652 8076 5661
rect 7104 5627 7156 5636
rect 7104 5593 7113 5627
rect 7113 5593 7147 5627
rect 7147 5593 7156 5627
rect 9956 5652 10008 5704
rect 10140 5652 10192 5704
rect 11060 5695 11112 5704
rect 7104 5584 7156 5593
rect 5356 5559 5408 5568
rect 5356 5525 5365 5559
rect 5365 5525 5399 5559
rect 5399 5525 5408 5559
rect 5356 5516 5408 5525
rect 5816 5516 5868 5568
rect 10508 5584 10560 5636
rect 11060 5661 11069 5695
rect 11069 5661 11103 5695
rect 11103 5661 11112 5695
rect 11060 5652 11112 5661
rect 12348 5652 12400 5704
rect 13084 5652 13136 5704
rect 13268 5695 13320 5704
rect 13268 5661 13277 5695
rect 13277 5661 13311 5695
rect 13311 5661 13320 5695
rect 13268 5652 13320 5661
rect 13452 5652 13504 5704
rect 13912 5720 13964 5772
rect 14372 5720 14424 5772
rect 13728 5695 13780 5704
rect 13728 5661 13737 5695
rect 13737 5661 13771 5695
rect 13771 5661 13780 5695
rect 13728 5652 13780 5661
rect 16396 5720 16448 5772
rect 11336 5627 11388 5636
rect 9956 5516 10008 5568
rect 11336 5593 11345 5627
rect 11345 5593 11379 5627
rect 11379 5593 11388 5627
rect 11336 5584 11388 5593
rect 12164 5516 12216 5568
rect 13084 5559 13136 5568
rect 13084 5525 13093 5559
rect 13093 5525 13127 5559
rect 13127 5525 13136 5559
rect 13084 5516 13136 5525
rect 13636 5516 13688 5568
rect 14372 5584 14424 5636
rect 16304 5695 16356 5704
rect 16304 5661 16313 5695
rect 16313 5661 16347 5695
rect 16347 5661 16356 5695
rect 16672 5695 16724 5704
rect 16304 5652 16356 5661
rect 16672 5661 16681 5695
rect 16681 5661 16715 5695
rect 16715 5661 16724 5695
rect 16672 5652 16724 5661
rect 18144 5720 18196 5772
rect 17500 5652 17552 5704
rect 17776 5652 17828 5704
rect 18512 5695 18564 5704
rect 18512 5661 18521 5695
rect 18521 5661 18555 5695
rect 18555 5661 18564 5695
rect 18512 5652 18564 5661
rect 17868 5584 17920 5636
rect 16212 5559 16264 5568
rect 16212 5525 16221 5559
rect 16221 5525 16255 5559
rect 16255 5525 16264 5559
rect 16212 5516 16264 5525
rect 17592 5516 17644 5568
rect 17684 5559 17736 5568
rect 17684 5525 17693 5559
rect 17693 5525 17727 5559
rect 17727 5525 17736 5559
rect 17684 5516 17736 5525
rect 6144 5414 6196 5466
rect 6208 5414 6260 5466
rect 6272 5414 6324 5466
rect 6336 5414 6388 5466
rect 6400 5414 6452 5466
rect 12443 5414 12495 5466
rect 12507 5414 12559 5466
rect 12571 5414 12623 5466
rect 12635 5414 12687 5466
rect 12699 5414 12751 5466
rect 4068 5312 4120 5364
rect 4896 5312 4948 5364
rect 4344 5244 4396 5296
rect 5632 5176 5684 5228
rect 7840 5176 7892 5228
rect 10968 5312 11020 5364
rect 11796 5312 11848 5364
rect 12348 5312 12400 5364
rect 9220 5244 9272 5296
rect 9956 5287 10008 5296
rect 9956 5253 9965 5287
rect 9965 5253 9999 5287
rect 9999 5253 10008 5287
rect 9956 5244 10008 5253
rect 10416 5244 10468 5296
rect 13452 5312 13504 5364
rect 13820 5312 13872 5364
rect 14740 5312 14792 5364
rect 17684 5312 17736 5364
rect 17868 5312 17920 5364
rect 14372 5244 14424 5296
rect 16028 5244 16080 5296
rect 3700 5108 3752 5160
rect 5816 5151 5868 5160
rect 5816 5117 5825 5151
rect 5825 5117 5859 5151
rect 5859 5117 5868 5151
rect 5816 5108 5868 5117
rect 6828 5108 6880 5160
rect 7656 5151 7708 5160
rect 7656 5117 7665 5151
rect 7665 5117 7699 5151
rect 7699 5117 7708 5151
rect 7656 5108 7708 5117
rect 9772 5151 9824 5160
rect 9772 5117 9781 5151
rect 9781 5117 9815 5151
rect 9815 5117 9824 5151
rect 9772 5108 9824 5117
rect 10600 5176 10652 5228
rect 11060 5176 11112 5228
rect 11520 5151 11572 5160
rect 11520 5117 11529 5151
rect 11529 5117 11563 5151
rect 11563 5117 11572 5151
rect 11520 5108 11572 5117
rect 13360 5176 13412 5228
rect 13544 5219 13596 5228
rect 13544 5185 13553 5219
rect 13553 5185 13587 5219
rect 13587 5185 13596 5219
rect 13544 5176 13596 5185
rect 16304 5219 16356 5228
rect 16304 5185 16313 5219
rect 16313 5185 16347 5219
rect 16347 5185 16356 5219
rect 16304 5176 16356 5185
rect 16948 5244 17000 5296
rect 12348 5108 12400 5160
rect 12440 5108 12492 5160
rect 16396 5151 16448 5160
rect 10784 5015 10836 5024
rect 10784 4981 10793 5015
rect 10793 4981 10827 5015
rect 10827 4981 10836 5015
rect 10784 4972 10836 4981
rect 11980 4972 12032 5024
rect 13360 5040 13412 5092
rect 16396 5117 16405 5151
rect 16405 5117 16439 5151
rect 16439 5117 16448 5151
rect 16396 5108 16448 5117
rect 17040 5151 17092 5160
rect 17040 5117 17049 5151
rect 17049 5117 17083 5151
rect 17083 5117 17092 5151
rect 17040 5108 17092 5117
rect 16764 5040 16816 5092
rect 17224 4972 17276 5024
rect 2995 4870 3047 4922
rect 3059 4870 3111 4922
rect 3123 4870 3175 4922
rect 3187 4870 3239 4922
rect 3251 4870 3303 4922
rect 9294 4870 9346 4922
rect 9358 4870 9410 4922
rect 9422 4870 9474 4922
rect 9486 4870 9538 4922
rect 9550 4870 9602 4922
rect 15592 4870 15644 4922
rect 15656 4870 15708 4922
rect 15720 4870 15772 4922
rect 15784 4870 15836 4922
rect 15848 4870 15900 4922
rect 7656 4768 7708 4820
rect 11520 4768 11572 4820
rect 12348 4768 12400 4820
rect 12532 4768 12584 4820
rect 12808 4768 12860 4820
rect 14280 4768 14332 4820
rect 14464 4811 14516 4820
rect 14464 4777 14473 4811
rect 14473 4777 14507 4811
rect 14507 4777 14516 4811
rect 14464 4768 14516 4777
rect 14556 4768 14608 4820
rect 17040 4768 17092 4820
rect 7380 4700 7432 4752
rect 8024 4743 8076 4752
rect 8024 4709 8033 4743
rect 8033 4709 8067 4743
rect 8067 4709 8076 4743
rect 8024 4700 8076 4709
rect 5540 4564 5592 4616
rect 8300 4564 8352 4616
rect 9036 4700 9088 4752
rect 8576 4675 8628 4684
rect 8576 4641 8585 4675
rect 8585 4641 8619 4675
rect 8619 4641 8628 4675
rect 8576 4632 8628 4641
rect 9956 4632 10008 4684
rect 10876 4632 10928 4684
rect 6000 4496 6052 4548
rect 7564 4496 7616 4548
rect 8208 4496 8260 4548
rect 8300 4428 8352 4480
rect 9220 4564 9272 4616
rect 11980 4607 12032 4616
rect 11980 4573 11989 4607
rect 11989 4573 12023 4607
rect 12023 4573 12032 4607
rect 11980 4564 12032 4573
rect 15384 4700 15436 4752
rect 13084 4632 13136 4684
rect 13360 4607 13412 4616
rect 13360 4573 13369 4607
rect 13369 4573 13403 4607
rect 13403 4573 13412 4607
rect 13360 4564 13412 4573
rect 13728 4564 13780 4616
rect 15200 4632 15252 4684
rect 16212 4632 16264 4684
rect 16764 4632 16816 4684
rect 12532 4539 12584 4548
rect 12532 4505 12541 4539
rect 12541 4505 12575 4539
rect 12575 4505 12584 4539
rect 14188 4564 14240 4616
rect 14924 4607 14976 4616
rect 14924 4573 14933 4607
rect 14933 4573 14967 4607
rect 14967 4573 14976 4607
rect 14924 4564 14976 4573
rect 15108 4607 15160 4616
rect 15108 4573 15117 4607
rect 15117 4573 15151 4607
rect 15151 4573 15160 4607
rect 15108 4564 15160 4573
rect 16672 4564 16724 4616
rect 17592 4607 17644 4616
rect 17592 4573 17601 4607
rect 17601 4573 17635 4607
rect 17635 4573 17644 4607
rect 17592 4564 17644 4573
rect 17960 4607 18012 4616
rect 17960 4573 17969 4607
rect 17969 4573 18003 4607
rect 18003 4573 18012 4607
rect 17960 4564 18012 4573
rect 18512 4607 18564 4616
rect 18512 4573 18521 4607
rect 18521 4573 18555 4607
rect 18555 4573 18564 4607
rect 18512 4564 18564 4573
rect 12532 4496 12584 4505
rect 8944 4471 8996 4480
rect 8944 4437 8953 4471
rect 8953 4437 8987 4471
rect 8987 4437 8996 4471
rect 8944 4428 8996 4437
rect 9128 4428 9180 4480
rect 12992 4471 13044 4480
rect 12992 4437 13001 4471
rect 13001 4437 13035 4471
rect 13035 4437 13044 4471
rect 12992 4428 13044 4437
rect 14004 4428 14056 4480
rect 14924 4428 14976 4480
rect 15108 4428 15160 4480
rect 16304 4428 16356 4480
rect 16948 4428 17000 4480
rect 6144 4326 6196 4378
rect 6208 4326 6260 4378
rect 6272 4326 6324 4378
rect 6336 4326 6388 4378
rect 6400 4326 6452 4378
rect 12443 4326 12495 4378
rect 12507 4326 12559 4378
rect 12571 4326 12623 4378
rect 12635 4326 12687 4378
rect 12699 4326 12751 4378
rect 6000 4224 6052 4276
rect 7380 4267 7432 4276
rect 7380 4233 7389 4267
rect 7389 4233 7423 4267
rect 7423 4233 7432 4267
rect 7380 4224 7432 4233
rect 10692 4224 10744 4276
rect 8852 4156 8904 4208
rect 9036 4199 9088 4208
rect 9036 4165 9045 4199
rect 9045 4165 9079 4199
rect 9079 4165 9088 4199
rect 9036 4156 9088 4165
rect 10600 4156 10652 4208
rect 10876 4199 10928 4208
rect 10876 4165 10885 4199
rect 10885 4165 10919 4199
rect 10919 4165 10928 4199
rect 10876 4156 10928 4165
rect 8484 4131 8536 4140
rect 7564 4063 7616 4072
rect 7564 4029 7573 4063
rect 7573 4029 7607 4063
rect 7607 4029 7616 4063
rect 7564 4020 7616 4029
rect 8484 4097 8493 4131
rect 8493 4097 8527 4131
rect 8527 4097 8536 4131
rect 8484 4088 8536 4097
rect 9680 4131 9732 4140
rect 9680 4097 9689 4131
rect 9689 4097 9723 4131
rect 9723 4097 9732 4131
rect 9680 4088 9732 4097
rect 10416 4088 10468 4140
rect 10692 4121 10744 4130
rect 10692 4087 10701 4121
rect 10701 4087 10735 4121
rect 10735 4087 10744 4121
rect 11060 4131 11112 4140
rect 10692 4078 10744 4087
rect 11060 4097 11069 4131
rect 11069 4097 11103 4131
rect 11103 4097 11112 4131
rect 11060 4088 11112 4097
rect 11520 4156 11572 4208
rect 8208 4020 8260 4072
rect 9220 4020 9272 4072
rect 9956 4063 10008 4072
rect 9956 4029 9965 4063
rect 9965 4029 9999 4063
rect 9999 4029 10008 4063
rect 9956 4020 10008 4029
rect 12440 4088 12492 4140
rect 12992 4156 13044 4208
rect 14464 4224 14516 4276
rect 16948 4224 17000 4276
rect 13452 4156 13504 4208
rect 15200 4156 15252 4208
rect 12808 4131 12860 4140
rect 12808 4097 12842 4131
rect 12842 4097 12860 4131
rect 12808 4088 12860 4097
rect 13084 4088 13136 4140
rect 18512 4131 18564 4140
rect 14004 4063 14056 4072
rect 14004 4029 14013 4063
rect 14013 4029 14047 4063
rect 14047 4029 14056 4063
rect 14004 4020 14056 4029
rect 8208 3884 8260 3936
rect 8944 3927 8996 3936
rect 8944 3893 8953 3927
rect 8953 3893 8987 3927
rect 8987 3893 8996 3927
rect 8944 3884 8996 3893
rect 12900 3884 12952 3936
rect 15200 3884 15252 3936
rect 18512 4097 18521 4131
rect 18521 4097 18555 4131
rect 18555 4097 18564 4131
rect 18512 4088 18564 4097
rect 17224 4020 17276 4072
rect 17960 4020 18012 4072
rect 18052 3884 18104 3936
rect 2995 3782 3047 3834
rect 3059 3782 3111 3834
rect 3123 3782 3175 3834
rect 3187 3782 3239 3834
rect 3251 3782 3303 3834
rect 9294 3782 9346 3834
rect 9358 3782 9410 3834
rect 9422 3782 9474 3834
rect 9486 3782 9538 3834
rect 9550 3782 9602 3834
rect 15592 3782 15644 3834
rect 15656 3782 15708 3834
rect 15720 3782 15772 3834
rect 15784 3782 15836 3834
rect 15848 3782 15900 3834
rect 5908 3680 5960 3732
rect 8484 3680 8536 3732
rect 10600 3680 10652 3732
rect 11060 3680 11112 3732
rect 5264 3655 5316 3664
rect 5264 3621 5273 3655
rect 5273 3621 5307 3655
rect 5307 3621 5316 3655
rect 5264 3612 5316 3621
rect 3332 3476 3384 3528
rect 5356 3519 5408 3528
rect 5356 3485 5365 3519
rect 5365 3485 5399 3519
rect 5399 3485 5408 3519
rect 5356 3476 5408 3485
rect 8944 3544 8996 3596
rect 8208 3519 8260 3528
rect 8208 3485 8217 3519
rect 8217 3485 8251 3519
rect 8251 3485 8260 3519
rect 8208 3476 8260 3485
rect 9772 3476 9824 3528
rect 11888 3476 11940 3528
rect 12532 3587 12584 3596
rect 12532 3553 12541 3587
rect 12541 3553 12575 3587
rect 12575 3553 12584 3587
rect 12532 3544 12584 3553
rect 12992 3680 13044 3732
rect 13268 3680 13320 3732
rect 15108 3680 15160 3732
rect 13544 3612 13596 3664
rect 13636 3612 13688 3664
rect 15384 3612 15436 3664
rect 17960 3544 18012 3596
rect 5540 3408 5592 3460
rect 5816 3408 5868 3460
rect 3240 3340 3292 3392
rect 3608 3340 3660 3392
rect 7012 3340 7064 3392
rect 8300 3340 8352 3392
rect 8576 3408 8628 3460
rect 12900 3476 12952 3528
rect 13360 3519 13412 3528
rect 13360 3485 13369 3519
rect 13369 3485 13403 3519
rect 13403 3485 13412 3519
rect 13360 3476 13412 3485
rect 13636 3519 13688 3528
rect 13636 3485 13645 3519
rect 13645 3485 13679 3519
rect 13679 3485 13688 3519
rect 13636 3476 13688 3485
rect 14464 3476 14516 3528
rect 13452 3408 13504 3460
rect 8852 3340 8904 3392
rect 14556 3340 14608 3392
rect 15016 3519 15068 3528
rect 15016 3485 15025 3519
rect 15025 3485 15059 3519
rect 15059 3485 15068 3519
rect 15200 3519 15252 3528
rect 15016 3476 15068 3485
rect 15200 3485 15209 3519
rect 15209 3485 15243 3519
rect 15243 3485 15252 3519
rect 15200 3476 15252 3485
rect 16948 3408 17000 3460
rect 18052 3408 18104 3460
rect 14924 3383 14976 3392
rect 14924 3349 14933 3383
rect 14933 3349 14967 3383
rect 14967 3349 14976 3383
rect 14924 3340 14976 3349
rect 16580 3340 16632 3392
rect 6144 3238 6196 3290
rect 6208 3238 6260 3290
rect 6272 3238 6324 3290
rect 6336 3238 6388 3290
rect 6400 3238 6452 3290
rect 12443 3238 12495 3290
rect 12507 3238 12559 3290
rect 12571 3238 12623 3290
rect 12635 3238 12687 3290
rect 12699 3238 12751 3290
rect 5816 3179 5868 3188
rect 5816 3145 5825 3179
rect 5825 3145 5859 3179
rect 5859 3145 5868 3179
rect 5816 3136 5868 3145
rect 5908 3136 5960 3188
rect 4344 3068 4396 3120
rect 3240 3043 3292 3052
rect 3240 3009 3249 3043
rect 3249 3009 3283 3043
rect 3283 3009 3292 3043
rect 3240 3000 3292 3009
rect 3608 3043 3660 3052
rect 3608 3009 3617 3043
rect 3617 3009 3651 3043
rect 3651 3009 3660 3043
rect 3608 3000 3660 3009
rect 4896 3000 4948 3052
rect 5632 3000 5684 3052
rect 5908 3000 5960 3052
rect 7012 3136 7064 3188
rect 8300 3136 8352 3188
rect 6460 3043 6512 3052
rect 6460 3009 6469 3043
rect 6469 3009 6503 3043
rect 6503 3009 6512 3043
rect 6460 3000 6512 3009
rect 9220 3136 9272 3188
rect 10416 3136 10468 3188
rect 11520 3136 11572 3188
rect 12808 3136 12860 3188
rect 13912 3136 13964 3188
rect 14832 3136 14884 3188
rect 6368 2932 6420 2984
rect 6552 2975 6604 2984
rect 6552 2941 6561 2975
rect 6561 2941 6595 2975
rect 6595 2941 6604 2975
rect 7012 3043 7064 3052
rect 6552 2932 6604 2941
rect 5356 2907 5408 2916
rect 5356 2873 5365 2907
rect 5365 2873 5399 2907
rect 5399 2873 5408 2907
rect 5356 2864 5408 2873
rect 6460 2864 6512 2916
rect 5908 2796 5960 2848
rect 7012 3009 7021 3043
rect 7021 3009 7055 3043
rect 7055 3009 7064 3043
rect 7012 3000 7064 3009
rect 13360 3068 13412 3120
rect 13636 3068 13688 3120
rect 8116 3043 8168 3052
rect 8116 3009 8125 3043
rect 8125 3009 8159 3043
rect 8159 3009 8168 3043
rect 8116 3000 8168 3009
rect 8852 3000 8904 3052
rect 12072 3043 12124 3052
rect 8668 2932 8720 2984
rect 8944 2932 8996 2984
rect 12072 3009 12081 3043
rect 12081 3009 12115 3043
rect 12115 3009 12124 3043
rect 12072 3000 12124 3009
rect 13084 3043 13136 3052
rect 13084 3009 13093 3043
rect 13093 3009 13127 3043
rect 13127 3009 13136 3043
rect 13084 3000 13136 3009
rect 12808 2932 12860 2984
rect 14372 3043 14424 3052
rect 13452 2932 13504 2984
rect 10048 2864 10100 2916
rect 13084 2864 13136 2916
rect 14372 3009 14381 3043
rect 14381 3009 14415 3043
rect 14415 3009 14424 3043
rect 14372 3000 14424 3009
rect 14556 3043 14608 3052
rect 14556 3009 14565 3043
rect 14565 3009 14599 3043
rect 14599 3009 14608 3043
rect 14556 3000 14608 3009
rect 14924 3068 14976 3120
rect 17592 3136 17644 3188
rect 16948 3068 17000 3120
rect 15016 3000 15068 3052
rect 14740 2932 14792 2984
rect 15384 3043 15436 3052
rect 15384 3009 15393 3043
rect 15393 3009 15427 3043
rect 15427 3009 15436 3043
rect 15384 3000 15436 3009
rect 17960 3000 18012 3052
rect 18420 3000 18472 3052
rect 18604 3000 18656 3052
rect 16028 2975 16080 2984
rect 16028 2941 16037 2975
rect 16037 2941 16071 2975
rect 16071 2941 16080 2975
rect 16028 2932 16080 2941
rect 16120 2975 16172 2984
rect 16120 2941 16129 2975
rect 16129 2941 16163 2975
rect 16163 2941 16172 2975
rect 16120 2932 16172 2941
rect 16396 2932 16448 2984
rect 15016 2864 15068 2916
rect 7932 2839 7984 2848
rect 7932 2805 7941 2839
rect 7941 2805 7975 2839
rect 7975 2805 7984 2839
rect 7932 2796 7984 2805
rect 9680 2796 9732 2848
rect 10968 2796 11020 2848
rect 13268 2839 13320 2848
rect 13268 2805 13277 2839
rect 13277 2805 13311 2839
rect 13311 2805 13320 2839
rect 13268 2796 13320 2805
rect 13360 2796 13412 2848
rect 13820 2796 13872 2848
rect 14280 2796 14332 2848
rect 15108 2796 15160 2848
rect 18328 2839 18380 2848
rect 18328 2805 18337 2839
rect 18337 2805 18371 2839
rect 18371 2805 18380 2839
rect 18328 2796 18380 2805
rect 2995 2694 3047 2746
rect 3059 2694 3111 2746
rect 3123 2694 3175 2746
rect 3187 2694 3239 2746
rect 3251 2694 3303 2746
rect 9294 2694 9346 2746
rect 9358 2694 9410 2746
rect 9422 2694 9474 2746
rect 9486 2694 9538 2746
rect 9550 2694 9602 2746
rect 15592 2694 15644 2746
rect 15656 2694 15708 2746
rect 15720 2694 15772 2746
rect 15784 2694 15836 2746
rect 15848 2694 15900 2746
rect 6000 2592 6052 2644
rect 5080 2456 5132 2508
rect 5632 2456 5684 2508
rect 9680 2592 9732 2644
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 5724 2431 5776 2440
rect 5724 2397 5733 2431
rect 5733 2397 5767 2431
rect 5767 2397 5776 2431
rect 5724 2388 5776 2397
rect 6000 2388 6052 2440
rect 6552 2524 6604 2576
rect 8024 2524 8076 2576
rect 6828 2431 6880 2440
rect 6828 2397 6837 2431
rect 6837 2397 6871 2431
rect 6871 2397 6880 2431
rect 7932 2456 7984 2508
rect 8668 2456 8720 2508
rect 9220 2499 9272 2508
rect 9220 2465 9229 2499
rect 9229 2465 9263 2499
rect 9263 2465 9272 2499
rect 11888 2592 11940 2644
rect 12072 2592 12124 2644
rect 13176 2592 13228 2644
rect 14372 2592 14424 2644
rect 16120 2592 16172 2644
rect 13360 2524 13412 2576
rect 17868 2524 17920 2576
rect 9220 2456 9272 2465
rect 6828 2388 6880 2397
rect 8392 2320 8444 2372
rect 9312 2388 9364 2440
rect 14004 2499 14056 2508
rect 14004 2465 14013 2499
rect 14013 2465 14047 2499
rect 14047 2465 14056 2499
rect 14004 2456 14056 2465
rect 16396 2499 16448 2508
rect 16396 2465 16405 2499
rect 16405 2465 16439 2499
rect 16439 2465 16448 2499
rect 16396 2456 16448 2465
rect 9588 2431 9640 2440
rect 9588 2397 9597 2431
rect 9597 2397 9631 2431
rect 9631 2397 9640 2431
rect 9588 2388 9640 2397
rect 10048 2431 10100 2440
rect 10048 2397 10057 2431
rect 10057 2397 10091 2431
rect 10091 2397 10100 2431
rect 10048 2388 10100 2397
rect 3608 2252 3660 2304
rect 7748 2252 7800 2304
rect 8208 2295 8260 2304
rect 8208 2261 8217 2295
rect 8217 2261 8251 2295
rect 8251 2261 8260 2295
rect 8208 2252 8260 2261
rect 8484 2252 8536 2304
rect 9128 2252 9180 2304
rect 9496 2252 9548 2304
rect 9864 2295 9916 2304
rect 9864 2261 9873 2295
rect 9873 2261 9907 2295
rect 9907 2261 9916 2295
rect 9864 2252 9916 2261
rect 13084 2431 13136 2440
rect 13084 2397 13093 2431
rect 13093 2397 13127 2431
rect 13127 2397 13136 2431
rect 13084 2388 13136 2397
rect 11796 2320 11848 2372
rect 12900 2320 12952 2372
rect 13360 2388 13412 2440
rect 13820 2431 13872 2440
rect 13820 2397 13829 2431
rect 13829 2397 13863 2431
rect 13863 2397 13872 2431
rect 13820 2388 13872 2397
rect 14280 2363 14332 2372
rect 14280 2329 14289 2363
rect 14289 2329 14323 2363
rect 14323 2329 14332 2363
rect 14280 2320 14332 2329
rect 15568 2320 15620 2372
rect 16488 2320 16540 2372
rect 16948 2320 17000 2372
rect 17684 2320 17736 2372
rect 13820 2252 13872 2304
rect 15108 2252 15160 2304
rect 17776 2252 17828 2304
rect 6144 2150 6196 2202
rect 6208 2150 6260 2202
rect 6272 2150 6324 2202
rect 6336 2150 6388 2202
rect 6400 2150 6452 2202
rect 12443 2150 12495 2202
rect 12507 2150 12559 2202
rect 12571 2150 12623 2202
rect 12635 2150 12687 2202
rect 12699 2150 12751 2202
rect 5080 2091 5132 2100
rect 5080 2057 5089 2091
rect 5089 2057 5123 2091
rect 5123 2057 5132 2091
rect 5080 2048 5132 2057
rect 5264 2091 5316 2100
rect 5264 2057 5273 2091
rect 5273 2057 5307 2091
rect 5307 2057 5316 2091
rect 5264 2048 5316 2057
rect 5724 2048 5776 2100
rect 3608 2023 3660 2032
rect 3608 1989 3617 2023
rect 3617 1989 3651 2023
rect 3651 1989 3660 2023
rect 3608 1980 3660 1989
rect 4896 1980 4948 2032
rect 3332 1955 3384 1964
rect 3332 1921 3341 1955
rect 3341 1921 3375 1955
rect 3375 1921 3384 1955
rect 3332 1912 3384 1921
rect 5448 1980 5500 2032
rect 8024 2048 8076 2100
rect 8944 2091 8996 2100
rect 7932 1980 7984 2032
rect 8944 2057 8953 2091
rect 8953 2057 8987 2091
rect 8987 2057 8996 2091
rect 8944 2048 8996 2057
rect 5816 1955 5868 1964
rect 5816 1921 5825 1955
rect 5825 1921 5859 1955
rect 5859 1921 5868 1955
rect 5816 1912 5868 1921
rect 5908 1912 5960 1964
rect 6552 1912 6604 1964
rect 7564 1912 7616 1964
rect 8116 1912 8168 1964
rect 8392 1955 8444 1964
rect 8392 1921 8401 1955
rect 8401 1921 8435 1955
rect 8435 1921 8444 1955
rect 8392 1912 8444 1921
rect 8668 1955 8720 1964
rect 8668 1921 8677 1955
rect 8677 1921 8711 1955
rect 8711 1921 8720 1955
rect 9128 1980 9180 2032
rect 9496 2048 9548 2100
rect 9864 1980 9916 2032
rect 11520 1980 11572 2032
rect 8668 1912 8720 1921
rect 6828 1844 6880 1896
rect 9312 1955 9364 1964
rect 9312 1921 9321 1955
rect 9321 1921 9355 1955
rect 9355 1921 9364 1955
rect 9312 1912 9364 1921
rect 9496 1955 9548 1964
rect 9496 1921 9505 1955
rect 9505 1921 9539 1955
rect 9539 1921 9548 1955
rect 9496 1912 9548 1921
rect 9772 1955 9824 1964
rect 9772 1921 9781 1955
rect 9781 1921 9815 1955
rect 9815 1921 9824 1955
rect 9772 1912 9824 1921
rect 9956 1912 10008 1964
rect 10968 1955 11020 1964
rect 10508 1844 10560 1896
rect 10968 1921 10977 1955
rect 10977 1921 11011 1955
rect 11011 1921 11020 1955
rect 10968 1912 11020 1921
rect 16580 2048 16632 2100
rect 16948 2048 17000 2100
rect 12072 1980 12124 2032
rect 14832 1980 14884 2032
rect 18328 1980 18380 2032
rect 11888 1844 11940 1896
rect 8484 1776 8536 1828
rect 6644 1708 6696 1760
rect 8300 1708 8352 1760
rect 8668 1708 8720 1760
rect 10048 1776 10100 1828
rect 12808 1912 12860 1964
rect 13084 1887 13136 1896
rect 13084 1853 13093 1887
rect 13093 1853 13127 1887
rect 13127 1853 13136 1887
rect 13544 1912 13596 1964
rect 14280 1955 14332 1964
rect 13084 1844 13136 1853
rect 13820 1844 13872 1896
rect 14280 1921 14289 1955
rect 14289 1921 14323 1955
rect 14323 1921 14332 1955
rect 14280 1912 14332 1921
rect 14924 1955 14976 1964
rect 14924 1921 14933 1955
rect 14933 1921 14967 1955
rect 14967 1921 14976 1955
rect 14924 1912 14976 1921
rect 15384 1912 15436 1964
rect 15108 1887 15160 1896
rect 15108 1853 15117 1887
rect 15117 1853 15151 1887
rect 15151 1853 15160 1887
rect 16948 1912 17000 1964
rect 18512 1955 18564 1964
rect 18512 1921 18521 1955
rect 18521 1921 18555 1955
rect 18555 1921 18564 1955
rect 18512 1912 18564 1921
rect 15108 1844 15160 1853
rect 16580 1887 16632 1896
rect 14188 1776 14240 1828
rect 15384 1776 15436 1828
rect 16304 1776 16356 1828
rect 16580 1853 16589 1887
rect 16589 1853 16623 1887
rect 16623 1853 16632 1887
rect 16580 1844 16632 1853
rect 17040 1776 17092 1828
rect 9220 1708 9272 1760
rect 9864 1708 9916 1760
rect 12808 1708 12860 1760
rect 13268 1751 13320 1760
rect 13268 1717 13277 1751
rect 13277 1717 13311 1751
rect 13311 1717 13320 1751
rect 13268 1708 13320 1717
rect 14832 1708 14884 1760
rect 15476 1708 15528 1760
rect 15936 1751 15988 1760
rect 15936 1717 15945 1751
rect 15945 1717 15979 1751
rect 15979 1717 15988 1751
rect 15936 1708 15988 1717
rect 2995 1606 3047 1658
rect 3059 1606 3111 1658
rect 3123 1606 3175 1658
rect 3187 1606 3239 1658
rect 3251 1606 3303 1658
rect 9294 1606 9346 1658
rect 9358 1606 9410 1658
rect 9422 1606 9474 1658
rect 9486 1606 9538 1658
rect 9550 1606 9602 1658
rect 15592 1606 15644 1658
rect 15656 1606 15708 1658
rect 15720 1606 15772 1658
rect 15784 1606 15836 1658
rect 15848 1606 15900 1658
rect 8484 1436 8536 1488
rect 14924 1504 14976 1556
rect 15016 1547 15068 1556
rect 15016 1513 15025 1547
rect 15025 1513 15059 1547
rect 15059 1513 15068 1547
rect 15016 1504 15068 1513
rect 16948 1504 17000 1556
rect 6920 1368 6972 1420
rect 8024 1368 8076 1420
rect 7564 1343 7616 1352
rect 7564 1309 7573 1343
rect 7573 1309 7607 1343
rect 7607 1309 7616 1343
rect 7564 1300 7616 1309
rect 7748 1300 7800 1352
rect 8760 1343 8812 1352
rect 8760 1309 8769 1343
rect 8769 1309 8803 1343
rect 8803 1309 8812 1343
rect 8760 1300 8812 1309
rect 9036 1300 9088 1352
rect 10416 1436 10468 1488
rect 10692 1368 10744 1420
rect 10968 1368 11020 1420
rect 14188 1436 14240 1488
rect 14464 1411 14516 1420
rect 14464 1377 14473 1411
rect 14473 1377 14507 1411
rect 14507 1377 14516 1411
rect 14464 1368 14516 1377
rect 15476 1368 15528 1420
rect 15936 1368 15988 1420
rect 16120 1411 16172 1420
rect 16120 1377 16129 1411
rect 16129 1377 16163 1411
rect 16163 1377 16172 1411
rect 16120 1368 16172 1377
rect 16580 1368 16632 1420
rect 17040 1368 17092 1420
rect 17776 1411 17828 1420
rect 17776 1377 17785 1411
rect 17785 1377 17819 1411
rect 17819 1377 17828 1411
rect 17776 1368 17828 1377
rect 7012 1232 7064 1284
rect 5540 1164 5592 1216
rect 6552 1164 6604 1216
rect 7472 1164 7524 1216
rect 8944 1164 8996 1216
rect 9128 1164 9180 1216
rect 9772 1164 9824 1216
rect 10600 1164 10652 1216
rect 11060 1207 11112 1216
rect 11060 1173 11069 1207
rect 11069 1173 11103 1207
rect 11103 1173 11112 1207
rect 11060 1164 11112 1173
rect 11888 1300 11940 1352
rect 14280 1300 14332 1352
rect 14832 1343 14884 1352
rect 14832 1309 14841 1343
rect 14841 1309 14875 1343
rect 14875 1309 14884 1343
rect 14832 1300 14884 1309
rect 15384 1343 15436 1352
rect 15384 1309 15393 1343
rect 15393 1309 15427 1343
rect 15427 1309 15436 1343
rect 15384 1300 15436 1309
rect 14740 1232 14792 1284
rect 16028 1232 16080 1284
rect 11888 1207 11940 1216
rect 11888 1173 11897 1207
rect 11897 1173 11931 1207
rect 11931 1173 11940 1207
rect 11888 1164 11940 1173
rect 15936 1164 15988 1216
rect 17960 1232 18012 1284
rect 16764 1207 16816 1216
rect 16764 1173 16773 1207
rect 16773 1173 16807 1207
rect 16807 1173 16816 1207
rect 16764 1164 16816 1173
rect 17408 1164 17460 1216
rect 6144 1062 6196 1114
rect 6208 1062 6260 1114
rect 6272 1062 6324 1114
rect 6336 1062 6388 1114
rect 6400 1062 6452 1114
rect 12443 1062 12495 1114
rect 12507 1062 12559 1114
rect 12571 1062 12623 1114
rect 12635 1062 12687 1114
rect 12699 1062 12751 1114
rect 6828 960 6880 1012
rect 7472 960 7524 1012
rect 6644 892 6696 944
rect 8208 892 8260 944
rect 8760 960 8812 1012
rect 9588 960 9640 1012
rect 10508 1003 10560 1012
rect 10508 969 10517 1003
rect 10517 969 10551 1003
rect 10551 969 10560 1003
rect 10508 960 10560 969
rect 11060 960 11112 1012
rect 12072 1003 12124 1012
rect 12072 969 12081 1003
rect 12081 969 12115 1003
rect 12115 969 12124 1003
rect 12072 960 12124 969
rect 14464 960 14516 1012
rect 16764 960 16816 1012
rect 17868 1003 17920 1012
rect 17868 969 17877 1003
rect 17877 969 17911 1003
rect 17911 969 17920 1003
rect 17868 960 17920 969
rect 17960 1003 18012 1012
rect 17960 969 17969 1003
rect 17969 969 18003 1003
rect 18003 969 18012 1003
rect 18420 1003 18472 1012
rect 17960 960 18012 969
rect 18420 969 18429 1003
rect 18429 969 18463 1003
rect 18463 969 18472 1003
rect 18420 960 18472 969
rect 8852 935 8904 944
rect 8852 901 8861 935
rect 8861 901 8895 935
rect 8895 901 8904 935
rect 8852 892 8904 901
rect 8944 892 8996 944
rect 6552 867 6604 876
rect 6552 833 6561 867
rect 6561 833 6595 867
rect 6595 833 6604 867
rect 7196 867 7248 876
rect 6552 824 6604 833
rect 7196 833 7205 867
rect 7205 833 7239 867
rect 7239 833 7248 867
rect 7196 824 7248 833
rect 9680 892 9732 944
rect 11152 892 11204 944
rect 9220 799 9272 808
rect 9220 765 9229 799
rect 9229 765 9263 799
rect 9263 765 9272 799
rect 9220 756 9272 765
rect 10140 867 10192 876
rect 10140 833 10149 867
rect 10149 833 10183 867
rect 10183 833 10192 867
rect 10140 824 10192 833
rect 10692 867 10744 876
rect 10692 833 10701 867
rect 10701 833 10735 867
rect 10735 833 10744 867
rect 10692 824 10744 833
rect 11796 892 11848 944
rect 13268 892 13320 944
rect 16856 892 16908 944
rect 9864 799 9916 808
rect 9864 765 9873 799
rect 9873 765 9907 799
rect 9907 765 9916 799
rect 9864 756 9916 765
rect 11060 756 11112 808
rect 14004 824 14056 876
rect 14740 824 14792 876
rect 15384 824 15436 876
rect 15936 867 15988 876
rect 15936 833 15945 867
rect 15945 833 15979 867
rect 15979 833 15988 867
rect 15936 824 15988 833
rect 18328 867 18380 876
rect 18328 833 18337 867
rect 18337 833 18371 867
rect 18371 833 18380 867
rect 18328 824 18380 833
rect 8024 688 8076 740
rect 17776 756 17828 808
rect 7748 620 7800 672
rect 9036 620 9088 672
rect 17132 620 17184 672
rect 2995 518 3047 570
rect 3059 518 3111 570
rect 3123 518 3175 570
rect 3187 518 3239 570
rect 3251 518 3303 570
rect 9294 518 9346 570
rect 9358 518 9410 570
rect 9422 518 9474 570
rect 9486 518 9538 570
rect 9550 518 9602 570
rect 15592 518 15644 570
rect 15656 518 15708 570
rect 15720 518 15772 570
rect 15784 518 15836 570
rect 15848 518 15900 570
rect 7564 416 7616 468
rect 11888 416 11940 468
rect 17408 459 17460 468
rect 17408 425 17417 459
rect 17417 425 17451 459
rect 17451 425 17460 459
rect 17408 416 17460 425
rect 18328 459 18380 468
rect 18328 425 18337 459
rect 18337 425 18371 459
rect 18371 425 18380 459
rect 18328 416 18380 425
rect 8392 323 8444 332
rect 8392 289 8401 323
rect 8401 289 8435 323
rect 8435 289 8444 323
rect 8392 280 8444 289
rect 9036 280 9088 332
rect 10140 323 10192 332
rect 10140 289 10149 323
rect 10149 289 10183 323
rect 10183 289 10192 323
rect 10140 280 10192 289
rect 7472 255 7524 264
rect 7472 221 7481 255
rect 7481 221 7515 255
rect 7515 221 7524 255
rect 7472 212 7524 221
rect 14740 280 14792 332
rect 17684 280 17736 332
rect 11060 255 11112 264
rect 11060 221 11069 255
rect 11069 221 11103 255
rect 11103 221 11112 255
rect 11060 212 11112 221
rect 11152 212 11204 264
rect 17132 255 17184 264
rect 17132 221 17141 255
rect 17141 221 17175 255
rect 17175 221 17184 255
rect 17132 212 17184 221
rect 18512 255 18564 264
rect 18512 221 18521 255
rect 18521 221 18555 255
rect 18555 221 18564 255
rect 18512 212 18564 221
rect 8208 144 8260 196
rect 6144 -26 6196 26
rect 6208 -26 6260 26
rect 6272 -26 6324 26
rect 6336 -26 6388 26
rect 6400 -26 6452 26
rect 12443 -26 12495 26
rect 12507 -26 12559 26
rect 12571 -26 12623 26
rect 12635 -26 12687 26
rect 12699 -26 12751 26
<< metal2 >>
rect 1398 11200 1454 12000
rect 4250 11200 4306 12000
rect 7102 11200 7158 12000
rect 9954 11200 10010 12000
rect 12806 11200 12862 12000
rect 15396 11206 15608 11234
rect 1412 9602 1440 11200
rect 1320 9586 1440 9602
rect 1308 9580 1440 9586
rect 1360 9574 1440 9580
rect 1308 9522 1360 9528
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2332 9178 2360 9454
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 572 8968 624 8974
rect 572 8910 624 8916
rect 388 8832 440 8838
rect 388 8774 440 8780
rect 400 8498 428 8774
rect 388 8492 440 8498
rect 388 8434 440 8440
rect 584 7410 612 8910
rect 2332 8566 2360 9114
rect 2700 8974 2728 9454
rect 2995 9276 3303 9296
rect 2995 9274 3001 9276
rect 3057 9274 3081 9276
rect 3137 9274 3161 9276
rect 3217 9274 3241 9276
rect 3297 9274 3303 9276
rect 3057 9222 3059 9274
rect 3239 9222 3241 9274
rect 2995 9220 3001 9222
rect 3057 9220 3081 9222
rect 3137 9220 3161 9222
rect 3217 9220 3241 9222
rect 3297 9220 3303 9222
rect 2995 9200 3303 9220
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2964 8900 3016 8906
rect 2964 8842 3016 8848
rect 2976 8634 3004 8842
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 1952 8560 2004 8566
rect 1952 8502 2004 8508
rect 2320 8560 2372 8566
rect 2320 8502 2372 8508
rect 756 8424 808 8430
rect 756 8366 808 8372
rect 768 8090 796 8366
rect 756 8084 808 8090
rect 756 8026 808 8032
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 1872 7546 1900 7822
rect 1860 7540 1912 7546
rect 1860 7482 1912 7488
rect 1964 7410 1992 8502
rect 3896 8498 3924 8774
rect 2964 8492 3016 8498
rect 2884 8452 2964 8480
rect 2412 8288 2464 8294
rect 2412 8230 2464 8236
rect 2320 8084 2372 8090
rect 2320 8026 2372 8032
rect 2332 7750 2360 8026
rect 2424 7886 2452 8230
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2320 7744 2372 7750
rect 2320 7686 2372 7692
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2516 7478 2544 7686
rect 2504 7472 2556 7478
rect 2504 7414 2556 7420
rect 2700 7410 2728 7822
rect 2884 7478 2912 8452
rect 3332 8492 3384 8498
rect 3016 8452 3332 8480
rect 2964 8434 3016 8440
rect 3332 8434 3384 8440
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 3792 8424 3844 8430
rect 3792 8366 3844 8372
rect 3332 8356 3384 8362
rect 3332 8298 3384 8304
rect 2995 8188 3303 8208
rect 2995 8186 3001 8188
rect 3057 8186 3081 8188
rect 3137 8186 3161 8188
rect 3217 8186 3241 8188
rect 3297 8186 3303 8188
rect 3057 8134 3059 8186
rect 3239 8134 3241 8186
rect 2995 8132 3001 8134
rect 3057 8132 3081 8134
rect 3137 8132 3161 8134
rect 3217 8132 3241 8134
rect 3297 8132 3303 8134
rect 2995 8112 3303 8132
rect 3344 8090 3372 8298
rect 3608 8288 3660 8294
rect 3608 8230 3660 8236
rect 3332 8084 3384 8090
rect 3332 8026 3384 8032
rect 3056 8016 3108 8022
rect 3056 7958 3108 7964
rect 3068 7546 3096 7958
rect 3620 7886 3648 8230
rect 3804 8090 3832 8366
rect 4172 8090 4200 8434
rect 3792 8084 3844 8090
rect 3712 8044 3792 8072
rect 3712 7954 3740 8044
rect 3792 8026 3844 8032
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 3700 7948 3752 7954
rect 3700 7890 3752 7896
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 4080 7546 4108 7822
rect 4172 7818 4200 8026
rect 4264 8022 4292 11200
rect 6144 9820 6452 9840
rect 6144 9818 6150 9820
rect 6206 9818 6230 9820
rect 6286 9818 6310 9820
rect 6366 9818 6390 9820
rect 6446 9818 6452 9820
rect 6206 9766 6208 9818
rect 6388 9766 6390 9818
rect 6144 9764 6150 9766
rect 6206 9764 6230 9766
rect 6286 9764 6310 9766
rect 6366 9764 6390 9766
rect 6446 9764 6452 9766
rect 6144 9744 6452 9764
rect 5632 9648 5684 9654
rect 5632 9590 5684 9596
rect 5644 9178 5672 9590
rect 5724 9512 5776 9518
rect 5724 9454 5776 9460
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5644 8974 5672 9114
rect 5736 9042 5764 9454
rect 7116 9450 7144 11200
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 7288 9512 7340 9518
rect 7288 9454 7340 9460
rect 7104 9444 7156 9450
rect 7104 9386 7156 9392
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 6736 8900 6788 8906
rect 6736 8842 6788 8848
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 4252 8016 4304 8022
rect 4252 7958 4304 7964
rect 4356 7886 4384 8774
rect 5460 8566 5488 8774
rect 6144 8732 6452 8752
rect 6144 8730 6150 8732
rect 6206 8730 6230 8732
rect 6286 8730 6310 8732
rect 6366 8730 6390 8732
rect 6446 8730 6452 8732
rect 6206 8678 6208 8730
rect 6388 8678 6390 8730
rect 6144 8676 6150 8678
rect 6206 8676 6230 8678
rect 6286 8676 6310 8678
rect 6366 8676 6390 8678
rect 6446 8676 6452 8678
rect 6144 8656 6452 8676
rect 6748 8634 6776 8842
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6460 8424 6512 8430
rect 6460 8366 6512 8372
rect 6472 8090 6500 8366
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 5552 7886 5580 8026
rect 6472 7954 6500 8026
rect 6368 7948 6420 7954
rect 6368 7890 6420 7896
rect 6460 7948 6512 7954
rect 6460 7890 6512 7896
rect 4344 7880 4396 7886
rect 4264 7840 4344 7868
rect 4160 7812 4212 7818
rect 4160 7754 4212 7760
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 2872 7472 2924 7478
rect 2872 7414 2924 7420
rect 572 7404 624 7410
rect 572 7346 624 7352
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 584 6322 612 7346
rect 1964 7274 1992 7346
rect 4172 7274 4200 7754
rect 4264 7478 4292 7840
rect 4344 7822 4396 7828
rect 5540 7880 5592 7886
rect 5908 7880 5960 7886
rect 5540 7822 5592 7828
rect 5630 7848 5686 7857
rect 6380 7857 6408 7890
rect 5908 7822 5960 7828
rect 6366 7848 6422 7857
rect 5630 7783 5686 7792
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 4252 7472 4304 7478
rect 4252 7414 4304 7420
rect 1952 7268 2004 7274
rect 1952 7210 2004 7216
rect 2596 7268 2648 7274
rect 2596 7210 2648 7216
rect 4160 7268 4212 7274
rect 4160 7210 4212 7216
rect 1676 6656 1728 6662
rect 1676 6598 1728 6604
rect 1688 6390 1716 6598
rect 2608 6458 2636 7210
rect 2995 7100 3303 7120
rect 2995 7098 3001 7100
rect 3057 7098 3081 7100
rect 3137 7098 3161 7100
rect 3217 7098 3241 7100
rect 3297 7098 3303 7100
rect 3057 7046 3059 7098
rect 3239 7046 3241 7098
rect 2995 7044 3001 7046
rect 3057 7044 3081 7046
rect 3137 7044 3161 7046
rect 3217 7044 3241 7046
rect 3297 7044 3303 7046
rect 2995 7024 3303 7044
rect 3608 6928 3660 6934
rect 3608 6870 3660 6876
rect 3620 6798 3648 6870
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 3608 6792 3660 6798
rect 3608 6734 3660 6740
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3068 6458 3096 6734
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 1676 6384 1728 6390
rect 1676 6326 1728 6332
rect 572 6316 624 6322
rect 572 6258 624 6264
rect 584 5778 612 6258
rect 572 5772 624 5778
rect 572 5714 624 5720
rect 2608 5642 2636 6394
rect 3252 6322 3280 6598
rect 3608 6384 3660 6390
rect 3608 6326 3660 6332
rect 3240 6316 3292 6322
rect 3292 6276 3464 6304
rect 3240 6258 3292 6264
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 2995 6012 3303 6032
rect 2995 6010 3001 6012
rect 3057 6010 3081 6012
rect 3137 6010 3161 6012
rect 3217 6010 3241 6012
rect 3297 6010 3303 6012
rect 3057 5958 3059 6010
rect 3239 5958 3241 6010
rect 2995 5956 3001 5958
rect 3057 5956 3081 5958
rect 3137 5956 3161 5958
rect 3217 5956 3241 5958
rect 3297 5956 3303 5958
rect 2995 5936 3303 5956
rect 3344 5846 3372 6054
rect 3332 5840 3384 5846
rect 3332 5782 3384 5788
rect 3332 5704 3384 5710
rect 3436 5692 3464 6276
rect 3620 5710 3648 6326
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 3804 5846 3832 6258
rect 3896 6186 3924 6734
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 4264 6458 4292 6598
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4356 6254 4384 7686
rect 4816 7410 4844 7686
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 5000 6866 5028 7142
rect 5460 7002 5488 7686
rect 5644 7410 5672 7783
rect 5920 7546 5948 7822
rect 6366 7783 6422 7792
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6144 7644 6452 7664
rect 6144 7642 6150 7644
rect 6206 7642 6230 7644
rect 6286 7642 6310 7644
rect 6366 7642 6390 7644
rect 6446 7642 6452 7644
rect 6206 7590 6208 7642
rect 6388 7590 6390 7642
rect 6144 7588 6150 7590
rect 6206 7588 6230 7590
rect 6286 7588 6310 7590
rect 6366 7588 6390 7590
rect 6446 7588 6452 7590
rect 6144 7568 6452 7588
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 6564 7478 6592 7686
rect 6552 7472 6604 7478
rect 6656 7449 6684 8434
rect 6748 7750 6776 8434
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6840 8090 6868 8230
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6748 7478 6776 7686
rect 6840 7546 6868 7822
rect 7104 7812 7156 7818
rect 7104 7754 7156 7760
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6736 7472 6788 7478
rect 6552 7414 6604 7420
rect 6642 7440 6698 7449
rect 5632 7404 5684 7410
rect 6736 7414 6788 7420
rect 6642 7375 6698 7384
rect 5632 7346 5684 7352
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 4988 6860 5040 6866
rect 4988 6802 5040 6808
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 5080 6792 5132 6798
rect 5080 6734 5132 6740
rect 5092 6322 5120 6734
rect 5368 6390 5396 6802
rect 5448 6724 5500 6730
rect 5448 6666 5500 6672
rect 5356 6384 5408 6390
rect 5356 6326 5408 6332
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 5080 6316 5132 6322
rect 5080 6258 5132 6264
rect 4252 6248 4304 6254
rect 4252 6190 4304 6196
rect 4344 6248 4396 6254
rect 4344 6190 4396 6196
rect 3884 6180 3936 6186
rect 3884 6122 3936 6128
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 4080 6066 4108 6122
rect 3988 6038 4108 6066
rect 3792 5840 3844 5846
rect 3792 5782 3844 5788
rect 3988 5778 4016 6038
rect 4264 5914 4292 6190
rect 4160 5908 4212 5914
rect 4160 5850 4212 5856
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 4172 5710 4200 5850
rect 4908 5710 4936 6258
rect 3384 5664 3464 5692
rect 3608 5704 3660 5710
rect 3332 5646 3384 5652
rect 3792 5704 3844 5710
rect 3608 5646 3660 5652
rect 3712 5652 3792 5658
rect 3712 5646 3844 5652
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 4896 5704 4948 5710
rect 4896 5646 4948 5652
rect 2596 5636 2648 5642
rect 2596 5578 2648 5584
rect 3712 5630 3832 5646
rect 4068 5636 4120 5642
rect 3712 5166 3740 5630
rect 4068 5578 4120 5584
rect 4080 5370 4108 5578
rect 4908 5370 4936 5646
rect 5368 5574 5396 6326
rect 5460 6322 5488 6666
rect 5644 6662 5672 7346
rect 6656 7342 6684 7375
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 6000 7268 6052 7274
rect 6000 7210 6052 7216
rect 5908 7200 5960 7206
rect 5908 7142 5960 7148
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5644 6458 5672 6598
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 5828 6118 5856 6734
rect 5920 6390 5948 7142
rect 6012 6798 6040 7210
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 6104 6934 6132 7142
rect 6092 6928 6144 6934
rect 6092 6870 6144 6876
rect 6552 6928 6604 6934
rect 6552 6870 6604 6876
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 6144 6556 6452 6576
rect 6144 6554 6150 6556
rect 6206 6554 6230 6556
rect 6286 6554 6310 6556
rect 6366 6554 6390 6556
rect 6446 6554 6452 6556
rect 6206 6502 6208 6554
rect 6388 6502 6390 6554
rect 6144 6500 6150 6502
rect 6206 6500 6230 6502
rect 6286 6500 6310 6502
rect 6366 6500 6390 6502
rect 6446 6500 6452 6502
rect 6144 6480 6452 6500
rect 5908 6384 5960 6390
rect 5908 6326 5960 6332
rect 6564 6254 6592 6870
rect 6840 6662 6868 7482
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 7024 7002 7052 7346
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 7116 6866 7144 7754
rect 7208 7546 7236 8978
rect 7300 8090 7328 9454
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 7852 7886 7880 8026
rect 8128 7886 8156 9318
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8220 8566 8248 8978
rect 8312 8974 8340 9522
rect 9232 9178 9260 9522
rect 9692 9382 9720 9522
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9294 9276 9602 9296
rect 9294 9274 9300 9276
rect 9356 9274 9380 9276
rect 9436 9274 9460 9276
rect 9516 9274 9540 9276
rect 9596 9274 9602 9276
rect 9356 9222 9358 9274
rect 9538 9222 9540 9274
rect 9294 9220 9300 9222
rect 9356 9220 9380 9222
rect 9436 9220 9460 9222
rect 9516 9220 9540 9222
rect 9596 9220 9602 9222
rect 9294 9200 9602 9220
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8404 8634 8432 8978
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 8864 8634 8892 8910
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 8956 8498 8984 8910
rect 9140 8888 9168 9114
rect 9680 9104 9732 9110
rect 9600 9064 9680 9092
rect 9220 8900 9272 8906
rect 9140 8860 9220 8888
rect 9220 8842 9272 8848
rect 9600 8634 9628 9064
rect 9680 9046 9732 9052
rect 9784 9042 9812 9522
rect 9968 9518 9996 11200
rect 12443 9820 12751 9840
rect 12443 9818 12449 9820
rect 12505 9818 12529 9820
rect 12585 9818 12609 9820
rect 12665 9818 12689 9820
rect 12745 9818 12751 9820
rect 12505 9766 12507 9818
rect 12687 9766 12689 9818
rect 12443 9764 12449 9766
rect 12505 9764 12529 9766
rect 12585 9764 12609 9766
rect 12665 9764 12689 9766
rect 12745 9764 12751 9766
rect 12443 9744 12751 9764
rect 10888 9710 11100 9738
rect 10048 9580 10100 9586
rect 10048 9522 10100 9528
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 10060 9110 10088 9522
rect 10888 9518 10916 9710
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10692 9444 10744 9450
rect 10692 9386 10744 9392
rect 10784 9444 10836 9450
rect 10784 9386 10836 9392
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10048 9104 10100 9110
rect 10048 9046 10100 9052
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10416 8900 10468 8906
rect 10416 8842 10468 8848
rect 10048 8832 10100 8838
rect 10048 8774 10100 8780
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8576 8288 8628 8294
rect 8576 8230 8628 8236
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 6656 5914 6684 6598
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 5632 5772 5684 5778
rect 5632 5714 5684 5720
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4896 5364 4948 5370
rect 4896 5306 4948 5312
rect 4344 5296 4396 5302
rect 4344 5238 4396 5244
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 2995 4924 3303 4944
rect 2995 4922 3001 4924
rect 3057 4922 3081 4924
rect 3137 4922 3161 4924
rect 3217 4922 3241 4924
rect 3297 4922 3303 4924
rect 3057 4870 3059 4922
rect 3239 4870 3241 4922
rect 2995 4868 3001 4870
rect 3057 4868 3081 4870
rect 3137 4868 3161 4870
rect 3217 4868 3241 4870
rect 3297 4868 3303 4870
rect 2995 4848 3303 4868
rect 2995 3836 3303 3856
rect 2995 3834 3001 3836
rect 3057 3834 3081 3836
rect 3137 3834 3161 3836
rect 3217 3834 3241 3836
rect 3297 3834 3303 3836
rect 3057 3782 3059 3834
rect 3239 3782 3241 3834
rect 2995 3780 3001 3782
rect 3057 3780 3081 3782
rect 3137 3780 3161 3782
rect 3217 3780 3241 3782
rect 3297 3780 3303 3782
rect 2995 3760 3303 3780
rect 3332 3528 3384 3534
rect 3332 3470 3384 3476
rect 3240 3392 3292 3398
rect 3240 3334 3292 3340
rect 3252 3058 3280 3334
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 2995 2748 3303 2768
rect 2995 2746 3001 2748
rect 3057 2746 3081 2748
rect 3137 2746 3161 2748
rect 3217 2746 3241 2748
rect 3297 2746 3303 2748
rect 3057 2694 3059 2746
rect 3239 2694 3241 2746
rect 2995 2692 3001 2694
rect 3057 2692 3081 2694
rect 3137 2692 3161 2694
rect 3217 2692 3241 2694
rect 3297 2692 3303 2694
rect 2995 2672 3303 2692
rect 3344 1970 3372 3470
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 3620 3058 3648 3334
rect 4356 3126 4384 5238
rect 5644 5234 5672 5714
rect 5816 5568 5868 5574
rect 5816 5510 5868 5516
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5828 5166 5856 5510
rect 6144 5468 6452 5488
rect 6144 5466 6150 5468
rect 6206 5466 6230 5468
rect 6286 5466 6310 5468
rect 6366 5466 6390 5468
rect 6446 5466 6452 5468
rect 6206 5414 6208 5466
rect 6388 5414 6390 5466
rect 6144 5412 6150 5414
rect 6206 5412 6230 5414
rect 6286 5412 6310 5414
rect 6366 5412 6390 5414
rect 6446 5412 6452 5414
rect 6144 5392 6452 5412
rect 6840 5166 6868 6258
rect 7116 5642 7144 6598
rect 7208 6322 7236 7482
rect 7300 7274 7328 7822
rect 7852 7449 7880 7822
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8390 7712 8446 7721
rect 8312 7478 8340 7686
rect 8390 7647 8446 7656
rect 8300 7472 8352 7478
rect 7838 7440 7894 7449
rect 8300 7414 8352 7420
rect 7838 7375 7894 7384
rect 8404 7342 8432 7647
rect 8588 7342 8616 8230
rect 8392 7336 8444 7342
rect 8392 7278 8444 7284
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 7288 7268 7340 7274
rect 7288 7210 7340 7216
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 8220 6866 8248 7142
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7380 6724 7432 6730
rect 7380 6666 7432 6672
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7392 6202 7420 6666
rect 7852 6458 7880 6734
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 8128 6458 8156 6598
rect 7840 6452 7892 6458
rect 7840 6394 7892 6400
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 7208 6186 7420 6202
rect 7196 6180 7420 6186
rect 7248 6174 7420 6180
rect 7196 6122 7248 6128
rect 7208 5778 7236 6122
rect 8128 5778 8156 6258
rect 8404 6118 8432 7278
rect 8588 7002 8616 7278
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 8496 6322 8524 6802
rect 8680 6390 8708 8366
rect 8956 7886 8984 8434
rect 9036 8424 9088 8430
rect 9036 8366 9088 8372
rect 9048 7954 9076 8366
rect 9036 7948 9088 7954
rect 9036 7890 9088 7896
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8772 7478 8800 7686
rect 8760 7472 8812 7478
rect 8760 7414 8812 7420
rect 8956 7410 8984 7822
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 9048 6662 9076 7890
rect 9140 7478 9168 8434
rect 9128 7472 9180 7478
rect 9128 7414 9180 7420
rect 9232 7342 9260 8434
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9294 8188 9602 8208
rect 9294 8186 9300 8188
rect 9356 8186 9380 8188
rect 9436 8186 9460 8188
rect 9516 8186 9540 8188
rect 9596 8186 9602 8188
rect 9356 8134 9358 8186
rect 9538 8134 9540 8186
rect 9294 8132 9300 8134
rect 9356 8132 9380 8134
rect 9436 8132 9460 8134
rect 9516 8132 9540 8134
rect 9596 8132 9602 8134
rect 9294 8112 9602 8132
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9312 7812 9364 7818
rect 9312 7754 9364 7760
rect 9324 7410 9352 7754
rect 9404 7744 9456 7750
rect 9402 7712 9404 7721
rect 9456 7712 9458 7721
rect 9402 7647 9458 7656
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9600 7342 9628 7822
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 9588 7336 9640 7342
rect 9588 7278 9640 7284
rect 9692 7274 9720 8366
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9784 7410 9812 8026
rect 9956 7744 10008 7750
rect 9956 7686 10008 7692
rect 9968 7546 9996 7686
rect 9956 7540 10008 7546
rect 9956 7482 10008 7488
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9956 7404 10008 7410
rect 9956 7346 10008 7352
rect 9680 7268 9732 7274
rect 9680 7210 9732 7216
rect 9294 7100 9602 7120
rect 9294 7098 9300 7100
rect 9356 7098 9380 7100
rect 9436 7098 9460 7100
rect 9516 7098 9540 7100
rect 9596 7098 9602 7100
rect 9356 7046 9358 7098
rect 9538 7046 9540 7098
rect 9294 7044 9300 7046
rect 9356 7044 9380 7046
rect 9436 7044 9460 7046
rect 9516 7044 9540 7046
rect 9596 7044 9602 7046
rect 9294 7024 9602 7044
rect 9784 7002 9812 7346
rect 9772 6996 9824 7002
rect 9772 6938 9824 6944
rect 9220 6724 9272 6730
rect 9220 6666 9272 6672
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 8668 6384 8720 6390
rect 8668 6326 8720 6332
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 7104 5636 7156 5642
rect 7104 5578 7156 5584
rect 7852 5234 7880 5646
rect 7840 5228 7892 5234
rect 7840 5170 7892 5176
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 7668 4826 7696 5102
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 8036 4758 8064 5646
rect 9232 5302 9260 6666
rect 9968 6202 9996 7346
rect 10060 6730 10088 8774
rect 10428 8634 10456 8842
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10428 8498 10456 8570
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 10152 7954 10180 8230
rect 10140 7948 10192 7954
rect 10140 7890 10192 7896
rect 10140 7336 10192 7342
rect 10140 7278 10192 7284
rect 10152 6934 10180 7278
rect 10520 7002 10548 8910
rect 10612 8566 10640 9318
rect 10704 8974 10732 9386
rect 10796 9042 10824 9386
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10980 8634 11008 9522
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 10600 8560 10652 8566
rect 10600 8502 10652 8508
rect 10876 8288 10928 8294
rect 10928 8248 11008 8276
rect 10876 8230 10928 8236
rect 10980 7342 11008 8248
rect 11072 8090 11100 9710
rect 11336 9716 11388 9722
rect 11336 9658 11388 9664
rect 11348 9518 11376 9658
rect 11428 9648 11480 9654
rect 11428 9590 11480 9596
rect 11612 9648 11664 9654
rect 11612 9590 11664 9596
rect 11440 9518 11468 9590
rect 11336 9512 11388 9518
rect 11336 9454 11388 9460
rect 11428 9512 11480 9518
rect 11428 9454 11480 9460
rect 11520 9104 11572 9110
rect 11518 9072 11520 9081
rect 11572 9072 11574 9081
rect 11152 9036 11204 9042
rect 11518 9007 11574 9016
rect 11152 8978 11204 8984
rect 11164 8498 11192 8978
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 11256 8498 11284 8910
rect 11520 8900 11572 8906
rect 11624 8888 11652 9590
rect 12820 9466 12848 11200
rect 13084 9648 13136 9654
rect 13084 9590 13136 9596
rect 14280 9648 14332 9654
rect 14280 9590 14332 9596
rect 12820 9450 12940 9466
rect 12820 9444 12952 9450
rect 12820 9438 12900 9444
rect 12900 9386 12952 9392
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11572 8860 11652 8888
rect 11520 8842 11572 8848
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 11164 7970 11192 8434
rect 11624 8362 11652 8860
rect 11612 8356 11664 8362
rect 11072 7942 11192 7970
rect 11532 8316 11612 8344
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10140 6928 10192 6934
rect 10140 6870 10192 6876
rect 10152 6798 10180 6870
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10048 6724 10100 6730
rect 10048 6666 10100 6672
rect 10230 6488 10286 6497
rect 10230 6423 10232 6432
rect 10284 6423 10286 6432
rect 10232 6394 10284 6400
rect 10244 6322 10272 6394
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 9968 6174 10548 6202
rect 9294 6012 9602 6032
rect 9294 6010 9300 6012
rect 9356 6010 9380 6012
rect 9436 6010 9460 6012
rect 9516 6010 9540 6012
rect 9596 6010 9602 6012
rect 9356 5958 9358 6010
rect 9538 5958 9540 6010
rect 9294 5956 9300 5958
rect 9356 5956 9380 5958
rect 9436 5956 9460 5958
rect 9516 5956 9540 5958
rect 9596 5956 9602 5958
rect 9294 5936 9602 5956
rect 9968 5710 9996 6174
rect 10520 6118 10548 6174
rect 10140 6112 10192 6118
rect 10140 6054 10192 6060
rect 10416 6112 10468 6118
rect 10416 6054 10468 6060
rect 10508 6112 10560 6118
rect 10508 6054 10560 6060
rect 10152 5710 10180 6054
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 9968 5302 9996 5510
rect 10428 5302 10456 6054
rect 10520 5794 10548 6054
rect 10796 5914 10824 6258
rect 10968 6248 11020 6254
rect 10968 6190 11020 6196
rect 10784 5908 10836 5914
rect 10784 5850 10836 5856
rect 10520 5766 10640 5794
rect 10508 5636 10560 5642
rect 10508 5578 10560 5584
rect 9220 5296 9272 5302
rect 9220 5238 9272 5244
rect 9956 5296 10008 5302
rect 9956 5238 10008 5244
rect 10416 5296 10468 5302
rect 10416 5238 10468 5244
rect 7380 4752 7432 4758
rect 7380 4694 7432 4700
rect 8024 4752 8076 4758
rect 8024 4694 8076 4700
rect 9036 4752 9088 4758
rect 9036 4694 9088 4700
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 4344 3120 4396 3126
rect 4344 3062 4396 3068
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 3608 2304 3660 2310
rect 3608 2246 3660 2252
rect 3620 2038 3648 2246
rect 4908 2038 4936 2994
rect 5080 2508 5132 2514
rect 5080 2450 5132 2456
rect 5092 2106 5120 2450
rect 5276 2106 5304 3606
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 5368 2922 5396 3470
rect 5552 3466 5580 4558
rect 6000 4548 6052 4554
rect 6000 4490 6052 4496
rect 6012 4282 6040 4490
rect 6144 4380 6452 4400
rect 6144 4378 6150 4380
rect 6206 4378 6230 4380
rect 6286 4378 6310 4380
rect 6366 4378 6390 4380
rect 6446 4378 6452 4380
rect 6206 4326 6208 4378
rect 6388 4326 6390 4378
rect 6144 4324 6150 4326
rect 6206 4324 6230 4326
rect 6286 4324 6310 4326
rect 6366 4324 6390 4326
rect 6446 4324 6452 4326
rect 6144 4304 6452 4324
rect 7392 4282 7420 4694
rect 8576 4684 8628 4690
rect 8496 4644 8576 4672
rect 8300 4616 8352 4622
rect 8496 4604 8524 4644
rect 8576 4626 8628 4632
rect 8352 4576 8524 4604
rect 8300 4558 8352 4564
rect 7564 4548 7616 4554
rect 7564 4490 7616 4496
rect 8208 4548 8260 4554
rect 8208 4490 8260 4496
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 7380 4276 7432 4282
rect 7380 4218 7432 4224
rect 7576 4078 7604 4490
rect 8220 4078 8248 4490
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 5908 3732 5960 3738
rect 5908 3674 5960 3680
rect 5540 3460 5592 3466
rect 5540 3402 5592 3408
rect 5816 3460 5868 3466
rect 5816 3402 5868 3408
rect 5356 2916 5408 2922
rect 5356 2858 5408 2864
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5080 2100 5132 2106
rect 5080 2042 5132 2048
rect 5264 2100 5316 2106
rect 5264 2042 5316 2048
rect 5460 2038 5488 2382
rect 3608 2032 3660 2038
rect 3608 1974 3660 1980
rect 4896 2032 4948 2038
rect 4896 1974 4948 1980
rect 5448 2032 5500 2038
rect 5448 1974 5500 1980
rect 3332 1964 3384 1970
rect 3332 1906 3384 1912
rect 2995 1660 3303 1680
rect 2995 1658 3001 1660
rect 3057 1658 3081 1660
rect 3137 1658 3161 1660
rect 3217 1658 3241 1660
rect 3297 1658 3303 1660
rect 3057 1606 3059 1658
rect 3239 1606 3241 1658
rect 2995 1604 3001 1606
rect 3057 1604 3081 1606
rect 3137 1604 3161 1606
rect 3217 1604 3241 1606
rect 3297 1604 3303 1606
rect 2995 1584 3303 1604
rect 4908 1465 4936 1974
rect 4894 1456 4950 1465
rect 4894 1391 4950 1400
rect 5552 1222 5580 3402
rect 5828 3194 5856 3402
rect 5920 3194 5948 3674
rect 8220 3534 8248 3878
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8312 3398 8340 4422
rect 8496 4146 8524 4576
rect 8944 4480 8996 4486
rect 8944 4422 8996 4428
rect 8956 4298 8984 4422
rect 8864 4270 8984 4298
rect 8864 4214 8892 4270
rect 9048 4214 9076 4694
rect 9232 4622 9260 5238
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 9294 4924 9602 4944
rect 9294 4922 9300 4924
rect 9356 4922 9380 4924
rect 9436 4922 9460 4924
rect 9516 4922 9540 4924
rect 9596 4922 9602 4924
rect 9356 4870 9358 4922
rect 9538 4870 9540 4922
rect 9294 4868 9300 4870
rect 9356 4868 9380 4870
rect 9436 4868 9460 4870
rect 9516 4868 9540 4870
rect 9596 4868 9602 4870
rect 9294 4848 9602 4868
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 8852 4208 8904 4214
rect 8852 4150 8904 4156
rect 9036 4208 9088 4214
rect 9036 4150 9088 4156
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 8496 3738 8524 4082
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8956 3602 8984 3878
rect 8944 3596 8996 3602
rect 8944 3538 8996 3544
rect 8576 3460 8628 3466
rect 8576 3402 8628 3408
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 6144 3292 6452 3312
rect 6144 3290 6150 3292
rect 6206 3290 6230 3292
rect 6286 3290 6310 3292
rect 6366 3290 6390 3292
rect 6446 3290 6452 3292
rect 6206 3238 6208 3290
rect 6388 3238 6390 3290
rect 6144 3236 6150 3238
rect 6206 3236 6230 3238
rect 6286 3236 6310 3238
rect 6366 3236 6390 3238
rect 6446 3236 6452 3238
rect 6144 3216 6452 3236
rect 7024 3194 7052 3334
rect 8312 3194 8340 3334
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5908 3188 5960 3194
rect 7012 3188 7064 3194
rect 5960 3148 6040 3176
rect 5908 3130 5960 3136
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 5644 2514 5672 2994
rect 5920 2854 5948 2994
rect 5908 2848 5960 2854
rect 5908 2790 5960 2796
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 5736 2106 5764 2382
rect 5724 2100 5776 2106
rect 5724 2042 5776 2048
rect 5920 1970 5948 2790
rect 6012 2650 6040 3148
rect 7012 3130 7064 3136
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 7024 3058 7052 3130
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 8116 3052 8168 3058
rect 8116 2994 8168 3000
rect 6368 2984 6420 2990
rect 6368 2926 6420 2932
rect 6380 2802 6408 2926
rect 6472 2922 6500 2994
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 6460 2916 6512 2922
rect 6460 2858 6512 2864
rect 6564 2802 6592 2926
rect 6380 2774 6592 2802
rect 7932 2848 7984 2854
rect 7932 2790 7984 2796
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 6552 2576 6604 2582
rect 6552 2518 6604 2524
rect 6000 2440 6052 2446
rect 6000 2382 6052 2388
rect 5816 1964 5868 1970
rect 5816 1906 5868 1912
rect 5908 1964 5960 1970
rect 5908 1906 5960 1912
rect 5828 1850 5856 1906
rect 6012 1850 6040 2382
rect 6144 2204 6452 2224
rect 6144 2202 6150 2204
rect 6206 2202 6230 2204
rect 6286 2202 6310 2204
rect 6366 2202 6390 2204
rect 6446 2202 6452 2204
rect 6206 2150 6208 2202
rect 6388 2150 6390 2202
rect 6144 2148 6150 2150
rect 6206 2148 6230 2150
rect 6286 2148 6310 2150
rect 6366 2148 6390 2150
rect 6446 2148 6452 2150
rect 6144 2128 6452 2148
rect 6564 1970 6592 2518
rect 7944 2514 7972 2790
rect 8024 2576 8076 2582
rect 8024 2518 8076 2524
rect 7932 2508 7984 2514
rect 7932 2450 7984 2456
rect 6828 2440 6880 2446
rect 6828 2382 6880 2388
rect 6552 1964 6604 1970
rect 6552 1906 6604 1912
rect 6840 1902 6868 2382
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 7564 1964 7616 1970
rect 7564 1906 7616 1912
rect 5828 1822 6040 1850
rect 6828 1896 6880 1902
rect 6828 1838 6880 1844
rect 6644 1760 6696 1766
rect 6644 1702 6696 1708
rect 5540 1216 5592 1222
rect 5540 1158 5592 1164
rect 6552 1216 6604 1222
rect 6552 1158 6604 1164
rect 6144 1116 6452 1136
rect 6144 1114 6150 1116
rect 6206 1114 6230 1116
rect 6286 1114 6310 1116
rect 6366 1114 6390 1116
rect 6446 1114 6452 1116
rect 6206 1062 6208 1114
rect 6388 1062 6390 1114
rect 6144 1060 6150 1062
rect 6206 1060 6230 1062
rect 6286 1060 6310 1062
rect 6366 1060 6390 1062
rect 6446 1060 6452 1062
rect 6144 1040 6452 1060
rect 6564 882 6592 1158
rect 6656 950 6684 1702
rect 6920 1420 6972 1426
rect 6920 1362 6972 1368
rect 6932 1306 6960 1362
rect 7576 1358 7604 1906
rect 7760 1358 7788 2246
rect 7944 2038 7972 2450
rect 8036 2106 8064 2518
rect 8024 2100 8076 2106
rect 8024 2042 8076 2048
rect 7932 2032 7984 2038
rect 8128 2009 8156 2994
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 8208 2304 8260 2310
rect 8208 2246 8260 2252
rect 7932 1974 7984 1980
rect 8114 2000 8170 2009
rect 8114 1935 8116 1944
rect 8168 1935 8170 1944
rect 8116 1906 8168 1912
rect 8128 1875 8156 1906
rect 8022 1864 8078 1873
rect 8022 1799 8078 1808
rect 8036 1426 8064 1799
rect 8220 1748 8248 2246
rect 8404 1970 8432 2314
rect 8484 2304 8536 2310
rect 8484 2246 8536 2252
rect 8392 1964 8444 1970
rect 8392 1906 8444 1912
rect 8496 1834 8524 2246
rect 8484 1828 8536 1834
rect 8484 1770 8536 1776
rect 8300 1760 8352 1766
rect 8220 1720 8300 1748
rect 8300 1702 8352 1708
rect 8312 1465 8340 1702
rect 8496 1494 8524 1770
rect 8484 1488 8536 1494
rect 8298 1456 8354 1465
rect 8024 1420 8076 1426
rect 8484 1430 8536 1436
rect 8298 1391 8354 1400
rect 8024 1362 8076 1368
rect 6840 1278 6960 1306
rect 7564 1352 7616 1358
rect 7564 1294 7616 1300
rect 7748 1352 7800 1358
rect 7748 1294 7800 1300
rect 7012 1284 7064 1290
rect 6840 1018 6868 1278
rect 7012 1226 7064 1232
rect 7024 1193 7052 1226
rect 7472 1216 7524 1222
rect 7010 1184 7066 1193
rect 7472 1158 7524 1164
rect 7010 1119 7066 1128
rect 7484 1018 7512 1158
rect 6828 1012 6880 1018
rect 6828 954 6880 960
rect 7472 1012 7524 1018
rect 7472 954 7524 960
rect 6644 944 6696 950
rect 6644 886 6696 892
rect 7194 912 7250 921
rect 6552 876 6604 882
rect 7194 847 7196 856
rect 6552 818 6604 824
rect 7248 847 7250 856
rect 7196 818 7248 824
rect 6564 785 6592 818
rect 6550 776 6606 785
rect 6550 711 6606 720
rect 2995 572 3303 592
rect 2995 570 3001 572
rect 3057 570 3081 572
rect 3137 570 3161 572
rect 3217 570 3241 572
rect 3297 570 3303 572
rect 3057 518 3059 570
rect 3239 518 3241 570
rect 2995 516 3001 518
rect 3057 516 3081 518
rect 3137 516 3161 518
rect 3217 516 3241 518
rect 3297 516 3303 518
rect 2995 496 3303 516
rect 7484 270 7512 954
rect 7576 474 7604 1294
rect 7760 678 7788 1294
rect 8036 746 8064 1362
rect 8588 1193 8616 3402
rect 8852 3392 8904 3398
rect 8852 3334 8904 3340
rect 8864 3058 8892 3334
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 8668 2984 8720 2990
rect 8668 2926 8720 2932
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 8680 2514 8708 2926
rect 8668 2508 8720 2514
rect 8668 2450 8720 2456
rect 8956 2106 8984 2926
rect 9140 2774 9168 4422
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9232 3194 9260 4014
rect 9294 3836 9602 3856
rect 9294 3834 9300 3836
rect 9356 3834 9380 3836
rect 9436 3834 9460 3836
rect 9516 3834 9540 3836
rect 9596 3834 9602 3836
rect 9356 3782 9358 3834
rect 9538 3782 9540 3834
rect 9294 3780 9300 3782
rect 9356 3780 9380 3782
rect 9436 3780 9460 3782
rect 9516 3780 9540 3782
rect 9596 3780 9602 3782
rect 9294 3760 9602 3780
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9048 2746 9168 2774
rect 9048 2394 9076 2746
rect 9232 2514 9260 3130
rect 9692 2854 9720 4082
rect 9784 3534 9812 5102
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 9968 4078 9996 4626
rect 10520 4604 10548 5578
rect 10612 5234 10640 5766
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 10796 5030 10824 5850
rect 10980 5370 11008 6190
rect 11072 5710 11100 7942
rect 11532 6662 11560 8316
rect 11612 8298 11664 8304
rect 11704 8288 11756 8294
rect 11704 8230 11756 8236
rect 11716 7886 11744 8230
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11808 7818 11836 9318
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 12808 9104 12860 9110
rect 12452 9052 12808 9058
rect 12452 9046 12860 9052
rect 12452 9030 12848 9046
rect 12452 8906 12480 9030
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 12440 8900 12492 8906
rect 12440 8842 12492 8848
rect 12443 8732 12751 8752
rect 12443 8730 12449 8732
rect 12505 8730 12529 8732
rect 12585 8730 12609 8732
rect 12665 8730 12689 8732
rect 12745 8730 12751 8732
rect 12505 8678 12507 8730
rect 12687 8678 12689 8730
rect 12443 8676 12449 8678
rect 12505 8676 12529 8678
rect 12585 8676 12609 8678
rect 12665 8676 12689 8678
rect 12745 8676 12751 8678
rect 12443 8656 12751 8676
rect 12440 8560 12492 8566
rect 12440 8502 12492 8508
rect 12716 8560 12768 8566
rect 12716 8502 12768 8508
rect 11980 8356 12032 8362
rect 11980 8298 12032 8304
rect 11992 7954 12020 8298
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 12176 7886 12204 8230
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 11796 7812 11848 7818
rect 11796 7754 11848 7760
rect 12452 7732 12480 8502
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12544 8090 12572 8434
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12728 7954 12756 8502
rect 12820 7954 12848 8910
rect 12900 8900 12952 8906
rect 12900 8842 12952 8848
rect 12716 7948 12768 7954
rect 12716 7890 12768 7896
rect 12808 7948 12860 7954
rect 12808 7890 12860 7896
rect 12360 7704 12480 7732
rect 12728 7732 12756 7890
rect 12728 7704 12848 7732
rect 12360 7528 12388 7704
rect 12443 7644 12751 7664
rect 12443 7642 12449 7644
rect 12505 7642 12529 7644
rect 12585 7642 12609 7644
rect 12665 7642 12689 7644
rect 12745 7642 12751 7644
rect 12505 7590 12507 7642
rect 12687 7590 12689 7642
rect 12443 7588 12449 7590
rect 12505 7588 12529 7590
rect 12585 7588 12609 7590
rect 12665 7588 12689 7590
rect 12745 7588 12751 7590
rect 12443 7568 12751 7588
rect 12360 7500 12480 7528
rect 12346 7440 12402 7449
rect 12346 7375 12402 7384
rect 11888 7336 11940 7342
rect 11888 7278 11940 7284
rect 11610 6896 11666 6905
rect 11610 6831 11612 6840
rect 11664 6831 11666 6840
rect 11612 6802 11664 6808
rect 11900 6798 11928 7278
rect 12360 7002 12388 7375
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12452 6866 12480 7500
rect 12716 7472 12768 7478
rect 12530 7440 12586 7449
rect 12820 7460 12848 7704
rect 12768 7432 12848 7460
rect 12716 7414 12768 7420
rect 12530 7375 12586 7384
rect 12544 7206 12572 7375
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12622 6896 12678 6905
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 12440 6860 12492 6866
rect 12622 6831 12678 6840
rect 12440 6802 12492 6808
rect 11888 6792 11940 6798
rect 11888 6734 11940 6740
rect 11612 6724 11664 6730
rect 11612 6666 11664 6672
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11520 6656 11572 6662
rect 11520 6598 11572 6604
rect 11256 6322 11284 6598
rect 11624 6458 11652 6666
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11808 6497 11836 6598
rect 11794 6488 11850 6497
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11704 6452 11756 6458
rect 11900 6458 11928 6734
rect 11794 6423 11850 6432
rect 11888 6452 11940 6458
rect 11704 6394 11756 6400
rect 11610 6352 11666 6361
rect 11244 6316 11296 6322
rect 11610 6287 11666 6296
rect 11244 6258 11296 6264
rect 11624 6254 11652 6287
rect 11612 6248 11664 6254
rect 11612 6190 11664 6196
rect 11716 5778 11744 6394
rect 11808 6304 11836 6423
rect 11888 6394 11940 6400
rect 11888 6316 11940 6322
rect 11808 6276 11888 6304
rect 11888 6258 11940 6264
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 11072 5234 11100 5646
rect 11336 5636 11388 5642
rect 11336 5578 11388 5584
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 10520 4576 10732 4604
rect 10704 4282 10732 4576
rect 10692 4276 10744 4282
rect 10692 4218 10744 4224
rect 10600 4208 10652 4214
rect 10600 4150 10652 4156
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 10428 3194 10456 4082
rect 10612 3738 10640 4150
rect 10704 4136 10732 4218
rect 10888 4214 10916 4626
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 11060 4140 11112 4146
rect 10692 4130 10744 4136
rect 11060 4082 11112 4088
rect 10692 4072 10744 4078
rect 11072 3738 11100 4082
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10048 2916 10100 2922
rect 10048 2858 10100 2864
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 9294 2748 9602 2768
rect 9294 2746 9300 2748
rect 9356 2746 9380 2748
rect 9436 2746 9460 2748
rect 9516 2746 9540 2748
rect 9596 2746 9602 2748
rect 9356 2694 9358 2746
rect 9538 2694 9540 2746
rect 9294 2692 9300 2694
rect 9356 2692 9380 2694
rect 9436 2692 9460 2694
rect 9516 2692 9540 2694
rect 9596 2692 9602 2694
rect 9294 2672 9602 2692
rect 9692 2650 9720 2790
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 10060 2446 10088 2858
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 9312 2440 9364 2446
rect 9048 2388 9312 2394
rect 9048 2382 9364 2388
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 10048 2440 10100 2446
rect 10048 2382 10100 2388
rect 9048 2366 9352 2382
rect 8944 2100 8996 2106
rect 8944 2042 8996 2048
rect 8668 1964 8720 1970
rect 8668 1906 8720 1912
rect 8680 1766 8708 1906
rect 8668 1760 8720 1766
rect 8668 1702 8720 1708
rect 9048 1358 9076 2366
rect 9128 2304 9180 2310
rect 9128 2246 9180 2252
rect 9496 2304 9548 2310
rect 9496 2246 9548 2252
rect 9140 2038 9168 2246
rect 9508 2106 9536 2246
rect 9496 2100 9548 2106
rect 9496 2042 9548 2048
rect 9128 2032 9180 2038
rect 9128 1974 9180 1980
rect 9312 1964 9364 1970
rect 9312 1906 9364 1912
rect 9496 1964 9548 1970
rect 9496 1906 9548 1912
rect 9324 1850 9352 1906
rect 9508 1873 9536 1906
rect 9140 1822 9352 1850
rect 9494 1864 9550 1873
rect 8760 1352 8812 1358
rect 8760 1294 8812 1300
rect 9036 1352 9088 1358
rect 9036 1294 9088 1300
rect 8206 1184 8262 1193
rect 8206 1119 8262 1128
rect 8574 1184 8630 1193
rect 8574 1119 8630 1128
rect 8220 950 8248 1119
rect 8772 1057 8800 1294
rect 9140 1222 9168 1822
rect 9494 1799 9550 1808
rect 9220 1760 9272 1766
rect 9600 1748 9628 2382
rect 9864 2304 9916 2310
rect 9864 2246 9916 2252
rect 9876 2038 9904 2246
rect 9864 2032 9916 2038
rect 9864 1974 9916 1980
rect 9954 2000 10010 2009
rect 9772 1964 9824 1970
rect 9954 1935 9956 1944
rect 9772 1906 9824 1912
rect 10008 1935 10010 1944
rect 9956 1906 10008 1912
rect 9600 1720 9720 1748
rect 9220 1702 9272 1708
rect 8944 1216 8996 1222
rect 8944 1158 8996 1164
rect 9128 1216 9180 1222
rect 9128 1158 9180 1164
rect 8758 1048 8814 1057
rect 8758 983 8760 992
rect 8812 983 8814 992
rect 8760 954 8812 960
rect 8208 944 8260 950
rect 8772 923 8800 954
rect 8956 950 8984 1158
rect 8852 944 8904 950
rect 8208 886 8260 892
rect 8852 886 8904 892
rect 8944 944 8996 950
rect 8944 886 8996 892
rect 8024 740 8076 746
rect 8024 682 8076 688
rect 7748 672 7800 678
rect 7748 614 7800 620
rect 7564 468 7616 474
rect 7564 410 7616 416
rect 7472 264 7524 270
rect 7472 206 7524 212
rect 8220 202 8248 886
rect 8390 776 8446 785
rect 8390 711 8446 720
rect 8404 338 8432 711
rect 8864 377 8892 886
rect 9232 814 9260 1702
rect 9294 1660 9602 1680
rect 9294 1658 9300 1660
rect 9356 1658 9380 1660
rect 9436 1658 9460 1660
rect 9516 1658 9540 1660
rect 9596 1658 9602 1660
rect 9356 1606 9358 1658
rect 9538 1606 9540 1658
rect 9294 1604 9300 1606
rect 9356 1604 9380 1606
rect 9436 1604 9460 1606
rect 9516 1604 9540 1606
rect 9596 1604 9602 1606
rect 9294 1584 9602 1604
rect 9692 1442 9720 1720
rect 9600 1414 9720 1442
rect 9600 1018 9628 1414
rect 9784 1222 9812 1906
rect 10060 1834 10088 2382
rect 10980 1970 11008 2790
rect 10968 1964 11020 1970
rect 10968 1906 11020 1912
rect 10508 1896 10560 1902
rect 10508 1838 10560 1844
rect 10048 1828 10100 1834
rect 10048 1770 10100 1776
rect 9864 1760 9916 1766
rect 9864 1702 9916 1708
rect 9772 1216 9824 1222
rect 9772 1158 9824 1164
rect 9588 1012 9640 1018
rect 9588 954 9640 960
rect 9680 944 9732 950
rect 9678 912 9680 921
rect 9732 912 9734 921
rect 9678 847 9734 856
rect 9876 814 9904 1702
rect 10416 1488 10468 1494
rect 10520 1442 10548 1838
rect 10468 1436 10548 1442
rect 10416 1430 10548 1436
rect 10428 1414 10548 1430
rect 10980 1426 11008 1906
rect 11348 1873 11376 5578
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11520 5160 11572 5166
rect 11520 5102 11572 5108
rect 11532 4826 11560 5102
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11520 4208 11572 4214
rect 11520 4150 11572 4156
rect 11532 3194 11560 4150
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 11532 2038 11560 3130
rect 11808 2378 11836 5306
rect 11900 4729 11928 6258
rect 11992 6118 12020 6802
rect 12164 6792 12216 6798
rect 12164 6734 12216 6740
rect 12072 6656 12124 6662
rect 12072 6598 12124 6604
rect 12084 6390 12112 6598
rect 12072 6384 12124 6390
rect 12072 6326 12124 6332
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 12176 5574 12204 6734
rect 12636 6730 12664 6831
rect 12624 6724 12676 6730
rect 12624 6666 12676 6672
rect 12820 6662 12848 7432
rect 12912 6882 12940 8842
rect 13004 8090 13032 9114
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 13096 7750 13124 9590
rect 13176 9376 13228 9382
rect 13176 9318 13228 9324
rect 13084 7744 13136 7750
rect 13084 7686 13136 7692
rect 12912 6866 13032 6882
rect 13188 6866 13216 9318
rect 14002 9072 14058 9081
rect 13268 9036 13320 9042
rect 14002 9007 14058 9016
rect 13268 8978 13320 8984
rect 13280 8430 13308 8978
rect 13728 8900 13780 8906
rect 13728 8842 13780 8848
rect 13740 8566 13768 8842
rect 13728 8560 13780 8566
rect 13728 8502 13780 8508
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 13280 8022 13308 8230
rect 13268 8016 13320 8022
rect 13268 7958 13320 7964
rect 13372 7886 13400 8434
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13372 7002 13400 7822
rect 13360 6996 13412 7002
rect 13360 6938 13412 6944
rect 12912 6860 13044 6866
rect 12912 6854 12992 6860
rect 12992 6802 13044 6808
rect 13176 6860 13228 6866
rect 13176 6802 13228 6808
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12268 6361 12296 6598
rect 12443 6556 12751 6576
rect 12443 6554 12449 6556
rect 12505 6554 12529 6556
rect 12585 6554 12609 6556
rect 12665 6554 12689 6556
rect 12745 6554 12751 6556
rect 12505 6502 12507 6554
rect 12687 6502 12689 6554
rect 12443 6500 12449 6502
rect 12505 6500 12529 6502
rect 12585 6500 12609 6502
rect 12665 6500 12689 6502
rect 12745 6500 12751 6502
rect 12443 6480 12751 6500
rect 12254 6352 12310 6361
rect 12254 6287 12310 6296
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 12348 5704 12400 5710
rect 12348 5646 12400 5652
rect 12164 5568 12216 5574
rect 12164 5510 12216 5516
rect 12176 5250 12204 5510
rect 12360 5370 12388 5646
rect 12443 5468 12751 5488
rect 12443 5466 12449 5468
rect 12505 5466 12529 5468
rect 12585 5466 12609 5468
rect 12665 5466 12689 5468
rect 12745 5466 12751 5468
rect 12505 5414 12507 5466
rect 12687 5414 12689 5466
rect 12443 5412 12449 5414
rect 12505 5412 12529 5414
rect 12585 5412 12609 5414
rect 12665 5412 12689 5414
rect 12745 5412 12751 5414
rect 12443 5392 12751 5412
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12176 5222 12480 5250
rect 12452 5166 12480 5222
rect 12348 5160 12400 5166
rect 12348 5102 12400 5108
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11886 4720 11942 4729
rect 11886 4655 11942 4664
rect 11992 4622 12020 4966
rect 12360 4826 12388 5102
rect 12820 4826 12848 6190
rect 12912 6118 12940 6734
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 13004 5914 13032 6802
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 13096 6390 13124 6598
rect 13084 6384 13136 6390
rect 13084 6326 13136 6332
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 13096 5710 13124 6326
rect 13360 6316 13412 6322
rect 13360 6258 13412 6264
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13280 5710 13308 5850
rect 13084 5704 13136 5710
rect 13084 5646 13136 5652
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12532 4820 12584 4826
rect 12532 4762 12584 4768
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 12360 4162 12388 4762
rect 12544 4554 12572 4762
rect 13096 4690 13124 5510
rect 13372 5234 13400 6258
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 13464 5370 13492 5646
rect 13452 5364 13504 5370
rect 13452 5306 13504 5312
rect 13556 5234 13584 8366
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 13832 7886 13860 8298
rect 14016 7886 14044 9007
rect 14188 8560 14240 8566
rect 14292 8548 14320 9590
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14476 9042 14504 9318
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 14464 9036 14516 9042
rect 14464 8978 14516 8984
rect 14476 8634 14504 8978
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14240 8520 14320 8548
rect 14188 8502 14240 8508
rect 14188 8356 14240 8362
rect 14188 8298 14240 8304
rect 14200 8090 14228 8298
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 13740 7478 13768 7822
rect 14292 7750 14320 8520
rect 14752 8362 14780 8774
rect 14740 8356 14792 8362
rect 14740 8298 14792 8304
rect 14648 7880 14700 7886
rect 14646 7848 14648 7857
rect 14700 7848 14702 7857
rect 14646 7783 14702 7792
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 14280 7744 14332 7750
rect 14280 7686 14332 7692
rect 13728 7472 13780 7478
rect 13728 7414 13780 7420
rect 13832 7342 13860 7686
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 14004 7336 14056 7342
rect 14004 7278 14056 7284
rect 14016 6769 14044 7278
rect 14108 7002 14136 7346
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 14002 6760 14058 6769
rect 14002 6695 14058 6704
rect 13636 6248 13688 6254
rect 13636 6190 13688 6196
rect 13648 5574 13676 6190
rect 13728 6180 13780 6186
rect 13728 6122 13780 6128
rect 13740 5710 13768 6122
rect 13912 5772 13964 5778
rect 14016 5760 14044 6695
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14108 6236 14136 6598
rect 14200 6390 14228 7482
rect 14280 7268 14332 7274
rect 14280 7210 14332 7216
rect 14292 6798 14320 7210
rect 14936 7206 14964 8910
rect 15304 8566 15332 9114
rect 15200 8560 15252 8566
rect 15200 8502 15252 8508
rect 15292 8560 15344 8566
rect 15292 8502 15344 8508
rect 15212 7478 15240 8502
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 15200 7472 15252 7478
rect 15200 7414 15252 7420
rect 14924 7200 14976 7206
rect 14924 7142 14976 7148
rect 15108 6996 15160 7002
rect 15108 6938 15160 6944
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14372 6656 14424 6662
rect 14372 6598 14424 6604
rect 14384 6390 14412 6598
rect 14188 6384 14240 6390
rect 14188 6326 14240 6332
rect 14372 6384 14424 6390
rect 14372 6326 14424 6332
rect 14108 6208 14228 6236
rect 14200 6118 14228 6208
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 13964 5732 14044 5760
rect 13912 5714 13964 5720
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13544 5228 13596 5234
rect 13544 5170 13596 5176
rect 13360 5092 13412 5098
rect 13360 5034 13412 5040
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 13372 4622 13400 5034
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 12532 4548 12584 4554
rect 12532 4490 12584 4496
rect 12992 4480 13044 4486
rect 12992 4422 13044 4428
rect 12443 4380 12751 4400
rect 12443 4378 12449 4380
rect 12505 4378 12529 4380
rect 12585 4378 12609 4380
rect 12665 4378 12689 4380
rect 12745 4378 12751 4380
rect 12505 4326 12507 4378
rect 12687 4326 12689 4378
rect 12443 4324 12449 4326
rect 12505 4324 12529 4326
rect 12585 4324 12609 4326
rect 12665 4324 12689 4326
rect 12745 4324 12751 4326
rect 12443 4304 12751 4324
rect 13004 4214 13032 4422
rect 12992 4208 13044 4214
rect 12360 4146 12480 4162
rect 12992 4150 13044 4156
rect 13452 4208 13504 4214
rect 13452 4150 13504 4156
rect 12360 4140 12492 4146
rect 12360 4134 12440 4140
rect 12440 4082 12492 4088
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 12820 4026 12848 4082
rect 12820 3998 13032 4026
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12532 3596 12584 3602
rect 12532 3538 12584 3544
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 12544 3482 12572 3538
rect 12912 3534 12940 3878
rect 13004 3738 13032 3998
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 12900 3528 12952 3534
rect 11900 2650 11928 3470
rect 12544 3454 12848 3482
rect 12900 3470 12952 3476
rect 12443 3292 12751 3312
rect 12443 3290 12449 3292
rect 12505 3290 12529 3292
rect 12585 3290 12609 3292
rect 12665 3290 12689 3292
rect 12745 3290 12751 3292
rect 12505 3238 12507 3290
rect 12687 3238 12689 3290
rect 12443 3236 12449 3238
rect 12505 3236 12529 3238
rect 12585 3236 12609 3238
rect 12665 3236 12689 3238
rect 12745 3236 12751 3238
rect 12443 3216 12751 3236
rect 12820 3194 12848 3454
rect 12808 3188 12860 3194
rect 12808 3130 12860 3136
rect 12820 3074 12848 3130
rect 12072 3052 12124 3058
rect 12820 3046 12940 3074
rect 13096 3058 13124 4082
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 12072 2994 12124 3000
rect 12084 2650 12112 2994
rect 12808 2984 12860 2990
rect 12808 2926 12860 2932
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 12072 2644 12124 2650
rect 12072 2586 12124 2592
rect 11796 2372 11848 2378
rect 11796 2314 11848 2320
rect 11520 2032 11572 2038
rect 11520 1974 11572 1980
rect 11334 1864 11390 1873
rect 11334 1799 11390 1808
rect 10520 1018 10548 1414
rect 10692 1420 10744 1426
rect 10692 1362 10744 1368
rect 10968 1420 11020 1426
rect 10968 1362 11020 1368
rect 10704 1306 10732 1362
rect 10612 1278 10732 1306
rect 10612 1222 10640 1278
rect 10600 1216 10652 1222
rect 10600 1158 10652 1164
rect 11060 1216 11112 1222
rect 11060 1158 11112 1164
rect 10690 1048 10746 1057
rect 10508 1012 10560 1018
rect 11072 1018 11100 1158
rect 10690 983 10746 992
rect 11060 1012 11112 1018
rect 10508 954 10560 960
rect 10704 882 10732 983
rect 11060 954 11112 960
rect 11808 950 11836 2314
rect 11900 1902 11928 2586
rect 12443 2204 12751 2224
rect 12443 2202 12449 2204
rect 12505 2202 12529 2204
rect 12585 2202 12609 2204
rect 12665 2202 12689 2204
rect 12745 2202 12751 2204
rect 12505 2150 12507 2202
rect 12687 2150 12689 2202
rect 12443 2148 12449 2150
rect 12505 2148 12529 2150
rect 12585 2148 12609 2150
rect 12665 2148 12689 2150
rect 12745 2148 12751 2150
rect 12443 2128 12751 2148
rect 12072 2032 12124 2038
rect 12072 1974 12124 1980
rect 11888 1896 11940 1902
rect 11888 1838 11940 1844
rect 11900 1358 11928 1838
rect 11888 1352 11940 1358
rect 11888 1294 11940 1300
rect 11888 1216 11940 1222
rect 11888 1158 11940 1164
rect 11152 944 11204 950
rect 11152 886 11204 892
rect 11796 944 11848 950
rect 11796 886 11848 892
rect 10140 876 10192 882
rect 10140 818 10192 824
rect 10692 876 10744 882
rect 10692 818 10744 824
rect 9220 808 9272 814
rect 9220 750 9272 756
rect 9864 808 9916 814
rect 9864 750 9916 756
rect 9036 672 9088 678
rect 9036 614 9088 620
rect 8850 368 8906 377
rect 8392 332 8444 338
rect 9048 338 9076 614
rect 9294 572 9602 592
rect 9294 570 9300 572
rect 9356 570 9380 572
rect 9436 570 9460 572
rect 9516 570 9540 572
rect 9596 570 9602 572
rect 9356 518 9358 570
rect 9538 518 9540 570
rect 9294 516 9300 518
rect 9356 516 9380 518
rect 9436 516 9460 518
rect 9516 516 9540 518
rect 9596 516 9602 518
rect 9294 496 9602 516
rect 10152 338 10180 818
rect 11060 808 11112 814
rect 11060 750 11112 756
rect 11072 377 11100 750
rect 11058 368 11114 377
rect 8850 303 8906 312
rect 9036 332 9088 338
rect 8392 274 8444 280
rect 9036 274 9088 280
rect 10140 332 10192 338
rect 11058 303 11114 312
rect 10140 274 10192 280
rect 11072 270 11100 303
rect 11164 270 11192 886
rect 11900 474 11928 1158
rect 12084 1018 12112 1974
rect 12820 1970 12848 2926
rect 12912 2378 12940 3046
rect 13084 3052 13136 3058
rect 13084 2994 13136 3000
rect 13084 2916 13136 2922
rect 13084 2858 13136 2864
rect 13096 2446 13124 2858
rect 13280 2854 13308 3674
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13372 3126 13400 3470
rect 13464 3466 13492 4150
rect 13556 3670 13584 5170
rect 13728 4616 13780 4622
rect 13832 4604 13860 5306
rect 14200 4622 14228 6054
rect 14280 5908 14332 5914
rect 14280 5850 14332 5856
rect 14292 4826 14320 5850
rect 14384 5778 14412 6326
rect 14372 5772 14424 5778
rect 14372 5714 14424 5720
rect 14372 5636 14424 5642
rect 14372 5578 14424 5584
rect 14384 5302 14412 5578
rect 14372 5296 14424 5302
rect 14372 5238 14424 5244
rect 14476 5114 14504 6802
rect 14740 6792 14792 6798
rect 14738 6760 14740 6769
rect 14924 6792 14976 6798
rect 14792 6760 14794 6769
rect 14648 6724 14700 6730
rect 14738 6695 14794 6704
rect 14922 6760 14924 6769
rect 14976 6760 14978 6769
rect 14922 6695 14978 6704
rect 14648 6666 14700 6672
rect 14660 5914 14688 6666
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 14752 5370 14780 6598
rect 14936 6254 14964 6695
rect 15120 6458 15148 6938
rect 15304 6730 15332 7686
rect 15292 6724 15344 6730
rect 15292 6666 15344 6672
rect 15016 6452 15068 6458
rect 15016 6394 15068 6400
rect 15108 6452 15160 6458
rect 15108 6394 15160 6400
rect 14924 6248 14976 6254
rect 14924 6190 14976 6196
rect 15028 6118 15056 6394
rect 15016 6112 15068 6118
rect 15016 6054 15068 6060
rect 14740 5364 14792 5370
rect 14740 5306 14792 5312
rect 14476 5086 14596 5114
rect 14568 4826 14596 5086
rect 14280 4820 14332 4826
rect 14280 4762 14332 4768
rect 14464 4820 14516 4826
rect 14464 4762 14516 4768
rect 14556 4820 14608 4826
rect 14556 4762 14608 4768
rect 13780 4576 13860 4604
rect 14188 4616 14240 4622
rect 13728 4558 13780 4564
rect 14188 4558 14240 4564
rect 14004 4480 14056 4486
rect 14004 4422 14056 4428
rect 14016 4078 14044 4422
rect 14476 4282 14504 4762
rect 14922 4720 14978 4729
rect 14922 4655 14978 4664
rect 14936 4622 14964 4655
rect 15120 4622 15148 6394
rect 15292 6248 15344 6254
rect 15292 6190 15344 6196
rect 15304 5846 15332 6190
rect 15292 5840 15344 5846
rect 15292 5782 15344 5788
rect 15396 4758 15424 11206
rect 15580 11098 15608 11206
rect 15658 11200 15714 12000
rect 17866 11248 17922 11257
rect 15672 11098 15700 11200
rect 18510 11200 18566 12000
rect 17866 11183 17922 11192
rect 15580 11070 15700 11098
rect 17774 9752 17830 9761
rect 17774 9687 17830 9696
rect 16856 9648 16908 9654
rect 16856 9590 16908 9596
rect 16488 9512 16540 9518
rect 16488 9454 16540 9460
rect 15476 9376 15528 9382
rect 15476 9318 15528 9324
rect 16028 9376 16080 9382
rect 16028 9318 16080 9324
rect 15488 9042 15516 9318
rect 15592 9276 15900 9296
rect 15592 9274 15598 9276
rect 15654 9274 15678 9276
rect 15734 9274 15758 9276
rect 15814 9274 15838 9276
rect 15894 9274 15900 9276
rect 15654 9222 15656 9274
rect 15836 9222 15838 9274
rect 15592 9220 15598 9222
rect 15654 9220 15678 9222
rect 15734 9220 15758 9222
rect 15814 9220 15838 9222
rect 15894 9220 15900 9222
rect 15592 9200 15900 9220
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 16040 8906 16068 9318
rect 16500 9178 16528 9454
rect 16868 9382 16896 9590
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16488 9172 16540 9178
rect 16488 9114 16540 9120
rect 16028 8900 16080 8906
rect 16028 8842 16080 8848
rect 15936 8356 15988 8362
rect 15936 8298 15988 8304
rect 15592 8188 15900 8208
rect 15592 8186 15598 8188
rect 15654 8186 15678 8188
rect 15734 8186 15758 8188
rect 15814 8186 15838 8188
rect 15894 8186 15900 8188
rect 15654 8134 15656 8186
rect 15836 8134 15838 8186
rect 15592 8132 15598 8134
rect 15654 8132 15678 8134
rect 15734 8132 15758 8134
rect 15814 8132 15838 8134
rect 15894 8132 15900 8134
rect 15592 8112 15900 8132
rect 15592 7100 15900 7120
rect 15592 7098 15598 7100
rect 15654 7098 15678 7100
rect 15734 7098 15758 7100
rect 15814 7098 15838 7100
rect 15894 7098 15900 7100
rect 15654 7046 15656 7098
rect 15836 7046 15838 7098
rect 15592 7044 15598 7046
rect 15654 7044 15678 7046
rect 15734 7044 15758 7046
rect 15814 7044 15838 7046
rect 15894 7044 15900 7046
rect 15592 7024 15900 7044
rect 15476 6316 15528 6322
rect 15476 6258 15528 6264
rect 15488 5914 15516 6258
rect 15948 6254 15976 8298
rect 16040 7886 16068 8842
rect 16868 8566 16896 9318
rect 17788 8974 17816 9687
rect 17880 9042 17908 11183
rect 18328 9580 18380 9586
rect 18328 9522 18380 9528
rect 18340 9178 18368 9522
rect 18328 9172 18380 9178
rect 18328 9114 18380 9120
rect 17868 9036 17920 9042
rect 17868 8978 17920 8984
rect 17776 8968 17828 8974
rect 17776 8910 17828 8916
rect 16856 8560 16908 8566
rect 16856 8502 16908 8508
rect 16488 8424 16540 8430
rect 16488 8366 16540 8372
rect 16856 8424 16908 8430
rect 16856 8366 16908 8372
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 16500 7954 16528 8366
rect 16488 7948 16540 7954
rect 16488 7890 16540 7896
rect 16028 7880 16080 7886
rect 16028 7822 16080 7828
rect 16764 7812 16816 7818
rect 16764 7754 16816 7760
rect 16396 7744 16448 7750
rect 16448 7704 16620 7732
rect 16396 7686 16448 7692
rect 16028 7336 16080 7342
rect 16028 7278 16080 7284
rect 16040 6866 16068 7278
rect 16592 6866 16620 7704
rect 16776 7478 16804 7754
rect 16764 7472 16816 7478
rect 16764 7414 16816 7420
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16684 6798 16712 7278
rect 16672 6792 16724 6798
rect 16592 6740 16672 6746
rect 16592 6734 16724 6740
rect 16592 6718 16712 6734
rect 16304 6656 16356 6662
rect 16304 6598 16356 6604
rect 16316 6390 16344 6598
rect 16304 6384 16356 6390
rect 16304 6326 16356 6332
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 15936 6248 15988 6254
rect 15936 6190 15988 6196
rect 15592 6012 15900 6032
rect 15592 6010 15598 6012
rect 15654 6010 15678 6012
rect 15734 6010 15758 6012
rect 15814 6010 15838 6012
rect 15894 6010 15900 6012
rect 15654 5958 15656 6010
rect 15836 5958 15838 6010
rect 15592 5956 15598 5958
rect 15654 5956 15678 5958
rect 15734 5956 15758 5958
rect 15814 5956 15838 5958
rect 15894 5956 15900 5958
rect 15592 5936 15900 5956
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 16040 5302 16068 6258
rect 16316 5914 16344 6326
rect 16304 5908 16356 5914
rect 16304 5850 16356 5856
rect 16592 5846 16620 6718
rect 16868 6662 16896 8366
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 16960 7206 16988 7890
rect 16948 7200 17000 7206
rect 16948 7142 17000 7148
rect 16960 6866 16988 7142
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17590 6760 17646 6769
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 17420 6458 17448 6598
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 17512 6322 17540 6734
rect 17590 6695 17646 6704
rect 17604 6322 17632 6695
rect 17500 6316 17552 6322
rect 17500 6258 17552 6264
rect 17592 6316 17644 6322
rect 17592 6258 17644 6264
rect 17224 6112 17276 6118
rect 17224 6054 17276 6060
rect 17236 5914 17264 6054
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 17224 5908 17276 5914
rect 17224 5850 17276 5856
rect 16580 5840 16632 5846
rect 16580 5782 16632 5788
rect 16396 5772 16448 5778
rect 16396 5714 16448 5720
rect 16304 5704 16356 5710
rect 16304 5646 16356 5652
rect 16212 5568 16264 5574
rect 16212 5510 16264 5516
rect 16028 5296 16080 5302
rect 16028 5238 16080 5244
rect 15592 4924 15900 4944
rect 15592 4922 15598 4924
rect 15654 4922 15678 4924
rect 15734 4922 15758 4924
rect 15814 4922 15838 4924
rect 15894 4922 15900 4924
rect 15654 4870 15656 4922
rect 15836 4870 15838 4922
rect 15592 4868 15598 4870
rect 15654 4868 15678 4870
rect 15734 4868 15758 4870
rect 15814 4868 15838 4870
rect 15894 4868 15900 4870
rect 15592 4848 15900 4868
rect 15384 4752 15436 4758
rect 15384 4694 15436 4700
rect 16224 4690 16252 5510
rect 16316 5234 16344 5646
rect 16304 5228 16356 5234
rect 16304 5170 16356 5176
rect 16408 5166 16436 5714
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 16396 5160 16448 5166
rect 16396 5102 16448 5108
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 16212 4684 16264 4690
rect 16212 4626 16264 4632
rect 14924 4616 14976 4622
rect 14924 4558 14976 4564
rect 15108 4616 15160 4622
rect 15108 4558 15160 4564
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 15108 4480 15160 4486
rect 15108 4422 15160 4428
rect 14464 4276 14516 4282
rect 14464 4218 14516 4224
rect 14004 4072 14056 4078
rect 14004 4014 14056 4020
rect 13544 3664 13596 3670
rect 13544 3606 13596 3612
rect 13636 3664 13688 3670
rect 13636 3606 13688 3612
rect 13648 3534 13676 3606
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13452 3460 13504 3466
rect 13452 3402 13504 3408
rect 13360 3120 13412 3126
rect 13360 3062 13412 3068
rect 13464 2990 13492 3402
rect 13648 3126 13676 3470
rect 13912 3188 13964 3194
rect 13912 3130 13964 3136
rect 13636 3120 13688 3126
rect 13636 3062 13688 3068
rect 13452 2984 13504 2990
rect 13452 2926 13504 2932
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 13360 2848 13412 2854
rect 13360 2790 13412 2796
rect 13176 2644 13228 2650
rect 13176 2586 13228 2592
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 12900 2372 12952 2378
rect 12900 2314 12952 2320
rect 12808 1964 12860 1970
rect 12808 1906 12860 1912
rect 12820 1766 12848 1906
rect 13084 1896 13136 1902
rect 13188 1884 13216 2586
rect 13372 2582 13400 2790
rect 13464 2774 13492 2926
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 13464 2746 13584 2774
rect 13360 2576 13412 2582
rect 13360 2518 13412 2524
rect 13372 2446 13400 2518
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 13556 1970 13584 2746
rect 13832 2446 13860 2790
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 13820 2304 13872 2310
rect 13924 2258 13952 3130
rect 14016 2514 14044 4014
rect 14476 3534 14504 4218
rect 14936 3890 14964 4422
rect 14936 3862 15056 3890
rect 15028 3534 15056 3862
rect 15120 3738 15148 4422
rect 15212 4214 15240 4626
rect 16684 4622 16712 5646
rect 16960 5302 16988 5850
rect 17512 5710 17540 6258
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 17604 5574 17632 6258
rect 17788 5710 17816 8366
rect 18524 8294 18552 11200
rect 18512 8288 18564 8294
rect 18512 8230 18564 8236
rect 18602 8256 18658 8265
rect 18602 8191 18658 8200
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18234 7848 18290 7857
rect 18234 7783 18290 7792
rect 18248 7750 18276 7783
rect 18144 7744 18196 7750
rect 18144 7686 18196 7692
rect 18236 7744 18288 7750
rect 18236 7686 18288 7692
rect 18156 7478 18184 7686
rect 18144 7472 18196 7478
rect 18144 7414 18196 7420
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 17972 6458 18000 6598
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 18156 5778 18184 6190
rect 18340 5914 18368 8026
rect 18616 7886 18644 8191
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18510 6760 18566 6769
rect 18510 6695 18566 6704
rect 18328 5908 18380 5914
rect 18328 5850 18380 5856
rect 18144 5772 18196 5778
rect 18144 5714 18196 5720
rect 18524 5710 18552 6695
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 18512 5704 18564 5710
rect 18512 5646 18564 5652
rect 17592 5568 17644 5574
rect 17592 5510 17644 5516
rect 17684 5568 17736 5574
rect 17684 5510 17736 5516
rect 17696 5370 17724 5510
rect 17684 5364 17736 5370
rect 17684 5306 17736 5312
rect 16948 5296 17000 5302
rect 16948 5238 17000 5244
rect 16764 5092 16816 5098
rect 16764 5034 16816 5040
rect 16776 4690 16804 5034
rect 16764 4684 16816 4690
rect 16764 4626 16816 4632
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16960 4486 16988 5238
rect 17040 5160 17092 5166
rect 17040 5102 17092 5108
rect 17052 4826 17080 5102
rect 17224 5024 17276 5030
rect 17224 4966 17276 4972
rect 17040 4820 17092 4826
rect 17040 4762 17092 4768
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 16948 4480 17000 4486
rect 16948 4422 17000 4428
rect 15200 4208 15252 4214
rect 15200 4150 15252 4156
rect 15200 3936 15252 3942
rect 15200 3878 15252 3884
rect 15108 3732 15160 3738
rect 15108 3674 15160 3680
rect 15212 3534 15240 3878
rect 15592 3836 15900 3856
rect 15592 3834 15598 3836
rect 15654 3834 15678 3836
rect 15734 3834 15758 3836
rect 15814 3834 15838 3836
rect 15894 3834 15900 3836
rect 15654 3782 15656 3834
rect 15836 3782 15838 3834
rect 15592 3780 15598 3782
rect 15654 3780 15678 3782
rect 15734 3780 15758 3782
rect 15814 3780 15838 3782
rect 15894 3780 15900 3782
rect 15592 3760 15900 3780
rect 15384 3664 15436 3670
rect 15384 3606 15436 3612
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 14556 3392 14608 3398
rect 14556 3334 14608 3340
rect 14924 3392 14976 3398
rect 14924 3334 14976 3340
rect 14568 3058 14596 3334
rect 14832 3188 14884 3194
rect 14832 3130 14884 3136
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14280 2848 14332 2854
rect 14280 2790 14332 2796
rect 14004 2508 14056 2514
rect 14004 2450 14056 2456
rect 13872 2252 13952 2258
rect 13820 2246 13952 2252
rect 13832 2230 13952 2246
rect 13544 1964 13596 1970
rect 13544 1906 13596 1912
rect 13832 1902 13860 2230
rect 13136 1856 13216 1884
rect 13820 1896 13872 1902
rect 13084 1838 13136 1844
rect 13820 1838 13872 1844
rect 12808 1760 12860 1766
rect 12808 1702 12860 1708
rect 13096 1465 13124 1838
rect 13268 1760 13320 1766
rect 13268 1702 13320 1708
rect 13082 1456 13138 1465
rect 13082 1391 13138 1400
rect 12443 1116 12751 1136
rect 12443 1114 12449 1116
rect 12505 1114 12529 1116
rect 12585 1114 12609 1116
rect 12665 1114 12689 1116
rect 12745 1114 12751 1116
rect 12505 1062 12507 1114
rect 12687 1062 12689 1114
rect 12443 1060 12449 1062
rect 12505 1060 12529 1062
rect 12585 1060 12609 1062
rect 12665 1060 12689 1062
rect 12745 1060 12751 1062
rect 12443 1040 12751 1060
rect 12072 1012 12124 1018
rect 12072 954 12124 960
rect 13280 950 13308 1702
rect 13268 944 13320 950
rect 13268 886 13320 892
rect 14016 882 14044 2450
rect 14292 2378 14320 2790
rect 14384 2650 14412 2994
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 14280 2372 14332 2378
rect 14280 2314 14332 2320
rect 14280 1964 14332 1970
rect 14280 1906 14332 1912
rect 14188 1828 14240 1834
rect 14188 1770 14240 1776
rect 14200 1494 14228 1770
rect 14188 1488 14240 1494
rect 14188 1430 14240 1436
rect 14292 1358 14320 1906
rect 14464 1420 14516 1426
rect 14464 1362 14516 1368
rect 14280 1352 14332 1358
rect 14280 1294 14332 1300
rect 14476 1018 14504 1362
rect 14752 1290 14780 2926
rect 14844 2038 14872 3130
rect 14936 3126 14964 3334
rect 14924 3120 14976 3126
rect 14924 3062 14976 3068
rect 15396 3058 15424 3606
rect 15016 3052 15068 3058
rect 15016 2994 15068 3000
rect 15384 3052 15436 3058
rect 15384 2994 15436 3000
rect 15028 2922 15056 2994
rect 15016 2916 15068 2922
rect 15016 2858 15068 2864
rect 14832 2032 14884 2038
rect 14832 1974 14884 1980
rect 14924 1964 14976 1970
rect 14924 1906 14976 1912
rect 14832 1760 14884 1766
rect 14832 1702 14884 1708
rect 14844 1358 14872 1702
rect 14936 1562 14964 1906
rect 15028 1562 15056 2858
rect 15108 2848 15160 2854
rect 15108 2790 15160 2796
rect 15120 2310 15148 2790
rect 15108 2304 15160 2310
rect 15108 2246 15160 2252
rect 15120 1902 15148 2246
rect 15396 1970 15424 2994
rect 16028 2984 16080 2990
rect 16028 2926 16080 2932
rect 16120 2984 16172 2990
rect 16120 2926 16172 2932
rect 15592 2748 15900 2768
rect 15592 2746 15598 2748
rect 15654 2746 15678 2748
rect 15734 2746 15758 2748
rect 15814 2746 15838 2748
rect 15894 2746 15900 2748
rect 15654 2694 15656 2746
rect 15836 2694 15838 2746
rect 15592 2692 15598 2694
rect 15654 2692 15678 2694
rect 15734 2692 15758 2694
rect 15814 2692 15838 2694
rect 15894 2692 15900 2694
rect 15592 2672 15900 2692
rect 15566 2408 15622 2417
rect 15566 2343 15568 2352
rect 15620 2343 15622 2352
rect 15568 2314 15620 2320
rect 15384 1964 15436 1970
rect 15384 1906 15436 1912
rect 15108 1896 15160 1902
rect 15108 1838 15160 1844
rect 15384 1828 15436 1834
rect 15384 1770 15436 1776
rect 14924 1556 14976 1562
rect 14924 1498 14976 1504
rect 15016 1556 15068 1562
rect 15016 1498 15068 1504
rect 15396 1358 15424 1770
rect 15476 1760 15528 1766
rect 15476 1702 15528 1708
rect 15936 1760 15988 1766
rect 15936 1702 15988 1708
rect 15488 1426 15516 1702
rect 15592 1660 15900 1680
rect 15592 1658 15598 1660
rect 15654 1658 15678 1660
rect 15734 1658 15758 1660
rect 15814 1658 15838 1660
rect 15894 1658 15900 1660
rect 15654 1606 15656 1658
rect 15836 1606 15838 1658
rect 15592 1604 15598 1606
rect 15654 1604 15678 1606
rect 15734 1604 15758 1606
rect 15814 1604 15838 1606
rect 15894 1604 15900 1606
rect 15592 1584 15900 1604
rect 15948 1426 15976 1702
rect 15476 1420 15528 1426
rect 15476 1362 15528 1368
rect 15936 1420 15988 1426
rect 15936 1362 15988 1368
rect 14832 1352 14884 1358
rect 14832 1294 14884 1300
rect 15384 1352 15436 1358
rect 15384 1294 15436 1300
rect 14740 1284 14792 1290
rect 14740 1226 14792 1232
rect 14464 1012 14516 1018
rect 14464 954 14516 960
rect 14752 882 14780 1226
rect 15396 882 15424 1294
rect 16040 1290 16068 2926
rect 16132 2650 16160 2926
rect 16120 2644 16172 2650
rect 16120 2586 16172 2592
rect 16132 1426 16160 2586
rect 16316 1834 16344 4422
rect 16960 4282 16988 4422
rect 16948 4276 17000 4282
rect 16948 4218 17000 4224
rect 16960 3466 16988 4218
rect 17236 4078 17264 4966
rect 17788 4729 17816 5646
rect 17868 5636 17920 5642
rect 17868 5578 17920 5584
rect 17880 5370 17908 5578
rect 17868 5364 17920 5370
rect 17868 5306 17920 5312
rect 18510 5264 18566 5273
rect 18510 5199 18566 5208
rect 17774 4720 17830 4729
rect 17774 4655 17830 4664
rect 18524 4622 18552 5199
rect 17592 4616 17644 4622
rect 17592 4558 17644 4564
rect 17960 4616 18012 4622
rect 17960 4558 18012 4564
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 16948 3460 17000 3466
rect 16948 3402 17000 3408
rect 16580 3392 16632 3398
rect 16580 3334 16632 3340
rect 16396 2984 16448 2990
rect 16396 2926 16448 2932
rect 16408 2514 16436 2926
rect 16396 2508 16448 2514
rect 16396 2450 16448 2456
rect 16488 2372 16540 2378
rect 16488 2314 16540 2320
rect 16500 1884 16528 2314
rect 16592 2106 16620 3334
rect 16960 3126 16988 3402
rect 17604 3194 17632 4558
rect 17972 4078 18000 4558
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 17972 3602 18000 4014
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 17960 3596 18012 3602
rect 17960 3538 18012 3544
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 16948 3120 17000 3126
rect 16948 3062 17000 3068
rect 16960 2417 16988 3062
rect 17972 3058 18000 3538
rect 18064 3466 18092 3878
rect 18524 3777 18552 4082
rect 18510 3768 18566 3777
rect 18510 3703 18566 3712
rect 18052 3460 18104 3466
rect 18052 3402 18104 3408
rect 17960 3052 18012 3058
rect 17960 2994 18012 3000
rect 17868 2576 17920 2582
rect 17868 2518 17920 2524
rect 16946 2408 17002 2417
rect 16946 2343 16948 2352
rect 17000 2343 17002 2352
rect 17684 2372 17736 2378
rect 16948 2314 17000 2320
rect 17684 2314 17736 2320
rect 16960 2106 16988 2314
rect 16580 2100 16632 2106
rect 16948 2100 17000 2106
rect 16580 2042 16632 2048
rect 16868 2060 16948 2088
rect 16580 1896 16632 1902
rect 16500 1856 16580 1884
rect 16580 1838 16632 1844
rect 16304 1828 16356 1834
rect 16304 1770 16356 1776
rect 16592 1426 16620 1838
rect 16120 1420 16172 1426
rect 16120 1362 16172 1368
rect 16580 1420 16632 1426
rect 16580 1362 16632 1368
rect 16028 1284 16080 1290
rect 16028 1226 16080 1232
rect 15936 1216 15988 1222
rect 15936 1158 15988 1164
rect 16764 1216 16816 1222
rect 16764 1158 16816 1164
rect 15948 882 15976 1158
rect 16776 1018 16804 1158
rect 16764 1012 16816 1018
rect 16764 954 16816 960
rect 16868 950 16896 2060
rect 16948 2042 17000 2048
rect 16948 1964 17000 1970
rect 16948 1906 17000 1912
rect 16960 1562 16988 1906
rect 17040 1828 17092 1834
rect 17040 1770 17092 1776
rect 16948 1556 17000 1562
rect 16948 1498 17000 1504
rect 17052 1426 17080 1770
rect 17040 1420 17092 1426
rect 17040 1362 17092 1368
rect 17408 1216 17460 1222
rect 17408 1158 17460 1164
rect 16856 944 16908 950
rect 16856 886 16908 892
rect 14004 876 14056 882
rect 14004 818 14056 824
rect 14740 876 14792 882
rect 14740 818 14792 824
rect 15384 876 15436 882
rect 15384 818 15436 824
rect 15936 876 15988 882
rect 15936 818 15988 824
rect 11888 468 11940 474
rect 11888 410 11940 416
rect 14752 338 14780 818
rect 17132 672 17184 678
rect 17132 614 17184 620
rect 15592 572 15900 592
rect 15592 570 15598 572
rect 15654 570 15678 572
rect 15734 570 15758 572
rect 15814 570 15838 572
rect 15894 570 15900 572
rect 15654 518 15656 570
rect 15836 518 15838 570
rect 15592 516 15598 518
rect 15654 516 15678 518
rect 15734 516 15758 518
rect 15814 516 15838 518
rect 15894 516 15900 518
rect 15592 496 15900 516
rect 14740 332 14792 338
rect 14740 274 14792 280
rect 17144 270 17172 614
rect 17420 474 17448 1158
rect 17408 468 17460 474
rect 17408 410 17460 416
rect 17696 338 17724 2314
rect 17776 2304 17828 2310
rect 17776 2246 17828 2252
rect 17788 1426 17816 2246
rect 17776 1420 17828 1426
rect 17776 1362 17828 1368
rect 17788 814 17816 1362
rect 17880 1018 17908 2518
rect 17960 1284 18012 1290
rect 18064 1272 18092 3402
rect 18420 3052 18472 3058
rect 18420 2994 18472 3000
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18328 2848 18380 2854
rect 18328 2790 18380 2796
rect 18340 2038 18368 2790
rect 18432 2774 18460 2994
rect 18432 2746 18552 2774
rect 18328 2032 18380 2038
rect 18328 1974 18380 1980
rect 18524 1970 18552 2746
rect 18616 2281 18644 2994
rect 18602 2272 18658 2281
rect 18602 2207 18658 2216
rect 18512 1964 18564 1970
rect 18512 1906 18564 1912
rect 18418 1864 18474 1873
rect 18418 1799 18474 1808
rect 18012 1244 18092 1272
rect 17960 1226 18012 1232
rect 17972 1018 18000 1226
rect 18432 1018 18460 1799
rect 17868 1012 17920 1018
rect 17868 954 17920 960
rect 17960 1012 18012 1018
rect 17960 954 18012 960
rect 18420 1012 18472 1018
rect 18420 954 18472 960
rect 18328 876 18380 882
rect 18328 818 18380 824
rect 17776 808 17828 814
rect 17776 750 17828 756
rect 18340 474 18368 818
rect 18510 776 18566 785
rect 18510 711 18566 720
rect 18328 468 18380 474
rect 18328 410 18380 416
rect 17684 332 17736 338
rect 17684 274 17736 280
rect 18524 270 18552 711
rect 11060 264 11112 270
rect 11060 206 11112 212
rect 11152 264 11204 270
rect 11152 206 11204 212
rect 17132 264 17184 270
rect 17132 206 17184 212
rect 18512 264 18564 270
rect 18512 206 18564 212
rect 8208 196 8260 202
rect 8208 138 8260 144
rect 6144 28 6452 48
rect 6144 26 6150 28
rect 6206 26 6230 28
rect 6286 26 6310 28
rect 6366 26 6390 28
rect 6446 26 6452 28
rect 6206 -26 6208 26
rect 6388 -26 6390 26
rect 6144 -28 6150 -26
rect 6206 -28 6230 -26
rect 6286 -28 6310 -26
rect 6366 -28 6390 -26
rect 6446 -28 6452 -26
rect 6144 -48 6452 -28
rect 12443 28 12751 48
rect 12443 26 12449 28
rect 12505 26 12529 28
rect 12585 26 12609 28
rect 12665 26 12689 28
rect 12745 26 12751 28
rect 12505 -26 12507 26
rect 12687 -26 12689 26
rect 12443 -28 12449 -26
rect 12505 -28 12529 -26
rect 12585 -28 12609 -26
rect 12665 -28 12689 -26
rect 12745 -28 12751 -26
rect 12443 -48 12751 -28
<< via2 >>
rect 3001 9274 3057 9276
rect 3081 9274 3137 9276
rect 3161 9274 3217 9276
rect 3241 9274 3297 9276
rect 3001 9222 3047 9274
rect 3047 9222 3057 9274
rect 3081 9222 3111 9274
rect 3111 9222 3123 9274
rect 3123 9222 3137 9274
rect 3161 9222 3175 9274
rect 3175 9222 3187 9274
rect 3187 9222 3217 9274
rect 3241 9222 3251 9274
rect 3251 9222 3297 9274
rect 3001 9220 3057 9222
rect 3081 9220 3137 9222
rect 3161 9220 3217 9222
rect 3241 9220 3297 9222
rect 3001 8186 3057 8188
rect 3081 8186 3137 8188
rect 3161 8186 3217 8188
rect 3241 8186 3297 8188
rect 3001 8134 3047 8186
rect 3047 8134 3057 8186
rect 3081 8134 3111 8186
rect 3111 8134 3123 8186
rect 3123 8134 3137 8186
rect 3161 8134 3175 8186
rect 3175 8134 3187 8186
rect 3187 8134 3217 8186
rect 3241 8134 3251 8186
rect 3251 8134 3297 8186
rect 3001 8132 3057 8134
rect 3081 8132 3137 8134
rect 3161 8132 3217 8134
rect 3241 8132 3297 8134
rect 6150 9818 6206 9820
rect 6230 9818 6286 9820
rect 6310 9818 6366 9820
rect 6390 9818 6446 9820
rect 6150 9766 6196 9818
rect 6196 9766 6206 9818
rect 6230 9766 6260 9818
rect 6260 9766 6272 9818
rect 6272 9766 6286 9818
rect 6310 9766 6324 9818
rect 6324 9766 6336 9818
rect 6336 9766 6366 9818
rect 6390 9766 6400 9818
rect 6400 9766 6446 9818
rect 6150 9764 6206 9766
rect 6230 9764 6286 9766
rect 6310 9764 6366 9766
rect 6390 9764 6446 9766
rect 6150 8730 6206 8732
rect 6230 8730 6286 8732
rect 6310 8730 6366 8732
rect 6390 8730 6446 8732
rect 6150 8678 6196 8730
rect 6196 8678 6206 8730
rect 6230 8678 6260 8730
rect 6260 8678 6272 8730
rect 6272 8678 6286 8730
rect 6310 8678 6324 8730
rect 6324 8678 6336 8730
rect 6336 8678 6366 8730
rect 6390 8678 6400 8730
rect 6400 8678 6446 8730
rect 6150 8676 6206 8678
rect 6230 8676 6286 8678
rect 6310 8676 6366 8678
rect 6390 8676 6446 8678
rect 5630 7792 5686 7848
rect 3001 7098 3057 7100
rect 3081 7098 3137 7100
rect 3161 7098 3217 7100
rect 3241 7098 3297 7100
rect 3001 7046 3047 7098
rect 3047 7046 3057 7098
rect 3081 7046 3111 7098
rect 3111 7046 3123 7098
rect 3123 7046 3137 7098
rect 3161 7046 3175 7098
rect 3175 7046 3187 7098
rect 3187 7046 3217 7098
rect 3241 7046 3251 7098
rect 3251 7046 3297 7098
rect 3001 7044 3057 7046
rect 3081 7044 3137 7046
rect 3161 7044 3217 7046
rect 3241 7044 3297 7046
rect 3001 6010 3057 6012
rect 3081 6010 3137 6012
rect 3161 6010 3217 6012
rect 3241 6010 3297 6012
rect 3001 5958 3047 6010
rect 3047 5958 3057 6010
rect 3081 5958 3111 6010
rect 3111 5958 3123 6010
rect 3123 5958 3137 6010
rect 3161 5958 3175 6010
rect 3175 5958 3187 6010
rect 3187 5958 3217 6010
rect 3241 5958 3251 6010
rect 3251 5958 3297 6010
rect 3001 5956 3057 5958
rect 3081 5956 3137 5958
rect 3161 5956 3217 5958
rect 3241 5956 3297 5958
rect 6366 7792 6422 7848
rect 6150 7642 6206 7644
rect 6230 7642 6286 7644
rect 6310 7642 6366 7644
rect 6390 7642 6446 7644
rect 6150 7590 6196 7642
rect 6196 7590 6206 7642
rect 6230 7590 6260 7642
rect 6260 7590 6272 7642
rect 6272 7590 6286 7642
rect 6310 7590 6324 7642
rect 6324 7590 6336 7642
rect 6336 7590 6366 7642
rect 6390 7590 6400 7642
rect 6400 7590 6446 7642
rect 6150 7588 6206 7590
rect 6230 7588 6286 7590
rect 6310 7588 6366 7590
rect 6390 7588 6446 7590
rect 6642 7384 6698 7440
rect 6150 6554 6206 6556
rect 6230 6554 6286 6556
rect 6310 6554 6366 6556
rect 6390 6554 6446 6556
rect 6150 6502 6196 6554
rect 6196 6502 6206 6554
rect 6230 6502 6260 6554
rect 6260 6502 6272 6554
rect 6272 6502 6286 6554
rect 6310 6502 6324 6554
rect 6324 6502 6336 6554
rect 6336 6502 6366 6554
rect 6390 6502 6400 6554
rect 6400 6502 6446 6554
rect 6150 6500 6206 6502
rect 6230 6500 6286 6502
rect 6310 6500 6366 6502
rect 6390 6500 6446 6502
rect 9300 9274 9356 9276
rect 9380 9274 9436 9276
rect 9460 9274 9516 9276
rect 9540 9274 9596 9276
rect 9300 9222 9346 9274
rect 9346 9222 9356 9274
rect 9380 9222 9410 9274
rect 9410 9222 9422 9274
rect 9422 9222 9436 9274
rect 9460 9222 9474 9274
rect 9474 9222 9486 9274
rect 9486 9222 9516 9274
rect 9540 9222 9550 9274
rect 9550 9222 9596 9274
rect 9300 9220 9356 9222
rect 9380 9220 9436 9222
rect 9460 9220 9516 9222
rect 9540 9220 9596 9222
rect 12449 9818 12505 9820
rect 12529 9818 12585 9820
rect 12609 9818 12665 9820
rect 12689 9818 12745 9820
rect 12449 9766 12495 9818
rect 12495 9766 12505 9818
rect 12529 9766 12559 9818
rect 12559 9766 12571 9818
rect 12571 9766 12585 9818
rect 12609 9766 12623 9818
rect 12623 9766 12635 9818
rect 12635 9766 12665 9818
rect 12689 9766 12699 9818
rect 12699 9766 12745 9818
rect 12449 9764 12505 9766
rect 12529 9764 12585 9766
rect 12609 9764 12665 9766
rect 12689 9764 12745 9766
rect 3001 4922 3057 4924
rect 3081 4922 3137 4924
rect 3161 4922 3217 4924
rect 3241 4922 3297 4924
rect 3001 4870 3047 4922
rect 3047 4870 3057 4922
rect 3081 4870 3111 4922
rect 3111 4870 3123 4922
rect 3123 4870 3137 4922
rect 3161 4870 3175 4922
rect 3175 4870 3187 4922
rect 3187 4870 3217 4922
rect 3241 4870 3251 4922
rect 3251 4870 3297 4922
rect 3001 4868 3057 4870
rect 3081 4868 3137 4870
rect 3161 4868 3217 4870
rect 3241 4868 3297 4870
rect 3001 3834 3057 3836
rect 3081 3834 3137 3836
rect 3161 3834 3217 3836
rect 3241 3834 3297 3836
rect 3001 3782 3047 3834
rect 3047 3782 3057 3834
rect 3081 3782 3111 3834
rect 3111 3782 3123 3834
rect 3123 3782 3137 3834
rect 3161 3782 3175 3834
rect 3175 3782 3187 3834
rect 3187 3782 3217 3834
rect 3241 3782 3251 3834
rect 3251 3782 3297 3834
rect 3001 3780 3057 3782
rect 3081 3780 3137 3782
rect 3161 3780 3217 3782
rect 3241 3780 3297 3782
rect 3001 2746 3057 2748
rect 3081 2746 3137 2748
rect 3161 2746 3217 2748
rect 3241 2746 3297 2748
rect 3001 2694 3047 2746
rect 3047 2694 3057 2746
rect 3081 2694 3111 2746
rect 3111 2694 3123 2746
rect 3123 2694 3137 2746
rect 3161 2694 3175 2746
rect 3175 2694 3187 2746
rect 3187 2694 3217 2746
rect 3241 2694 3251 2746
rect 3251 2694 3297 2746
rect 3001 2692 3057 2694
rect 3081 2692 3137 2694
rect 3161 2692 3217 2694
rect 3241 2692 3297 2694
rect 6150 5466 6206 5468
rect 6230 5466 6286 5468
rect 6310 5466 6366 5468
rect 6390 5466 6446 5468
rect 6150 5414 6196 5466
rect 6196 5414 6206 5466
rect 6230 5414 6260 5466
rect 6260 5414 6272 5466
rect 6272 5414 6286 5466
rect 6310 5414 6324 5466
rect 6324 5414 6336 5466
rect 6336 5414 6366 5466
rect 6390 5414 6400 5466
rect 6400 5414 6446 5466
rect 6150 5412 6206 5414
rect 6230 5412 6286 5414
rect 6310 5412 6366 5414
rect 6390 5412 6446 5414
rect 8390 7656 8446 7712
rect 7838 7384 7894 7440
rect 9300 8186 9356 8188
rect 9380 8186 9436 8188
rect 9460 8186 9516 8188
rect 9540 8186 9596 8188
rect 9300 8134 9346 8186
rect 9346 8134 9356 8186
rect 9380 8134 9410 8186
rect 9410 8134 9422 8186
rect 9422 8134 9436 8186
rect 9460 8134 9474 8186
rect 9474 8134 9486 8186
rect 9486 8134 9516 8186
rect 9540 8134 9550 8186
rect 9550 8134 9596 8186
rect 9300 8132 9356 8134
rect 9380 8132 9436 8134
rect 9460 8132 9516 8134
rect 9540 8132 9596 8134
rect 9402 7692 9404 7712
rect 9404 7692 9456 7712
rect 9456 7692 9458 7712
rect 9402 7656 9458 7692
rect 9300 7098 9356 7100
rect 9380 7098 9436 7100
rect 9460 7098 9516 7100
rect 9540 7098 9596 7100
rect 9300 7046 9346 7098
rect 9346 7046 9356 7098
rect 9380 7046 9410 7098
rect 9410 7046 9422 7098
rect 9422 7046 9436 7098
rect 9460 7046 9474 7098
rect 9474 7046 9486 7098
rect 9486 7046 9516 7098
rect 9540 7046 9550 7098
rect 9550 7046 9596 7098
rect 9300 7044 9356 7046
rect 9380 7044 9436 7046
rect 9460 7044 9516 7046
rect 9540 7044 9596 7046
rect 11518 9052 11520 9072
rect 11520 9052 11572 9072
rect 11572 9052 11574 9072
rect 11518 9016 11574 9052
rect 10230 6452 10286 6488
rect 10230 6432 10232 6452
rect 10232 6432 10284 6452
rect 10284 6432 10286 6452
rect 9300 6010 9356 6012
rect 9380 6010 9436 6012
rect 9460 6010 9516 6012
rect 9540 6010 9596 6012
rect 9300 5958 9346 6010
rect 9346 5958 9356 6010
rect 9380 5958 9410 6010
rect 9410 5958 9422 6010
rect 9422 5958 9436 6010
rect 9460 5958 9474 6010
rect 9474 5958 9486 6010
rect 9486 5958 9516 6010
rect 9540 5958 9550 6010
rect 9550 5958 9596 6010
rect 9300 5956 9356 5958
rect 9380 5956 9436 5958
rect 9460 5956 9516 5958
rect 9540 5956 9596 5958
rect 6150 4378 6206 4380
rect 6230 4378 6286 4380
rect 6310 4378 6366 4380
rect 6390 4378 6446 4380
rect 6150 4326 6196 4378
rect 6196 4326 6206 4378
rect 6230 4326 6260 4378
rect 6260 4326 6272 4378
rect 6272 4326 6286 4378
rect 6310 4326 6324 4378
rect 6324 4326 6336 4378
rect 6336 4326 6366 4378
rect 6390 4326 6400 4378
rect 6400 4326 6446 4378
rect 6150 4324 6206 4326
rect 6230 4324 6286 4326
rect 6310 4324 6366 4326
rect 6390 4324 6446 4326
rect 3001 1658 3057 1660
rect 3081 1658 3137 1660
rect 3161 1658 3217 1660
rect 3241 1658 3297 1660
rect 3001 1606 3047 1658
rect 3047 1606 3057 1658
rect 3081 1606 3111 1658
rect 3111 1606 3123 1658
rect 3123 1606 3137 1658
rect 3161 1606 3175 1658
rect 3175 1606 3187 1658
rect 3187 1606 3217 1658
rect 3241 1606 3251 1658
rect 3251 1606 3297 1658
rect 3001 1604 3057 1606
rect 3081 1604 3137 1606
rect 3161 1604 3217 1606
rect 3241 1604 3297 1606
rect 4894 1400 4950 1456
rect 9300 4922 9356 4924
rect 9380 4922 9436 4924
rect 9460 4922 9516 4924
rect 9540 4922 9596 4924
rect 9300 4870 9346 4922
rect 9346 4870 9356 4922
rect 9380 4870 9410 4922
rect 9410 4870 9422 4922
rect 9422 4870 9436 4922
rect 9460 4870 9474 4922
rect 9474 4870 9486 4922
rect 9486 4870 9516 4922
rect 9540 4870 9550 4922
rect 9550 4870 9596 4922
rect 9300 4868 9356 4870
rect 9380 4868 9436 4870
rect 9460 4868 9516 4870
rect 9540 4868 9596 4870
rect 6150 3290 6206 3292
rect 6230 3290 6286 3292
rect 6310 3290 6366 3292
rect 6390 3290 6446 3292
rect 6150 3238 6196 3290
rect 6196 3238 6206 3290
rect 6230 3238 6260 3290
rect 6260 3238 6272 3290
rect 6272 3238 6286 3290
rect 6310 3238 6324 3290
rect 6324 3238 6336 3290
rect 6336 3238 6366 3290
rect 6390 3238 6400 3290
rect 6400 3238 6446 3290
rect 6150 3236 6206 3238
rect 6230 3236 6286 3238
rect 6310 3236 6366 3238
rect 6390 3236 6446 3238
rect 6150 2202 6206 2204
rect 6230 2202 6286 2204
rect 6310 2202 6366 2204
rect 6390 2202 6446 2204
rect 6150 2150 6196 2202
rect 6196 2150 6206 2202
rect 6230 2150 6260 2202
rect 6260 2150 6272 2202
rect 6272 2150 6286 2202
rect 6310 2150 6324 2202
rect 6324 2150 6336 2202
rect 6336 2150 6366 2202
rect 6390 2150 6400 2202
rect 6400 2150 6446 2202
rect 6150 2148 6206 2150
rect 6230 2148 6286 2150
rect 6310 2148 6366 2150
rect 6390 2148 6446 2150
rect 6150 1114 6206 1116
rect 6230 1114 6286 1116
rect 6310 1114 6366 1116
rect 6390 1114 6446 1116
rect 6150 1062 6196 1114
rect 6196 1062 6206 1114
rect 6230 1062 6260 1114
rect 6260 1062 6272 1114
rect 6272 1062 6286 1114
rect 6310 1062 6324 1114
rect 6324 1062 6336 1114
rect 6336 1062 6366 1114
rect 6390 1062 6400 1114
rect 6400 1062 6446 1114
rect 6150 1060 6206 1062
rect 6230 1060 6286 1062
rect 6310 1060 6366 1062
rect 6390 1060 6446 1062
rect 8114 1964 8170 2000
rect 8114 1944 8116 1964
rect 8116 1944 8168 1964
rect 8168 1944 8170 1964
rect 8022 1808 8078 1864
rect 8298 1400 8354 1456
rect 7010 1128 7066 1184
rect 7194 876 7250 912
rect 7194 856 7196 876
rect 7196 856 7248 876
rect 7248 856 7250 876
rect 6550 720 6606 776
rect 3001 570 3057 572
rect 3081 570 3137 572
rect 3161 570 3217 572
rect 3241 570 3297 572
rect 3001 518 3047 570
rect 3047 518 3057 570
rect 3081 518 3111 570
rect 3111 518 3123 570
rect 3123 518 3137 570
rect 3161 518 3175 570
rect 3175 518 3187 570
rect 3187 518 3217 570
rect 3241 518 3251 570
rect 3251 518 3297 570
rect 3001 516 3057 518
rect 3081 516 3137 518
rect 3161 516 3217 518
rect 3241 516 3297 518
rect 9300 3834 9356 3836
rect 9380 3834 9436 3836
rect 9460 3834 9516 3836
rect 9540 3834 9596 3836
rect 9300 3782 9346 3834
rect 9346 3782 9356 3834
rect 9380 3782 9410 3834
rect 9410 3782 9422 3834
rect 9422 3782 9436 3834
rect 9460 3782 9474 3834
rect 9474 3782 9486 3834
rect 9486 3782 9516 3834
rect 9540 3782 9550 3834
rect 9550 3782 9596 3834
rect 9300 3780 9356 3782
rect 9380 3780 9436 3782
rect 9460 3780 9516 3782
rect 9540 3780 9596 3782
rect 12449 8730 12505 8732
rect 12529 8730 12585 8732
rect 12609 8730 12665 8732
rect 12689 8730 12745 8732
rect 12449 8678 12495 8730
rect 12495 8678 12505 8730
rect 12529 8678 12559 8730
rect 12559 8678 12571 8730
rect 12571 8678 12585 8730
rect 12609 8678 12623 8730
rect 12623 8678 12635 8730
rect 12635 8678 12665 8730
rect 12689 8678 12699 8730
rect 12699 8678 12745 8730
rect 12449 8676 12505 8678
rect 12529 8676 12585 8678
rect 12609 8676 12665 8678
rect 12689 8676 12745 8678
rect 12449 7642 12505 7644
rect 12529 7642 12585 7644
rect 12609 7642 12665 7644
rect 12689 7642 12745 7644
rect 12449 7590 12495 7642
rect 12495 7590 12505 7642
rect 12529 7590 12559 7642
rect 12559 7590 12571 7642
rect 12571 7590 12585 7642
rect 12609 7590 12623 7642
rect 12623 7590 12635 7642
rect 12635 7590 12665 7642
rect 12689 7590 12699 7642
rect 12699 7590 12745 7642
rect 12449 7588 12505 7590
rect 12529 7588 12585 7590
rect 12609 7588 12665 7590
rect 12689 7588 12745 7590
rect 12346 7384 12402 7440
rect 11610 6860 11666 6896
rect 11610 6840 11612 6860
rect 11612 6840 11664 6860
rect 11664 6840 11666 6860
rect 12530 7384 12586 7440
rect 12622 6840 12678 6896
rect 11794 6432 11850 6488
rect 11610 6296 11666 6352
rect 9300 2746 9356 2748
rect 9380 2746 9436 2748
rect 9460 2746 9516 2748
rect 9540 2746 9596 2748
rect 9300 2694 9346 2746
rect 9346 2694 9356 2746
rect 9380 2694 9410 2746
rect 9410 2694 9422 2746
rect 9422 2694 9436 2746
rect 9460 2694 9474 2746
rect 9474 2694 9486 2746
rect 9486 2694 9516 2746
rect 9540 2694 9550 2746
rect 9550 2694 9596 2746
rect 9300 2692 9356 2694
rect 9380 2692 9436 2694
rect 9460 2692 9516 2694
rect 9540 2692 9596 2694
rect 8206 1128 8262 1184
rect 8574 1128 8630 1184
rect 9494 1808 9550 1864
rect 9954 1964 10010 2000
rect 9954 1944 9956 1964
rect 9956 1944 10008 1964
rect 10008 1944 10010 1964
rect 8758 1012 8814 1048
rect 8758 992 8760 1012
rect 8760 992 8812 1012
rect 8812 992 8814 1012
rect 8390 720 8446 776
rect 9300 1658 9356 1660
rect 9380 1658 9436 1660
rect 9460 1658 9516 1660
rect 9540 1658 9596 1660
rect 9300 1606 9346 1658
rect 9346 1606 9356 1658
rect 9380 1606 9410 1658
rect 9410 1606 9422 1658
rect 9422 1606 9436 1658
rect 9460 1606 9474 1658
rect 9474 1606 9486 1658
rect 9486 1606 9516 1658
rect 9540 1606 9550 1658
rect 9550 1606 9596 1658
rect 9300 1604 9356 1606
rect 9380 1604 9436 1606
rect 9460 1604 9516 1606
rect 9540 1604 9596 1606
rect 9678 892 9680 912
rect 9680 892 9732 912
rect 9732 892 9734 912
rect 9678 856 9734 892
rect 14002 9016 14058 9072
rect 12449 6554 12505 6556
rect 12529 6554 12585 6556
rect 12609 6554 12665 6556
rect 12689 6554 12745 6556
rect 12449 6502 12495 6554
rect 12495 6502 12505 6554
rect 12529 6502 12559 6554
rect 12559 6502 12571 6554
rect 12571 6502 12585 6554
rect 12609 6502 12623 6554
rect 12623 6502 12635 6554
rect 12635 6502 12665 6554
rect 12689 6502 12699 6554
rect 12699 6502 12745 6554
rect 12449 6500 12505 6502
rect 12529 6500 12585 6502
rect 12609 6500 12665 6502
rect 12689 6500 12745 6502
rect 12254 6296 12310 6352
rect 12449 5466 12505 5468
rect 12529 5466 12585 5468
rect 12609 5466 12665 5468
rect 12689 5466 12745 5468
rect 12449 5414 12495 5466
rect 12495 5414 12505 5466
rect 12529 5414 12559 5466
rect 12559 5414 12571 5466
rect 12571 5414 12585 5466
rect 12609 5414 12623 5466
rect 12623 5414 12635 5466
rect 12635 5414 12665 5466
rect 12689 5414 12699 5466
rect 12699 5414 12745 5466
rect 12449 5412 12505 5414
rect 12529 5412 12585 5414
rect 12609 5412 12665 5414
rect 12689 5412 12745 5414
rect 11886 4664 11942 4720
rect 14646 7828 14648 7848
rect 14648 7828 14700 7848
rect 14700 7828 14702 7848
rect 14646 7792 14702 7828
rect 14002 6704 14058 6760
rect 12449 4378 12505 4380
rect 12529 4378 12585 4380
rect 12609 4378 12665 4380
rect 12689 4378 12745 4380
rect 12449 4326 12495 4378
rect 12495 4326 12505 4378
rect 12529 4326 12559 4378
rect 12559 4326 12571 4378
rect 12571 4326 12585 4378
rect 12609 4326 12623 4378
rect 12623 4326 12635 4378
rect 12635 4326 12665 4378
rect 12689 4326 12699 4378
rect 12699 4326 12745 4378
rect 12449 4324 12505 4326
rect 12529 4324 12585 4326
rect 12609 4324 12665 4326
rect 12689 4324 12745 4326
rect 12449 3290 12505 3292
rect 12529 3290 12585 3292
rect 12609 3290 12665 3292
rect 12689 3290 12745 3292
rect 12449 3238 12495 3290
rect 12495 3238 12505 3290
rect 12529 3238 12559 3290
rect 12559 3238 12571 3290
rect 12571 3238 12585 3290
rect 12609 3238 12623 3290
rect 12623 3238 12635 3290
rect 12635 3238 12665 3290
rect 12689 3238 12699 3290
rect 12699 3238 12745 3290
rect 12449 3236 12505 3238
rect 12529 3236 12585 3238
rect 12609 3236 12665 3238
rect 12689 3236 12745 3238
rect 11334 1808 11390 1864
rect 10690 992 10746 1048
rect 12449 2202 12505 2204
rect 12529 2202 12585 2204
rect 12609 2202 12665 2204
rect 12689 2202 12745 2204
rect 12449 2150 12495 2202
rect 12495 2150 12505 2202
rect 12529 2150 12559 2202
rect 12559 2150 12571 2202
rect 12571 2150 12585 2202
rect 12609 2150 12623 2202
rect 12623 2150 12635 2202
rect 12635 2150 12665 2202
rect 12689 2150 12699 2202
rect 12699 2150 12745 2202
rect 12449 2148 12505 2150
rect 12529 2148 12585 2150
rect 12609 2148 12665 2150
rect 12689 2148 12745 2150
rect 8850 312 8906 368
rect 9300 570 9356 572
rect 9380 570 9436 572
rect 9460 570 9516 572
rect 9540 570 9596 572
rect 9300 518 9346 570
rect 9346 518 9356 570
rect 9380 518 9410 570
rect 9410 518 9422 570
rect 9422 518 9436 570
rect 9460 518 9474 570
rect 9474 518 9486 570
rect 9486 518 9516 570
rect 9540 518 9550 570
rect 9550 518 9596 570
rect 9300 516 9356 518
rect 9380 516 9436 518
rect 9460 516 9516 518
rect 9540 516 9596 518
rect 11058 312 11114 368
rect 14738 6740 14740 6760
rect 14740 6740 14792 6760
rect 14792 6740 14794 6760
rect 14738 6704 14794 6740
rect 14922 6740 14924 6760
rect 14924 6740 14976 6760
rect 14976 6740 14978 6760
rect 14922 6704 14978 6740
rect 14922 4664 14978 4720
rect 17866 11192 17922 11248
rect 17774 9696 17830 9752
rect 15598 9274 15654 9276
rect 15678 9274 15734 9276
rect 15758 9274 15814 9276
rect 15838 9274 15894 9276
rect 15598 9222 15644 9274
rect 15644 9222 15654 9274
rect 15678 9222 15708 9274
rect 15708 9222 15720 9274
rect 15720 9222 15734 9274
rect 15758 9222 15772 9274
rect 15772 9222 15784 9274
rect 15784 9222 15814 9274
rect 15838 9222 15848 9274
rect 15848 9222 15894 9274
rect 15598 9220 15654 9222
rect 15678 9220 15734 9222
rect 15758 9220 15814 9222
rect 15838 9220 15894 9222
rect 15598 8186 15654 8188
rect 15678 8186 15734 8188
rect 15758 8186 15814 8188
rect 15838 8186 15894 8188
rect 15598 8134 15644 8186
rect 15644 8134 15654 8186
rect 15678 8134 15708 8186
rect 15708 8134 15720 8186
rect 15720 8134 15734 8186
rect 15758 8134 15772 8186
rect 15772 8134 15784 8186
rect 15784 8134 15814 8186
rect 15838 8134 15848 8186
rect 15848 8134 15894 8186
rect 15598 8132 15654 8134
rect 15678 8132 15734 8134
rect 15758 8132 15814 8134
rect 15838 8132 15894 8134
rect 15598 7098 15654 7100
rect 15678 7098 15734 7100
rect 15758 7098 15814 7100
rect 15838 7098 15894 7100
rect 15598 7046 15644 7098
rect 15644 7046 15654 7098
rect 15678 7046 15708 7098
rect 15708 7046 15720 7098
rect 15720 7046 15734 7098
rect 15758 7046 15772 7098
rect 15772 7046 15784 7098
rect 15784 7046 15814 7098
rect 15838 7046 15848 7098
rect 15848 7046 15894 7098
rect 15598 7044 15654 7046
rect 15678 7044 15734 7046
rect 15758 7044 15814 7046
rect 15838 7044 15894 7046
rect 15598 6010 15654 6012
rect 15678 6010 15734 6012
rect 15758 6010 15814 6012
rect 15838 6010 15894 6012
rect 15598 5958 15644 6010
rect 15644 5958 15654 6010
rect 15678 5958 15708 6010
rect 15708 5958 15720 6010
rect 15720 5958 15734 6010
rect 15758 5958 15772 6010
rect 15772 5958 15784 6010
rect 15784 5958 15814 6010
rect 15838 5958 15848 6010
rect 15848 5958 15894 6010
rect 15598 5956 15654 5958
rect 15678 5956 15734 5958
rect 15758 5956 15814 5958
rect 15838 5956 15894 5958
rect 17590 6704 17646 6760
rect 15598 4922 15654 4924
rect 15678 4922 15734 4924
rect 15758 4922 15814 4924
rect 15838 4922 15894 4924
rect 15598 4870 15644 4922
rect 15644 4870 15654 4922
rect 15678 4870 15708 4922
rect 15708 4870 15720 4922
rect 15720 4870 15734 4922
rect 15758 4870 15772 4922
rect 15772 4870 15784 4922
rect 15784 4870 15814 4922
rect 15838 4870 15848 4922
rect 15848 4870 15894 4922
rect 15598 4868 15654 4870
rect 15678 4868 15734 4870
rect 15758 4868 15814 4870
rect 15838 4868 15894 4870
rect 18602 8200 18658 8256
rect 18234 7792 18290 7848
rect 18510 6704 18566 6760
rect 15598 3834 15654 3836
rect 15678 3834 15734 3836
rect 15758 3834 15814 3836
rect 15838 3834 15894 3836
rect 15598 3782 15644 3834
rect 15644 3782 15654 3834
rect 15678 3782 15708 3834
rect 15708 3782 15720 3834
rect 15720 3782 15734 3834
rect 15758 3782 15772 3834
rect 15772 3782 15784 3834
rect 15784 3782 15814 3834
rect 15838 3782 15848 3834
rect 15848 3782 15894 3834
rect 15598 3780 15654 3782
rect 15678 3780 15734 3782
rect 15758 3780 15814 3782
rect 15838 3780 15894 3782
rect 13082 1400 13138 1456
rect 12449 1114 12505 1116
rect 12529 1114 12585 1116
rect 12609 1114 12665 1116
rect 12689 1114 12745 1116
rect 12449 1062 12495 1114
rect 12495 1062 12505 1114
rect 12529 1062 12559 1114
rect 12559 1062 12571 1114
rect 12571 1062 12585 1114
rect 12609 1062 12623 1114
rect 12623 1062 12635 1114
rect 12635 1062 12665 1114
rect 12689 1062 12699 1114
rect 12699 1062 12745 1114
rect 12449 1060 12505 1062
rect 12529 1060 12585 1062
rect 12609 1060 12665 1062
rect 12689 1060 12745 1062
rect 15598 2746 15654 2748
rect 15678 2746 15734 2748
rect 15758 2746 15814 2748
rect 15838 2746 15894 2748
rect 15598 2694 15644 2746
rect 15644 2694 15654 2746
rect 15678 2694 15708 2746
rect 15708 2694 15720 2746
rect 15720 2694 15734 2746
rect 15758 2694 15772 2746
rect 15772 2694 15784 2746
rect 15784 2694 15814 2746
rect 15838 2694 15848 2746
rect 15848 2694 15894 2746
rect 15598 2692 15654 2694
rect 15678 2692 15734 2694
rect 15758 2692 15814 2694
rect 15838 2692 15894 2694
rect 15566 2372 15622 2408
rect 15566 2352 15568 2372
rect 15568 2352 15620 2372
rect 15620 2352 15622 2372
rect 15598 1658 15654 1660
rect 15678 1658 15734 1660
rect 15758 1658 15814 1660
rect 15838 1658 15894 1660
rect 15598 1606 15644 1658
rect 15644 1606 15654 1658
rect 15678 1606 15708 1658
rect 15708 1606 15720 1658
rect 15720 1606 15734 1658
rect 15758 1606 15772 1658
rect 15772 1606 15784 1658
rect 15784 1606 15814 1658
rect 15838 1606 15848 1658
rect 15848 1606 15894 1658
rect 15598 1604 15654 1606
rect 15678 1604 15734 1606
rect 15758 1604 15814 1606
rect 15838 1604 15894 1606
rect 18510 5208 18566 5264
rect 17774 4664 17830 4720
rect 18510 3712 18566 3768
rect 16946 2372 17002 2408
rect 16946 2352 16948 2372
rect 16948 2352 17000 2372
rect 17000 2352 17002 2372
rect 15598 570 15654 572
rect 15678 570 15734 572
rect 15758 570 15814 572
rect 15838 570 15894 572
rect 15598 518 15644 570
rect 15644 518 15654 570
rect 15678 518 15708 570
rect 15708 518 15720 570
rect 15720 518 15734 570
rect 15758 518 15772 570
rect 15772 518 15784 570
rect 15784 518 15814 570
rect 15838 518 15848 570
rect 15848 518 15894 570
rect 15598 516 15654 518
rect 15678 516 15734 518
rect 15758 516 15814 518
rect 15838 516 15894 518
rect 18602 2216 18658 2272
rect 18418 1808 18474 1864
rect 18510 720 18566 776
rect 6150 26 6206 28
rect 6230 26 6286 28
rect 6310 26 6366 28
rect 6390 26 6446 28
rect 6150 -26 6196 26
rect 6196 -26 6206 26
rect 6230 -26 6260 26
rect 6260 -26 6272 26
rect 6272 -26 6286 26
rect 6310 -26 6324 26
rect 6324 -26 6336 26
rect 6336 -26 6366 26
rect 6390 -26 6400 26
rect 6400 -26 6446 26
rect 6150 -28 6206 -26
rect 6230 -28 6286 -26
rect 6310 -28 6366 -26
rect 6390 -28 6446 -26
rect 12449 26 12505 28
rect 12529 26 12585 28
rect 12609 26 12665 28
rect 12689 26 12745 28
rect 12449 -26 12495 26
rect 12495 -26 12505 26
rect 12529 -26 12559 26
rect 12559 -26 12571 26
rect 12571 -26 12585 26
rect 12609 -26 12623 26
rect 12623 -26 12635 26
rect 12635 -26 12665 26
rect 12689 -26 12699 26
rect 12699 -26 12745 26
rect 12449 -28 12505 -26
rect 12529 -28 12585 -26
rect 12609 -28 12665 -26
rect 12689 -28 12745 -26
<< metal3 >>
rect 17861 11250 17927 11253
rect 19200 11250 20000 11280
rect 17861 11248 20000 11250
rect 17861 11192 17866 11248
rect 17922 11192 20000 11248
rect 17861 11190 20000 11192
rect 17861 11187 17927 11190
rect 19200 11160 20000 11190
rect 6138 9824 6458 9825
rect 6138 9760 6146 9824
rect 6210 9760 6226 9824
rect 6290 9760 6306 9824
rect 6370 9760 6386 9824
rect 6450 9760 6458 9824
rect 6138 9759 6458 9760
rect 12437 9824 12757 9825
rect 12437 9760 12445 9824
rect 12509 9760 12525 9824
rect 12589 9760 12605 9824
rect 12669 9760 12685 9824
rect 12749 9760 12757 9824
rect 12437 9759 12757 9760
rect 17769 9754 17835 9757
rect 19200 9754 20000 9784
rect 17769 9752 20000 9754
rect 17769 9696 17774 9752
rect 17830 9696 20000 9752
rect 17769 9694 20000 9696
rect 17769 9691 17835 9694
rect 19200 9664 20000 9694
rect 2989 9280 3309 9281
rect 2989 9216 2997 9280
rect 3061 9216 3077 9280
rect 3141 9216 3157 9280
rect 3221 9216 3237 9280
rect 3301 9216 3309 9280
rect 2989 9215 3309 9216
rect 9288 9280 9608 9281
rect 9288 9216 9296 9280
rect 9360 9216 9376 9280
rect 9440 9216 9456 9280
rect 9520 9216 9536 9280
rect 9600 9216 9608 9280
rect 9288 9215 9608 9216
rect 15586 9280 15906 9281
rect 15586 9216 15594 9280
rect 15658 9216 15674 9280
rect 15738 9216 15754 9280
rect 15818 9216 15834 9280
rect 15898 9216 15906 9280
rect 15586 9215 15906 9216
rect 11513 9074 11579 9077
rect 13997 9074 14063 9077
rect 11513 9072 14063 9074
rect 11513 9016 11518 9072
rect 11574 9016 14002 9072
rect 14058 9016 14063 9072
rect 11513 9014 14063 9016
rect 11513 9011 11579 9014
rect 13997 9011 14063 9014
rect 6138 8736 6458 8737
rect 6138 8672 6146 8736
rect 6210 8672 6226 8736
rect 6290 8672 6306 8736
rect 6370 8672 6386 8736
rect 6450 8672 6458 8736
rect 6138 8671 6458 8672
rect 12437 8736 12757 8737
rect 12437 8672 12445 8736
rect 12509 8672 12525 8736
rect 12589 8672 12605 8736
rect 12669 8672 12685 8736
rect 12749 8672 12757 8736
rect 12437 8671 12757 8672
rect 18597 8258 18663 8261
rect 19200 8258 20000 8288
rect 18597 8256 20000 8258
rect 18597 8200 18602 8256
rect 18658 8200 20000 8256
rect 18597 8198 20000 8200
rect 18597 8195 18663 8198
rect 2989 8192 3309 8193
rect 2989 8128 2997 8192
rect 3061 8128 3077 8192
rect 3141 8128 3157 8192
rect 3221 8128 3237 8192
rect 3301 8128 3309 8192
rect 2989 8127 3309 8128
rect 9288 8192 9608 8193
rect 9288 8128 9296 8192
rect 9360 8128 9376 8192
rect 9440 8128 9456 8192
rect 9520 8128 9536 8192
rect 9600 8128 9608 8192
rect 9288 8127 9608 8128
rect 15586 8192 15906 8193
rect 15586 8128 15594 8192
rect 15658 8128 15674 8192
rect 15738 8128 15754 8192
rect 15818 8128 15834 8192
rect 15898 8128 15906 8192
rect 19200 8168 20000 8198
rect 15586 8127 15906 8128
rect 5625 7850 5691 7853
rect 6361 7850 6427 7853
rect 14641 7850 14707 7853
rect 18229 7850 18295 7853
rect 5625 7848 8448 7850
rect 5625 7792 5630 7848
rect 5686 7792 6366 7848
rect 6422 7792 8448 7848
rect 5625 7790 8448 7792
rect 5625 7787 5691 7790
rect 6361 7787 6427 7790
rect 8388 7717 8448 7790
rect 14641 7848 18295 7850
rect 14641 7792 14646 7848
rect 14702 7792 18234 7848
rect 18290 7792 18295 7848
rect 14641 7790 18295 7792
rect 14641 7787 14707 7790
rect 18229 7787 18295 7790
rect 8385 7714 8451 7717
rect 9397 7714 9463 7717
rect 8385 7712 9463 7714
rect 8385 7656 8390 7712
rect 8446 7656 9402 7712
rect 9458 7656 9463 7712
rect 8385 7654 9463 7656
rect 8385 7651 8451 7654
rect 9397 7651 9463 7654
rect 6138 7648 6458 7649
rect 6138 7584 6146 7648
rect 6210 7584 6226 7648
rect 6290 7584 6306 7648
rect 6370 7584 6386 7648
rect 6450 7584 6458 7648
rect 6138 7583 6458 7584
rect 12437 7648 12757 7649
rect 12437 7584 12445 7648
rect 12509 7584 12525 7648
rect 12589 7584 12605 7648
rect 12669 7584 12685 7648
rect 12749 7584 12757 7648
rect 12437 7583 12757 7584
rect 6637 7442 6703 7445
rect 7833 7442 7899 7445
rect 6637 7440 7899 7442
rect 6637 7384 6642 7440
rect 6698 7384 7838 7440
rect 7894 7384 7899 7440
rect 6637 7382 7899 7384
rect 6637 7379 6703 7382
rect 7833 7379 7899 7382
rect 12341 7442 12407 7445
rect 12525 7442 12591 7445
rect 12341 7440 12591 7442
rect 12341 7384 12346 7440
rect 12402 7384 12530 7440
rect 12586 7384 12591 7440
rect 12341 7382 12591 7384
rect 12341 7379 12407 7382
rect 12525 7379 12591 7382
rect 2989 7104 3309 7105
rect 2989 7040 2997 7104
rect 3061 7040 3077 7104
rect 3141 7040 3157 7104
rect 3221 7040 3237 7104
rect 3301 7040 3309 7104
rect 2989 7039 3309 7040
rect 9288 7104 9608 7105
rect 9288 7040 9296 7104
rect 9360 7040 9376 7104
rect 9440 7040 9456 7104
rect 9520 7040 9536 7104
rect 9600 7040 9608 7104
rect 9288 7039 9608 7040
rect 15586 7104 15906 7105
rect 15586 7040 15594 7104
rect 15658 7040 15674 7104
rect 15738 7040 15754 7104
rect 15818 7040 15834 7104
rect 15898 7040 15906 7104
rect 15586 7039 15906 7040
rect 11605 6898 11671 6901
rect 12617 6898 12683 6901
rect 11605 6896 12683 6898
rect 11605 6840 11610 6896
rect 11666 6840 12622 6896
rect 12678 6840 12683 6896
rect 11605 6838 12683 6840
rect 11605 6835 11671 6838
rect 12617 6835 12683 6838
rect 13997 6762 14063 6765
rect 14733 6762 14799 6765
rect 13997 6760 14799 6762
rect 13997 6704 14002 6760
rect 14058 6704 14738 6760
rect 14794 6704 14799 6760
rect 13997 6702 14799 6704
rect 13997 6699 14063 6702
rect 14733 6699 14799 6702
rect 14917 6762 14983 6765
rect 17585 6762 17651 6765
rect 14917 6760 17651 6762
rect 14917 6704 14922 6760
rect 14978 6704 17590 6760
rect 17646 6704 17651 6760
rect 14917 6702 17651 6704
rect 14917 6699 14983 6702
rect 17585 6699 17651 6702
rect 18505 6762 18571 6765
rect 19200 6762 20000 6792
rect 18505 6760 20000 6762
rect 18505 6704 18510 6760
rect 18566 6704 20000 6760
rect 18505 6702 20000 6704
rect 18505 6699 18571 6702
rect 19200 6672 20000 6702
rect 6138 6560 6458 6561
rect 6138 6496 6146 6560
rect 6210 6496 6226 6560
rect 6290 6496 6306 6560
rect 6370 6496 6386 6560
rect 6450 6496 6458 6560
rect 6138 6495 6458 6496
rect 12437 6560 12757 6561
rect 12437 6496 12445 6560
rect 12509 6496 12525 6560
rect 12589 6496 12605 6560
rect 12669 6496 12685 6560
rect 12749 6496 12757 6560
rect 12437 6495 12757 6496
rect 10225 6490 10291 6493
rect 11789 6490 11855 6493
rect 10225 6488 11855 6490
rect 10225 6432 10230 6488
rect 10286 6432 11794 6488
rect 11850 6432 11855 6488
rect 10225 6430 11855 6432
rect 10225 6427 10291 6430
rect 11789 6427 11855 6430
rect 11605 6354 11671 6357
rect 12249 6354 12315 6357
rect 11605 6352 12315 6354
rect 11605 6296 11610 6352
rect 11666 6296 12254 6352
rect 12310 6296 12315 6352
rect 11605 6294 12315 6296
rect 11605 6291 11671 6294
rect 12249 6291 12315 6294
rect 2989 6016 3309 6017
rect 2989 5952 2997 6016
rect 3061 5952 3077 6016
rect 3141 5952 3157 6016
rect 3221 5952 3237 6016
rect 3301 5952 3309 6016
rect 2989 5951 3309 5952
rect 9288 6016 9608 6017
rect 9288 5952 9296 6016
rect 9360 5952 9376 6016
rect 9440 5952 9456 6016
rect 9520 5952 9536 6016
rect 9600 5952 9608 6016
rect 9288 5951 9608 5952
rect 15586 6016 15906 6017
rect 15586 5952 15594 6016
rect 15658 5952 15674 6016
rect 15738 5952 15754 6016
rect 15818 5952 15834 6016
rect 15898 5952 15906 6016
rect 15586 5951 15906 5952
rect 6138 5472 6458 5473
rect 6138 5408 6146 5472
rect 6210 5408 6226 5472
rect 6290 5408 6306 5472
rect 6370 5408 6386 5472
rect 6450 5408 6458 5472
rect 6138 5407 6458 5408
rect 12437 5472 12757 5473
rect 12437 5408 12445 5472
rect 12509 5408 12525 5472
rect 12589 5408 12605 5472
rect 12669 5408 12685 5472
rect 12749 5408 12757 5472
rect 12437 5407 12757 5408
rect 18505 5266 18571 5269
rect 19200 5266 20000 5296
rect 18505 5264 20000 5266
rect 18505 5208 18510 5264
rect 18566 5208 20000 5264
rect 18505 5206 20000 5208
rect 18505 5203 18571 5206
rect 19200 5176 20000 5206
rect 2989 4928 3309 4929
rect 2989 4864 2997 4928
rect 3061 4864 3077 4928
rect 3141 4864 3157 4928
rect 3221 4864 3237 4928
rect 3301 4864 3309 4928
rect 2989 4863 3309 4864
rect 9288 4928 9608 4929
rect 9288 4864 9296 4928
rect 9360 4864 9376 4928
rect 9440 4864 9456 4928
rect 9520 4864 9536 4928
rect 9600 4864 9608 4928
rect 9288 4863 9608 4864
rect 15586 4928 15906 4929
rect 15586 4864 15594 4928
rect 15658 4864 15674 4928
rect 15738 4864 15754 4928
rect 15818 4864 15834 4928
rect 15898 4864 15906 4928
rect 15586 4863 15906 4864
rect 11881 4722 11947 4725
rect 14917 4722 14983 4725
rect 17769 4722 17835 4725
rect 11881 4720 17835 4722
rect 11881 4664 11886 4720
rect 11942 4664 14922 4720
rect 14978 4664 17774 4720
rect 17830 4664 17835 4720
rect 11881 4662 17835 4664
rect 11881 4659 11947 4662
rect 14917 4659 14983 4662
rect 17769 4659 17835 4662
rect 6138 4384 6458 4385
rect 6138 4320 6146 4384
rect 6210 4320 6226 4384
rect 6290 4320 6306 4384
rect 6370 4320 6386 4384
rect 6450 4320 6458 4384
rect 6138 4319 6458 4320
rect 12437 4384 12757 4385
rect 12437 4320 12445 4384
rect 12509 4320 12525 4384
rect 12589 4320 12605 4384
rect 12669 4320 12685 4384
rect 12749 4320 12757 4384
rect 12437 4319 12757 4320
rect 2989 3840 3309 3841
rect 2989 3776 2997 3840
rect 3061 3776 3077 3840
rect 3141 3776 3157 3840
rect 3221 3776 3237 3840
rect 3301 3776 3309 3840
rect 2989 3775 3309 3776
rect 9288 3840 9608 3841
rect 9288 3776 9296 3840
rect 9360 3776 9376 3840
rect 9440 3776 9456 3840
rect 9520 3776 9536 3840
rect 9600 3776 9608 3840
rect 9288 3775 9608 3776
rect 15586 3840 15906 3841
rect 15586 3776 15594 3840
rect 15658 3776 15674 3840
rect 15738 3776 15754 3840
rect 15818 3776 15834 3840
rect 15898 3776 15906 3840
rect 15586 3775 15906 3776
rect 18505 3770 18571 3773
rect 19200 3770 20000 3800
rect 18505 3768 20000 3770
rect 18505 3712 18510 3768
rect 18566 3712 20000 3768
rect 18505 3710 20000 3712
rect 18505 3707 18571 3710
rect 19200 3680 20000 3710
rect 6138 3296 6458 3297
rect 6138 3232 6146 3296
rect 6210 3232 6226 3296
rect 6290 3232 6306 3296
rect 6370 3232 6386 3296
rect 6450 3232 6458 3296
rect 6138 3231 6458 3232
rect 12437 3296 12757 3297
rect 12437 3232 12445 3296
rect 12509 3232 12525 3296
rect 12589 3232 12605 3296
rect 12669 3232 12685 3296
rect 12749 3232 12757 3296
rect 12437 3231 12757 3232
rect 2989 2752 3309 2753
rect 2989 2688 2997 2752
rect 3061 2688 3077 2752
rect 3141 2688 3157 2752
rect 3221 2688 3237 2752
rect 3301 2688 3309 2752
rect 2989 2687 3309 2688
rect 9288 2752 9608 2753
rect 9288 2688 9296 2752
rect 9360 2688 9376 2752
rect 9440 2688 9456 2752
rect 9520 2688 9536 2752
rect 9600 2688 9608 2752
rect 9288 2687 9608 2688
rect 15586 2752 15906 2753
rect 15586 2688 15594 2752
rect 15658 2688 15674 2752
rect 15738 2688 15754 2752
rect 15818 2688 15834 2752
rect 15898 2688 15906 2752
rect 15586 2687 15906 2688
rect 15561 2410 15627 2413
rect 16941 2410 17007 2413
rect 15561 2408 17007 2410
rect 15561 2352 15566 2408
rect 15622 2352 16946 2408
rect 17002 2352 17007 2408
rect 15561 2350 17007 2352
rect 15561 2347 15627 2350
rect 16941 2347 17007 2350
rect 18597 2274 18663 2277
rect 19200 2274 20000 2304
rect 18597 2272 20000 2274
rect 18597 2216 18602 2272
rect 18658 2216 20000 2272
rect 18597 2214 20000 2216
rect 18597 2211 18663 2214
rect 6138 2208 6458 2209
rect 6138 2144 6146 2208
rect 6210 2144 6226 2208
rect 6290 2144 6306 2208
rect 6370 2144 6386 2208
rect 6450 2144 6458 2208
rect 6138 2143 6458 2144
rect 12437 2208 12757 2209
rect 12437 2144 12445 2208
rect 12509 2144 12525 2208
rect 12589 2144 12605 2208
rect 12669 2144 12685 2208
rect 12749 2144 12757 2208
rect 19200 2184 20000 2214
rect 12437 2143 12757 2144
rect 8109 2002 8175 2005
rect 9949 2002 10015 2005
rect 8109 2000 10015 2002
rect 8109 1944 8114 2000
rect 8170 1944 9954 2000
rect 10010 1944 10015 2000
rect 8109 1942 10015 1944
rect 8109 1939 8175 1942
rect 9949 1939 10015 1942
rect 8017 1866 8083 1869
rect 9489 1866 9555 1869
rect 8017 1864 9555 1866
rect 8017 1808 8022 1864
rect 8078 1808 9494 1864
rect 9550 1808 9555 1864
rect 8017 1806 9555 1808
rect 8017 1803 8083 1806
rect 9489 1803 9555 1806
rect 11329 1866 11395 1869
rect 18413 1866 18479 1869
rect 11329 1864 18479 1866
rect 11329 1808 11334 1864
rect 11390 1808 18418 1864
rect 18474 1808 18479 1864
rect 11329 1806 18479 1808
rect 11329 1803 11395 1806
rect 18413 1803 18479 1806
rect 2989 1664 3309 1665
rect 2989 1600 2997 1664
rect 3061 1600 3077 1664
rect 3141 1600 3157 1664
rect 3221 1600 3237 1664
rect 3301 1600 3309 1664
rect 2989 1599 3309 1600
rect 9288 1664 9608 1665
rect 9288 1600 9296 1664
rect 9360 1600 9376 1664
rect 9440 1600 9456 1664
rect 9520 1600 9536 1664
rect 9600 1600 9608 1664
rect 9288 1599 9608 1600
rect 15586 1664 15906 1665
rect 15586 1600 15594 1664
rect 15658 1600 15674 1664
rect 15738 1600 15754 1664
rect 15818 1600 15834 1664
rect 15898 1600 15906 1664
rect 15586 1599 15906 1600
rect 4889 1458 4955 1461
rect 8293 1458 8359 1461
rect 13077 1458 13143 1461
rect 4889 1456 5642 1458
rect 4889 1400 4894 1456
rect 4950 1400 5642 1456
rect 4889 1398 5642 1400
rect 4889 1395 4955 1398
rect 5582 1322 5642 1398
rect 8293 1456 13143 1458
rect 8293 1400 8298 1456
rect 8354 1400 13082 1456
rect 13138 1400 13143 1456
rect 8293 1398 13143 1400
rect 8293 1395 8359 1398
rect 13077 1395 13143 1398
rect 5582 1262 6746 1322
rect 6686 1186 6746 1262
rect 7005 1186 7071 1189
rect 8201 1186 8267 1189
rect 8569 1186 8635 1189
rect 6686 1184 8635 1186
rect 6686 1128 7010 1184
rect 7066 1128 8206 1184
rect 8262 1128 8574 1184
rect 8630 1128 8635 1184
rect 6686 1126 8635 1128
rect 7005 1123 7071 1126
rect 8201 1123 8267 1126
rect 8569 1123 8635 1126
rect 6138 1120 6458 1121
rect 6138 1056 6146 1120
rect 6210 1056 6226 1120
rect 6290 1056 6306 1120
rect 6370 1056 6386 1120
rect 6450 1056 6458 1120
rect 6138 1055 6458 1056
rect 12437 1120 12757 1121
rect 12437 1056 12445 1120
rect 12509 1056 12525 1120
rect 12589 1056 12605 1120
rect 12669 1056 12685 1120
rect 12749 1056 12757 1120
rect 12437 1055 12757 1056
rect 8753 1050 8819 1053
rect 10685 1050 10751 1053
rect 8753 1048 10751 1050
rect 8753 992 8758 1048
rect 8814 992 10690 1048
rect 10746 992 10751 1048
rect 8753 990 10751 992
rect 8753 987 8819 990
rect 10685 987 10751 990
rect 7189 914 7255 917
rect 9673 914 9739 917
rect 7189 912 9739 914
rect 7189 856 7194 912
rect 7250 856 9678 912
rect 9734 856 9739 912
rect 7189 854 9739 856
rect 7189 851 7255 854
rect 9673 851 9739 854
rect 6545 778 6611 781
rect 8385 778 8451 781
rect 6545 776 8451 778
rect 6545 720 6550 776
rect 6606 720 8390 776
rect 8446 720 8451 776
rect 6545 718 8451 720
rect 6545 715 6611 718
rect 8385 715 8451 718
rect 18505 778 18571 781
rect 19200 778 20000 808
rect 18505 776 20000 778
rect 18505 720 18510 776
rect 18566 720 20000 776
rect 18505 718 20000 720
rect 18505 715 18571 718
rect 19200 688 20000 718
rect 2989 576 3309 577
rect 2989 512 2997 576
rect 3061 512 3077 576
rect 3141 512 3157 576
rect 3221 512 3237 576
rect 3301 512 3309 576
rect 2989 511 3309 512
rect 9288 576 9608 577
rect 9288 512 9296 576
rect 9360 512 9376 576
rect 9440 512 9456 576
rect 9520 512 9536 576
rect 9600 512 9608 576
rect 9288 511 9608 512
rect 15586 576 15906 577
rect 15586 512 15594 576
rect 15658 512 15674 576
rect 15738 512 15754 576
rect 15818 512 15834 576
rect 15898 512 15906 576
rect 15586 511 15906 512
rect 8845 370 8911 373
rect 11053 370 11119 373
rect 8845 368 11119 370
rect 8845 312 8850 368
rect 8906 312 11058 368
rect 11114 312 11119 368
rect 8845 310 11119 312
rect 8845 307 8911 310
rect 11053 307 11119 310
rect 6138 32 6458 33
rect 6138 -32 6146 32
rect 6210 -32 6226 32
rect 6290 -32 6306 32
rect 6370 -32 6386 32
rect 6450 -32 6458 32
rect 6138 -33 6458 -32
rect 12437 32 12757 33
rect 12437 -32 12445 32
rect 12509 -32 12525 32
rect 12589 -32 12605 32
rect 12669 -32 12685 32
rect 12749 -32 12757 32
rect 12437 -33 12757 -32
<< via3 >>
rect 6146 9820 6210 9824
rect 6146 9764 6150 9820
rect 6150 9764 6206 9820
rect 6206 9764 6210 9820
rect 6146 9760 6210 9764
rect 6226 9820 6290 9824
rect 6226 9764 6230 9820
rect 6230 9764 6286 9820
rect 6286 9764 6290 9820
rect 6226 9760 6290 9764
rect 6306 9820 6370 9824
rect 6306 9764 6310 9820
rect 6310 9764 6366 9820
rect 6366 9764 6370 9820
rect 6306 9760 6370 9764
rect 6386 9820 6450 9824
rect 6386 9764 6390 9820
rect 6390 9764 6446 9820
rect 6446 9764 6450 9820
rect 6386 9760 6450 9764
rect 12445 9820 12509 9824
rect 12445 9764 12449 9820
rect 12449 9764 12505 9820
rect 12505 9764 12509 9820
rect 12445 9760 12509 9764
rect 12525 9820 12589 9824
rect 12525 9764 12529 9820
rect 12529 9764 12585 9820
rect 12585 9764 12589 9820
rect 12525 9760 12589 9764
rect 12605 9820 12669 9824
rect 12605 9764 12609 9820
rect 12609 9764 12665 9820
rect 12665 9764 12669 9820
rect 12605 9760 12669 9764
rect 12685 9820 12749 9824
rect 12685 9764 12689 9820
rect 12689 9764 12745 9820
rect 12745 9764 12749 9820
rect 12685 9760 12749 9764
rect 2997 9276 3061 9280
rect 2997 9220 3001 9276
rect 3001 9220 3057 9276
rect 3057 9220 3061 9276
rect 2997 9216 3061 9220
rect 3077 9276 3141 9280
rect 3077 9220 3081 9276
rect 3081 9220 3137 9276
rect 3137 9220 3141 9276
rect 3077 9216 3141 9220
rect 3157 9276 3221 9280
rect 3157 9220 3161 9276
rect 3161 9220 3217 9276
rect 3217 9220 3221 9276
rect 3157 9216 3221 9220
rect 3237 9276 3301 9280
rect 3237 9220 3241 9276
rect 3241 9220 3297 9276
rect 3297 9220 3301 9276
rect 3237 9216 3301 9220
rect 9296 9276 9360 9280
rect 9296 9220 9300 9276
rect 9300 9220 9356 9276
rect 9356 9220 9360 9276
rect 9296 9216 9360 9220
rect 9376 9276 9440 9280
rect 9376 9220 9380 9276
rect 9380 9220 9436 9276
rect 9436 9220 9440 9276
rect 9376 9216 9440 9220
rect 9456 9276 9520 9280
rect 9456 9220 9460 9276
rect 9460 9220 9516 9276
rect 9516 9220 9520 9276
rect 9456 9216 9520 9220
rect 9536 9276 9600 9280
rect 9536 9220 9540 9276
rect 9540 9220 9596 9276
rect 9596 9220 9600 9276
rect 9536 9216 9600 9220
rect 15594 9276 15658 9280
rect 15594 9220 15598 9276
rect 15598 9220 15654 9276
rect 15654 9220 15658 9276
rect 15594 9216 15658 9220
rect 15674 9276 15738 9280
rect 15674 9220 15678 9276
rect 15678 9220 15734 9276
rect 15734 9220 15738 9276
rect 15674 9216 15738 9220
rect 15754 9276 15818 9280
rect 15754 9220 15758 9276
rect 15758 9220 15814 9276
rect 15814 9220 15818 9276
rect 15754 9216 15818 9220
rect 15834 9276 15898 9280
rect 15834 9220 15838 9276
rect 15838 9220 15894 9276
rect 15894 9220 15898 9276
rect 15834 9216 15898 9220
rect 6146 8732 6210 8736
rect 6146 8676 6150 8732
rect 6150 8676 6206 8732
rect 6206 8676 6210 8732
rect 6146 8672 6210 8676
rect 6226 8732 6290 8736
rect 6226 8676 6230 8732
rect 6230 8676 6286 8732
rect 6286 8676 6290 8732
rect 6226 8672 6290 8676
rect 6306 8732 6370 8736
rect 6306 8676 6310 8732
rect 6310 8676 6366 8732
rect 6366 8676 6370 8732
rect 6306 8672 6370 8676
rect 6386 8732 6450 8736
rect 6386 8676 6390 8732
rect 6390 8676 6446 8732
rect 6446 8676 6450 8732
rect 6386 8672 6450 8676
rect 12445 8732 12509 8736
rect 12445 8676 12449 8732
rect 12449 8676 12505 8732
rect 12505 8676 12509 8732
rect 12445 8672 12509 8676
rect 12525 8732 12589 8736
rect 12525 8676 12529 8732
rect 12529 8676 12585 8732
rect 12585 8676 12589 8732
rect 12525 8672 12589 8676
rect 12605 8732 12669 8736
rect 12605 8676 12609 8732
rect 12609 8676 12665 8732
rect 12665 8676 12669 8732
rect 12605 8672 12669 8676
rect 12685 8732 12749 8736
rect 12685 8676 12689 8732
rect 12689 8676 12745 8732
rect 12745 8676 12749 8732
rect 12685 8672 12749 8676
rect 2997 8188 3061 8192
rect 2997 8132 3001 8188
rect 3001 8132 3057 8188
rect 3057 8132 3061 8188
rect 2997 8128 3061 8132
rect 3077 8188 3141 8192
rect 3077 8132 3081 8188
rect 3081 8132 3137 8188
rect 3137 8132 3141 8188
rect 3077 8128 3141 8132
rect 3157 8188 3221 8192
rect 3157 8132 3161 8188
rect 3161 8132 3217 8188
rect 3217 8132 3221 8188
rect 3157 8128 3221 8132
rect 3237 8188 3301 8192
rect 3237 8132 3241 8188
rect 3241 8132 3297 8188
rect 3297 8132 3301 8188
rect 3237 8128 3301 8132
rect 9296 8188 9360 8192
rect 9296 8132 9300 8188
rect 9300 8132 9356 8188
rect 9356 8132 9360 8188
rect 9296 8128 9360 8132
rect 9376 8188 9440 8192
rect 9376 8132 9380 8188
rect 9380 8132 9436 8188
rect 9436 8132 9440 8188
rect 9376 8128 9440 8132
rect 9456 8188 9520 8192
rect 9456 8132 9460 8188
rect 9460 8132 9516 8188
rect 9516 8132 9520 8188
rect 9456 8128 9520 8132
rect 9536 8188 9600 8192
rect 9536 8132 9540 8188
rect 9540 8132 9596 8188
rect 9596 8132 9600 8188
rect 9536 8128 9600 8132
rect 15594 8188 15658 8192
rect 15594 8132 15598 8188
rect 15598 8132 15654 8188
rect 15654 8132 15658 8188
rect 15594 8128 15658 8132
rect 15674 8188 15738 8192
rect 15674 8132 15678 8188
rect 15678 8132 15734 8188
rect 15734 8132 15738 8188
rect 15674 8128 15738 8132
rect 15754 8188 15818 8192
rect 15754 8132 15758 8188
rect 15758 8132 15814 8188
rect 15814 8132 15818 8188
rect 15754 8128 15818 8132
rect 15834 8188 15898 8192
rect 15834 8132 15838 8188
rect 15838 8132 15894 8188
rect 15894 8132 15898 8188
rect 15834 8128 15898 8132
rect 6146 7644 6210 7648
rect 6146 7588 6150 7644
rect 6150 7588 6206 7644
rect 6206 7588 6210 7644
rect 6146 7584 6210 7588
rect 6226 7644 6290 7648
rect 6226 7588 6230 7644
rect 6230 7588 6286 7644
rect 6286 7588 6290 7644
rect 6226 7584 6290 7588
rect 6306 7644 6370 7648
rect 6306 7588 6310 7644
rect 6310 7588 6366 7644
rect 6366 7588 6370 7644
rect 6306 7584 6370 7588
rect 6386 7644 6450 7648
rect 6386 7588 6390 7644
rect 6390 7588 6446 7644
rect 6446 7588 6450 7644
rect 6386 7584 6450 7588
rect 12445 7644 12509 7648
rect 12445 7588 12449 7644
rect 12449 7588 12505 7644
rect 12505 7588 12509 7644
rect 12445 7584 12509 7588
rect 12525 7644 12589 7648
rect 12525 7588 12529 7644
rect 12529 7588 12585 7644
rect 12585 7588 12589 7644
rect 12525 7584 12589 7588
rect 12605 7644 12669 7648
rect 12605 7588 12609 7644
rect 12609 7588 12665 7644
rect 12665 7588 12669 7644
rect 12605 7584 12669 7588
rect 12685 7644 12749 7648
rect 12685 7588 12689 7644
rect 12689 7588 12745 7644
rect 12745 7588 12749 7644
rect 12685 7584 12749 7588
rect 2997 7100 3061 7104
rect 2997 7044 3001 7100
rect 3001 7044 3057 7100
rect 3057 7044 3061 7100
rect 2997 7040 3061 7044
rect 3077 7100 3141 7104
rect 3077 7044 3081 7100
rect 3081 7044 3137 7100
rect 3137 7044 3141 7100
rect 3077 7040 3141 7044
rect 3157 7100 3221 7104
rect 3157 7044 3161 7100
rect 3161 7044 3217 7100
rect 3217 7044 3221 7100
rect 3157 7040 3221 7044
rect 3237 7100 3301 7104
rect 3237 7044 3241 7100
rect 3241 7044 3297 7100
rect 3297 7044 3301 7100
rect 3237 7040 3301 7044
rect 9296 7100 9360 7104
rect 9296 7044 9300 7100
rect 9300 7044 9356 7100
rect 9356 7044 9360 7100
rect 9296 7040 9360 7044
rect 9376 7100 9440 7104
rect 9376 7044 9380 7100
rect 9380 7044 9436 7100
rect 9436 7044 9440 7100
rect 9376 7040 9440 7044
rect 9456 7100 9520 7104
rect 9456 7044 9460 7100
rect 9460 7044 9516 7100
rect 9516 7044 9520 7100
rect 9456 7040 9520 7044
rect 9536 7100 9600 7104
rect 9536 7044 9540 7100
rect 9540 7044 9596 7100
rect 9596 7044 9600 7100
rect 9536 7040 9600 7044
rect 15594 7100 15658 7104
rect 15594 7044 15598 7100
rect 15598 7044 15654 7100
rect 15654 7044 15658 7100
rect 15594 7040 15658 7044
rect 15674 7100 15738 7104
rect 15674 7044 15678 7100
rect 15678 7044 15734 7100
rect 15734 7044 15738 7100
rect 15674 7040 15738 7044
rect 15754 7100 15818 7104
rect 15754 7044 15758 7100
rect 15758 7044 15814 7100
rect 15814 7044 15818 7100
rect 15754 7040 15818 7044
rect 15834 7100 15898 7104
rect 15834 7044 15838 7100
rect 15838 7044 15894 7100
rect 15894 7044 15898 7100
rect 15834 7040 15898 7044
rect 6146 6556 6210 6560
rect 6146 6500 6150 6556
rect 6150 6500 6206 6556
rect 6206 6500 6210 6556
rect 6146 6496 6210 6500
rect 6226 6556 6290 6560
rect 6226 6500 6230 6556
rect 6230 6500 6286 6556
rect 6286 6500 6290 6556
rect 6226 6496 6290 6500
rect 6306 6556 6370 6560
rect 6306 6500 6310 6556
rect 6310 6500 6366 6556
rect 6366 6500 6370 6556
rect 6306 6496 6370 6500
rect 6386 6556 6450 6560
rect 6386 6500 6390 6556
rect 6390 6500 6446 6556
rect 6446 6500 6450 6556
rect 6386 6496 6450 6500
rect 12445 6556 12509 6560
rect 12445 6500 12449 6556
rect 12449 6500 12505 6556
rect 12505 6500 12509 6556
rect 12445 6496 12509 6500
rect 12525 6556 12589 6560
rect 12525 6500 12529 6556
rect 12529 6500 12585 6556
rect 12585 6500 12589 6556
rect 12525 6496 12589 6500
rect 12605 6556 12669 6560
rect 12605 6500 12609 6556
rect 12609 6500 12665 6556
rect 12665 6500 12669 6556
rect 12605 6496 12669 6500
rect 12685 6556 12749 6560
rect 12685 6500 12689 6556
rect 12689 6500 12745 6556
rect 12745 6500 12749 6556
rect 12685 6496 12749 6500
rect 2997 6012 3061 6016
rect 2997 5956 3001 6012
rect 3001 5956 3057 6012
rect 3057 5956 3061 6012
rect 2997 5952 3061 5956
rect 3077 6012 3141 6016
rect 3077 5956 3081 6012
rect 3081 5956 3137 6012
rect 3137 5956 3141 6012
rect 3077 5952 3141 5956
rect 3157 6012 3221 6016
rect 3157 5956 3161 6012
rect 3161 5956 3217 6012
rect 3217 5956 3221 6012
rect 3157 5952 3221 5956
rect 3237 6012 3301 6016
rect 3237 5956 3241 6012
rect 3241 5956 3297 6012
rect 3297 5956 3301 6012
rect 3237 5952 3301 5956
rect 9296 6012 9360 6016
rect 9296 5956 9300 6012
rect 9300 5956 9356 6012
rect 9356 5956 9360 6012
rect 9296 5952 9360 5956
rect 9376 6012 9440 6016
rect 9376 5956 9380 6012
rect 9380 5956 9436 6012
rect 9436 5956 9440 6012
rect 9376 5952 9440 5956
rect 9456 6012 9520 6016
rect 9456 5956 9460 6012
rect 9460 5956 9516 6012
rect 9516 5956 9520 6012
rect 9456 5952 9520 5956
rect 9536 6012 9600 6016
rect 9536 5956 9540 6012
rect 9540 5956 9596 6012
rect 9596 5956 9600 6012
rect 9536 5952 9600 5956
rect 15594 6012 15658 6016
rect 15594 5956 15598 6012
rect 15598 5956 15654 6012
rect 15654 5956 15658 6012
rect 15594 5952 15658 5956
rect 15674 6012 15738 6016
rect 15674 5956 15678 6012
rect 15678 5956 15734 6012
rect 15734 5956 15738 6012
rect 15674 5952 15738 5956
rect 15754 6012 15818 6016
rect 15754 5956 15758 6012
rect 15758 5956 15814 6012
rect 15814 5956 15818 6012
rect 15754 5952 15818 5956
rect 15834 6012 15898 6016
rect 15834 5956 15838 6012
rect 15838 5956 15894 6012
rect 15894 5956 15898 6012
rect 15834 5952 15898 5956
rect 6146 5468 6210 5472
rect 6146 5412 6150 5468
rect 6150 5412 6206 5468
rect 6206 5412 6210 5468
rect 6146 5408 6210 5412
rect 6226 5468 6290 5472
rect 6226 5412 6230 5468
rect 6230 5412 6286 5468
rect 6286 5412 6290 5468
rect 6226 5408 6290 5412
rect 6306 5468 6370 5472
rect 6306 5412 6310 5468
rect 6310 5412 6366 5468
rect 6366 5412 6370 5468
rect 6306 5408 6370 5412
rect 6386 5468 6450 5472
rect 6386 5412 6390 5468
rect 6390 5412 6446 5468
rect 6446 5412 6450 5468
rect 6386 5408 6450 5412
rect 12445 5468 12509 5472
rect 12445 5412 12449 5468
rect 12449 5412 12505 5468
rect 12505 5412 12509 5468
rect 12445 5408 12509 5412
rect 12525 5468 12589 5472
rect 12525 5412 12529 5468
rect 12529 5412 12585 5468
rect 12585 5412 12589 5468
rect 12525 5408 12589 5412
rect 12605 5468 12669 5472
rect 12605 5412 12609 5468
rect 12609 5412 12665 5468
rect 12665 5412 12669 5468
rect 12605 5408 12669 5412
rect 12685 5468 12749 5472
rect 12685 5412 12689 5468
rect 12689 5412 12745 5468
rect 12745 5412 12749 5468
rect 12685 5408 12749 5412
rect 2997 4924 3061 4928
rect 2997 4868 3001 4924
rect 3001 4868 3057 4924
rect 3057 4868 3061 4924
rect 2997 4864 3061 4868
rect 3077 4924 3141 4928
rect 3077 4868 3081 4924
rect 3081 4868 3137 4924
rect 3137 4868 3141 4924
rect 3077 4864 3141 4868
rect 3157 4924 3221 4928
rect 3157 4868 3161 4924
rect 3161 4868 3217 4924
rect 3217 4868 3221 4924
rect 3157 4864 3221 4868
rect 3237 4924 3301 4928
rect 3237 4868 3241 4924
rect 3241 4868 3297 4924
rect 3297 4868 3301 4924
rect 3237 4864 3301 4868
rect 9296 4924 9360 4928
rect 9296 4868 9300 4924
rect 9300 4868 9356 4924
rect 9356 4868 9360 4924
rect 9296 4864 9360 4868
rect 9376 4924 9440 4928
rect 9376 4868 9380 4924
rect 9380 4868 9436 4924
rect 9436 4868 9440 4924
rect 9376 4864 9440 4868
rect 9456 4924 9520 4928
rect 9456 4868 9460 4924
rect 9460 4868 9516 4924
rect 9516 4868 9520 4924
rect 9456 4864 9520 4868
rect 9536 4924 9600 4928
rect 9536 4868 9540 4924
rect 9540 4868 9596 4924
rect 9596 4868 9600 4924
rect 9536 4864 9600 4868
rect 15594 4924 15658 4928
rect 15594 4868 15598 4924
rect 15598 4868 15654 4924
rect 15654 4868 15658 4924
rect 15594 4864 15658 4868
rect 15674 4924 15738 4928
rect 15674 4868 15678 4924
rect 15678 4868 15734 4924
rect 15734 4868 15738 4924
rect 15674 4864 15738 4868
rect 15754 4924 15818 4928
rect 15754 4868 15758 4924
rect 15758 4868 15814 4924
rect 15814 4868 15818 4924
rect 15754 4864 15818 4868
rect 15834 4924 15898 4928
rect 15834 4868 15838 4924
rect 15838 4868 15894 4924
rect 15894 4868 15898 4924
rect 15834 4864 15898 4868
rect 6146 4380 6210 4384
rect 6146 4324 6150 4380
rect 6150 4324 6206 4380
rect 6206 4324 6210 4380
rect 6146 4320 6210 4324
rect 6226 4380 6290 4384
rect 6226 4324 6230 4380
rect 6230 4324 6286 4380
rect 6286 4324 6290 4380
rect 6226 4320 6290 4324
rect 6306 4380 6370 4384
rect 6306 4324 6310 4380
rect 6310 4324 6366 4380
rect 6366 4324 6370 4380
rect 6306 4320 6370 4324
rect 6386 4380 6450 4384
rect 6386 4324 6390 4380
rect 6390 4324 6446 4380
rect 6446 4324 6450 4380
rect 6386 4320 6450 4324
rect 12445 4380 12509 4384
rect 12445 4324 12449 4380
rect 12449 4324 12505 4380
rect 12505 4324 12509 4380
rect 12445 4320 12509 4324
rect 12525 4380 12589 4384
rect 12525 4324 12529 4380
rect 12529 4324 12585 4380
rect 12585 4324 12589 4380
rect 12525 4320 12589 4324
rect 12605 4380 12669 4384
rect 12605 4324 12609 4380
rect 12609 4324 12665 4380
rect 12665 4324 12669 4380
rect 12605 4320 12669 4324
rect 12685 4380 12749 4384
rect 12685 4324 12689 4380
rect 12689 4324 12745 4380
rect 12745 4324 12749 4380
rect 12685 4320 12749 4324
rect 2997 3836 3061 3840
rect 2997 3780 3001 3836
rect 3001 3780 3057 3836
rect 3057 3780 3061 3836
rect 2997 3776 3061 3780
rect 3077 3836 3141 3840
rect 3077 3780 3081 3836
rect 3081 3780 3137 3836
rect 3137 3780 3141 3836
rect 3077 3776 3141 3780
rect 3157 3836 3221 3840
rect 3157 3780 3161 3836
rect 3161 3780 3217 3836
rect 3217 3780 3221 3836
rect 3157 3776 3221 3780
rect 3237 3836 3301 3840
rect 3237 3780 3241 3836
rect 3241 3780 3297 3836
rect 3297 3780 3301 3836
rect 3237 3776 3301 3780
rect 9296 3836 9360 3840
rect 9296 3780 9300 3836
rect 9300 3780 9356 3836
rect 9356 3780 9360 3836
rect 9296 3776 9360 3780
rect 9376 3836 9440 3840
rect 9376 3780 9380 3836
rect 9380 3780 9436 3836
rect 9436 3780 9440 3836
rect 9376 3776 9440 3780
rect 9456 3836 9520 3840
rect 9456 3780 9460 3836
rect 9460 3780 9516 3836
rect 9516 3780 9520 3836
rect 9456 3776 9520 3780
rect 9536 3836 9600 3840
rect 9536 3780 9540 3836
rect 9540 3780 9596 3836
rect 9596 3780 9600 3836
rect 9536 3776 9600 3780
rect 15594 3836 15658 3840
rect 15594 3780 15598 3836
rect 15598 3780 15654 3836
rect 15654 3780 15658 3836
rect 15594 3776 15658 3780
rect 15674 3836 15738 3840
rect 15674 3780 15678 3836
rect 15678 3780 15734 3836
rect 15734 3780 15738 3836
rect 15674 3776 15738 3780
rect 15754 3836 15818 3840
rect 15754 3780 15758 3836
rect 15758 3780 15814 3836
rect 15814 3780 15818 3836
rect 15754 3776 15818 3780
rect 15834 3836 15898 3840
rect 15834 3780 15838 3836
rect 15838 3780 15894 3836
rect 15894 3780 15898 3836
rect 15834 3776 15898 3780
rect 6146 3292 6210 3296
rect 6146 3236 6150 3292
rect 6150 3236 6206 3292
rect 6206 3236 6210 3292
rect 6146 3232 6210 3236
rect 6226 3292 6290 3296
rect 6226 3236 6230 3292
rect 6230 3236 6286 3292
rect 6286 3236 6290 3292
rect 6226 3232 6290 3236
rect 6306 3292 6370 3296
rect 6306 3236 6310 3292
rect 6310 3236 6366 3292
rect 6366 3236 6370 3292
rect 6306 3232 6370 3236
rect 6386 3292 6450 3296
rect 6386 3236 6390 3292
rect 6390 3236 6446 3292
rect 6446 3236 6450 3292
rect 6386 3232 6450 3236
rect 12445 3292 12509 3296
rect 12445 3236 12449 3292
rect 12449 3236 12505 3292
rect 12505 3236 12509 3292
rect 12445 3232 12509 3236
rect 12525 3292 12589 3296
rect 12525 3236 12529 3292
rect 12529 3236 12585 3292
rect 12585 3236 12589 3292
rect 12525 3232 12589 3236
rect 12605 3292 12669 3296
rect 12605 3236 12609 3292
rect 12609 3236 12665 3292
rect 12665 3236 12669 3292
rect 12605 3232 12669 3236
rect 12685 3292 12749 3296
rect 12685 3236 12689 3292
rect 12689 3236 12745 3292
rect 12745 3236 12749 3292
rect 12685 3232 12749 3236
rect 2997 2748 3061 2752
rect 2997 2692 3001 2748
rect 3001 2692 3057 2748
rect 3057 2692 3061 2748
rect 2997 2688 3061 2692
rect 3077 2748 3141 2752
rect 3077 2692 3081 2748
rect 3081 2692 3137 2748
rect 3137 2692 3141 2748
rect 3077 2688 3141 2692
rect 3157 2748 3221 2752
rect 3157 2692 3161 2748
rect 3161 2692 3217 2748
rect 3217 2692 3221 2748
rect 3157 2688 3221 2692
rect 3237 2748 3301 2752
rect 3237 2692 3241 2748
rect 3241 2692 3297 2748
rect 3297 2692 3301 2748
rect 3237 2688 3301 2692
rect 9296 2748 9360 2752
rect 9296 2692 9300 2748
rect 9300 2692 9356 2748
rect 9356 2692 9360 2748
rect 9296 2688 9360 2692
rect 9376 2748 9440 2752
rect 9376 2692 9380 2748
rect 9380 2692 9436 2748
rect 9436 2692 9440 2748
rect 9376 2688 9440 2692
rect 9456 2748 9520 2752
rect 9456 2692 9460 2748
rect 9460 2692 9516 2748
rect 9516 2692 9520 2748
rect 9456 2688 9520 2692
rect 9536 2748 9600 2752
rect 9536 2692 9540 2748
rect 9540 2692 9596 2748
rect 9596 2692 9600 2748
rect 9536 2688 9600 2692
rect 15594 2748 15658 2752
rect 15594 2692 15598 2748
rect 15598 2692 15654 2748
rect 15654 2692 15658 2748
rect 15594 2688 15658 2692
rect 15674 2748 15738 2752
rect 15674 2692 15678 2748
rect 15678 2692 15734 2748
rect 15734 2692 15738 2748
rect 15674 2688 15738 2692
rect 15754 2748 15818 2752
rect 15754 2692 15758 2748
rect 15758 2692 15814 2748
rect 15814 2692 15818 2748
rect 15754 2688 15818 2692
rect 15834 2748 15898 2752
rect 15834 2692 15838 2748
rect 15838 2692 15894 2748
rect 15894 2692 15898 2748
rect 15834 2688 15898 2692
rect 6146 2204 6210 2208
rect 6146 2148 6150 2204
rect 6150 2148 6206 2204
rect 6206 2148 6210 2204
rect 6146 2144 6210 2148
rect 6226 2204 6290 2208
rect 6226 2148 6230 2204
rect 6230 2148 6286 2204
rect 6286 2148 6290 2204
rect 6226 2144 6290 2148
rect 6306 2204 6370 2208
rect 6306 2148 6310 2204
rect 6310 2148 6366 2204
rect 6366 2148 6370 2204
rect 6306 2144 6370 2148
rect 6386 2204 6450 2208
rect 6386 2148 6390 2204
rect 6390 2148 6446 2204
rect 6446 2148 6450 2204
rect 6386 2144 6450 2148
rect 12445 2204 12509 2208
rect 12445 2148 12449 2204
rect 12449 2148 12505 2204
rect 12505 2148 12509 2204
rect 12445 2144 12509 2148
rect 12525 2204 12589 2208
rect 12525 2148 12529 2204
rect 12529 2148 12585 2204
rect 12585 2148 12589 2204
rect 12525 2144 12589 2148
rect 12605 2204 12669 2208
rect 12605 2148 12609 2204
rect 12609 2148 12665 2204
rect 12665 2148 12669 2204
rect 12605 2144 12669 2148
rect 12685 2204 12749 2208
rect 12685 2148 12689 2204
rect 12689 2148 12745 2204
rect 12745 2148 12749 2204
rect 12685 2144 12749 2148
rect 2997 1660 3061 1664
rect 2997 1604 3001 1660
rect 3001 1604 3057 1660
rect 3057 1604 3061 1660
rect 2997 1600 3061 1604
rect 3077 1660 3141 1664
rect 3077 1604 3081 1660
rect 3081 1604 3137 1660
rect 3137 1604 3141 1660
rect 3077 1600 3141 1604
rect 3157 1660 3221 1664
rect 3157 1604 3161 1660
rect 3161 1604 3217 1660
rect 3217 1604 3221 1660
rect 3157 1600 3221 1604
rect 3237 1660 3301 1664
rect 3237 1604 3241 1660
rect 3241 1604 3297 1660
rect 3297 1604 3301 1660
rect 3237 1600 3301 1604
rect 9296 1660 9360 1664
rect 9296 1604 9300 1660
rect 9300 1604 9356 1660
rect 9356 1604 9360 1660
rect 9296 1600 9360 1604
rect 9376 1660 9440 1664
rect 9376 1604 9380 1660
rect 9380 1604 9436 1660
rect 9436 1604 9440 1660
rect 9376 1600 9440 1604
rect 9456 1660 9520 1664
rect 9456 1604 9460 1660
rect 9460 1604 9516 1660
rect 9516 1604 9520 1660
rect 9456 1600 9520 1604
rect 9536 1660 9600 1664
rect 9536 1604 9540 1660
rect 9540 1604 9596 1660
rect 9596 1604 9600 1660
rect 9536 1600 9600 1604
rect 15594 1660 15658 1664
rect 15594 1604 15598 1660
rect 15598 1604 15654 1660
rect 15654 1604 15658 1660
rect 15594 1600 15658 1604
rect 15674 1660 15738 1664
rect 15674 1604 15678 1660
rect 15678 1604 15734 1660
rect 15734 1604 15738 1660
rect 15674 1600 15738 1604
rect 15754 1660 15818 1664
rect 15754 1604 15758 1660
rect 15758 1604 15814 1660
rect 15814 1604 15818 1660
rect 15754 1600 15818 1604
rect 15834 1660 15898 1664
rect 15834 1604 15838 1660
rect 15838 1604 15894 1660
rect 15894 1604 15898 1660
rect 15834 1600 15898 1604
rect 6146 1116 6210 1120
rect 6146 1060 6150 1116
rect 6150 1060 6206 1116
rect 6206 1060 6210 1116
rect 6146 1056 6210 1060
rect 6226 1116 6290 1120
rect 6226 1060 6230 1116
rect 6230 1060 6286 1116
rect 6286 1060 6290 1116
rect 6226 1056 6290 1060
rect 6306 1116 6370 1120
rect 6306 1060 6310 1116
rect 6310 1060 6366 1116
rect 6366 1060 6370 1116
rect 6306 1056 6370 1060
rect 6386 1116 6450 1120
rect 6386 1060 6390 1116
rect 6390 1060 6446 1116
rect 6446 1060 6450 1116
rect 6386 1056 6450 1060
rect 12445 1116 12509 1120
rect 12445 1060 12449 1116
rect 12449 1060 12505 1116
rect 12505 1060 12509 1116
rect 12445 1056 12509 1060
rect 12525 1116 12589 1120
rect 12525 1060 12529 1116
rect 12529 1060 12585 1116
rect 12585 1060 12589 1116
rect 12525 1056 12589 1060
rect 12605 1116 12669 1120
rect 12605 1060 12609 1116
rect 12609 1060 12665 1116
rect 12665 1060 12669 1116
rect 12605 1056 12669 1060
rect 12685 1116 12749 1120
rect 12685 1060 12689 1116
rect 12689 1060 12745 1116
rect 12745 1060 12749 1116
rect 12685 1056 12749 1060
rect 2997 572 3061 576
rect 2997 516 3001 572
rect 3001 516 3057 572
rect 3057 516 3061 572
rect 2997 512 3061 516
rect 3077 572 3141 576
rect 3077 516 3081 572
rect 3081 516 3137 572
rect 3137 516 3141 572
rect 3077 512 3141 516
rect 3157 572 3221 576
rect 3157 516 3161 572
rect 3161 516 3217 572
rect 3217 516 3221 572
rect 3157 512 3221 516
rect 3237 572 3301 576
rect 3237 516 3241 572
rect 3241 516 3297 572
rect 3297 516 3301 572
rect 3237 512 3301 516
rect 9296 572 9360 576
rect 9296 516 9300 572
rect 9300 516 9356 572
rect 9356 516 9360 572
rect 9296 512 9360 516
rect 9376 572 9440 576
rect 9376 516 9380 572
rect 9380 516 9436 572
rect 9436 516 9440 572
rect 9376 512 9440 516
rect 9456 572 9520 576
rect 9456 516 9460 572
rect 9460 516 9516 572
rect 9516 516 9520 572
rect 9456 512 9520 516
rect 9536 572 9600 576
rect 9536 516 9540 572
rect 9540 516 9596 572
rect 9596 516 9600 572
rect 9536 512 9600 516
rect 15594 572 15658 576
rect 15594 516 15598 572
rect 15598 516 15654 572
rect 15654 516 15658 572
rect 15594 512 15658 516
rect 15674 572 15738 576
rect 15674 516 15678 572
rect 15678 516 15734 572
rect 15734 516 15738 572
rect 15674 512 15738 516
rect 15754 572 15818 576
rect 15754 516 15758 572
rect 15758 516 15814 572
rect 15814 516 15818 572
rect 15754 512 15818 516
rect 15834 572 15898 576
rect 15834 516 15838 572
rect 15838 516 15894 572
rect 15894 516 15898 572
rect 15834 512 15898 516
rect 6146 28 6210 32
rect 6146 -28 6150 28
rect 6150 -28 6206 28
rect 6206 -28 6210 28
rect 6146 -32 6210 -28
rect 6226 28 6290 32
rect 6226 -28 6230 28
rect 6230 -28 6286 28
rect 6286 -28 6290 28
rect 6226 -32 6290 -28
rect 6306 28 6370 32
rect 6306 -28 6310 28
rect 6310 -28 6366 28
rect 6366 -28 6370 28
rect 6306 -32 6370 -28
rect 6386 28 6450 32
rect 6386 -28 6390 28
rect 6390 -28 6446 28
rect 6446 -28 6450 28
rect 6386 -32 6450 -28
rect 12445 28 12509 32
rect 12445 -28 12449 28
rect 12449 -28 12505 28
rect 12505 -28 12509 28
rect 12445 -32 12509 -28
rect 12525 28 12589 32
rect 12525 -28 12529 28
rect 12529 -28 12585 28
rect 12585 -28 12589 28
rect 12525 -32 12589 -28
rect 12605 28 12669 32
rect 12605 -28 12609 28
rect 12609 -28 12665 28
rect 12665 -28 12669 28
rect 12605 -32 12669 -28
rect 12685 28 12749 32
rect 12685 -28 12689 28
rect 12689 -28 12745 28
rect 12745 -28 12749 28
rect 12685 -32 12749 -28
<< metal4 >>
rect 2989 9280 3309 9840
rect 2989 9216 2997 9280
rect 3061 9216 3077 9280
rect 3141 9216 3157 9280
rect 3221 9216 3237 9280
rect 3301 9216 3309 9280
rect 2989 8256 3309 9216
rect 2989 8192 3031 8256
rect 3267 8192 3309 8256
rect 2989 8128 2997 8192
rect 3301 8128 3309 8192
rect 2989 8020 3031 8128
rect 3267 8020 3309 8128
rect 2989 7104 3309 8020
rect 2989 7040 2997 7104
rect 3061 7040 3077 7104
rect 3141 7040 3157 7104
rect 3221 7040 3237 7104
rect 3301 7040 3309 7104
rect 2989 6016 3309 7040
rect 2989 5952 2997 6016
rect 3061 5952 3077 6016
rect 3141 5952 3157 6016
rect 3221 5952 3237 6016
rect 3301 5952 3309 6016
rect 2989 4982 3309 5952
rect 2989 4928 3031 4982
rect 3267 4928 3309 4982
rect 2989 4864 2997 4928
rect 3301 4864 3309 4928
rect 2989 4746 3031 4864
rect 3267 4746 3309 4864
rect 2989 3840 3309 4746
rect 2989 3776 2997 3840
rect 3061 3776 3077 3840
rect 3141 3776 3157 3840
rect 3221 3776 3237 3840
rect 3301 3776 3309 3840
rect 2989 2752 3309 3776
rect 2989 2688 2997 2752
rect 3061 2688 3077 2752
rect 3141 2688 3157 2752
rect 3221 2688 3237 2752
rect 3301 2688 3309 2752
rect 2989 1707 3309 2688
rect 2989 1664 3031 1707
rect 3267 1664 3309 1707
rect 2989 1600 2997 1664
rect 3301 1600 3309 1664
rect 2989 1471 3031 1600
rect 3267 1471 3309 1600
rect 2989 576 3309 1471
rect 2989 512 2997 576
rect 3061 512 3077 576
rect 3141 512 3157 576
rect 3221 512 3237 576
rect 3301 512 3309 576
rect 2989 -48 3309 512
rect 6138 9824 6458 9840
rect 6138 9760 6146 9824
rect 6210 9760 6226 9824
rect 6290 9760 6306 9824
rect 6370 9760 6386 9824
rect 6450 9760 6458 9824
rect 6138 8736 6458 9760
rect 6138 8672 6146 8736
rect 6210 8672 6226 8736
rect 6290 8672 6306 8736
rect 6370 8672 6386 8736
rect 6450 8672 6458 8736
rect 6138 7648 6458 8672
rect 6138 7584 6146 7648
rect 6210 7584 6226 7648
rect 6290 7584 6306 7648
rect 6370 7584 6386 7648
rect 6450 7584 6458 7648
rect 6138 6619 6458 7584
rect 6138 6560 6180 6619
rect 6416 6560 6458 6619
rect 6138 6496 6146 6560
rect 6450 6496 6458 6560
rect 6138 6383 6180 6496
rect 6416 6383 6458 6496
rect 6138 5472 6458 6383
rect 6138 5408 6146 5472
rect 6210 5408 6226 5472
rect 6290 5408 6306 5472
rect 6370 5408 6386 5472
rect 6450 5408 6458 5472
rect 6138 4384 6458 5408
rect 6138 4320 6146 4384
rect 6210 4320 6226 4384
rect 6290 4320 6306 4384
rect 6370 4320 6386 4384
rect 6450 4320 6458 4384
rect 6138 3344 6458 4320
rect 6138 3296 6180 3344
rect 6416 3296 6458 3344
rect 6138 3232 6146 3296
rect 6450 3232 6458 3296
rect 6138 3108 6180 3232
rect 6416 3108 6458 3232
rect 6138 2208 6458 3108
rect 6138 2144 6146 2208
rect 6210 2144 6226 2208
rect 6290 2144 6306 2208
rect 6370 2144 6386 2208
rect 6450 2144 6458 2208
rect 6138 1120 6458 2144
rect 6138 1056 6146 1120
rect 6210 1056 6226 1120
rect 6290 1056 6306 1120
rect 6370 1056 6386 1120
rect 6450 1056 6458 1120
rect 6138 32 6458 1056
rect 6138 -32 6146 32
rect 6210 -32 6226 32
rect 6290 -32 6306 32
rect 6370 -32 6386 32
rect 6450 -32 6458 32
rect 6138 -48 6458 -32
rect 9287 9280 9608 9840
rect 9287 9216 9296 9280
rect 9360 9216 9376 9280
rect 9440 9216 9456 9280
rect 9520 9216 9536 9280
rect 9600 9216 9608 9280
rect 9287 8256 9608 9216
rect 9287 8192 9330 8256
rect 9566 8192 9608 8256
rect 9287 8128 9296 8192
rect 9600 8128 9608 8192
rect 9287 8020 9330 8128
rect 9566 8020 9608 8128
rect 9287 7104 9608 8020
rect 9287 7040 9296 7104
rect 9360 7040 9376 7104
rect 9440 7040 9456 7104
rect 9520 7040 9536 7104
rect 9600 7040 9608 7104
rect 9287 6016 9608 7040
rect 9287 5952 9296 6016
rect 9360 5952 9376 6016
rect 9440 5952 9456 6016
rect 9520 5952 9536 6016
rect 9600 5952 9608 6016
rect 9287 4982 9608 5952
rect 9287 4928 9330 4982
rect 9566 4928 9608 4982
rect 9287 4864 9296 4928
rect 9600 4864 9608 4928
rect 9287 4746 9330 4864
rect 9566 4746 9608 4864
rect 9287 3840 9608 4746
rect 9287 3776 9296 3840
rect 9360 3776 9376 3840
rect 9440 3776 9456 3840
rect 9520 3776 9536 3840
rect 9600 3776 9608 3840
rect 9287 2752 9608 3776
rect 9287 2688 9296 2752
rect 9360 2688 9376 2752
rect 9440 2688 9456 2752
rect 9520 2688 9536 2752
rect 9600 2688 9608 2752
rect 9287 1707 9608 2688
rect 9287 1664 9330 1707
rect 9566 1664 9608 1707
rect 9287 1600 9296 1664
rect 9600 1600 9608 1664
rect 9287 1471 9330 1600
rect 9566 1471 9608 1600
rect 9287 576 9608 1471
rect 9287 512 9296 576
rect 9360 512 9376 576
rect 9440 512 9456 576
rect 9520 512 9536 576
rect 9600 512 9608 576
rect 9287 -48 9608 512
rect 12437 9824 12757 9840
rect 12437 9760 12445 9824
rect 12509 9760 12525 9824
rect 12589 9760 12605 9824
rect 12669 9760 12685 9824
rect 12749 9760 12757 9824
rect 12437 8736 12757 9760
rect 12437 8672 12445 8736
rect 12509 8672 12525 8736
rect 12589 8672 12605 8736
rect 12669 8672 12685 8736
rect 12749 8672 12757 8736
rect 12437 7648 12757 8672
rect 12437 7584 12445 7648
rect 12509 7584 12525 7648
rect 12589 7584 12605 7648
rect 12669 7584 12685 7648
rect 12749 7584 12757 7648
rect 12437 6619 12757 7584
rect 12437 6560 12479 6619
rect 12715 6560 12757 6619
rect 12437 6496 12445 6560
rect 12749 6496 12757 6560
rect 12437 6383 12479 6496
rect 12715 6383 12757 6496
rect 12437 5472 12757 6383
rect 12437 5408 12445 5472
rect 12509 5408 12525 5472
rect 12589 5408 12605 5472
rect 12669 5408 12685 5472
rect 12749 5408 12757 5472
rect 12437 4384 12757 5408
rect 12437 4320 12445 4384
rect 12509 4320 12525 4384
rect 12589 4320 12605 4384
rect 12669 4320 12685 4384
rect 12749 4320 12757 4384
rect 12437 3344 12757 4320
rect 12437 3296 12479 3344
rect 12715 3296 12757 3344
rect 12437 3232 12445 3296
rect 12749 3232 12757 3296
rect 12437 3108 12479 3232
rect 12715 3108 12757 3232
rect 12437 2208 12757 3108
rect 12437 2144 12445 2208
rect 12509 2144 12525 2208
rect 12589 2144 12605 2208
rect 12669 2144 12685 2208
rect 12749 2144 12757 2208
rect 12437 1120 12757 2144
rect 12437 1056 12445 1120
rect 12509 1056 12525 1120
rect 12589 1056 12605 1120
rect 12669 1056 12685 1120
rect 12749 1056 12757 1120
rect 12437 32 12757 1056
rect 12437 -32 12445 32
rect 12509 -32 12525 32
rect 12589 -32 12605 32
rect 12669 -32 12685 32
rect 12749 -32 12757 32
rect 12437 -48 12757 -32
rect 15586 9280 15906 9840
rect 15586 9216 15594 9280
rect 15658 9216 15674 9280
rect 15738 9216 15754 9280
rect 15818 9216 15834 9280
rect 15898 9216 15906 9280
rect 15586 8256 15906 9216
rect 15586 8192 15628 8256
rect 15864 8192 15906 8256
rect 15586 8128 15594 8192
rect 15898 8128 15906 8192
rect 15586 8020 15628 8128
rect 15864 8020 15906 8128
rect 15586 7104 15906 8020
rect 15586 7040 15594 7104
rect 15658 7040 15674 7104
rect 15738 7040 15754 7104
rect 15818 7040 15834 7104
rect 15898 7040 15906 7104
rect 15586 6016 15906 7040
rect 15586 5952 15594 6016
rect 15658 5952 15674 6016
rect 15738 5952 15754 6016
rect 15818 5952 15834 6016
rect 15898 5952 15906 6016
rect 15586 4982 15906 5952
rect 15586 4928 15628 4982
rect 15864 4928 15906 4982
rect 15586 4864 15594 4928
rect 15898 4864 15906 4928
rect 15586 4746 15628 4864
rect 15864 4746 15906 4864
rect 15586 3840 15906 4746
rect 15586 3776 15594 3840
rect 15658 3776 15674 3840
rect 15738 3776 15754 3840
rect 15818 3776 15834 3840
rect 15898 3776 15906 3840
rect 15586 2752 15906 3776
rect 15586 2688 15594 2752
rect 15658 2688 15674 2752
rect 15738 2688 15754 2752
rect 15818 2688 15834 2752
rect 15898 2688 15906 2752
rect 15586 1707 15906 2688
rect 15586 1664 15628 1707
rect 15864 1664 15906 1707
rect 15586 1600 15594 1664
rect 15898 1600 15906 1664
rect 15586 1471 15628 1600
rect 15864 1471 15906 1600
rect 15586 576 15906 1471
rect 15586 512 15594 576
rect 15658 512 15674 576
rect 15738 512 15754 576
rect 15818 512 15834 576
rect 15898 512 15906 576
rect 15586 -48 15906 512
<< via4 >>
rect 3031 8192 3267 8256
rect 3031 8128 3061 8192
rect 3061 8128 3077 8192
rect 3077 8128 3141 8192
rect 3141 8128 3157 8192
rect 3157 8128 3221 8192
rect 3221 8128 3237 8192
rect 3237 8128 3267 8192
rect 3031 8020 3267 8128
rect 3031 4928 3267 4982
rect 3031 4864 3061 4928
rect 3061 4864 3077 4928
rect 3077 4864 3141 4928
rect 3141 4864 3157 4928
rect 3157 4864 3221 4928
rect 3221 4864 3237 4928
rect 3237 4864 3267 4928
rect 3031 4746 3267 4864
rect 3031 1664 3267 1707
rect 3031 1600 3061 1664
rect 3061 1600 3077 1664
rect 3077 1600 3141 1664
rect 3141 1600 3157 1664
rect 3157 1600 3221 1664
rect 3221 1600 3237 1664
rect 3237 1600 3267 1664
rect 3031 1471 3267 1600
rect 6180 6560 6416 6619
rect 6180 6496 6210 6560
rect 6210 6496 6226 6560
rect 6226 6496 6290 6560
rect 6290 6496 6306 6560
rect 6306 6496 6370 6560
rect 6370 6496 6386 6560
rect 6386 6496 6416 6560
rect 6180 6383 6416 6496
rect 6180 3296 6416 3344
rect 6180 3232 6210 3296
rect 6210 3232 6226 3296
rect 6226 3232 6290 3296
rect 6290 3232 6306 3296
rect 6306 3232 6370 3296
rect 6370 3232 6386 3296
rect 6386 3232 6416 3296
rect 6180 3108 6416 3232
rect 9330 8192 9566 8256
rect 9330 8128 9360 8192
rect 9360 8128 9376 8192
rect 9376 8128 9440 8192
rect 9440 8128 9456 8192
rect 9456 8128 9520 8192
rect 9520 8128 9536 8192
rect 9536 8128 9566 8192
rect 9330 8020 9566 8128
rect 9330 4928 9566 4982
rect 9330 4864 9360 4928
rect 9360 4864 9376 4928
rect 9376 4864 9440 4928
rect 9440 4864 9456 4928
rect 9456 4864 9520 4928
rect 9520 4864 9536 4928
rect 9536 4864 9566 4928
rect 9330 4746 9566 4864
rect 9330 1664 9566 1707
rect 9330 1600 9360 1664
rect 9360 1600 9376 1664
rect 9376 1600 9440 1664
rect 9440 1600 9456 1664
rect 9456 1600 9520 1664
rect 9520 1600 9536 1664
rect 9536 1600 9566 1664
rect 9330 1471 9566 1600
rect 12479 6560 12715 6619
rect 12479 6496 12509 6560
rect 12509 6496 12525 6560
rect 12525 6496 12589 6560
rect 12589 6496 12605 6560
rect 12605 6496 12669 6560
rect 12669 6496 12685 6560
rect 12685 6496 12715 6560
rect 12479 6383 12715 6496
rect 12479 3296 12715 3344
rect 12479 3232 12509 3296
rect 12509 3232 12525 3296
rect 12525 3232 12589 3296
rect 12589 3232 12605 3296
rect 12605 3232 12669 3296
rect 12669 3232 12685 3296
rect 12685 3232 12715 3296
rect 12479 3108 12715 3232
rect 15628 8192 15864 8256
rect 15628 8128 15658 8192
rect 15658 8128 15674 8192
rect 15674 8128 15738 8192
rect 15738 8128 15754 8192
rect 15754 8128 15818 8192
rect 15818 8128 15834 8192
rect 15834 8128 15864 8192
rect 15628 8020 15864 8128
rect 15628 4928 15864 4982
rect 15628 4864 15658 4928
rect 15658 4864 15674 4928
rect 15674 4864 15738 4928
rect 15738 4864 15754 4928
rect 15754 4864 15818 4928
rect 15818 4864 15834 4928
rect 15834 4864 15864 4928
rect 15628 4746 15864 4864
rect 15628 1664 15864 1707
rect 15628 1600 15658 1664
rect 15658 1600 15674 1664
rect 15674 1600 15738 1664
rect 15738 1600 15754 1664
rect 15754 1600 15818 1664
rect 15818 1600 15834 1664
rect 15834 1600 15864 1664
rect 15628 1471 15864 1600
<< metal5 >>
rect 0 8256 18860 8298
rect 0 8020 3031 8256
rect 3267 8020 9330 8256
rect 9566 8020 15628 8256
rect 15864 8020 18860 8256
rect 0 7978 18860 8020
rect 0 6619 18860 6661
rect 0 6383 6180 6619
rect 6416 6383 12479 6619
rect 12715 6383 18860 6619
rect 0 6341 18860 6383
rect 0 4982 18860 5024
rect 0 4746 3031 4982
rect 3267 4746 9330 4982
rect 9566 4746 15628 4982
rect 15864 4746 18860 4982
rect 0 4704 18860 4746
rect 0 3344 18860 3386
rect 0 3108 6180 3344
rect 6416 3108 12479 3344
rect 12715 3108 18860 3344
rect 0 3066 18860 3108
rect 0 1707 18860 1749
rect 0 1471 3031 1707
rect 3267 1471 9330 1707
rect 9566 1471 15628 1707
rect 15864 1471 18860 1707
rect 0 1429 18860 1471
use sky130_fd_sc_hd__decap_12  FILLER_0_15 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1380 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1636915332
transform 1 0 276 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1636915332
transform 1 0 1380 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1636915332
transform 1 0 276 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 0 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1636915332
transform 1 0 0 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2484 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 1636915332
transform 1 0 2668 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 1636915332
transform 1 0 3772 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1636915332
transform 1 0 2484 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1636915332
transform 1 0 3588 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2576 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1636915332
transform 1 0 5152 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1636915332
transform 1 0 5152 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_57 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5244 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1636915332
transform 1 0 5060 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 4692 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1636915332
transform 1 0 4876 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _338_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 6256 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334__6 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 6532 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_65
timestamp 1636915332
transform 1 0 5980 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69
timestamp 1636915332
transform 1 0 6348 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__dfstp_1  _441_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 6808 0 -1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57
timestamp 1636915332
transform 1 0 5244 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 7084 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1636915332
transform 1 0 7544 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 7820 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_95
timestamp 1636915332
transform 1 0 8740 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1636915332
transform 1 0 7728 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _312_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 8832 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp 1636915332
transform -1 0 7544 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _442_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 8372 0 1 0
box -38 -48 1878 592
use sky130_fd_sc_hd__o21ai_1  _336_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 9568 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _333_
timestamp 1636915332
transform -1 0 9568 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1636915332
transform -1 0 10212 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1636915332
transform 1 0 10212 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1636915332
transform 1 0 10212 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _357_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 10396 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _356_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 11040 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _355_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 11960 0 -1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_2  _308_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 10396 0 -1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1636915332
transform 1 0 10304 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1636915332
transform 1 0 10304 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_123
timestamp 1636915332
transform 1 0 11316 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_135
timestamp 1636915332
transform 1 0 12420 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1636915332
transform 1 0 12788 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1636915332
transform 1 0 12972 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_130
timestamp 1636915332
transform 1 0 11960 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1636915332
transform 1 0 12880 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _453_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 13892 0 -1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_0_153
timestamp 1636915332
transform 1 0 14076 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1636915332
transform 1 0 15180 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_169
timestamp 1636915332
transform 1 0 15548 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_151
timestamp 1636915332
transform 1 0 13892 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1636915332
transform 1 0 15272 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1636915332
transform 1 0 15456 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1636915332
transform 1 0 15456 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _360_
timestamp 1636915332
transform 1 0 14996 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _452_
timestamp 1636915332
transform 1 0 15548 0 -1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_0_181
timestamp 1636915332
transform 1 0 16652 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp 1636915332
transform 1 0 17572 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1636915332
transform 1 0 17940 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1636915332
transform 1 0 18124 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1636915332
transform 1 0 18032 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  _359_
timestamp 1636915332
transform 1 0 16928 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _404_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 17480 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1636915332
transform -1 0 18860 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1636915332
transform -1 0 18860 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1636915332
transform 1 0 18308 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 18308 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1636915332
transform 1 0 1380 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1636915332
transform 1 0 276 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1636915332
transform 1 0 0 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1636915332
transform 1 0 2484 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1636915332
transform 1 0 2668 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1636915332
transform 1 0 3772 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1636915332
transform 1 0 2576 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_53
timestamp 1636915332
transform 1 0 4876 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtn_1  _440_
timestamp 1636915332
transform 1 0 5428 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1636915332
transform 1 0 7636 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1636915332
transform 1 0 7728 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _311_
timestamp 1636915332
transform 1 0 8740 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _331_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 7820 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _339_
timestamp 1636915332
transform -1 0 7636 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _407_
timestamp 1636915332
transform 1 0 9016 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _381_
timestamp 1636915332
transform 1 0 10672 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _382_
timestamp 1636915332
transform 1 0 9844 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_2_134
timestamp 1636915332
transform 1 0 12328 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1636915332
transform 1 0 12972 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1636915332
transform 1 0 12880 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _406_
timestamp 1636915332
transform 1 0 11500 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_153
timestamp 1636915332
transform 1 0 14076 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_168
timestamp 1636915332
transform 1 0 15456 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _275_
timestamp 1636915332
transform -1 0 15456 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _276_
timestamp 1636915332
transform -1 0 15180 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _290_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 15640 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _361_
timestamp 1636915332
transform 1 0 14168 0 1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_2_197
timestamp 1636915332
transform 1 0 18124 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1636915332
transform 1 0 18032 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _401_
timestamp 1636915332
transform 1 0 17204 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _405_
timestamp 1636915332
transform 1 0 16376 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_201
timestamp 1636915332
transform 1 0 18492 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1636915332
transform -1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1636915332
transform 1 0 1380 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1636915332
transform 1 0 276 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1636915332
transform 1 0 0 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_27
timestamp 1636915332
transform 1 0 2484 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_35
timestamp 1636915332
transform 1 0 3220 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtn_1  _448_
timestamp 1636915332
transform 1 0 3312 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_3_69
timestamp 1636915332
transform 1 0 6348 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1636915332
transform 1 0 5152 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _293_
timestamp 1636915332
transform 1 0 5796 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1636915332
transform -1 0 6348 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _302_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 5796 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _386_
timestamp 1636915332
transform 1 0 6440 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _286_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 8556 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _309_
timestamp 1636915332
transform -1 0 8924 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _316_
timestamp 1636915332
transform -1 0 9292 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _385_
timestamp 1636915332
transform 1 0 7268 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_107
timestamp 1636915332
transform 1 0 9844 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1636915332
transform 1 0 10212 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1636915332
transform 1 0 10396 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_122
timestamp 1636915332
transform 1 0 11224 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1636915332
transform 1 0 10304 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_2  _282_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 11224 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _283_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 11316 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _332_
timestamp 1636915332
transform 1 0 9292 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _335_
timestamp 1636915332
transform -1 0 9844 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_127
timestamp 1636915332
transform 1 0 11684 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_145
timestamp 1636915332
transform 1 0 13340 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _287_
timestamp 1636915332
transform 1 0 12236 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _288_
timestamp 1636915332
transform 1 0 12604 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _399_
timestamp 1636915332
transform 1 0 13432 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1636915332
transform 1 0 15364 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1636915332
transform 1 0 15456 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _274_
timestamp 1636915332
transform 1 0 14260 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _289_
timestamp 1636915332
transform -1 0 15916 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _398_
timestamp 1636915332
transform 1 0 14536 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _402_
timestamp 1636915332
transform 1 0 15916 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_1  _427_
timestamp 1636915332
transform -1 0 18584 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1636915332
transform -1 0 18860 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1636915332
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1636915332
transform 1 0 276 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1636915332
transform 1 0 0 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1636915332
transform 1 0 2484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1636915332
transform 1 0 2668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_41
timestamp 1636915332
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_49
timestamp 1636915332
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1636915332
transform 1 0 2576 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_58
timestamp 1636915332
transform 1 0 5336 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_71
timestamp 1636915332
transform 1 0 6532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1636915332
transform -1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _295_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5428 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _296_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5980 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _304_
timestamp 1636915332
transform -1 0 5336 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_75
timestamp 1636915332
transform 1 0 6900 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1636915332
transform 1 0 7728 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _281_
timestamp 1636915332
transform 1 0 8648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _314_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 9568 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _330_
timestamp 1636915332
transform 1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _397_
timestamp 1636915332
transform 1 0 7820 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_110
timestamp 1636915332
transform 1 0 10120 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_114
timestamp 1636915332
transform 1 0 10488 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__o21bai_1  _315_
timestamp 1636915332
transform -1 0 10120 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__dfstp_1  _454_
timestamp 1636915332
transform 1 0 10580 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_4_136
timestamp 1636915332
transform 1 0 12512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1636915332
transform 1 0 12880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1636915332
transform 1 0 12604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _279_
timestamp 1636915332
transform 1 0 12972 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _285_
timestamp 1636915332
transform -1 0 13892 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_151
timestamp 1636915332
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _443_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 13984 0 1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1636915332
transform 1 0 18032 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _358_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_2  _451_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 16100 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_4_201
timestamp 1636915332
transform 1 0 18492 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1636915332
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1636915332
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1636915332
transform 1 0 276 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1636915332
transform 1 0 0 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_27
timestamp 1636915332
transform 1 0 2484 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dfstp_1  _449_
timestamp 1636915332
transform 1 0 3220 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_5_73
timestamp 1636915332
transform 1 0 6716 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1636915332
transform 1 0 5152 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1636915332
transform 1 0 6164 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1636915332
transform -1 0 5520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _299_
timestamp 1636915332
transform 1 0 6440 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2ai_1  _300_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 6164 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _313_
timestamp 1636915332
transform 1 0 6808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_77
timestamp 1636915332
transform 1 0 7084 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_85
timestamp 1636915332
transform 1 0 7820 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_89
timestamp 1636915332
transform 1 0 8188 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  _306_
timestamp 1636915332
transform 1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _447_
timestamp 1636915332
transform 1 0 8372 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_5_116
timestamp 1636915332
transform 1 0 10672 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1636915332
transform 1 0 10304 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1636915332
transform -1 0 10672 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_128
timestamp 1636915332
transform 1 0 11776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_136
timestamp 1636915332
transform 1 0 12512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _278_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 12880 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _284_
timestamp 1636915332
transform 1 0 13432 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _349_
timestamp 1636915332
transform 1 0 11868 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_5_152
timestamp 1636915332
transform 1 0 13984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_160
timestamp 1636915332
transform 1 0 14720 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_169
timestamp 1636915332
transform 1 0 15548 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1636915332
transform 1 0 15456 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _291_
timestamp 1636915332
transform 1 0 15088 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _292_
timestamp 1636915332
transform 1 0 15640 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _329_
timestamp 1636915332
transform 1 0 14168 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1636915332
transform 1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _428_
timestamp 1636915332
transform -1 0 18308 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1636915332
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1636915332
transform 1 0 18308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1636915332
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1636915332
transform 1 0 276 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1636915332
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1636915332
transform 1 0 276 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1636915332
transform 1 0 0 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1636915332
transform 1 0 0 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1636915332
transform 1 0 2484 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_29
timestamp 1636915332
transform 1 0 2668 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_35
timestamp 1636915332
transform 1 0 3220 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_39
timestamp 1636915332
transform 1 0 3588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1636915332
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1636915332
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1636915332
transform 1 0 2576 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _301__4
timestamp 1636915332
transform -1 0 3588 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_51
timestamp 1636915332
transform 1 0 4692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1636915332
transform 1 0 4692 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1636915332
transform 1 0 5060 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1636915332
transform 1 0 5244 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_72
timestamp 1636915332
transform 1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1636915332
transform 1 0 5152 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _303_
timestamp 1636915332
transform -1 0 5428 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _320_
timestamp 1636915332
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _450_
timestamp 1636915332
transform 1 0 5428 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_6_79
timestamp 1636915332
transform 1 0 7268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1636915332
transform 1 0 7636 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1636915332
transform 1 0 7728 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _319_
timestamp 1636915332
transform 1 0 6900 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _321_
timestamp 1636915332
transform 1 0 8004 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _322_
timestamp 1636915332
transform -1 0 8004 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_2  _444_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 7820 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_pll_clk
timestamp 1636915332
transform -1 0 9200 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _400_
timestamp 1636915332
transform 1 0 9292 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _305__5
timestamp 1636915332
transform -1 0 10028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1636915332
transform 1 0 10120 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_100
timestamp 1636915332
transform 1 0 9200 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_109
timestamp 1636915332
transform 1 0 10028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _364_
timestamp 1636915332
transform -1 0 11684 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _362_
timestamp 1636915332
transform -1 0 11316 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _341_
timestamp 1636915332
transform 1 0 10396 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1636915332
transform 1 0 10304 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_123
timestamp 1636915332
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _416_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 10304 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_127
timestamp 1636915332
transform 1 0 11684 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1636915332
transform 1 0 12880 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _326_
timestamp 1636915332
transform 1 0 12604 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _327_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 11776 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _328_
timestamp 1636915332
transform 1 0 12236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_2  _350_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 11868 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_2  _351_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 12972 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _415_
timestamp 1636915332
transform 1 0 12512 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_6_150
timestamp 1636915332
transform 1 0 13800 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_166
timestamp 1636915332
transform 1 0 15272 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_172
timestamp 1636915332
transform 1 0 15824 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1636915332
transform 1 0 15456 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _323_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 14352 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _325_
timestamp 1636915332
transform -1 0 15272 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _414_
timestamp 1636915332
transform 1 0 13984 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_4  _430_
timestamp 1636915332
transform 1 0 15916 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _432_
timestamp 1636915332
transform -1 0 17664 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_6_197
timestamp 1636915332
transform 1 0 18124 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_192
timestamp 1636915332
transform 1 0 17664 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_198
timestamp 1636915332
transform 1 0 18216 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1636915332
transform 1 0 18032 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_201
timestamp 1636915332
transform 1 0 18492 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1636915332
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1636915332
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1636915332
transform 1 0 18308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1636915332
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1636915332
transform 1 0 276 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1636915332
transform 1 0 0 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1636915332
transform 1 0 2484 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1636915332
transform 1 0 2668 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1636915332
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1636915332
transform 1 0 2576 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_53
timestamp 1636915332
transform 1 0 4876 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_61
timestamp 1636915332
transform 1 0 5612 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_1  _445_
timestamp 1636915332
transform 1 0 5796 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1636915332
transform 1 0 7636 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_89
timestamp 1636915332
transform 1 0 8188 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1636915332
transform 1 0 7728 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_1  _317_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 8188 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _363_
timestamp 1636915332
transform 1 0 8280 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _403_
timestamp 1636915332
transform 1 0 8924 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_pll_clk OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 11592 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1636915332
transform 1 0 12880 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _273_
timestamp 1636915332
transform -1 0 12880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _342_
timestamp 1636915332
transform -1 0 12236 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _411_
timestamp 1636915332
transform 1 0 12972 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_pll_clk
timestamp 1636915332
transform 1 0 12236 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1636915332
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _324_
timestamp 1636915332
transform 1 0 14352 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _348_
timestamp 1636915332
transform 1 0 13800 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _352_
timestamp 1636915332
transform 1 0 14904 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _377_
timestamp 1636915332
transform 1 0 15180 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dfstp_4  _431_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 18032 0 1 4352
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1636915332
transform 1 0 18124 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1636915332
transform 1 0 18032 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1636915332
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1636915332
transform 1 0 18308 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1636915332
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1636915332
transform 1 0 276 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1636915332
transform 1 0 0 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_27
timestamp 1636915332
transform 1 0 2484 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_33
timestamp 1636915332
transform 1 0 3036 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _457_
timestamp 1636915332
transform 1 0 3128 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1636915332
transform 1 0 5060 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1636915332
transform 1 0 5244 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_61
timestamp 1636915332
transform 1 0 5612 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_69
timestamp 1636915332
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1636915332
transform 1 0 5152 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _367_
timestamp 1636915332
transform 1 0 5704 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_9_77
timestamp 1636915332
transform 1 0 7084 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _318_
timestamp 1636915332
transform 1 0 7360 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _446_
timestamp 1636915332
transform -1 0 9844 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_9_107
timestamp 1636915332
transform 1 0 9844 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_119
timestamp 1636915332
transform 1 0 10948 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1636915332
transform 1 0 10304 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _208_
timestamp 1636915332
transform -1 0 10948 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _210_
timestamp 1636915332
transform 1 0 9936 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _439_
timestamp 1636915332
transform 1 0 11132 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_9_145
timestamp 1636915332
transform 1 0 13340 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1636915332
transform 1 0 13064 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _429_
timestamp 1636915332
transform 1 0 13524 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1636915332
transform 1 0 15364 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_169
timestamp 1636915332
transform 1 0 15548 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1636915332
transform 1 0 15456 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  _373_
timestamp 1636915332
transform 1 0 16100 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _470_
timestamp 1636915332
transform 1 0 16744 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1636915332
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1636915332
transform 1 0 276 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_7
timestamp 1636915332
transform 1 0 644 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1636915332
transform 1 0 0 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _458_
timestamp 1636915332
transform 1 0 736 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_10_29
timestamp 1636915332
transform 1 0 2668 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_33
timestamp 1636915332
transform 1 0 3036 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_38
timestamp 1636915332
transform 1 0 3496 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_49
timestamp 1636915332
transform 1 0 4508 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1636915332
transform 1 0 2576 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1636915332
transform -1 0 4508 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _261_
timestamp 1636915332
transform -1 0 3496 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _262__3
timestamp 1636915332
transform -1 0 4232 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _264_
timestamp 1636915332
transform 1 0 3588 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_70
timestamp 1636915332
transform 1 0 6440 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__nor3b_2  _249_
timestamp 1636915332
transform -1 0 5520 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_1  _365_
timestamp 1636915332
transform 1 0 5796 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _366_
timestamp 1636915332
transform -1 0 5796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _408_
timestamp 1636915332
transform 1 0 6624 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_10_81
timestamp 1636915332
transform 1 0 7452 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1636915332
transform 1 0 7728 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _340_
timestamp 1636915332
transform -1 0 8096 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _418_
timestamp 1636915332
transform 1 0 8096 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _417_
timestamp 1636915332
transform -1 0 11040 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _424_
timestamp 1636915332
transform 1 0 11040 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_10_141
timestamp 1636915332
transform 1 0 12972 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_148
timestamp 1636915332
transform 1 0 13616 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1636915332
transform 1 0 12880 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _205_
timestamp 1636915332
transform -1 0 13984 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _271_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 13064 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_172
timestamp 1636915332
transform 1 0 15824 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_1  _376_
timestamp 1636915332
transform -1 0 16284 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _469_
timestamp 1636915332
transform 1 0 13984 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1636915332
transform 1 0 18124 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1636915332
transform 1 0 18032 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__nor3b_2  _268_
timestamp 1636915332
transform 1 0 16284 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _410_
timestamp 1636915332
transform 1 0 17204 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1636915332
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1636915332
transform 1 0 18308 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1636915332
transform 1 0 276 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1636915332
transform 1 0 0 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _456_
timestamp 1636915332
transform 1 0 1380 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__nand3_1  _253_
timestamp 1636915332
transform 1 0 3496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _260_
timestamp 1636915332
transform -1 0 3496 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _384_
timestamp 1636915332
transform 1 0 3864 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1636915332
transform 1 0 4968 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_60
timestamp 1636915332
transform 1 0 5520 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1636915332
transform 1 0 5152 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1636915332
transform -1 0 4968 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _263_
timestamp 1636915332
transform -1 0 5520 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _395_
timestamp 1636915332
transform 1 0 6440 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _396_
timestamp 1636915332
transform 1 0 5612 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_11_79
timestamp 1636915332
transform 1 0 7268 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_85
timestamp 1636915332
transform 1 0 7820 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_89
timestamp 1636915332
transform 1 0 8188 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _246__2
timestamp 1636915332
transform -1 0 8188 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1636915332
transform -1 0 8556 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _419_
timestamp 1636915332
transform 1 0 8556 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1636915332
transform 1 0 10304 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _209_
timestamp 1636915332
transform -1 0 10948 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _211_
timestamp 1636915332
transform -1 0 10304 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _218_
timestamp 1636915332
transform -1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_125
timestamp 1636915332
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__and2_1  _212_
timestamp 1636915332
transform 1 0 11684 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__dfstp_1  _455_
timestamp 1636915332
transform 1 0 12144 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_11_157
timestamp 1636915332
transform 1 0 14444 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1636915332
transform 1 0 15456 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _204_
timestamp 1636915332
transform 1 0 14628 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_1  _468_
timestamp 1636915332
transform 1 0 15548 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_pll_clk90
timestamp 1636915332
transform 1 0 14076 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _387_
timestamp 1636915332
transform 1 0 17480 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1636915332
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1636915332
transform 1 0 18308 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1636915332
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1636915332
transform 1 0 276 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1636915332
transform 1 0 0 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1636915332
transform 1 0 2484 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_29
timestamp 1636915332
transform 1 0 2668 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1636915332
transform 1 0 2576 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _259_
timestamp 1636915332
transform 1 0 3956 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1636915332
transform -1 0 3956 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _266_
timestamp 1636915332
transform 1 0 3036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _267_
timestamp 1636915332
transform -1 0 3680 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_62
timestamp 1636915332
transform 1 0 5704 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o21bai_1  _256_
timestamp 1636915332
transform -1 0 6348 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _383_
timestamp 1636915332
transform 1 0 4876 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _409_
timestamp 1636915332
transform 1 0 6348 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1636915332
transform 1 0 7544 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1636915332
transform 1 0 7728 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _250_
timestamp 1636915332
transform -1 0 7544 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _459_
timestamp 1636915332
transform 1 0 7820 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_12_106
timestamp 1636915332
transform 1 0 9752 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _467_
timestamp 1636915332
transform -1 0 11960 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1636915332
transform 1 0 12880 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _213_
timestamp 1636915332
transform -1 0 12512 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _214_
timestamp 1636915332
transform -1 0 12880 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _412_
timestamp 1636915332
transform -1 0 13800 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_163
timestamp 1636915332
transform 1 0 14996 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _272_
timestamp 1636915332
transform 1 0 14628 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _413_
timestamp 1636915332
transform 1 0 13800 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_2  _437_
timestamp 1636915332
transform -1 0 17020 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1636915332
transform 1 0 17848 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1636915332
transform 1 0 18032 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _206_
timestamp 1636915332
transform 1 0 17020 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_2  _372_
timestamp 1636915332
transform 1 0 18124 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_201
timestamp 1636915332
transform 1 0 18492 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1636915332
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1636915332
transform 1 0 276 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_15
timestamp 1636915332
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1636915332
transform 1 0 276 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1636915332
transform 1 0 0 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1636915332
transform 1 0 0 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _240_
timestamp 1636915332
transform 1 0 1748 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _244_
timestamp 1636915332
transform 1 0 2024 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtn_1  _462_
timestamp 1636915332
transform 1 0 552 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__nor2_1  _254_
timestamp 1636915332
transform -1 0 3036 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2ai_1  _241_
timestamp 1636915332
transform 1 0 2668 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1636915332
transform -1 0 2760 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1636915332
transform 1 0 2576 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1636915332
transform 1 0 2392 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_26
timestamp 1636915332
transform 1 0 2392 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__and2b_1  _243_
timestamp 1636915332
transform -1 0 4048 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _236_
timestamp 1636915332
transform 1 0 3312 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_37
timestamp 1636915332
transform 1 0 3404 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_33
timestamp 1636915332
transform 1 0 3036 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _237_
timestamp 1636915332
transform -1 0 4416 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_48
timestamp 1636915332
transform 1 0 4416 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_44
timestamp 1636915332
transform 1 0 4048 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _390_
timestamp 1636915332
transform 1 0 5060 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _258_
timestamp 1636915332
transform 1 0 4876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _255_
timestamp 1636915332
transform -1 0 5980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _247_
timestamp 1636915332
transform 1 0 4784 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _216_
timestamp 1636915332
transform -1 0 4876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1636915332
transform 1 0 5152 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1636915332
transform 1 0 5244 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  _225_
timestamp 1636915332
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _224_
timestamp 1636915332
transform 1 0 5980 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _217_
timestamp 1636915332
transform 1 0 5888 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _215_
timestamp 1636915332
transform -1 0 6716 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _257_
timestamp 1636915332
transform 1 0 6716 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_73
timestamp 1636915332
transform 1 0 6716 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_pll_clk90
timestamp 1636915332
transform -1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _233_
timestamp 1636915332
transform -1 0 7728 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1636915332
transform 1 0 7728 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_81
timestamp 1636915332
transform 1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _380_
timestamp 1636915332
transform 1 0 7912 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _379_
timestamp 1636915332
transform 1 0 8464 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_1  _232_
timestamp 1636915332
transform -1 0 8188 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_89
timestamp 1636915332
transform 1 0 8188 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_85
timestamp 1636915332
transform 1 0 7820 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _368_
timestamp 1636915332
transform -1 0 9108 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _230_
timestamp 1636915332
transform 1 0 9108 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_101
timestamp 1636915332
transform 1 0 9292 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1636915332
transform 1 0 10304 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _343_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 11316 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _369_
timestamp 1636915332
transform -1 0 11868 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _391_
timestamp 1636915332
transform 1 0 10396 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _392_
timestamp 1636915332
transform 1 0 9476 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_pll_clk90
timestamp 1636915332
transform -1 0 11316 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_13_129
timestamp 1636915332
transform 1 0 11868 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1636915332
transform 1 0 12880 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _394_
timestamp 1636915332
transform 1 0 12972 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_1  _466_
timestamp 1636915332
transform 1 0 11960 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 12144 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1636915332
transform 1 0 15364 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_154
timestamp 1636915332
transform 1 0 14168 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1636915332
transform 1 0 15456 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _227_
timestamp 1636915332
transform -1 0 14168 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _353_
timestamp 1636915332
transform -1 0 16192 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2ai_2  _354_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 13892 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dfstp_1  _434_
timestamp 1636915332
transform 1 0 14260 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_ext_clk
timestamp 1636915332
transform -1 0 15364 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_176
timestamp 1636915332
transform 1 0 16192 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1636915332
transform 1 0 18124 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1636915332
transform 1 0 18032 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _433_
timestamp 1636915332
transform 1 0 16192 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _436_
timestamp 1636915332
transform -1 0 18492 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_1  FILLER_13_201
timestamp 1636915332
transform 1 0 18492 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1636915332
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1636915332
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1636915332
transform 1 0 18308 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1636915332
transform 1 0 276 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1636915332
transform 1 0 0 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _461_
timestamp 1636915332
transform 1 0 368 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_15_28
timestamp 1636915332
transform 1 0 2576 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_46
timestamp 1636915332
transform 1 0 4232 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _234_
timestamp 1636915332
transform -1 0 3956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1636915332
transform -1 0 4232 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1636915332
transform -1 0 2576 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _245_
timestamp 1636915332
transform -1 0 3680 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1636915332
transform 1 0 4968 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1636915332
transform 1 0 5244 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1636915332
transform 1 0 5152 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _228_
timestamp 1636915332
transform 1 0 5428 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _229_
timestamp 1636915332
transform 1 0 5796 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _389_
timestamp 1636915332
transform 1 0 6532 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_15_80
timestamp 1636915332
transform 1 0 7360 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _370_
timestamp 1636915332
transform 1 0 8924 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _388_
timestamp 1636915332
transform 1 0 8096 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_100
timestamp 1636915332
transform 1 0 9200 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1636915332
transform 1 0 10396 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1636915332
transform 1 0 10304 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_1  _231_
timestamp 1636915332
transform -1 0 10028 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1636915332
transform -1 0 10304 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _420_
timestamp 1636915332
transform 1 0 10488 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__nand3b_1  _223_
timestamp 1636915332
transform 1 0 11960 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ext_clk
timestamp 1636915332
transform 1 0 12512 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_15_156
timestamp 1636915332
transform 1 0 14352 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1636915332
transform 1 0 15364 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_172
timestamp 1636915332
transform 1 0 15824 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1636915332
transform 1 0 15456 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _207_
timestamp 1636915332
transform -1 0 15824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _393_
timestamp 1636915332
transform 1 0 14536 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_178
timestamp 1636915332
transform 1 0 16376 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _438_
timestamp 1636915332
transform 1 0 16468 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1636915332
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_20
timestamp 1636915332
transform 1 0 1840 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1636915332
transform 1 0 276 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_8
timestamp 1636915332
transform 1 0 736 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1636915332
transform 1 0 0 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _242__1
timestamp 1636915332
transform -1 0 736 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_49
timestamp 1636915332
transform 1 0 4508 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1636915332
transform 1 0 2576 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtn_1  _460_
timestamp 1636915332
transform 1 0 2668 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _465_
timestamp 1636915332
transform -1 0 7084 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1636915332
transform 1 0 7084 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1636915332
transform 1 0 7636 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1636915332
transform 1 0 7728 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _371_
timestamp 1636915332
transform 1 0 7820 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__dfstp_1  _464_
timestamp 1636915332
transform 1 0 8464 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_16_113
timestamp 1636915332
transform 1 0 10396 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o21bai_1  _226_
timestamp 1636915332
transform -1 0 11040 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _435_
timestamp 1636915332
transform -1 0 12880 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1636915332
transform 1 0 12880 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _425_
timestamp 1636915332
transform 1 0 12972 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1636915332
transform -1 0 15088 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _422_
timestamp 1636915332
transform 1 0 15088 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_8  FILLER_16_185
timestamp 1636915332
transform 1 0 17020 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1636915332
transform 1 0 18124 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1636915332
transform 1 0 18032 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1636915332
transform 1 0 17756 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1636915332
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1636915332
transform 1 0 18308 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_11
timestamp 1636915332
transform 1 0 1012 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1636915332
transform 1 0 276 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1636915332
transform 1 0 0 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  input3 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1104 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_17_29
timestamp 1636915332
transform 1 0 2668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_41
timestamp 1636915332
transform 1 0 3772 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1636915332
transform 1 0 2576 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1636915332
transform 1 0 4876 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_57
timestamp 1636915332
transform 1 0 5244 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1636915332
transform 1 0 5152 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _463_
timestamp 1636915332
transform 1 0 5796 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_17_88
timestamp 1636915332
transform 1 0 8096 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_17_97
timestamp 1636915332
transform 1 0 8924 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1636915332
transform 1 0 7728 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _219_
timestamp 1636915332
transform 1 0 8648 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output10
timestamp 1636915332
transform 1 0 7820 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1636915332
transform 1 0 10120 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1636915332
transform 1 0 10304 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1636915332
transform -1 0 10120 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _221_
timestamp 1636915332
transform -1 0 9844 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _344_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 10396 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _426_
timestamp 1636915332
transform 1 0 11040 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_ext_clk
timestamp 1636915332
transform 1 0 10672 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output12
timestamp 1636915332
transform -1 0 9476 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_145
timestamp 1636915332
transform 1 0 13340 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1636915332
transform 1 0 12880 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _423_
timestamp 1636915332
transform 1 0 13524 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  output11 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 13340 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_172
timestamp 1636915332
transform 1 0 15824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1636915332
transform 1 0 15456 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _378__13 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 15824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1636915332
transform 1 0 18032 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _375_
timestamp 1636915332
transform 1 0 18124 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _421_
timestamp 1636915332
transform 1 0 16100 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_17_200
timestamp 1636915332
transform 1 0 18400 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1636915332
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
<< labels >>
rlabel metal5 s 0 3066 18860 3386 6 VGND
port 0 nsew ground input
rlabel metal5 s 0 6341 18860 6661 6 VGND
port 0 nsew ground input
rlabel metal4 s 6138 -48 6458 9840 6 VGND
port 0 nsew ground input
rlabel metal4 s 12437 -48 12757 9840 6 VGND
port 0 nsew ground input
rlabel metal5 s 0 1429 18860 1749 6 VPWR
port 1 nsew power input
rlabel metal5 s 0 4704 18860 5024 6 VPWR
port 1 nsew power input
rlabel metal5 s 0 7978 18860 8298 6 VPWR
port 1 nsew power input
rlabel metal4 s 2989 -48 3309 9840 6 VPWR
port 1 nsew power input
rlabel metal4 s 9287 -48 9607 9840 6 VPWR
port 1 nsew power input
rlabel metal4 s 15586 -48 15906 9840 6 VPWR
port 1 nsew power input
rlabel metal2 s 7102 11200 7158 12000 6 core_clk
port 2 nsew signal tristate
rlabel metal2 s 4250 11200 4306 12000 6 ext_clk
port 3 nsew signal input
rlabel metal3 s 19200 688 20000 808 6 ext_clk_sel
port 4 nsew signal input
rlabel metal3 s 19200 11160 20000 11280 6 ext_reset
port 5 nsew signal input
rlabel metal2 s 15658 11200 15714 12000 6 pll_clk
port 6 nsew signal input
rlabel metal2 s 18510 11200 18566 12000 6 pll_clk90
port 7 nsew signal input
rlabel metal2 s 1398 11200 1454 12000 6 resetb
port 8 nsew signal input
rlabel metal2 s 12806 11200 12862 12000 6 resetb_sync
port 9 nsew signal tristate
rlabel metal3 s 19200 6672 20000 6792 6 sel2[0]
port 10 nsew signal input
rlabel metal3 s 19200 8168 20000 8288 6 sel2[1]
port 11 nsew signal input
rlabel metal3 s 19200 9664 20000 9784 6 sel2[2]
port 12 nsew signal input
rlabel metal3 s 19200 2184 20000 2304 6 sel[0]
port 13 nsew signal input
rlabel metal3 s 19200 3680 20000 3800 6 sel[1]
port 14 nsew signal input
rlabel metal3 s 19200 5176 20000 5296 6 sel[2]
port 15 nsew signal input
rlabel metal2 s 9954 11200 10010 12000 6 user_clk
port 16 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 20000 12000
<< end >>
