magic
tech sky130A
magscale 1 2
timestamp 1637447660
<< error_p >>
rect 30830 218031 31584 218032
rect 30830 216955 30831 218031
rect 31583 216955 31584 218031
rect 30830 216954 31584 216955
rect 37368 216463 38130 216464
rect 37368 215381 37369 216463
rect 38129 215381 38130 216463
rect 37368 215380 38130 215381
<< metal3 >>
rect 6032 221346 55470 221382
rect 6032 221338 54256 221346
rect 6032 220224 6162 221338
rect 6862 220248 54256 221338
rect 55338 220248 55470 221346
rect 6862 220224 55470 220248
rect 6032 220182 55470 220224
rect 7246 219742 53826 219782
rect 7246 218628 7360 219742
rect 8060 219728 53826 219742
rect 8060 218630 52662 219728
rect 53744 218630 53826 219728
rect 8060 218628 53826 218630
rect 7246 218582 53826 218628
rect 17838 218068 31672 218100
rect 17838 216936 17896 218068
rect 18646 218032 31672 218068
rect 18646 216954 30830 218032
rect 31584 216954 31672 218032
rect 18646 216936 31672 216954
rect 17838 216900 31672 216936
rect 19032 216470 38262 216500
rect 19032 215338 19100 216470
rect 19850 216464 38262 216470
rect 19850 215380 37368 216464
rect 38130 215380 38262 216464
rect 19850 215338 38262 215380
rect 19032 215300 38262 215338
<< via3 >>
rect 6162 220224 6862 221338
rect 54256 220248 55338 221346
rect 7360 218628 8060 219742
rect 52662 218630 53744 219728
rect 17896 216936 18646 218068
rect 30830 216954 31584 218032
rect 19100 215338 19850 216470
rect 37368 215380 38130 216464
<< metal4 >>
rect 6116 221338 6916 221470
rect 6116 220224 6162 221338
rect 6862 220224 6916 221338
rect 6116 211884 6916 220224
rect 54194 221346 55400 221388
rect 54194 220248 54256 221346
rect 55338 220248 55400 221346
rect 54194 220174 55400 220248
rect 6116 211606 6126 211884
rect 6898 211606 6916 211884
rect 6116 208518 6916 211606
rect 6116 208240 6130 208518
rect 6906 208240 6916 208518
rect 6116 205138 6916 208240
rect 7316 219742 8116 219842
rect 7316 218628 7360 219742
rect 8060 218628 8116 219742
rect 7316 213586 8116 218628
rect 52590 219728 53796 219788
rect 52590 218630 52662 219728
rect 53744 218630 53796 219728
rect 52590 218574 53796 218630
rect 7316 213288 7328 213586
rect 8102 213288 8116 213586
rect 7316 210196 8116 213288
rect 7316 209918 7330 210196
rect 8102 209918 8116 210196
rect 7316 206826 8116 209918
rect 7316 206528 7326 206826
rect 8100 206528 8116 206826
rect 7316 206476 8116 206528
rect 17880 218068 18680 218110
rect 17880 216936 17896 218068
rect 18646 217338 18680 218068
rect 18656 217056 18680 217338
rect 18646 216936 18680 217056
rect 17880 212534 18680 216936
rect 17880 212246 17896 212534
rect 18668 212246 18680 212534
rect 17880 209152 18680 212246
rect 17880 208864 17890 209152
rect 18662 208864 18680 209152
rect 17880 205770 18680 208864
rect 17880 205482 17892 205770
rect 18664 205482 18680 205770
rect 17880 205422 18680 205482
rect 19080 216634 19880 216732
rect 19080 215338 19100 216634
rect 19856 216352 19880 216634
rect 19850 215338 19880 216352
rect 19080 210844 19880 215338
rect 19080 210556 19092 210844
rect 19864 210556 19880 210844
rect 19080 207464 19880 210556
rect 19080 207176 19096 207464
rect 19868 207176 19880 207464
rect 6116 204840 6132 205138
rect 6906 204840 6916 205138
rect 6116 204746 6916 204840
rect 19080 204084 19880 207176
rect 19080 203796 19096 204084
rect 19868 203796 19880 204084
rect 19080 203748 19880 203796
<< via4 >>
rect 54256 220248 55338 221346
rect 6126 211606 6898 211884
rect 6130 208240 6906 208518
rect 52662 218630 53744 219728
rect 7328 213288 8102 213586
rect 7330 209918 8102 210196
rect 7326 206528 8100 206826
rect 17900 217056 18646 217338
rect 18646 217056 18656 217338
rect 17896 212246 18668 212534
rect 17890 208864 18662 209152
rect 17892 205482 18664 205770
rect 19100 216470 19856 216634
rect 19100 216352 19850 216470
rect 19850 216352 19856 216470
rect 19092 210556 19864 210844
rect 19096 207176 19868 207464
rect 6132 204840 6906 205138
rect 19096 203796 19868 204084
<< metal5 >>
rect 54224 221346 55376 221378
rect 54224 220248 54256 221346
rect 55338 220248 55376 221346
rect 54224 220198 55376 220248
rect 52630 219728 53782 219772
rect 52630 218630 52662 219728
rect 53744 218630 53782 219728
rect 52630 218592 53782 218630
rect 17856 217356 18695 217379
rect 14320 217338 18695 217356
rect 14320 217056 17900 217338
rect 18656 217056 18695 217338
rect 14320 217036 18695 217056
rect 17856 217018 18695 217036
rect 19062 216656 19901 216670
rect 14320 216634 19932 216656
rect 14320 216352 19100 216634
rect 19856 216352 19932 216634
rect 14320 216336 19932 216352
rect 19062 216309 19901 216336
rect 7289 213598 8128 213619
rect 7270 213586 8592 213598
rect 7270 213288 7328 213586
rect 8102 213288 8592 213586
rect 7270 213278 8592 213288
rect 7289 213258 8128 213278
rect 17859 212550 18701 212568
rect 17434 212534 18718 212550
rect 17434 212246 17896 212534
rect 18668 212246 18718 212534
rect 17434 212230 18718 212246
rect 17859 212208 18701 212230
rect 6098 211908 6937 211940
rect 6058 211884 8592 211908
rect 6058 211606 6126 211884
rect 6898 211606 8592 211884
rect 6058 211588 8592 211606
rect 6098 211579 6937 211588
rect 19066 210860 19908 210873
rect 17434 210844 19910 210860
rect 17434 210556 19092 210844
rect 19864 210556 19910 210844
rect 17434 210540 19910 210556
rect 19066 210524 19908 210540
rect 7307 210218 8146 210241
rect 7276 210196 8592 210218
rect 7276 209918 7330 210196
rect 8102 209918 8592 210196
rect 7276 209898 8592 209918
rect 7307 209880 8146 209898
rect 17867 209170 18709 209178
rect 17434 209152 18709 209170
rect 17434 208864 17890 209152
rect 18662 208864 18709 209152
rect 17434 208850 18709 208864
rect 17867 208829 18709 208850
rect 6044 208528 6939 208554
rect 6044 208518 8592 208528
rect 6044 208240 6130 208518
rect 6906 208240 8592 208518
rect 6044 208208 8592 208240
rect 6044 208206 6939 208208
rect 19063 207480 19905 207495
rect 17434 207464 19910 207480
rect 17434 207176 19096 207464
rect 19868 207176 19910 207464
rect 17434 207160 19910 207176
rect 19063 207146 19905 207160
rect 7287 206838 8182 206853
rect 7287 206826 8624 206838
rect 7287 206528 7326 206826
rect 8100 206528 8624 206826
rect 7287 206518 8624 206528
rect 7287 206502 8182 206518
rect 17863 205790 18705 205805
rect 17434 205770 18712 205790
rect 17434 205482 17892 205770
rect 18664 205482 18712 205770
rect 17434 205470 18712 205482
rect 17863 205456 18705 205470
rect 6095 205148 6990 205170
rect 6095 205138 8624 205148
rect 6095 204840 6132 205138
rect 6906 204840 8624 205138
rect 6095 204828 8624 204840
rect 6095 204808 6990 204828
rect 19072 204100 19914 204115
rect 17434 204084 19914 204100
rect 17434 203796 19096 204084
rect 19868 203796 19914 204084
rect 17434 203780 19914 203796
rect 19072 203766 19914 203780
<< end >>
