magic
tech sky130A
magscale 1 2
timestamp 1648835380
<< metal1 >>
rect 146938 1007088 146944 1007140
rect 146996 1007128 147002 1007140
rect 154574 1007128 154580 1007140
rect 146996 1007100 154580 1007128
rect 146996 1007088 147002 1007100
rect 154574 1007088 154580 1007100
rect 154632 1007088 154638 1007140
rect 195422 1006952 195428 1007004
rect 195480 1006992 195486 1007004
rect 203886 1006992 203892 1007004
rect 195480 1006964 203892 1006992
rect 195480 1006952 195486 1006964
rect 203886 1006952 203892 1006964
rect 203944 1006952 203950 1007004
rect 300302 1006952 300308 1007004
rect 300360 1006992 300366 1007004
rect 308950 1006992 308956 1007004
rect 300360 1006964 308956 1006992
rect 300360 1006952 300366 1006964
rect 308950 1006952 308956 1006964
rect 309008 1006952 309014 1007004
rect 426342 1006884 426348 1006936
rect 426400 1006924 426406 1006936
rect 429562 1006924 429568 1006936
rect 426400 1006896 429568 1006924
rect 426400 1006884 426406 1006896
rect 429562 1006884 429568 1006896
rect 429620 1006884 429626 1006936
rect 261018 1006816 261024 1006868
rect 261076 1006856 261082 1006868
rect 268378 1006856 268384 1006868
rect 261076 1006828 268384 1006856
rect 261076 1006816 261082 1006828
rect 268378 1006816 268384 1006828
rect 268436 1006816 268442 1006868
rect 427170 1006816 427176 1006868
rect 427228 1006856 427234 1006868
rect 440878 1006856 440884 1006868
rect 427228 1006828 440884 1006856
rect 427228 1006816 427234 1006828
rect 440878 1006816 440884 1006828
rect 440936 1006816 440942 1006868
rect 425146 1006748 425152 1006800
rect 425204 1006788 425210 1006800
rect 469858 1006788 469864 1006800
rect 425204 1006760 469864 1006788
rect 425204 1006748 425210 1006760
rect 469858 1006748 469864 1006760
rect 469916 1006748 469922 1006800
rect 427538 1006680 427544 1006732
rect 427596 1006720 427602 1006732
rect 443638 1006720 443644 1006732
rect 427596 1006692 443644 1006720
rect 427596 1006680 427602 1006692
rect 443638 1006680 443644 1006692
rect 443696 1006680 443702 1006732
rect 427998 1006612 428004 1006664
rect 428056 1006652 428062 1006664
rect 448606 1006652 448612 1006664
rect 428056 1006624 448612 1006652
rect 428056 1006612 428062 1006624
rect 448606 1006612 448612 1006624
rect 448664 1006612 448670 1006664
rect 197998 1006544 198004 1006596
rect 198056 1006584 198062 1006596
rect 203518 1006584 203524 1006596
rect 198056 1006556 203524 1006584
rect 198056 1006544 198062 1006556
rect 203518 1006544 203524 1006556
rect 203576 1006544 203582 1006596
rect 429562 1006544 429568 1006596
rect 429620 1006584 429626 1006596
rect 441614 1006584 441620 1006596
rect 429620 1006556 441620 1006584
rect 429620 1006544 429626 1006556
rect 441614 1006544 441620 1006556
rect 441672 1006544 441678 1006596
rect 95878 1006476 95884 1006528
rect 95936 1006516 95942 1006528
rect 103606 1006516 103612 1006528
rect 95936 1006488 103612 1006516
rect 95936 1006476 95942 1006488
rect 103606 1006476 103612 1006488
rect 103664 1006476 103670 1006528
rect 145742 1006476 145748 1006528
rect 145800 1006516 145806 1006528
rect 145800 1006488 151814 1006516
rect 145800 1006476 145806 1006488
rect 94498 1006408 94504 1006460
rect 94556 1006448 94562 1006460
rect 103146 1006448 103152 1006460
rect 94556 1006420 103152 1006448
rect 94556 1006408 94562 1006420
rect 103146 1006408 103152 1006420
rect 103204 1006408 103210 1006460
rect 144178 1006408 144184 1006460
rect 144236 1006448 144242 1006460
rect 151630 1006448 151636 1006460
rect 144236 1006420 151636 1006448
rect 144236 1006408 144242 1006420
rect 151630 1006408 151636 1006420
rect 151688 1006408 151694 1006460
rect 151786 1006448 151814 1006488
rect 423490 1006476 423496 1006528
rect 423548 1006516 423554 1006528
rect 446398 1006516 446404 1006528
rect 423548 1006488 446404 1006516
rect 423548 1006476 423554 1006488
rect 446398 1006476 446404 1006488
rect 446456 1006476 446462 1006528
rect 154114 1006448 154120 1006460
rect 151786 1006420 154120 1006448
rect 154114 1006408 154120 1006420
rect 154172 1006408 154178 1006460
rect 428458 1006408 428464 1006460
rect 428516 1006448 428522 1006460
rect 457438 1006448 457444 1006460
rect 428516 1006420 457444 1006448
rect 428516 1006408 428522 1006420
rect 457438 1006408 457444 1006420
rect 457496 1006408 457502 1006460
rect 508682 1006408 508688 1006460
rect 508740 1006448 508746 1006460
rect 515398 1006448 515404 1006460
rect 508740 1006420 515404 1006448
rect 508740 1006408 508746 1006420
rect 515398 1006408 515404 1006420
rect 515456 1006408 515462 1006460
rect 100110 1006340 100116 1006392
rect 100168 1006380 100174 1006392
rect 104342 1006380 104348 1006392
rect 100168 1006352 104348 1006380
rect 100168 1006340 100174 1006352
rect 104342 1006340 104348 1006352
rect 104400 1006340 104406 1006392
rect 150434 1006340 150440 1006392
rect 150492 1006380 150498 1006392
rect 177298 1006380 177304 1006392
rect 150492 1006352 177304 1006380
rect 150492 1006340 150498 1006352
rect 177298 1006340 177304 1006352
rect 177356 1006340 177362 1006392
rect 253308 1006352 267734 1006380
rect 93302 1006272 93308 1006324
rect 93360 1006312 93366 1006324
rect 100662 1006312 100668 1006324
rect 93360 1006284 100668 1006312
rect 93360 1006272 93366 1006284
rect 100662 1006272 100668 1006284
rect 100720 1006272 100726 1006324
rect 108850 1006312 108856 1006324
rect 103486 1006284 108856 1006312
rect 93118 1006204 93124 1006256
rect 93176 1006244 93182 1006256
rect 101950 1006244 101956 1006256
rect 93176 1006216 101956 1006244
rect 93176 1006204 93182 1006216
rect 101950 1006204 101956 1006216
rect 102008 1006204 102014 1006256
rect 102778 1006204 102784 1006256
rect 102836 1006244 102842 1006256
rect 103486 1006244 103514 1006284
rect 108850 1006272 108856 1006284
rect 108908 1006272 108914 1006324
rect 195146 1006272 195152 1006324
rect 195204 1006312 195210 1006324
rect 204714 1006312 204720 1006324
rect 195204 1006284 204720 1006312
rect 195204 1006272 195210 1006284
rect 204714 1006272 204720 1006284
rect 204772 1006272 204778 1006324
rect 228358 1006312 228364 1006324
rect 205652 1006284 228364 1006312
rect 102836 1006216 103514 1006244
rect 102836 1006204 102842 1006216
rect 108482 1006204 108488 1006256
rect 108540 1006244 108546 1006256
rect 113818 1006244 113824 1006256
rect 108540 1006216 113824 1006244
rect 108540 1006204 108546 1006216
rect 113818 1006204 113824 1006216
rect 113876 1006204 113882 1006256
rect 97258 1006136 97264 1006188
rect 97316 1006176 97322 1006188
rect 104802 1006176 104808 1006188
rect 97316 1006148 104808 1006176
rect 97316 1006136 97322 1006148
rect 104802 1006136 104808 1006148
rect 104860 1006136 104866 1006188
rect 145558 1006136 145564 1006188
rect 145616 1006176 145622 1006188
rect 156138 1006176 156144 1006188
rect 145616 1006148 156144 1006176
rect 145616 1006136 145622 1006148
rect 156138 1006136 156144 1006148
rect 156196 1006136 156202 1006188
rect 196618 1006136 196624 1006188
rect 196676 1006176 196682 1006188
rect 205542 1006176 205548 1006188
rect 196676 1006148 205548 1006176
rect 196676 1006136 196682 1006148
rect 205542 1006136 205548 1006148
rect 205600 1006136 205606 1006188
rect 98270 1006068 98276 1006120
rect 98328 1006108 98334 1006120
rect 99098 1006108 99104 1006120
rect 98328 1006080 99104 1006108
rect 98328 1006068 98334 1006080
rect 99098 1006068 99104 1006080
rect 99156 1006068 99162 1006120
rect 149698 1006068 149704 1006120
rect 149756 1006108 149762 1006120
rect 150434 1006108 150440 1006120
rect 149756 1006080 150440 1006108
rect 149756 1006068 149762 1006080
rect 150434 1006068 150440 1006080
rect 150492 1006068 150498 1006120
rect 157426 1006108 157432 1006120
rect 151786 1006080 157432 1006108
rect 99116 1006040 99144 1006068
rect 126238 1006040 126244 1006052
rect 99116 1006012 126244 1006040
rect 126238 1006000 126244 1006012
rect 126296 1006000 126302 1006052
rect 145650 1006000 145656 1006052
rect 145708 1006040 145714 1006052
rect 151786 1006040 151814 1006080
rect 157426 1006068 157432 1006080
rect 157484 1006068 157490 1006120
rect 159082 1006068 159088 1006120
rect 159140 1006108 159146 1006120
rect 166258 1006108 166264 1006120
rect 159140 1006080 166264 1006108
rect 159140 1006068 159146 1006080
rect 166258 1006068 166264 1006080
rect 166316 1006068 166322 1006120
rect 195238 1006068 195244 1006120
rect 195296 1006108 195302 1006120
rect 204346 1006108 204352 1006120
rect 195296 1006080 204352 1006108
rect 195296 1006068 195302 1006080
rect 204346 1006068 204352 1006080
rect 204404 1006068 204410 1006120
rect 205652 1006108 205680 1006284
rect 228358 1006272 228364 1006284
rect 228416 1006272 228422 1006324
rect 253308 1006256 253336 1006352
rect 254670 1006272 254676 1006324
rect 254728 1006312 254734 1006324
rect 258166 1006312 258172 1006324
rect 254728 1006284 258172 1006312
rect 254728 1006272 254734 1006284
rect 258166 1006272 258172 1006284
rect 258224 1006272 258230 1006324
rect 267706 1006312 267734 1006352
rect 301498 1006340 301504 1006392
rect 301556 1006380 301562 1006392
rect 310146 1006380 310152 1006392
rect 301556 1006352 310152 1006380
rect 301556 1006340 301562 1006352
rect 310146 1006340 310152 1006352
rect 310204 1006340 310210 1006392
rect 425974 1006340 425980 1006392
rect 426032 1006380 426038 1006392
rect 451918 1006380 451924 1006392
rect 426032 1006352 451924 1006380
rect 426032 1006340 426038 1006352
rect 451918 1006340 451924 1006352
rect 451976 1006340 451982 1006392
rect 551922 1006340 551928 1006392
rect 551980 1006380 551986 1006392
rect 574738 1006380 574744 1006392
rect 551980 1006352 574744 1006380
rect 551980 1006340 551986 1006352
rect 574738 1006340 574744 1006352
rect 574796 1006340 574802 1006392
rect 280798 1006312 280804 1006324
rect 267706 1006284 280804 1006312
rect 280798 1006272 280804 1006284
rect 280856 1006272 280862 1006324
rect 300210 1006272 300216 1006324
rect 300268 1006312 300274 1006324
rect 308122 1006312 308128 1006324
rect 300268 1006284 308128 1006312
rect 300268 1006272 300274 1006284
rect 308122 1006272 308128 1006284
rect 308180 1006272 308186 1006324
rect 423858 1006272 423864 1006324
rect 423916 1006312 423922 1006324
rect 454678 1006312 454684 1006324
rect 423916 1006284 454684 1006312
rect 423916 1006272 423922 1006284
rect 454678 1006272 454684 1006284
rect 454736 1006272 454742 1006324
rect 501322 1006272 501328 1006324
rect 501380 1006312 501386 1006324
rect 517514 1006312 517520 1006324
rect 501380 1006284 517520 1006312
rect 501380 1006272 501386 1006284
rect 517514 1006272 517520 1006284
rect 517572 1006272 517578 1006324
rect 553946 1006272 553952 1006324
rect 554004 1006312 554010 1006324
rect 563790 1006312 563796 1006324
rect 554004 1006284 563796 1006312
rect 554004 1006272 554010 1006284
rect 563790 1006272 563796 1006284
rect 563848 1006272 563854 1006324
rect 252462 1006204 252468 1006256
rect 252520 1006244 252526 1006256
rect 253290 1006244 253296 1006256
rect 252520 1006216 253296 1006244
rect 252520 1006204 252526 1006216
rect 253290 1006204 253296 1006216
rect 253348 1006204 253354 1006256
rect 300118 1006204 300124 1006256
rect 300176 1006244 300182 1006256
rect 300176 1006216 306374 1006244
rect 300176 1006204 300182 1006216
rect 250438 1006136 250444 1006188
rect 250496 1006176 250502 1006188
rect 256510 1006176 256516 1006188
rect 250496 1006148 256516 1006176
rect 250496 1006136 250502 1006148
rect 256510 1006136 256516 1006148
rect 256568 1006136 256574 1006188
rect 298738 1006136 298744 1006188
rect 298796 1006176 298802 1006188
rect 306098 1006176 306104 1006188
rect 298796 1006148 306104 1006176
rect 298796 1006136 298802 1006148
rect 306098 1006136 306104 1006148
rect 306156 1006136 306162 1006188
rect 204824 1006080 205680 1006108
rect 145708 1006012 151814 1006040
rect 145708 1006000 145714 1006012
rect 154482 1006000 154488 1006052
rect 154540 1006040 154546 1006052
rect 160646 1006040 160652 1006052
rect 154540 1006012 160652 1006040
rect 154540 1006000 154546 1006012
rect 160646 1006000 160652 1006012
rect 160704 1006000 160710 1006052
rect 201034 1006000 201040 1006052
rect 201092 1006040 201098 1006052
rect 201862 1006040 201868 1006052
rect 201092 1006012 201868 1006040
rect 201092 1006000 201098 1006012
rect 201862 1006000 201868 1006012
rect 201920 1006040 201926 1006052
rect 204824 1006040 204852 1006080
rect 209590 1006068 209596 1006120
rect 209648 1006108 209654 1006120
rect 216030 1006108 216036 1006120
rect 209648 1006080 216036 1006108
rect 209648 1006068 209654 1006080
rect 216030 1006068 216036 1006080
rect 216088 1006068 216094 1006120
rect 247678 1006068 247684 1006120
rect 247736 1006108 247742 1006120
rect 258534 1006108 258540 1006120
rect 247736 1006080 258540 1006108
rect 247736 1006068 247742 1006080
rect 258534 1006068 258540 1006080
rect 258592 1006068 258598 1006120
rect 263042 1006068 263048 1006120
rect 263100 1006108 263106 1006120
rect 269758 1006108 269764 1006120
rect 263100 1006080 269764 1006108
rect 263100 1006068 263106 1006080
rect 269758 1006068 269764 1006080
rect 269816 1006068 269822 1006120
rect 298922 1006068 298928 1006120
rect 298980 1006108 298986 1006120
rect 305638 1006108 305644 1006120
rect 298980 1006080 305644 1006108
rect 298980 1006068 298986 1006080
rect 305638 1006068 305644 1006080
rect 305696 1006068 305702 1006120
rect 201920 1006012 204852 1006040
rect 201920 1006000 201926 1006012
rect 204898 1006000 204904 1006052
rect 204956 1006040 204962 1006052
rect 208762 1006040 208768 1006052
rect 204956 1006012 208768 1006040
rect 204956 1006000 204962 1006012
rect 208762 1006000 208768 1006012
rect 208820 1006000 208826 1006052
rect 249058 1006000 249064 1006052
rect 249116 1006040 249122 1006052
rect 255314 1006040 255320 1006052
rect 249116 1006012 255320 1006040
rect 249116 1006000 249122 1006012
rect 255314 1006000 255320 1006012
rect 255372 1006000 255378 1006052
rect 257338 1006000 257344 1006052
rect 257396 1006040 257402 1006052
rect 258994 1006040 259000 1006052
rect 257396 1006012 259000 1006040
rect 257396 1006000 257402 1006012
rect 258994 1006000 259000 1006012
rect 259052 1006000 259058 1006052
rect 262674 1006000 262680 1006052
rect 262732 1006040 262738 1006052
rect 268470 1006040 268476 1006052
rect 262732 1006012 268476 1006040
rect 262732 1006000 262738 1006012
rect 268470 1006000 268476 1006012
rect 268528 1006000 268534 1006052
rect 303522 1006000 303528 1006052
rect 303580 1006040 303586 1006052
rect 304074 1006040 304080 1006052
rect 303580 1006012 304080 1006040
rect 303580 1006000 303586 1006012
rect 304074 1006000 304080 1006012
rect 304132 1006040 304138 1006052
rect 304902 1006040 304908 1006052
rect 304132 1006012 304908 1006040
rect 304132 1006000 304138 1006012
rect 304902 1006000 304908 1006012
rect 304960 1006000 304966 1006052
rect 306346 1006040 306374 1006216
rect 357342 1006204 357348 1006256
rect 357400 1006244 357406 1006256
rect 374638 1006244 374644 1006256
rect 357400 1006216 374644 1006244
rect 357400 1006204 357406 1006216
rect 374638 1006204 374644 1006216
rect 374696 1006204 374702 1006256
rect 430022 1006204 430028 1006256
rect 430080 1006244 430086 1006256
rect 468478 1006244 468484 1006256
rect 430080 1006216 468484 1006244
rect 430080 1006204 430086 1006216
rect 468478 1006204 468484 1006216
rect 468536 1006204 468542 1006256
rect 505830 1006204 505836 1006256
rect 505888 1006244 505894 1006256
rect 514754 1006244 514760 1006256
rect 505888 1006216 514760 1006244
rect 505888 1006204 505894 1006216
rect 514754 1006204 514760 1006216
rect 514812 1006204 514818 1006256
rect 555970 1006204 555976 1006256
rect 556028 1006244 556034 1006256
rect 570598 1006244 570604 1006256
rect 556028 1006216 570604 1006244
rect 556028 1006204 556034 1006216
rect 570598 1006204 570604 1006216
rect 570656 1006204 570662 1006256
rect 361390 1006136 361396 1006188
rect 361448 1006176 361454 1006188
rect 369210 1006176 369216 1006188
rect 361448 1006148 369216 1006176
rect 361448 1006136 361454 1006148
rect 369210 1006136 369216 1006148
rect 369268 1006136 369274 1006188
rect 424686 1006136 424692 1006188
rect 424744 1006176 424750 1006188
rect 460198 1006176 460204 1006188
rect 424744 1006148 460204 1006176
rect 424744 1006136 424750 1006148
rect 460198 1006136 460204 1006148
rect 460256 1006136 460262 1006188
rect 520826 1006176 520832 1006188
rect 508240 1006148 520832 1006176
rect 358538 1006068 358544 1006120
rect 358596 1006108 358602 1006120
rect 371878 1006108 371884 1006120
rect 358596 1006080 371884 1006108
rect 358596 1006068 358602 1006080
rect 371878 1006068 371884 1006080
rect 371936 1006068 371942 1006120
rect 425514 1006068 425520 1006120
rect 425572 1006108 425578 1006120
rect 464982 1006108 464988 1006120
rect 425572 1006080 464988 1006108
rect 425572 1006068 425578 1006080
rect 464982 1006068 464988 1006080
rect 465040 1006068 465046 1006120
rect 498102 1006068 498108 1006120
rect 498160 1006108 498166 1006120
rect 499666 1006108 499672 1006120
rect 498160 1006080 499672 1006108
rect 498160 1006068 498166 1006080
rect 499666 1006068 499672 1006080
rect 499724 1006068 499730 1006120
rect 504542 1006068 504548 1006120
rect 504600 1006108 504606 1006120
rect 508240 1006108 508268 1006148
rect 520826 1006136 520832 1006148
rect 520884 1006136 520890 1006188
rect 557166 1006136 557172 1006188
rect 557224 1006176 557230 1006188
rect 557224 1006148 560708 1006176
rect 557224 1006136 557230 1006148
rect 522298 1006108 522304 1006120
rect 504600 1006080 508268 1006108
rect 514726 1006080 522304 1006108
rect 504600 1006068 504606 1006080
rect 306466 1006040 306472 1006052
rect 306346 1006012 306472 1006040
rect 306466 1006000 306472 1006012
rect 306524 1006000 306530 1006052
rect 307018 1006000 307024 1006052
rect 307076 1006040 307082 1006052
rect 310606 1006040 310612 1006052
rect 307076 1006012 310612 1006040
rect 307076 1006000 307082 1006012
rect 310606 1006000 310612 1006012
rect 310664 1006000 310670 1006052
rect 314654 1006000 314660 1006052
rect 314712 1006040 314718 1006052
rect 330478 1006040 330484 1006052
rect 314712 1006012 330484 1006040
rect 314712 1006000 314718 1006012
rect 330478 1006000 330484 1006012
rect 330536 1006000 330542 1006052
rect 353110 1006000 353116 1006052
rect 353168 1006040 353174 1006052
rect 354490 1006040 354496 1006052
rect 353168 1006012 354496 1006040
rect 353168 1006000 353174 1006012
rect 354490 1006000 354496 1006012
rect 354548 1006000 354554 1006052
rect 356054 1006000 356060 1006052
rect 356112 1006040 356118 1006052
rect 360838 1006040 360844 1006052
rect 356112 1006012 360844 1006040
rect 356112 1006000 356118 1006012
rect 360838 1006000 360844 1006012
rect 360896 1006000 360902 1006052
rect 420730 1006000 420736 1006052
rect 420788 1006040 420794 1006052
rect 422662 1006040 422668 1006052
rect 420788 1006012 422668 1006040
rect 420788 1006000 420794 1006012
rect 422662 1006000 422668 1006012
rect 422720 1006000 422726 1006052
rect 505370 1006000 505376 1006052
rect 505428 1006040 505434 1006052
rect 514726 1006040 514754 1006080
rect 522298 1006068 522304 1006080
rect 522356 1006068 522362 1006120
rect 549162 1006068 549168 1006120
rect 549220 1006108 549226 1006120
rect 550266 1006108 550272 1006120
rect 549220 1006080 550272 1006108
rect 549220 1006068 549226 1006080
rect 550266 1006068 550272 1006080
rect 550324 1006108 550330 1006120
rect 551094 1006108 551100 1006120
rect 550324 1006080 551100 1006108
rect 550324 1006068 550330 1006080
rect 551094 1006068 551100 1006080
rect 551152 1006068 551158 1006120
rect 556798 1006068 556804 1006120
rect 556856 1006108 556862 1006120
rect 560680 1006108 560708 1006148
rect 573358 1006108 573364 1006120
rect 556856 1006080 560616 1006108
rect 560680 1006080 573364 1006108
rect 556856 1006068 556862 1006080
rect 505428 1006012 514754 1006040
rect 505428 1006000 505434 1006012
rect 553118 1006000 553124 1006052
rect 553176 1006040 553182 1006052
rect 556706 1006040 556712 1006052
rect 553176 1006012 556712 1006040
rect 553176 1006000 553182 1006012
rect 556706 1006000 556712 1006012
rect 556764 1006000 556770 1006052
rect 560588 1006040 560616 1006080
rect 573358 1006068 573364 1006080
rect 573416 1006068 573422 1006120
rect 563698 1006040 563704 1006052
rect 560588 1006012 563704 1006040
rect 563698 1006000 563704 1006012
rect 563756 1006000 563762 1006052
rect 143718 1005388 143724 1005440
rect 143776 1005428 143782 1005440
rect 152550 1005428 152556 1005440
rect 143776 1005400 152556 1005428
rect 143776 1005388 143782 1005400
rect 152550 1005388 152556 1005400
rect 152608 1005388 152614 1005440
rect 428826 1005388 428832 1005440
rect 428884 1005428 428890 1005440
rect 448514 1005428 448520 1005440
rect 428884 1005400 448520 1005428
rect 428884 1005388 428890 1005400
rect 448514 1005388 448520 1005400
rect 448572 1005388 448578 1005440
rect 360562 1005320 360568 1005372
rect 360620 1005360 360626 1005372
rect 380158 1005360 380164 1005372
rect 360620 1005332 380164 1005360
rect 360620 1005320 360626 1005332
rect 380158 1005320 380164 1005332
rect 380216 1005320 380222 1005372
rect 432874 1005320 432880 1005372
rect 432932 1005360 432938 1005372
rect 462314 1005360 462320 1005372
rect 432932 1005332 462320 1005360
rect 432932 1005320 432938 1005332
rect 462314 1005320 462320 1005332
rect 462372 1005320 462378 1005372
rect 509878 1005320 509884 1005372
rect 509936 1005360 509942 1005372
rect 520918 1005360 520924 1005372
rect 509936 1005332 520924 1005360
rect 509936 1005320 509942 1005332
rect 520918 1005320 520924 1005332
rect 520976 1005320 520982 1005372
rect 215202 1005252 215208 1005304
rect 215260 1005292 215266 1005304
rect 219434 1005292 219440 1005304
rect 215260 1005264 219440 1005292
rect 215260 1005252 215266 1005264
rect 219434 1005252 219440 1005264
rect 219492 1005252 219498 1005304
rect 356514 1005252 356520 1005304
rect 356572 1005292 356578 1005304
rect 377398 1005292 377404 1005304
rect 356572 1005264 377404 1005292
rect 356572 1005252 356578 1005264
rect 377398 1005252 377404 1005264
rect 377456 1005252 377462 1005304
rect 432506 1005252 432512 1005304
rect 432564 1005292 432570 1005304
rect 467098 1005292 467104 1005304
rect 432564 1005264 467104 1005292
rect 432564 1005252 432570 1005264
rect 467098 1005252 467104 1005264
rect 467156 1005252 467162 1005304
rect 502886 1005252 502892 1005304
rect 502944 1005292 502950 1005304
rect 517606 1005292 517612 1005304
rect 502944 1005264 517612 1005292
rect 502944 1005252 502950 1005264
rect 517606 1005252 517612 1005264
rect 517664 1005252 517670 1005304
rect 564342 1005252 564348 1005304
rect 564400 1005292 564406 1005304
rect 571978 1005292 571984 1005304
rect 564400 1005264 571984 1005292
rect 564400 1005252 564406 1005264
rect 571978 1005252 571984 1005264
rect 572036 1005252 572042 1005304
rect 149698 1004912 149704 1004964
rect 149756 1004952 149762 1004964
rect 152918 1004952 152924 1004964
rect 149756 1004924 152924 1004952
rect 149756 1004912 149762 1004924
rect 152918 1004912 152924 1004924
rect 152976 1004912 152982 1004964
rect 160646 1004912 160652 1004964
rect 160704 1004952 160710 1004964
rect 162854 1004952 162860 1004964
rect 160704 1004924 162860 1004952
rect 160704 1004912 160710 1004924
rect 162854 1004912 162860 1004924
rect 162912 1004912 162918 1004964
rect 208394 1004844 208400 1004896
rect 208452 1004884 208458 1004896
rect 209774 1004884 209780 1004896
rect 208452 1004856 209780 1004884
rect 208452 1004844 208458 1004856
rect 209774 1004844 209780 1004856
rect 209832 1004844 209838 1004896
rect 304442 1004844 304448 1004896
rect 304500 1004884 304506 1004896
rect 307294 1004884 307300 1004896
rect 304500 1004856 307300 1004884
rect 304500 1004844 304506 1004856
rect 307294 1004844 307300 1004856
rect 307352 1004844 307358 1004896
rect 363414 1004844 363420 1004896
rect 363472 1004884 363478 1004896
rect 366358 1004884 366364 1004896
rect 363472 1004856 366364 1004884
rect 363472 1004844 363478 1004856
rect 366358 1004844 366364 1004856
rect 366416 1004844 366422 1004896
rect 151078 1004776 151084 1004828
rect 151136 1004816 151142 1004828
rect 153746 1004816 153752 1004828
rect 151136 1004788 153752 1004816
rect 151136 1004776 151142 1004788
rect 153746 1004776 153752 1004788
rect 153804 1004776 153810 1004828
rect 159450 1004776 159456 1004828
rect 159508 1004816 159514 1004828
rect 161474 1004816 161480 1004828
rect 159508 1004788 161480 1004816
rect 159508 1004776 159514 1004788
rect 161474 1004776 161480 1004788
rect 161532 1004776 161538 1004828
rect 304258 1004776 304264 1004828
rect 304316 1004816 304322 1004828
rect 306926 1004816 306932 1004828
rect 304316 1004788 306932 1004816
rect 304316 1004776 304322 1004788
rect 306926 1004776 306932 1004788
rect 306984 1004776 306990 1004828
rect 361758 1004776 361764 1004828
rect 361816 1004816 361822 1004828
rect 364978 1004816 364984 1004828
rect 361816 1004788 364984 1004816
rect 361816 1004776 361822 1004788
rect 364978 1004776 364984 1004788
rect 365036 1004776 365042 1004828
rect 499206 1004776 499212 1004828
rect 499264 1004816 499270 1004828
rect 501690 1004816 501696 1004828
rect 499264 1004788 501696 1004816
rect 499264 1004776 499270 1004788
rect 501690 1004776 501696 1004788
rect 501748 1004776 501754 1004828
rect 150342 1004708 150348 1004760
rect 150400 1004748 150406 1004760
rect 152090 1004748 152096 1004760
rect 150400 1004720 152096 1004748
rect 150400 1004708 150406 1004720
rect 152090 1004708 152096 1004720
rect 152148 1004708 152154 1004760
rect 160278 1004708 160284 1004760
rect 160336 1004748 160342 1004760
rect 163498 1004748 163504 1004760
rect 160336 1004720 163504 1004748
rect 160336 1004708 160342 1004720
rect 163498 1004708 163504 1004720
rect 163556 1004708 163562 1004760
rect 208762 1004708 208768 1004760
rect 208820 1004748 208826 1004760
rect 211798 1004748 211804 1004760
rect 208820 1004720 211804 1004748
rect 208820 1004708 208826 1004720
rect 211798 1004708 211804 1004720
rect 211856 1004708 211862 1004760
rect 305822 1004708 305828 1004760
rect 305880 1004748 305886 1004760
rect 308582 1004748 308588 1004760
rect 305880 1004720 308588 1004748
rect 305880 1004708 305886 1004720
rect 308582 1004708 308588 1004720
rect 308640 1004708 308646 1004760
rect 364242 1004708 364248 1004760
rect 364300 1004748 364306 1004760
rect 366542 1004748 366548 1004760
rect 364300 1004720 366548 1004748
rect 364300 1004708 364306 1004720
rect 366542 1004708 366548 1004720
rect 366600 1004708 366606 1004760
rect 499482 1004708 499488 1004760
rect 499540 1004748 499546 1004760
rect 499540 1004720 499712 1004748
rect 499540 1004708 499546 1004720
rect 94590 1004640 94596 1004692
rect 94648 1004680 94654 1004692
rect 103146 1004680 103152 1004692
rect 94648 1004652 103152 1004680
rect 94648 1004640 94654 1004652
rect 103146 1004640 103152 1004652
rect 103204 1004640 103210 1004692
rect 151262 1004640 151268 1004692
rect 151320 1004680 151326 1004692
rect 153286 1004680 153292 1004692
rect 151320 1004652 153292 1004680
rect 151320 1004640 151326 1004652
rect 153286 1004640 153292 1004652
rect 153344 1004640 153350 1004692
rect 159818 1004640 159824 1004692
rect 159876 1004680 159882 1004692
rect 162118 1004680 162124 1004692
rect 159876 1004652 162124 1004680
rect 159876 1004640 159882 1004652
rect 162118 1004640 162124 1004652
rect 162176 1004640 162182 1004692
rect 199378 1004640 199384 1004692
rect 199436 1004680 199442 1004692
rect 202322 1004680 202328 1004692
rect 199436 1004652 202328 1004680
rect 199436 1004640 199442 1004652
rect 202322 1004640 202328 1004652
rect 202380 1004640 202386 1004692
rect 305638 1004640 305644 1004692
rect 305696 1004680 305702 1004692
rect 307754 1004680 307760 1004692
rect 305696 1004652 307760 1004680
rect 305696 1004640 305702 1004652
rect 307754 1004640 307760 1004652
rect 307812 1004640 307818 1004692
rect 354582 1004640 354588 1004692
rect 354640 1004680 354646 1004692
rect 354640 1004640 354674 1004680
rect 362586 1004640 362592 1004692
rect 362644 1004680 362650 1004692
rect 365162 1004680 365168 1004692
rect 362644 1004652 365168 1004680
rect 362644 1004640 362650 1004652
rect 365162 1004640 365168 1004652
rect 365220 1004640 365226 1004692
rect 354646 1004612 354674 1004640
rect 356514 1004612 356520 1004624
rect 354646 1004584 356520 1004612
rect 356514 1004572 356520 1004584
rect 356572 1004572 356578 1004624
rect 499684 1004612 499712 1004720
rect 500494 1004708 500500 1004760
rect 500552 1004748 500558 1004760
rect 504358 1004748 504364 1004760
rect 500552 1004720 504364 1004748
rect 500552 1004708 500558 1004720
rect 504358 1004708 504364 1004720
rect 504416 1004708 504422 1004760
rect 556338 1004708 556344 1004760
rect 556396 1004748 556402 1004760
rect 559742 1004748 559748 1004760
rect 556396 1004720 559748 1004748
rect 556396 1004708 556402 1004720
rect 559742 1004708 559748 1004720
rect 559800 1004708 559806 1004760
rect 557626 1004640 557632 1004692
rect 557684 1004680 557690 1004692
rect 559558 1004680 559564 1004692
rect 557684 1004652 559564 1004680
rect 557684 1004640 557690 1004652
rect 559558 1004640 559564 1004652
rect 559616 1004640 559622 1004692
rect 500494 1004612 500500 1004624
rect 499684 1004584 500500 1004612
rect 500494 1004572 500500 1004584
rect 500552 1004572 500558 1004624
rect 499390 1004504 499396 1004556
rect 499448 1004544 499454 1004556
rect 501322 1004544 501328 1004556
rect 499448 1004516 501328 1004544
rect 499448 1004504 499454 1004516
rect 501322 1004504 501328 1004516
rect 501380 1004504 501386 1004556
rect 514754 1004096 514760 1004148
rect 514812 1004136 514818 1004148
rect 517974 1004136 517980 1004148
rect 514812 1004108 517980 1004136
rect 514812 1004096 514818 1004108
rect 517974 1004096 517980 1004108
rect 518032 1004096 518038 1004148
rect 358078 1003892 358084 1003944
rect 358136 1003932 358142 1003944
rect 378318 1003932 378324 1003944
rect 358136 1003904 378324 1003932
rect 358136 1003892 358142 1003904
rect 378318 1003892 378324 1003904
rect 378376 1003892 378382 1003944
rect 448606 1003892 448612 1003944
rect 448664 1003932 448670 1003944
rect 464798 1003932 464804 1003944
rect 448664 1003904 464804 1003932
rect 448664 1003892 448670 1003904
rect 464798 1003892 464804 1003904
rect 464856 1003892 464862 1003944
rect 499482 1003484 499488 1003536
rect 499540 1003524 499546 1003536
rect 500954 1003524 500960 1003536
rect 499540 1003496 500960 1003524
rect 499540 1003484 499546 1003496
rect 500954 1003484 500960 1003496
rect 501012 1003484 501018 1003536
rect 253658 1002640 253664 1002652
rect 246592 1002612 253664 1002640
rect 207198 1002572 207204 1002584
rect 195072 1002544 207204 1002572
rect 106826 1002328 106832 1002380
rect 106884 1002368 106890 1002380
rect 109862 1002368 109868 1002380
rect 106884 1002340 109868 1002368
rect 106884 1002328 106890 1002340
rect 109862 1002328 109868 1002340
rect 109920 1002328 109926 1002380
rect 106182 1002260 106188 1002312
rect 106240 1002300 106246 1002312
rect 108482 1002300 108488 1002312
rect 106240 1002272 108488 1002300
rect 106240 1002260 106246 1002272
rect 108482 1002260 108488 1002272
rect 108540 1002260 108546 1002312
rect 97350 1002192 97356 1002244
rect 97408 1002232 97414 1002244
rect 100294 1002232 100300 1002244
rect 97408 1002204 100300 1002232
rect 97408 1002192 97414 1002204
rect 100294 1002192 100300 1002204
rect 100352 1002192 100358 1002244
rect 105998 1002192 106004 1002244
rect 106056 1002232 106062 1002244
rect 108298 1002232 108304 1002244
rect 106056 1002204 108304 1002232
rect 106056 1002192 106062 1002204
rect 108298 1002192 108304 1002204
rect 108356 1002192 108362 1002244
rect 95970 1002124 95976 1002176
rect 96028 1002164 96034 1002176
rect 99466 1002164 99472 1002176
rect 96028 1002136 99472 1002164
rect 96028 1002124 96034 1002136
rect 99466 1002124 99472 1002136
rect 99524 1002124 99530 1002176
rect 107654 1002124 107660 1002176
rect 107712 1002164 107718 1002176
rect 109678 1002164 109684 1002176
rect 107712 1002136 109684 1002164
rect 107712 1002124 107718 1002136
rect 109678 1002124 109684 1002136
rect 109736 1002124 109742 1002176
rect 158254 1002124 158260 1002176
rect 158312 1002164 158318 1002176
rect 161106 1002164 161112 1002176
rect 158312 1002136 161112 1002164
rect 158312 1002124 158318 1002136
rect 161106 1002124 161112 1002136
rect 161164 1002124 161170 1002176
rect 98822 1002056 98828 1002108
rect 98880 1002096 98886 1002108
rect 101490 1002096 101496 1002108
rect 98880 1002068 101496 1002096
rect 98880 1002056 98886 1002068
rect 101490 1002056 101496 1002068
rect 101548 1002056 101554 1002108
rect 105630 1002056 105636 1002108
rect 105688 1002096 105694 1002108
rect 107746 1002096 107752 1002108
rect 105688 1002068 107752 1002096
rect 105688 1002056 105694 1002068
rect 107746 1002056 107752 1002068
rect 107804 1002056 107810 1002108
rect 144086 1002056 144092 1002108
rect 144144 1002096 144150 1002108
rect 150342 1002096 150348 1002108
rect 144144 1002068 150348 1002096
rect 144144 1002056 144150 1002068
rect 150342 1002056 150348 1002068
rect 150400 1002056 150406 1002108
rect 155770 1002056 155776 1002108
rect 155828 1002096 155834 1002108
rect 157334 1002096 157340 1002108
rect 155828 1002068 157340 1002096
rect 155828 1002056 155834 1002068
rect 157334 1002056 157340 1002068
rect 157392 1002056 157398 1002108
rect 157426 1002056 157432 1002108
rect 157484 1002096 157490 1002108
rect 159358 1002096 159364 1002108
rect 157484 1002068 159364 1002096
rect 157484 1002056 157490 1002068
rect 159358 1002056 159364 1002068
rect 159416 1002056 159422 1002108
rect 98638 1001988 98644 1002040
rect 98696 1002028 98702 1002040
rect 101122 1002028 101128 1002040
rect 98696 1002000 101128 1002028
rect 98696 1001988 98702 1002000
rect 101122 1001988 101128 1002000
rect 101180 1001988 101186 1002040
rect 104342 1001988 104348 1002040
rect 104400 1002028 104406 1002040
rect 106642 1002028 106648 1002040
rect 104400 1002000 106648 1002028
rect 104400 1001988 104406 1002000
rect 106642 1001988 106648 1002000
rect 106700 1001988 106706 1002040
rect 107194 1001988 107200 1002040
rect 107252 1002028 107258 1002040
rect 109034 1002028 109040 1002040
rect 107252 1002000 109040 1002028
rect 107252 1001988 107258 1002000
rect 109034 1001988 109040 1002000
rect 109092 1001988 109098 1002040
rect 148318 1001988 148324 1002040
rect 148376 1002028 148382 1002040
rect 151722 1002028 151728 1002040
rect 148376 1002000 151728 1002028
rect 148376 1001988 148382 1002000
rect 151722 1001988 151728 1002000
rect 151780 1001988 151786 1002040
rect 158622 1001988 158628 1002040
rect 158680 1002028 158686 1002040
rect 160186 1002028 160192 1002040
rect 158680 1002000 160192 1002028
rect 158680 1001988 158686 1002000
rect 160186 1001988 160192 1002000
rect 160244 1001988 160250 1002040
rect 97534 1001920 97540 1001972
rect 97592 1001960 97598 1001972
rect 99926 1001960 99932 1001972
rect 97592 1001932 99932 1001960
rect 97592 1001920 97598 1001932
rect 99926 1001920 99932 1001932
rect 99984 1001920 99990 1001972
rect 100018 1001920 100024 1001972
rect 100076 1001960 100082 1001972
rect 102318 1001960 102324 1001972
rect 100076 1001932 102324 1001960
rect 100076 1001920 100082 1001932
rect 102318 1001920 102324 1001932
rect 102376 1001920 102382 1001972
rect 106458 1001920 106464 1001972
rect 106516 1001960 106522 1001972
rect 107930 1001960 107936 1001972
rect 106516 1001932 107936 1001960
rect 106516 1001920 106522 1001932
rect 107930 1001920 107936 1001932
rect 107988 1001920 107994 1001972
rect 108022 1001920 108028 1001972
rect 108080 1001960 108086 1001972
rect 110506 1001960 110512 1001972
rect 108080 1001932 110512 1001960
rect 108080 1001920 108086 1001932
rect 110506 1001920 110512 1001932
rect 110564 1001920 110570 1001972
rect 148502 1001920 148508 1001972
rect 148560 1001960 148566 1001972
rect 150894 1001960 150900 1001972
rect 148560 1001932 150900 1001960
rect 148560 1001920 148566 1001932
rect 150894 1001920 150900 1001932
rect 150952 1001920 150958 1001972
rect 156966 1001920 156972 1001972
rect 157024 1001960 157030 1001972
rect 158714 1001960 158720 1001972
rect 157024 1001932 158720 1001960
rect 157024 1001920 157030 1001932
rect 158714 1001920 158720 1001932
rect 158772 1001920 158778 1001972
rect 195072 1001620 195100 1002544
rect 207198 1002532 207204 1002544
rect 207256 1002532 207262 1002584
rect 210418 1002192 210424 1002244
rect 210476 1002232 210482 1002244
rect 213178 1002232 213184 1002244
rect 210476 1002204 213184 1002232
rect 210476 1002192 210482 1002204
rect 213178 1002192 213184 1002204
rect 213236 1002192 213242 1002244
rect 210050 1002124 210056 1002176
rect 210108 1002164 210114 1002176
rect 212534 1002164 212540 1002176
rect 210108 1002136 212540 1002164
rect 210108 1002124 210114 1002136
rect 212534 1002124 212540 1002136
rect 212592 1002124 212598 1002176
rect 202138 1002056 202144 1002108
rect 202196 1002096 202202 1002108
rect 205174 1002096 205180 1002108
rect 202196 1002068 205180 1002096
rect 202196 1002056 202202 1002068
rect 205174 1002056 205180 1002068
rect 205232 1002056 205238 1002108
rect 206738 1002056 206744 1002108
rect 206796 1002096 206802 1002108
rect 208394 1002096 208400 1002108
rect 206796 1002068 208400 1002096
rect 206796 1002056 206802 1002068
rect 208394 1002056 208400 1002068
rect 208452 1002056 208458 1002108
rect 211246 1002056 211252 1002108
rect 211304 1002096 211310 1002108
rect 213362 1002096 213368 1002108
rect 211304 1002068 213368 1002096
rect 211304 1002056 211310 1002068
rect 213362 1002056 213368 1002068
rect 213420 1002056 213426 1002108
rect 200758 1001988 200764 1002040
rect 200816 1002028 200822 1002040
rect 202690 1002028 202696 1002040
rect 200816 1002000 202696 1002028
rect 200816 1001988 200822 1002000
rect 202690 1001988 202696 1002000
rect 202748 1001988 202754 1002040
rect 211706 1001988 211712 1002040
rect 211764 1002028 211770 1002040
rect 215938 1002028 215944 1002040
rect 211764 1002000 215944 1002028
rect 211764 1001988 211770 1002000
rect 215938 1001988 215944 1002000
rect 215996 1001988 216002 1002040
rect 200942 1001920 200948 1001972
rect 201000 1001960 201006 1001972
rect 203058 1001960 203064 1001972
rect 201000 1001932 203064 1001960
rect 201000 1001920 201006 1001932
rect 203058 1001920 203064 1001932
rect 203116 1001920 203122 1001972
rect 203518 1001920 203524 1001972
rect 203576 1001960 203582 1001972
rect 205910 1001960 205916 1001972
rect 203576 1001932 205916 1001960
rect 203576 1001920 203582 1001932
rect 205910 1001920 205916 1001932
rect 205968 1001920 205974 1001972
rect 212074 1001920 212080 1001972
rect 212132 1001960 212138 1001972
rect 213914 1001960 213920 1001972
rect 212132 1001932 213920 1001960
rect 212132 1001920 212138 1001932
rect 213914 1001920 213920 1001932
rect 213972 1001920 213978 1001972
rect 246592 1001904 246620 1002612
rect 253658 1002600 253664 1002612
rect 253716 1002600 253722 1002652
rect 552750 1002600 552756 1002652
rect 552808 1002640 552814 1002652
rect 565906 1002640 565912 1002652
rect 552808 1002612 565912 1002640
rect 552808 1002600 552814 1002612
rect 565906 1002600 565912 1002612
rect 565964 1002600 565970 1002652
rect 246666 1002532 246672 1002584
rect 246724 1002572 246730 1002584
rect 254946 1002572 254952 1002584
rect 246724 1002544 254952 1002572
rect 246724 1002532 246730 1002544
rect 254946 1002532 254952 1002544
rect 255004 1002532 255010 1002584
rect 552290 1002532 552296 1002584
rect 552348 1002572 552354 1002584
rect 568666 1002572 568672 1002584
rect 552348 1002544 568672 1002572
rect 552348 1002532 552354 1002544
rect 568666 1002532 568672 1002544
rect 568724 1002532 568730 1002584
rect 559190 1002260 559196 1002312
rect 559248 1002300 559254 1002312
rect 562318 1002300 562324 1002312
rect 559248 1002272 562324 1002300
rect 559248 1002260 559254 1002272
rect 562318 1002260 562324 1002272
rect 562376 1002260 562382 1002312
rect 260190 1002192 260196 1002244
rect 260248 1002232 260254 1002244
rect 262858 1002232 262864 1002244
rect 260248 1002204 262864 1002232
rect 260248 1002192 260254 1002204
rect 262858 1002192 262864 1002204
rect 262916 1002192 262922 1002244
rect 559650 1002192 559656 1002244
rect 559708 1002232 559714 1002244
rect 561766 1002232 561772 1002244
rect 559708 1002204 561772 1002232
rect 559708 1002192 559714 1002204
rect 561766 1002192 561772 1002204
rect 561824 1002192 561830 1002244
rect 253198 1002124 253204 1002176
rect 253256 1002164 253262 1002176
rect 256142 1002164 256148 1002176
rect 253256 1002136 256148 1002164
rect 253256 1002124 253262 1002136
rect 256142 1002124 256148 1002136
rect 256200 1002124 256206 1002176
rect 261846 1002124 261852 1002176
rect 261904 1002164 261910 1002176
rect 264238 1002164 264244 1002176
rect 261904 1002136 264244 1002164
rect 261904 1002124 261910 1002136
rect 264238 1002124 264244 1002136
rect 264296 1002124 264302 1002176
rect 558454 1002124 558460 1002176
rect 558512 1002164 558518 1002176
rect 560938 1002164 560944 1002176
rect 558512 1002136 560944 1002164
rect 558512 1002124 558518 1002136
rect 560938 1002124 560944 1002136
rect 560996 1002124 561002 1002176
rect 561306 1002124 561312 1002176
rect 561364 1002164 561370 1002176
rect 566458 1002164 566464 1002176
rect 561364 1002136 566464 1002164
rect 561364 1002124 561370 1002136
rect 566458 1002124 566464 1002136
rect 566516 1002124 566522 1002176
rect 253382 1002056 253388 1002108
rect 253440 1002096 253446 1002108
rect 255682 1002096 255688 1002108
rect 253440 1002068 255688 1002096
rect 253440 1002056 253446 1002068
rect 255682 1002056 255688 1002068
rect 255740 1002056 255746 1002108
rect 261478 1002056 261484 1002108
rect 261536 1002096 261542 1002108
rect 263594 1002096 263600 1002108
rect 261536 1002068 263600 1002096
rect 261536 1002056 261542 1002068
rect 263594 1002056 263600 1002068
rect 263652 1002056 263658 1002108
rect 502518 1002056 502524 1002108
rect 502576 1002096 502582 1002108
rect 505094 1002096 505100 1002108
rect 502576 1002068 505100 1002096
rect 502576 1002056 502582 1002068
rect 505094 1002056 505100 1002068
rect 505152 1002056 505158 1002108
rect 553210 1002056 553216 1002108
rect 553268 1002096 553274 1002108
rect 554774 1002096 554780 1002108
rect 553268 1002068 554780 1002096
rect 553268 1002056 553274 1002068
rect 554774 1002056 554780 1002068
rect 554832 1002056 554838 1002108
rect 560018 1002056 560024 1002108
rect 560076 1002096 560082 1002108
rect 562502 1002096 562508 1002108
rect 560076 1002068 562508 1002096
rect 560076 1002056 560082 1002068
rect 562502 1002056 562508 1002068
rect 562560 1002056 562566 1002108
rect 251910 1001988 251916 1002040
rect 251968 1002028 251974 1002040
rect 254486 1002028 254492 1002040
rect 251968 1002000 254492 1002028
rect 251968 1001988 251974 1002000
rect 254486 1001988 254492 1002000
rect 254544 1001988 254550 1002040
rect 254578 1001988 254584 1002040
rect 254636 1002028 254642 1002040
rect 256970 1002028 256976 1002040
rect 254636 1002000 256976 1002028
rect 254636 1001988 254642 1002000
rect 256970 1001988 256976 1002000
rect 257028 1001988 257034 1002040
rect 260650 1001988 260656 1002040
rect 260708 1002028 260714 1002040
rect 262214 1002028 262220 1002040
rect 260708 1002000 262220 1002028
rect 260708 1001988 260714 1002000
rect 262214 1001988 262220 1002000
rect 262272 1001988 262278 1002040
rect 311434 1001988 311440 1002040
rect 311492 1002028 311498 1002040
rect 313366 1002028 313372 1002040
rect 311492 1002000 313372 1002028
rect 311492 1001988 311498 1002000
rect 313366 1001988 313372 1002000
rect 313424 1001988 313430 1002040
rect 357066 1001988 357072 1002040
rect 357124 1002028 357130 1002040
rect 358906 1002028 358912 1002040
rect 357124 1002000 358912 1002028
rect 357124 1001988 357130 1002000
rect 358906 1001988 358912 1002000
rect 358964 1001988 358970 1002040
rect 361022 1001988 361028 1002040
rect 361080 1002028 361086 1002040
rect 363598 1002028 363604 1002040
rect 361080 1002000 363604 1002028
rect 361080 1001988 361086 1002000
rect 363598 1001988 363604 1002000
rect 363656 1001988 363662 1002040
rect 365070 1001988 365076 1002040
rect 365128 1002028 365134 1002040
rect 370498 1002028 370504 1002040
rect 365128 1002000 370504 1002028
rect 365128 1001988 365134 1002000
rect 370498 1001988 370504 1002000
rect 370556 1001988 370562 1002040
rect 500862 1001988 500868 1002040
rect 500920 1002028 500926 1002040
rect 503346 1002028 503352 1002040
rect 500920 1002000 503352 1002028
rect 500920 1001988 500926 1002000
rect 503346 1001988 503352 1002000
rect 503404 1001988 503410 1002040
rect 551738 1001988 551744 1002040
rect 551796 1002028 551802 1002040
rect 553946 1002028 553952 1002040
rect 551796 1002000 553952 1002028
rect 551796 1001988 551802 1002000
rect 553946 1001988 553952 1002000
rect 554004 1001988 554010 1002040
rect 557994 1001988 558000 1002040
rect 558052 1002028 558058 1002040
rect 560386 1002028 560392 1002040
rect 558052 1002000 560392 1002028
rect 558052 1001988 558058 1002000
rect 560386 1001988 560392 1002000
rect 560444 1001988 560450 1002040
rect 560846 1001988 560852 1002040
rect 560904 1002028 560910 1002040
rect 565078 1002028 565084 1002040
rect 560904 1002000 565084 1002028
rect 560904 1001988 560910 1002000
rect 565078 1001988 565084 1002000
rect 565136 1001988 565142 1002040
rect 249150 1001920 249156 1001972
rect 249208 1001960 249214 1001972
rect 254118 1001960 254124 1001972
rect 249208 1001932 254124 1001960
rect 249208 1001920 249214 1001932
rect 254118 1001920 254124 1001932
rect 254176 1001920 254182 1001972
rect 254762 1001920 254768 1001972
rect 254820 1001960 254826 1001972
rect 257798 1001960 257804 1001972
rect 254820 1001932 257804 1001960
rect 254820 1001920 254826 1001932
rect 257798 1001920 257804 1001932
rect 257856 1001920 257862 1001972
rect 259822 1001920 259828 1001972
rect 259880 1001960 259886 1001972
rect 260926 1001960 260932 1001972
rect 259880 1001932 260932 1001960
rect 259880 1001920 259886 1001932
rect 260926 1001920 260932 1001932
rect 260984 1001920 260990 1001972
rect 263502 1001920 263508 1001972
rect 263560 1001960 263566 1001972
rect 265618 1001960 265624 1001972
rect 263560 1001932 265624 1001960
rect 263560 1001920 263566 1001932
rect 265618 1001920 265624 1001932
rect 265676 1001920 265682 1001972
rect 302878 1001920 302884 1001972
rect 302936 1001960 302942 1001972
rect 305270 1001960 305276 1001972
rect 302936 1001932 305276 1001960
rect 302936 1001920 302942 1001932
rect 305270 1001920 305276 1001932
rect 305328 1001920 305334 1001972
rect 310146 1001920 310152 1001972
rect 310204 1001960 310210 1001972
rect 311894 1001960 311900 1001972
rect 310204 1001932 311900 1001960
rect 310204 1001920 310210 1001932
rect 311894 1001920 311900 1001932
rect 311952 1001920 311958 1001972
rect 355778 1001920 355784 1001972
rect 355836 1001960 355842 1001972
rect 358538 1001960 358544 1001972
rect 355836 1001932 358544 1001960
rect 355836 1001920 355842 1001932
rect 358538 1001920 358544 1001932
rect 358596 1001920 358602 1001972
rect 358722 1001920 358728 1001972
rect 358780 1001960 358786 1001972
rect 359366 1001960 359372 1001972
rect 358780 1001932 359372 1001960
rect 358780 1001920 358786 1001932
rect 359366 1001920 359372 1001932
rect 359424 1001920 359430 1001972
rect 360194 1001920 360200 1001972
rect 360252 1001960 360258 1001972
rect 362218 1001960 362224 1001972
rect 360252 1001932 362224 1001960
rect 360252 1001920 360258 1001932
rect 362218 1001920 362224 1001932
rect 362276 1001920 362282 1001972
rect 365438 1001920 365444 1001972
rect 365496 1001960 365502 1001972
rect 367738 1001960 367744 1001972
rect 365496 1001932 367744 1001960
rect 365496 1001920 365502 1001932
rect 367738 1001920 367744 1001932
rect 367796 1001920 367802 1001972
rect 420730 1001920 420736 1001972
rect 420788 1001960 420794 1001972
rect 421466 1001960 421472 1001972
rect 420788 1001932 421472 1001960
rect 420788 1001920 420794 1001932
rect 421466 1001920 421472 1001932
rect 421524 1001920 421530 1001972
rect 424318 1001920 424324 1001972
rect 424376 1001960 424382 1001972
rect 425698 1001960 425704 1001972
rect 424376 1001932 425704 1001960
rect 424376 1001920 424382 1001932
rect 425698 1001920 425704 1001932
rect 425756 1001920 425762 1001972
rect 464982 1001920 464988 1001972
rect 465040 1001960 465046 1001972
rect 472526 1001960 472532 1001972
rect 465040 1001932 472532 1001960
rect 465040 1001920 465046 1001932
rect 472526 1001920 472532 1001932
rect 472584 1001920 472590 1001972
rect 502150 1001920 502156 1001972
rect 502208 1001960 502214 1001972
rect 502886 1001960 502892 1001972
rect 502208 1001932 502892 1001960
rect 502208 1001920 502214 1001932
rect 502886 1001920 502892 1001932
rect 502944 1001920 502950 1001972
rect 505002 1001920 505008 1001972
rect 505060 1001960 505066 1001972
rect 506658 1001960 506664 1001972
rect 505060 1001932 506664 1001960
rect 505060 1001920 505066 1001932
rect 506658 1001920 506664 1001932
rect 506716 1001920 506722 1001972
rect 550542 1001920 550548 1001972
rect 550600 1001960 550606 1001972
rect 553118 1001960 553124 1001972
rect 550600 1001932 553124 1001960
rect 550600 1001920 550606 1001932
rect 553118 1001920 553124 1001932
rect 553176 1001920 553182 1001972
rect 558822 1001920 558828 1001972
rect 558880 1001960 558886 1001972
rect 560294 1001960 560300 1001972
rect 558880 1001932 560300 1001960
rect 558880 1001920 558886 1001932
rect 560294 1001920 560300 1001932
rect 560352 1001920 560358 1001972
rect 560478 1001920 560484 1001972
rect 560536 1001960 560542 1001972
rect 563054 1001960 563060 1001972
rect 560536 1001932 563060 1001960
rect 560536 1001920 560542 1001932
rect 563054 1001920 563060 1001932
rect 563112 1001920 563118 1001972
rect 195146 1001852 195152 1001904
rect 195204 1001892 195210 1001904
rect 195330 1001892 195336 1001904
rect 195204 1001864 195336 1001892
rect 195204 1001852 195210 1001864
rect 195330 1001852 195336 1001864
rect 195388 1001852 195394 1001904
rect 206922 1001852 206928 1001904
rect 206980 1001892 206986 1001904
rect 207566 1001892 207572 1001904
rect 206980 1001864 207572 1001892
rect 206980 1001852 206986 1001864
rect 207566 1001852 207572 1001864
rect 207624 1001852 207630 1001904
rect 246574 1001852 246580 1001904
rect 246632 1001852 246638 1001904
rect 195146 1001620 195152 1001632
rect 195072 1001592 195152 1001620
rect 195146 1001580 195152 1001592
rect 195204 1001580 195210 1001632
rect 247034 1001240 247040 1001292
rect 247092 1001280 247098 1001292
rect 251910 1001280 251916 1001292
rect 247092 1001252 251916 1001280
rect 247092 1001240 247098 1001252
rect 251910 1001240 251916 1001252
rect 251968 1001240 251974 1001292
rect 92290 1001172 92296 1001224
rect 92348 1001212 92354 1001224
rect 95970 1001212 95976 1001224
rect 92348 1001184 95976 1001212
rect 92348 1001172 92354 1001184
rect 95970 1001172 95976 1001184
rect 96028 1001172 96034 1001224
rect 247126 1001172 247132 1001224
rect 247184 1001212 247190 1001224
rect 253382 1001212 253388 1001224
rect 247184 1001184 253388 1001212
rect 247184 1001172 247190 1001184
rect 253382 1001172 253388 1001184
rect 253440 1001172 253446 1001224
rect 425698 1001172 425704 1001224
rect 425756 1001212 425762 1001224
rect 438762 1001212 438768 1001224
rect 425756 1001184 438768 1001212
rect 425756 1001172 425762 1001184
rect 438762 1001172 438768 1001184
rect 438820 1001172 438826 1001224
rect 251542 1000560 251548 1000612
rect 251600 1000600 251606 1000612
rect 254670 1000600 254676 1000612
rect 251600 1000572 254676 1000600
rect 251600 1000560 251606 1000572
rect 254670 1000560 254676 1000572
rect 254728 1000560 254734 1000612
rect 250438 1000492 250444 1000544
rect 250496 1000532 250502 1000544
rect 253198 1000532 253204 1000544
rect 250496 1000504 253204 1000532
rect 250496 1000492 250502 1000504
rect 253198 1000492 253204 1000504
rect 253256 1000492 253262 1000544
rect 612734 1000492 612740 1000544
rect 612792 1000532 612798 1000544
rect 625522 1000532 625528 1000544
rect 612792 1000504 625528 1000532
rect 612792 1000492 612798 1000504
rect 625522 1000492 625528 1000504
rect 625580 1000492 625586 1000544
rect 197354 1000356 197360 1000408
rect 197412 1000396 197418 1000408
rect 200942 1000396 200948 1000408
rect 197412 1000368 200948 1000396
rect 197412 1000356 197418 1000368
rect 200942 1000356 200948 1000368
rect 201000 1000356 201006 1000408
rect 563790 1000084 563796 1000136
rect 563848 1000124 563854 1000136
rect 565814 1000124 565820 1000136
rect 563848 1000096 565820 1000124
rect 563848 1000084 563854 1000096
rect 565814 1000084 565820 1000096
rect 565872 1000084 565878 1000136
rect 565906 1000016 565912 1000068
rect 565964 1000056 565970 1000068
rect 568758 1000056 568764 1000068
rect 565964 1000028 568764 1000056
rect 565964 1000016 565970 1000028
rect 568758 1000016 568764 1000028
rect 568816 1000016 568822 1000068
rect 426342 999744 426348 999796
rect 426400 999784 426406 999796
rect 446306 999784 446312 999796
rect 426400 999756 446312 999784
rect 426400 999744 426406 999756
rect 446306 999744 446312 999756
rect 446364 999744 446370 999796
rect 499390 999744 499396 999796
rect 499448 999784 499454 999796
rect 504266 999784 504272 999796
rect 499448 999756 504272 999784
rect 499448 999744 499454 999756
rect 504266 999744 504272 999756
rect 504324 999744 504330 999796
rect 505094 999744 505100 999796
rect 505152 999784 505158 999796
rect 515950 999784 515956 999796
rect 505152 999756 515956 999784
rect 505152 999744 505158 999756
rect 515950 999744 515956 999756
rect 516008 999744 516014 999796
rect 551738 999744 551744 999796
rect 551796 999784 551802 999796
rect 562226 999784 562232 999796
rect 551796 999756 562232 999784
rect 551796 999744 551802 999756
rect 562226 999744 562232 999756
rect 562284 999744 562290 999796
rect 563698 999744 563704 999796
rect 563756 999784 563762 999796
rect 572714 999784 572720 999796
rect 563756 999756 572720 999784
rect 563756 999744 563762 999756
rect 572714 999744 572720 999756
rect 572772 999744 572778 999796
rect 95970 999676 95976 999728
rect 96028 999716 96034 999728
rect 98822 999716 98828 999728
rect 96028 999688 98828 999716
rect 96028 999676 96034 999688
rect 98822 999676 98828 999688
rect 98880 999676 98886 999728
rect 94774 999336 94780 999388
rect 94832 999376 94838 999388
rect 97534 999376 97540 999388
rect 94832 999348 97540 999376
rect 94832 999336 94838 999348
rect 97534 999336 97540 999348
rect 97592 999336 97598 999388
rect 251358 999132 251364 999184
rect 251416 999172 251422 999184
rect 254762 999172 254768 999184
rect 251416 999144 254768 999172
rect 251416 999132 251422 999144
rect 254762 999132 254768 999144
rect 254820 999132 254826 999184
rect 298186 999132 298192 999184
rect 298244 999172 298250 999184
rect 327534 999172 327540 999184
rect 298244 999144 327540 999172
rect 298244 999132 298250 999144
rect 327534 999132 327540 999144
rect 327592 999132 327598 999184
rect 618162 999132 618168 999184
rect 618220 999172 618226 999184
rect 625430 999172 625436 999184
rect 618220 999144 625436 999172
rect 618220 999132 618226 999144
rect 625430 999132 625436 999144
rect 625488 999132 625494 999184
rect 92290 999064 92296 999116
rect 92348 999104 92354 999116
rect 94590 999104 94596 999116
rect 92348 999076 94596 999104
rect 92348 999064 92354 999076
rect 94590 999064 94596 999076
rect 94648 999064 94654 999116
rect 446398 999064 446404 999116
rect 446456 999104 446462 999116
rect 448606 999104 448612 999116
rect 446456 999076 448612 999104
rect 446456 999064 446462 999076
rect 448606 999064 448612 999076
rect 448664 999064 448670 999116
rect 357342 998724 357348 998776
rect 357400 998764 357406 998776
rect 360194 998764 360200 998776
rect 357400 998736 360200 998764
rect 357400 998724 357406 998736
rect 360194 998724 360200 998736
rect 360252 998724 360258 998776
rect 464798 998724 464804 998776
rect 464856 998764 464862 998776
rect 472434 998764 472440 998776
rect 464856 998736 472440 998764
rect 464856 998724 464862 998736
rect 472434 998724 472440 998736
rect 472492 998724 472498 998776
rect 360838 998588 360844 998640
rect 360896 998628 360902 998640
rect 367370 998628 367376 998640
rect 360896 998600 367376 998628
rect 360896 998588 360902 998600
rect 367370 998588 367376 998600
rect 367428 998588 367434 998640
rect 380158 998588 380164 998640
rect 380216 998628 380222 998640
rect 383562 998628 383568 998640
rect 380216 998600 383568 998628
rect 380216 998588 380222 998600
rect 383562 998588 383568 998600
rect 383620 998588 383626 998640
rect 550542 998588 550548 998640
rect 550600 998628 550606 998640
rect 556154 998628 556160 998640
rect 550600 998600 556160 998628
rect 550600 998588 550606 998600
rect 556154 998588 556160 998600
rect 556212 998588 556218 998640
rect 358722 998520 358728 998572
rect 358780 998560 358786 998572
rect 372430 998560 372436 998572
rect 358780 998532 372436 998560
rect 358780 998520 358786 998532
rect 372430 998520 372436 998532
rect 372488 998520 372494 998572
rect 472342 998560 472348 998572
rect 451246 998532 472348 998560
rect 355778 998452 355784 998504
rect 355836 998492 355842 998504
rect 383378 998492 383384 998504
rect 355836 998464 383384 998492
rect 355836 998452 355842 998464
rect 383378 998452 383384 998464
rect 383436 998452 383442 998504
rect 448514 998452 448520 998504
rect 448572 998492 448578 998504
rect 451246 998492 451274 998532
rect 472342 998520 472348 998532
rect 472400 998520 472406 998572
rect 448572 998464 451274 998492
rect 448572 998452 448578 998464
rect 500862 998452 500868 998504
rect 500920 998492 500926 998504
rect 513282 998492 513288 998504
rect 500920 998464 513288 998492
rect 500920 998452 500926 998464
rect 513282 998452 513288 998464
rect 513340 998452 513346 998504
rect 517606 998452 517612 998504
rect 517664 998492 517670 998504
rect 523862 998492 523868 998504
rect 517664 998464 523868 998492
rect 517664 998452 517670 998464
rect 523862 998452 523868 998464
rect 523920 998452 523926 998504
rect 92382 998384 92388 998436
rect 92440 998424 92446 998436
rect 100110 998424 100116 998436
rect 92440 998396 100116 998424
rect 92440 998384 92446 998396
rect 100110 998384 100116 998396
rect 100168 998384 100174 998436
rect 195974 998384 195980 998436
rect 196032 998424 196038 998436
rect 206278 998424 206284 998436
rect 196032 998396 206284 998424
rect 196032 998384 196038 998396
rect 206278 998384 206284 998396
rect 206336 998384 206342 998436
rect 246758 998384 246764 998436
rect 246816 998424 246822 998436
rect 254578 998424 254584 998436
rect 246816 998396 254584 998424
rect 246816 998384 246822 998396
rect 254578 998384 254584 998396
rect 254636 998384 254642 998436
rect 354582 998384 354588 998436
rect 354640 998424 354646 998436
rect 383562 998424 383568 998436
rect 354640 998396 383568 998424
rect 354640 998384 354646 998396
rect 383562 998384 383568 998396
rect 383620 998384 383626 998436
rect 441614 998384 441620 998436
rect 441672 998424 441678 998436
rect 441672 998396 451274 998424
rect 441672 998384 441678 998396
rect 369210 998316 369216 998368
rect 369268 998356 369274 998368
rect 372338 998356 372344 998368
rect 369268 998328 372344 998356
rect 369268 998316 369274 998328
rect 372338 998316 372344 998328
rect 372396 998316 372402 998368
rect 451246 998356 451274 998396
rect 502150 998384 502156 998436
rect 502208 998424 502214 998436
rect 516042 998424 516048 998436
rect 502208 998396 516048 998424
rect 502208 998384 502214 998396
rect 516042 998384 516048 998396
rect 516100 998384 516106 998436
rect 517514 998384 517520 998436
rect 517572 998424 517578 998436
rect 523770 998424 523776 998436
rect 517572 998396 523776 998424
rect 517572 998384 517578 998396
rect 523770 998384 523776 998396
rect 523828 998384 523834 998436
rect 472618 998356 472624 998368
rect 451246 998328 472624 998356
rect 472618 998316 472624 998328
rect 472676 998316 472682 998368
rect 202414 998248 202420 998300
rect 202472 998288 202478 998300
rect 206922 998288 206928 998300
rect 202472 998260 206928 998288
rect 202472 998248 202478 998260
rect 206922 998248 206928 998260
rect 206980 998248 206986 998300
rect 506658 998248 506664 998300
rect 506716 998288 506722 998300
rect 516686 998288 516692 998300
rect 506716 998260 516692 998288
rect 506716 998248 506722 998260
rect 516686 998248 516692 998260
rect 516744 998248 516750 998300
rect 430850 998112 430856 998164
rect 430908 998152 430914 998164
rect 436738 998152 436744 998164
rect 430908 998124 436744 998152
rect 430908 998112 430914 998124
rect 436738 998112 436744 998124
rect 436796 998112 436802 998164
rect 429654 998044 429660 998096
rect 429712 998084 429718 998096
rect 431954 998084 431960 998096
rect 429712 998056 431960 998084
rect 429712 998044 429718 998056
rect 431954 998044 431960 998056
rect 432012 998044 432018 998096
rect 507026 998044 507032 998096
rect 507084 998084 507090 998096
rect 510062 998084 510068 998096
rect 507084 998056 510068 998084
rect 507084 998044 507090 998056
rect 510062 998044 510068 998056
rect 510120 998044 510126 998096
rect 195422 997976 195428 998028
rect 195480 998016 195486 998028
rect 199378 998016 199384 998028
rect 195480 997988 199384 998016
rect 195480 997976 195486 997988
rect 199378 997976 199384 997988
rect 199436 997976 199442 998028
rect 428458 997976 428464 998028
rect 428516 998016 428522 998028
rect 430850 998016 430856 998028
rect 428516 997988 430856 998016
rect 428516 997976 428522 997988
rect 430850 997976 430856 997988
rect 430908 997976 430914 998028
rect 431678 997976 431684 998028
rect 431736 998016 431742 998028
rect 433978 998016 433984 998028
rect 431736 997988 433984 998016
rect 431736 997976 431742 997988
rect 433978 997976 433984 997988
rect 434036 997976 434042 998028
rect 508222 997976 508228 998028
rect 508280 998016 508286 998028
rect 510890 998016 510896 998028
rect 508280 997988 510896 998016
rect 508280 997976 508286 997988
rect 510890 997976 510896 997988
rect 510948 997976 510954 998028
rect 614114 997976 614120 998028
rect 614172 998016 614178 998028
rect 625614 998016 625620 998028
rect 614172 997988 625620 998016
rect 614172 997976 614178 997988
rect 625614 997976 625620 997988
rect 625672 997976 625678 998028
rect 312170 997908 312176 997960
rect 312228 997948 312234 997960
rect 314930 997948 314936 997960
rect 312228 997920 314936 997948
rect 312228 997908 312234 997920
rect 314930 997908 314936 997920
rect 314988 997908 314994 997960
rect 430390 997908 430396 997960
rect 430448 997948 430454 997960
rect 432138 997948 432144 997960
rect 430448 997920 432144 997948
rect 430448 997908 430454 997920
rect 432138 997908 432144 997920
rect 432196 997908 432202 997960
rect 507854 997908 507860 997960
rect 507912 997948 507918 997960
rect 509878 997948 509884 997960
rect 507912 997920 509884 997948
rect 507912 997908 507918 997920
rect 509878 997908 509884 997920
rect 509936 997908 509942 997960
rect 625706 997948 625712 997960
rect 620112 997920 625712 997948
rect 313826 997840 313832 997892
rect 313884 997880 313890 997892
rect 316034 997880 316040 997892
rect 313884 997852 316040 997880
rect 313884 997840 313890 997852
rect 316034 997840 316040 997852
rect 316092 997840 316098 997892
rect 429194 997840 429200 997892
rect 429252 997880 429258 997892
rect 431218 997880 431224 997892
rect 429252 997852 431224 997880
rect 429252 997840 429258 997852
rect 431218 997840 431224 997852
rect 431276 997840 431282 997892
rect 432046 997840 432052 997892
rect 432104 997880 432110 997892
rect 433426 997880 433432 997892
rect 432104 997852 433432 997880
rect 432104 997840 432110 997852
rect 433426 997840 433432 997852
rect 433484 997840 433490 997892
rect 506198 997840 506204 997892
rect 506256 997880 506262 997892
rect 508498 997880 508504 997892
rect 506256 997852 508504 997880
rect 506256 997840 506262 997852
rect 508498 997840 508504 997852
rect 508556 997840 508562 997892
rect 509050 997840 509056 997892
rect 509108 997880 509114 997892
rect 510706 997880 510712 997892
rect 509108 997852 510712 997880
rect 509108 997840 509114 997852
rect 510706 997840 510712 997852
rect 510764 997840 510770 997892
rect 143718 997772 143724 997824
rect 143776 997812 143782 997824
rect 145742 997812 145748 997824
rect 143776 997784 145748 997812
rect 143776 997772 143782 997784
rect 145742 997772 145748 997784
rect 145800 997772 145806 997824
rect 195330 997772 195336 997824
rect 195388 997812 195394 997824
rect 196618 997812 196624 997824
rect 195388 997784 196624 997812
rect 195388 997772 195394 997784
rect 196618 997772 196624 997784
rect 196676 997772 196682 997824
rect 246850 997772 246856 997824
rect 246908 997812 246914 997824
rect 279326 997812 279332 997824
rect 246908 997784 279332 997812
rect 246908 997772 246914 997784
rect 279326 997772 279332 997784
rect 279384 997772 279390 997824
rect 303246 997772 303252 997824
rect 303304 997812 303310 997824
rect 305822 997812 305828 997824
rect 303304 997784 305828 997812
rect 303304 997772 303310 997784
rect 305822 997772 305828 997784
rect 305880 997772 305886 997824
rect 312998 997772 313004 997824
rect 313056 997812 313062 997824
rect 314746 997812 314752 997824
rect 313056 997784 314752 997812
rect 313056 997772 313062 997784
rect 314746 997772 314752 997784
rect 314804 997772 314810 997824
rect 315114 997772 315120 997824
rect 315172 997812 315178 997824
rect 319438 997812 319444 997824
rect 315172 997784 319444 997812
rect 315172 997772 315178 997784
rect 319438 997772 319444 997784
rect 319496 997772 319502 997824
rect 400122 997772 400128 997824
rect 400180 997812 400186 997824
rect 400180 997784 437520 997812
rect 400180 997772 400186 997784
rect 143810 997704 143816 997756
rect 143868 997744 143874 997756
rect 161474 997744 161480 997756
rect 143868 997716 161480 997744
rect 143868 997704 143874 997716
rect 161474 997704 161480 997716
rect 161532 997704 161538 997756
rect 195238 997704 195244 997756
rect 195296 997744 195302 997756
rect 211246 997744 211252 997756
rect 195296 997716 211252 997744
rect 195296 997704 195302 997716
rect 211246 997704 211252 997716
rect 211304 997704 211310 997756
rect 246574 997704 246580 997756
rect 246632 997744 246638 997756
rect 261846 997744 261852 997756
rect 246632 997716 261852 997744
rect 246632 997704 246638 997716
rect 261846 997704 261852 997716
rect 261904 997704 261910 997756
rect 298370 997704 298376 997756
rect 298428 997744 298434 997756
rect 316034 997744 316040 997756
rect 298428 997716 316040 997744
rect 298428 997704 298434 997716
rect 316034 997704 316040 997716
rect 316092 997704 316098 997756
rect 399938 997704 399944 997756
rect 399996 997744 400002 997756
rect 433426 997744 433432 997756
rect 399996 997716 433432 997744
rect 399996 997704 400002 997716
rect 433426 997704 433432 997716
rect 433484 997704 433490 997756
rect 437492 997744 437520 997784
rect 507394 997772 507400 997824
rect 507452 997812 507458 997824
rect 509234 997812 509240 997824
rect 507452 997784 509240 997812
rect 507452 997772 507458 997784
rect 509234 997772 509240 997784
rect 509292 997772 509298 997824
rect 509510 997772 509516 997824
rect 509568 997812 509574 997824
rect 514018 997812 514024 997824
rect 509568 997784 514024 997812
rect 509568 997772 509574 997784
rect 514018 997772 514024 997784
rect 514076 997772 514082 997824
rect 540330 997772 540336 997824
rect 540388 997812 540394 997824
rect 575566 997812 575572 997824
rect 540388 997784 575572 997812
rect 540388 997772 540394 997784
rect 575566 997772 575572 997784
rect 575624 997772 575630 997824
rect 607122 997772 607128 997824
rect 607180 997812 607186 997824
rect 620112 997812 620140 997920
rect 625706 997908 625712 997920
rect 625764 997908 625770 997960
rect 625798 997812 625804 997824
rect 607180 997784 620140 997812
rect 620296 997784 625804 997812
rect 607180 997772 607186 997784
rect 440234 997744 440240 997756
rect 437492 997716 440240 997744
rect 440234 997704 440240 997716
rect 440292 997704 440298 997756
rect 488902 997704 488908 997756
rect 488960 997744 488966 997756
rect 510706 997744 510712 997756
rect 488960 997716 510712 997744
rect 488960 997704 488966 997716
rect 510706 997704 510712 997716
rect 510764 997704 510770 997756
rect 559742 997704 559748 997756
rect 559800 997744 559806 997756
rect 620296 997744 620324 997784
rect 625798 997772 625804 997784
rect 625856 997772 625862 997824
rect 559800 997716 620324 997744
rect 559800 997704 559806 997716
rect 143902 997636 143908 997688
rect 143960 997676 143966 997688
rect 155770 997676 155776 997688
rect 143960 997648 155776 997676
rect 143960 997636 143966 997648
rect 155770 997636 155776 997648
rect 155828 997636 155834 997688
rect 400030 997636 400036 997688
rect 400088 997676 400094 997688
rect 432046 997676 432052 997688
rect 400088 997648 432052 997676
rect 400088 997636 400094 997648
rect 432046 997636 432052 997648
rect 432104 997636 432110 997688
rect 540882 997636 540888 997688
rect 540940 997676 540946 997688
rect 563054 997676 563060 997688
rect 540940 997648 563060 997676
rect 540940 997636 540946 997648
rect 563054 997636 563060 997648
rect 563112 997636 563118 997688
rect 565814 997636 565820 997688
rect 565872 997676 565878 997688
rect 623682 997676 623688 997688
rect 565872 997648 623688 997676
rect 565872 997636 565878 997648
rect 623682 997636 623688 997648
rect 623740 997636 623746 997688
rect 554314 997568 554320 997620
rect 554372 997608 554378 997620
rect 607122 997608 607128 997620
rect 554372 997580 607128 997608
rect 554372 997568 554378 997580
rect 607122 997568 607128 997580
rect 607180 997568 607186 997620
rect 92658 997500 92664 997552
rect 92716 997540 92722 997552
rect 95970 997540 95976 997552
rect 92716 997512 95976 997540
rect 92716 997500 92722 997512
rect 95970 997500 95976 997512
rect 96028 997500 96034 997552
rect 554682 997500 554688 997552
rect 554740 997540 554746 997552
rect 561490 997540 561496 997552
rect 554740 997512 561496 997540
rect 554740 997500 554746 997512
rect 561490 997500 561496 997512
rect 561548 997500 561554 997552
rect 562226 997500 562232 997552
rect 562284 997540 562290 997552
rect 614114 997540 614120 997552
rect 562284 997512 614120 997540
rect 562284 997500 562290 997512
rect 614114 997500 614120 997512
rect 614172 997500 614178 997552
rect 553210 997432 553216 997484
rect 553268 997472 553274 997484
rect 561582 997472 561588 997484
rect 553268 997444 561588 997472
rect 553268 997432 553274 997444
rect 561582 997432 561588 997444
rect 561640 997432 561646 997484
rect 568758 997432 568764 997484
rect 568816 997472 568822 997484
rect 618162 997472 618168 997484
rect 568816 997444 618168 997472
rect 568816 997432 568822 997444
rect 618162 997432 618168 997444
rect 618220 997432 618226 997484
rect 154574 997364 154580 997416
rect 154632 997404 154638 997416
rect 157334 997404 157340 997416
rect 154632 997376 157340 997404
rect 154632 997364 154638 997376
rect 157334 997364 157340 997376
rect 157392 997364 157398 997416
rect 573358 997364 573364 997416
rect 573416 997404 573422 997416
rect 612734 997404 612740 997416
rect 573416 997376 612740 997404
rect 573416 997364 573422 997376
rect 612734 997364 612740 997376
rect 612792 997364 612798 997416
rect 215754 997296 215760 997348
rect 215812 997336 215818 997348
rect 218882 997336 218888 997348
rect 215812 997308 218888 997336
rect 215812 997296 215818 997308
rect 218882 997296 218888 997308
rect 218940 997296 218946 997348
rect 369210 997296 369216 997348
rect 369268 997336 369274 997348
rect 372338 997336 372344 997348
rect 369268 997308 372344 997336
rect 369268 997296 369274 997308
rect 372338 997296 372344 997308
rect 372396 997296 372402 997348
rect 113818 997228 113824 997280
rect 113876 997268 113882 997280
rect 116118 997268 116124 997280
rect 113876 997240 116124 997268
rect 113876 997228 113882 997240
rect 116118 997228 116124 997240
rect 116176 997228 116182 997280
rect 164418 997228 164424 997280
rect 164476 997268 164482 997280
rect 167546 997268 167552 997280
rect 164476 997240 167552 997268
rect 164476 997228 164482 997240
rect 167546 997228 167552 997240
rect 167604 997228 167610 997280
rect 268470 997228 268476 997280
rect 268528 997268 268534 997280
rect 270310 997268 270316 997280
rect 268528 997240 270316 997268
rect 268528 997228 268534 997240
rect 270310 997228 270316 997240
rect 270368 997228 270374 997280
rect 436554 997228 436560 997280
rect 436612 997268 436618 997280
rect 439682 997268 439688 997280
rect 436612 997240 439688 997268
rect 436612 997228 436618 997240
rect 439682 997228 439688 997240
rect 439740 997228 439746 997280
rect 515398 997228 515404 997280
rect 515456 997268 515462 997280
rect 516686 997268 516692 997280
rect 515456 997240 516692 997268
rect 515456 997228 515462 997240
rect 516686 997228 516692 997240
rect 516744 997228 516750 997280
rect 564986 997228 564992 997280
rect 565044 997268 565050 997280
rect 568114 997268 568120 997280
rect 565044 997240 568120 997268
rect 565044 997228 565050 997240
rect 568114 997228 568120 997240
rect 568172 997228 568178 997280
rect 572714 997228 572720 997280
rect 572772 997268 572778 997280
rect 572772 997240 581684 997268
rect 572772 997228 572778 997240
rect 575198 997160 575204 997212
rect 575256 997200 575262 997212
rect 580902 997200 580908 997212
rect 575256 997172 580908 997200
rect 575256 997160 575262 997172
rect 580902 997160 580908 997172
rect 580960 997160 580966 997212
rect 581656 997200 581684 997240
rect 585134 997228 585140 997280
rect 585192 997268 585198 997280
rect 590930 997268 590936 997280
rect 585192 997240 590936 997268
rect 585192 997228 585198 997240
rect 590930 997228 590936 997240
rect 590988 997228 590994 997280
rect 620278 997200 620284 997212
rect 581656 997172 620284 997200
rect 620278 997160 620284 997172
rect 620336 997160 620342 997212
rect 92474 997092 92480 997144
rect 92532 997132 92538 997144
rect 97350 997132 97356 997144
rect 92532 997104 97356 997132
rect 92532 997092 92538 997104
rect 97350 997092 97356 997104
rect 97408 997092 97414 997144
rect 112990 997092 112996 997144
rect 113048 997132 113054 997144
rect 116118 997132 116124 997144
rect 113048 997104 116124 997132
rect 113048 997092 113054 997104
rect 116118 997092 116124 997104
rect 116176 997092 116182 997144
rect 164418 997092 164424 997144
rect 164476 997132 164482 997144
rect 167546 997132 167552 997144
rect 164476 997104 167552 997132
rect 164476 997092 164482 997104
rect 167546 997092 167552 997104
rect 167604 997092 167610 997144
rect 195238 997092 195244 997144
rect 195296 997132 195302 997144
rect 197998 997132 198004 997144
rect 195296 997104 198004 997132
rect 195296 997092 195302 997104
rect 197998 997092 198004 997104
rect 198056 997092 198062 997144
rect 200206 997092 200212 997144
rect 200264 997132 200270 997144
rect 204898 997132 204904 997144
rect 200264 997104 204904 997132
rect 200264 997092 200270 997104
rect 204898 997092 204904 997104
rect 204956 997092 204962 997144
rect 319438 997092 319444 997144
rect 319496 997132 319502 997144
rect 332594 997132 332600 997144
rect 319496 997104 332600 997132
rect 319496 997092 319502 997104
rect 332594 997092 332600 997104
rect 332652 997092 332658 997144
rect 556706 997092 556712 997144
rect 556764 997132 556770 997144
rect 605926 997132 605932 997144
rect 556764 997104 605932 997132
rect 556764 997092 556770 997104
rect 605926 997092 605932 997104
rect 605984 997092 605990 997144
rect 92566 997024 92572 997076
rect 92624 997064 92630 997076
rect 100018 997064 100024 997076
rect 92624 997036 100024 997064
rect 92624 997024 92630 997036
rect 100018 997024 100024 997036
rect 100076 997024 100082 997076
rect 327534 997024 327540 997076
rect 327592 997064 327598 997076
rect 367830 997064 367836 997076
rect 327592 997036 367836 997064
rect 327592 997024 327598 997036
rect 367830 997024 367836 997036
rect 367888 997024 367894 997076
rect 570598 997024 570604 997076
rect 570656 997064 570662 997076
rect 622394 997064 622400 997076
rect 570656 997036 622400 997064
rect 570656 997024 570662 997036
rect 622394 997024 622400 997036
rect 622452 997024 622458 997076
rect 365162 996956 365168 997008
rect 365220 996996 365226 997008
rect 372338 996996 372344 997008
rect 365220 996968 372344 996996
rect 365220 996956 365226 996968
rect 372338 996956 372344 996968
rect 372396 996956 372402 997008
rect 564986 996888 564992 996940
rect 565044 996928 565050 996940
rect 568114 996928 568120 996940
rect 565044 996900 568120 996928
rect 565044 996888 565050 996900
rect 568114 996888 568120 996900
rect 568172 996888 568178 996940
rect 575474 996820 575480 996872
rect 575532 996860 575538 996872
rect 580718 996860 580724 996872
rect 575532 996832 580724 996860
rect 575532 996820 575538 996832
rect 580718 996820 580724 996832
rect 580776 996820 580782 996872
rect 585502 996820 585508 996872
rect 585560 996860 585566 996872
rect 590562 996860 590568 996872
rect 585560 996832 590568 996860
rect 585560 996820 585566 996832
rect 590562 996820 590568 996832
rect 590620 996820 590626 996872
rect 298278 996616 298284 996668
rect 298336 996656 298342 996668
rect 300210 996656 300216 996668
rect 298336 996628 300216 996656
rect 298336 996616 298342 996628
rect 300210 996616 300216 996628
rect 300268 996616 300274 996668
rect 144822 996344 144828 996396
rect 144880 996384 144886 996396
rect 149698 996384 149704 996396
rect 144880 996356 149704 996384
rect 144880 996344 144886 996356
rect 149698 996344 149704 996356
rect 149756 996344 149762 996396
rect 299014 996344 299020 996396
rect 299072 996384 299078 996396
rect 301498 996384 301504 996396
rect 299072 996356 301504 996384
rect 299072 996344 299078 996356
rect 301498 996344 301504 996356
rect 301556 996344 301562 996396
rect 159358 996140 159364 996192
rect 159416 996180 159422 996192
rect 209774 996180 209780 996192
rect 159416 996152 209780 996180
rect 159416 996140 159422 996152
rect 209774 996140 209780 996152
rect 209832 996140 209838 996192
rect 213178 996140 213184 996192
rect 213236 996180 213242 996192
rect 263594 996180 263600 996192
rect 213236 996152 263600 996180
rect 213236 996140 213242 996152
rect 263594 996140 263600 996152
rect 263652 996140 263658 996192
rect 264238 996140 264244 996192
rect 264296 996180 264302 996192
rect 314746 996180 314752 996192
rect 264296 996152 314752 996180
rect 264296 996140 264302 996152
rect 314746 996140 314752 996152
rect 314804 996140 314810 996192
rect 431218 996140 431224 996192
rect 431276 996180 431282 996192
rect 506566 996180 506572 996192
rect 431276 996152 506572 996180
rect 431276 996140 431282 996152
rect 506566 996140 506572 996152
rect 506624 996140 506630 996192
rect 508498 996140 508504 996192
rect 508556 996180 508562 996192
rect 560386 996180 560392 996192
rect 508556 996152 560392 996180
rect 508556 996140 508562 996152
rect 560386 996140 560392 996152
rect 560444 996140 560450 996192
rect 108298 996072 108304 996124
rect 108356 996112 108362 996124
rect 158714 996112 158720 996124
rect 108356 996084 158720 996112
rect 108356 996072 108362 996084
rect 158714 996072 158720 996084
rect 158772 996072 158778 996124
rect 211798 996072 211804 996124
rect 211856 996112 211862 996124
rect 260926 996112 260932 996124
rect 211856 996084 260932 996112
rect 211856 996072 211862 996084
rect 260926 996072 260932 996084
rect 260984 996072 260990 996124
rect 262858 996072 262864 996124
rect 262916 996112 262922 996124
rect 313366 996112 313372 996124
rect 262916 996084 313372 996112
rect 262916 996072 262922 996084
rect 313366 996072 313372 996084
rect 313424 996072 313430 996124
rect 366358 996072 366364 996124
rect 366416 996112 366422 996124
rect 428458 996112 428464 996124
rect 366416 996084 428464 996112
rect 366416 996072 366422 996084
rect 428458 996072 428464 996084
rect 428516 996072 428522 996124
rect 509878 996072 509884 996124
rect 509936 996112 509942 996124
rect 561766 996112 561772 996124
rect 509936 996084 561772 996112
rect 509936 996072 509942 996084
rect 561766 996072 561772 996084
rect 561824 996072 561830 996124
rect 109678 996004 109684 996056
rect 109736 996044 109742 996056
rect 160186 996044 160192 996056
rect 109736 996016 160192 996044
rect 109736 996004 109742 996016
rect 160186 996004 160192 996016
rect 160244 996004 160250 996056
rect 166258 996004 166264 996056
rect 166316 996044 166322 996056
rect 212534 996044 212540 996056
rect 166316 996016 212540 996044
rect 166316 996004 166322 996016
rect 212534 996004 212540 996016
rect 212592 996004 212598 996056
rect 216030 996004 216036 996056
rect 216088 996044 216094 996056
rect 262214 996044 262220 996056
rect 216088 996016 262220 996044
rect 216088 996004 216094 996016
rect 262214 996004 262220 996016
rect 262272 996004 262278 996056
rect 268378 996004 268384 996056
rect 268436 996044 268442 996056
rect 314930 996044 314936 996056
rect 268436 996016 314936 996044
rect 268436 996004 268442 996016
rect 314930 996004 314936 996016
rect 314988 996004 314994 996056
rect 367370 996004 367376 996056
rect 367428 996044 367434 996056
rect 381538 996044 381544 996056
rect 367428 996016 381544 996044
rect 367428 996004 367434 996016
rect 381538 996004 381544 996016
rect 381596 996004 381602 996056
rect 468478 996004 468484 996056
rect 468536 996044 468542 996056
rect 509234 996044 509240 996056
rect 468536 996016 509240 996044
rect 468536 996004 468542 996016
rect 509234 996004 509240 996016
rect 509292 996004 509298 996056
rect 510062 996004 510068 996056
rect 510120 996044 510126 996056
rect 560294 996044 560300 996056
rect 510120 996016 560300 996044
rect 510120 996004 510126 996016
rect 560294 996004 560300 996016
rect 560352 996004 560358 996056
rect 144086 995976 144092 995988
rect 137572 995948 144092 995976
rect 89622 995800 89628 995852
rect 89680 995840 89686 995852
rect 92382 995840 92388 995852
rect 89680 995812 92388 995840
rect 89680 995800 89686 995812
rect 92382 995800 92388 995812
rect 92440 995800 92446 995852
rect 137370 995800 137376 995852
rect 137428 995840 137434 995852
rect 137572 995840 137600 995948
rect 144086 995936 144092 995948
rect 144144 995936 144150 995988
rect 307018 995976 307024 995988
rect 287026 995948 307024 995976
rect 143994 995908 144000 995920
rect 137940 995880 144000 995908
rect 137940 995852 137968 995880
rect 143994 995868 144000 995880
rect 144052 995868 144058 995920
rect 195422 995908 195428 995920
rect 189460 995880 195428 995908
rect 189460 995852 189488 995880
rect 195422 995868 195428 995880
rect 195480 995868 195486 995920
rect 137428 995812 137600 995840
rect 137428 995800 137434 995812
rect 137922 995800 137928 995852
rect 137980 995800 137986 995852
rect 139210 995800 139216 995852
rect 139268 995840 139274 995852
rect 139268 995812 142568 995840
rect 139268 995800 139274 995812
rect 91554 995732 91560 995784
rect 91612 995772 91618 995784
rect 92290 995772 92296 995784
rect 91612 995744 92296 995772
rect 91612 995732 91618 995744
rect 92290 995732 92296 995744
rect 92348 995732 92354 995784
rect 141050 995732 141056 995784
rect 141108 995772 141114 995784
rect 142540 995772 142568 995812
rect 142890 995800 142896 995852
rect 142948 995840 142954 995852
rect 143718 995840 143724 995852
rect 142948 995812 143724 995840
rect 142948 995800 142954 995812
rect 143718 995800 143724 995812
rect 143776 995800 143782 995852
rect 189442 995800 189448 995852
rect 189500 995800 189506 995852
rect 194318 995800 194324 995852
rect 194376 995840 194382 995852
rect 195330 995840 195336 995852
rect 194376 995812 195336 995840
rect 194376 995800 194382 995812
rect 195330 995800 195336 995812
rect 195388 995800 195394 995852
rect 240870 995800 240876 995852
rect 240928 995840 240934 995852
rect 246482 995840 246488 995852
rect 240928 995812 246488 995840
rect 240928 995800 240934 995812
rect 246482 995800 246488 995812
rect 246540 995800 246546 995852
rect 284386 995800 284392 995852
rect 284444 995840 284450 995852
rect 287026 995840 287054 995948
rect 307018 995936 307024 995948
rect 307076 995936 307082 995988
rect 364978 995936 364984 995988
rect 365036 995976 365042 995988
rect 382090 995976 382096 995988
rect 365036 995948 382096 995976
rect 365036 995936 365042 995948
rect 382090 995936 382096 995948
rect 382148 995936 382154 995988
rect 382274 995936 382280 995988
rect 382332 995976 382338 995988
rect 431954 995976 431960 995988
rect 382332 995948 431960 995976
rect 382332 995936 382338 995948
rect 431954 995936 431960 995948
rect 432012 995936 432018 995988
rect 436738 995936 436744 995988
rect 436796 995976 436802 995988
rect 510890 995976 510896 995988
rect 436796 995948 510896 995976
rect 436796 995936 436802 995948
rect 510890 995936 510896 995948
rect 510948 995936 510954 995988
rect 625430 995936 625436 995988
rect 625488 995976 625494 995988
rect 625488 995948 631456 995976
rect 625488 995936 625494 995948
rect 381538 995868 381544 995920
rect 381596 995908 381602 995920
rect 381596 995880 393314 995908
rect 381596 995868 381602 995880
rect 284444 995812 287054 995840
rect 284444 995800 284450 995812
rect 294874 995800 294880 995852
rect 294932 995840 294938 995852
rect 298186 995840 298192 995852
rect 294932 995812 298192 995840
rect 294932 995800 294938 995812
rect 298186 995800 298192 995812
rect 298244 995800 298250 995852
rect 383378 995800 383384 995852
rect 383436 995840 383442 995852
rect 385034 995840 385040 995852
rect 383436 995812 385040 995840
rect 383436 995800 383442 995812
rect 385034 995800 385040 995812
rect 385092 995800 385098 995852
rect 393286 995840 393314 995880
rect 523862 995868 523868 995920
rect 523920 995908 523926 995920
rect 523920 995880 528554 995908
rect 523920 995868 523926 995880
rect 528526 995852 528554 995880
rect 625890 995868 625896 995920
rect 625948 995908 625954 995920
rect 625948 995880 630904 995908
rect 625948 995868 625954 995880
rect 630876 995852 630904 995880
rect 393590 995840 393596 995852
rect 393286 995812 393596 995840
rect 393590 995800 393596 995812
rect 393648 995800 393654 995852
rect 396626 995800 396632 995852
rect 396684 995840 396690 995852
rect 400122 995840 400128 995852
rect 396684 995812 400128 995840
rect 396684 995800 396690 995812
rect 400122 995800 400128 995812
rect 400180 995800 400186 995852
rect 472526 995800 472532 995852
rect 472584 995840 472590 995852
rect 477678 995840 477684 995852
rect 472584 995812 477684 995840
rect 472584 995800 472590 995812
rect 477678 995800 477684 995812
rect 477736 995800 477742 995852
rect 520826 995800 520832 995852
rect 520884 995840 520890 995852
rect 527910 995840 527916 995852
rect 520884 995812 527916 995840
rect 520884 995800 520890 995812
rect 527910 995800 527916 995812
rect 527968 995800 527974 995852
rect 528526 995812 528560 995852
rect 528554 995800 528560 995812
rect 528612 995800 528618 995852
rect 536834 995800 536840 995852
rect 536892 995840 536898 995852
rect 540330 995840 540336 995852
rect 536892 995812 540336 995840
rect 536892 995800 536898 995812
rect 540330 995800 540336 995812
rect 540388 995800 540394 995852
rect 625798 995800 625804 995852
rect 625856 995840 625862 995852
rect 626534 995840 626540 995852
rect 625856 995812 626540 995840
rect 625856 995800 625862 995812
rect 626534 995800 626540 995812
rect 626592 995800 626598 995852
rect 630858 995800 630864 995852
rect 630916 995800 630922 995852
rect 631428 995840 631456 995948
rect 631502 995840 631508 995852
rect 631428 995812 631508 995840
rect 631502 995800 631508 995812
rect 631560 995800 631566 995852
rect 143626 995772 143632 995784
rect 141108 995744 142154 995772
rect 142540 995744 143632 995772
rect 141108 995732 141114 995744
rect 86586 995664 86592 995716
rect 86644 995704 86650 995716
rect 92198 995704 92204 995716
rect 86644 995676 92204 995704
rect 86644 995664 86650 995676
rect 92198 995664 92204 995676
rect 92256 995664 92262 995716
rect 142126 995704 142154 995744
rect 143626 995732 143632 995744
rect 143684 995732 143690 995784
rect 192478 995732 192484 995784
rect 192536 995772 192542 995784
rect 195146 995772 195152 995784
rect 192536 995744 195152 995772
rect 192536 995732 192542 995744
rect 195146 995732 195152 995744
rect 195204 995732 195210 995784
rect 240042 995732 240048 995784
rect 240100 995772 240106 995784
rect 246666 995772 246672 995784
rect 240100 995744 246672 995772
rect 240100 995732 240106 995744
rect 246666 995732 246672 995744
rect 246724 995732 246730 995784
rect 297266 995732 297272 995784
rect 297324 995772 297330 995784
rect 298002 995772 298008 995784
rect 297324 995744 298008 995772
rect 297324 995732 297330 995744
rect 298002 995732 298008 995744
rect 298060 995732 298066 995784
rect 383654 995732 383660 995784
rect 383712 995772 383718 995784
rect 384390 995772 384396 995784
rect 383712 995744 384396 995772
rect 383712 995732 383718 995744
rect 384390 995732 384396 995744
rect 384448 995732 384454 995784
rect 472618 995732 472624 995784
rect 472676 995772 472682 995784
rect 473998 995772 474004 995784
rect 472676 995744 474004 995772
rect 472676 995732 472682 995744
rect 473998 995732 474004 995744
rect 474056 995732 474062 995784
rect 516042 995732 516048 995784
rect 516100 995772 516106 995784
rect 516686 995772 516692 995784
rect 516100 995744 516692 995772
rect 516100 995732 516106 995744
rect 516686 995732 516692 995744
rect 516744 995732 516750 995784
rect 524046 995732 524052 995784
rect 524104 995772 524110 995784
rect 524782 995772 524788 995784
rect 524104 995744 524788 995772
rect 524104 995732 524110 995744
rect 524782 995732 524788 995744
rect 524840 995732 524846 995784
rect 625706 995732 625712 995784
rect 625764 995772 625770 995784
rect 627178 995772 627184 995784
rect 625764 995744 627184 995772
rect 625764 995732 625770 995744
rect 627178 995732 627184 995744
rect 627236 995732 627242 995784
rect 143902 995704 143908 995716
rect 142126 995676 143908 995704
rect 143902 995664 143908 995676
rect 143960 995664 143966 995716
rect 190638 995664 190644 995716
rect 190696 995704 190702 995716
rect 195698 995704 195704 995716
rect 190696 995676 195704 995704
rect 190696 995664 190702 995676
rect 195698 995664 195704 995676
rect 195756 995664 195762 995716
rect 245562 995664 245568 995716
rect 245620 995704 245626 995716
rect 246758 995704 246764 995716
rect 245620 995676 246764 995704
rect 245620 995664 245626 995676
rect 246758 995664 246764 995676
rect 246816 995664 246822 995716
rect 383470 995664 383476 995716
rect 383528 995704 383534 995716
rect 385678 995704 385684 995716
rect 383528 995676 385684 995704
rect 383528 995664 383534 995676
rect 385678 995664 385684 995676
rect 385736 995664 385742 995716
rect 472434 995664 472440 995716
rect 472492 995704 472498 995716
rect 473354 995704 473360 995716
rect 472492 995676 473360 995704
rect 472492 995664 472498 995676
rect 473354 995664 473360 995676
rect 473412 995664 473418 995716
rect 523770 995664 523776 995716
rect 523828 995704 523834 995716
rect 529750 995704 529756 995716
rect 523828 995676 529756 995704
rect 523828 995664 523834 995676
rect 529750 995664 529756 995676
rect 529808 995664 529814 995716
rect 625614 995664 625620 995716
rect 625672 995704 625678 995716
rect 630214 995704 630220 995716
rect 625672 995676 630220 995704
rect 625672 995664 625678 995676
rect 630214 995664 630220 995676
rect 630272 995664 630278 995716
rect 55858 995596 55864 995648
rect 55916 995636 55922 995648
rect 107746 995636 107752 995648
rect 55916 995608 107752 995636
rect 55916 995596 55922 995608
rect 107746 995596 107752 995608
rect 107804 995596 107810 995648
rect 243262 995596 243268 995648
rect 243320 995636 243326 995648
rect 246850 995636 246856 995648
rect 243320 995608 246856 995636
rect 243320 995596 243326 995608
rect 246850 995596 246856 995608
rect 246908 995596 246914 995648
rect 279326 995596 279332 995648
rect 279384 995636 279390 995648
rect 316402 995636 316408 995648
rect 279384 995608 316408 995636
rect 279384 995596 279390 995608
rect 316402 995596 316408 995608
rect 316460 995596 316466 995648
rect 472710 995596 472716 995648
rect 472768 995636 472774 995648
rect 476390 995636 476396 995648
rect 472768 995608 476396 995636
rect 472768 995596 472774 995608
rect 476390 995596 476396 995608
rect 476448 995596 476454 995648
rect 515950 995596 515956 995648
rect 516008 995636 516014 995648
rect 516686 995636 516692 995648
rect 516008 995608 516692 995636
rect 516008 995596 516014 995608
rect 516686 995596 516692 995608
rect 516744 995596 516750 995648
rect 559558 995596 559564 995648
rect 559616 995636 559622 995648
rect 661678 995636 661684 995648
rect 559616 995608 661684 995636
rect 559616 995596 559622 995608
rect 661678 995596 661684 995608
rect 661736 995596 661742 995648
rect 472342 995528 472348 995580
rect 472400 995568 472406 995580
rect 474734 995568 474740 995580
rect 472400 995540 474740 995568
rect 472400 995528 472406 995540
rect 474734 995528 474740 995540
rect 474792 995528 474798 995580
rect 625522 995528 625528 995580
rect 625580 995568 625586 995580
rect 627914 995568 627920 995580
rect 625580 995540 627920 995568
rect 625580 995528 625586 995540
rect 627914 995528 627920 995540
rect 627972 995528 627978 995580
rect 369210 995460 369216 995512
rect 369268 995500 369274 995512
rect 372338 995500 372344 995512
rect 369268 995472 372344 995500
rect 369268 995460 369274 995472
rect 372338 995460 372344 995472
rect 372396 995460 372402 995512
rect 513282 995460 513288 995512
rect 513340 995500 513346 995512
rect 516686 995500 516692 995512
rect 513340 995472 516692 995500
rect 513340 995460 513346 995472
rect 516686 995460 516692 995472
rect 516744 995460 516750 995512
rect 370774 995324 370780 995376
rect 370832 995364 370838 995376
rect 372338 995364 372344 995376
rect 370832 995336 372344 995364
rect 370832 995324 370838 995336
rect 372338 995324 372344 995336
rect 372396 995324 372402 995376
rect 438762 995324 438768 995376
rect 438820 995364 438826 995376
rect 439682 995364 439688 995376
rect 438820 995336 439688 995364
rect 438820 995324 438826 995336
rect 439682 995324 439688 995336
rect 439740 995324 439746 995376
rect 515214 995324 515220 995376
rect 515272 995364 515278 995376
rect 516686 995364 516692 995376
rect 515272 995336 516692 995364
rect 515272 995324 515278 995336
rect 516686 995324 516692 995336
rect 516744 995324 516750 995376
rect 522298 995256 522304 995308
rect 522356 995296 522362 995308
rect 537386 995296 537392 995308
rect 522356 995268 537392 995296
rect 522356 995256 522362 995268
rect 537386 995256 537392 995268
rect 537444 995256 537450 995308
rect 81342 995188 81348 995240
rect 81400 995228 81406 995240
rect 92658 995228 92664 995240
rect 81400 995200 92664 995228
rect 81400 995188 81406 995200
rect 92658 995188 92664 995200
rect 92716 995188 92722 995240
rect 183508 995188 183514 995240
rect 183566 995228 183572 995240
rect 195514 995228 195520 995240
rect 183566 995200 195520 995228
rect 183566 995188 183572 995200
rect 195514 995188 195520 995200
rect 195572 995188 195578 995240
rect 239260 995188 239266 995240
rect 239318 995228 239324 995240
rect 249150 995228 249156 995240
rect 239318 995200 249156 995228
rect 239318 995188 239324 995200
rect 249150 995188 249156 995200
rect 249208 995188 249214 995240
rect 370774 995188 370780 995240
rect 370832 995228 370838 995240
rect 372338 995228 372344 995240
rect 370832 995200 372344 995228
rect 370832 995188 370838 995200
rect 372338 995188 372344 995200
rect 372396 995188 372402 995240
rect 509206 995200 518894 995228
rect 77662 995120 77668 995172
rect 77720 995160 77726 995172
rect 92566 995160 92572 995172
rect 77720 995132 92572 995160
rect 77720 995120 77726 995132
rect 92566 995120 92572 995132
rect 92624 995120 92630 995172
rect 133414 995120 133420 995172
rect 133472 995160 133478 995172
rect 144178 995160 144184 995172
rect 133472 995132 144184 995160
rect 133472 995120 133478 995132
rect 144178 995120 144184 995132
rect 144236 995120 144242 995172
rect 180150 995120 180156 995172
rect 180208 995160 180214 995172
rect 195974 995160 195980 995172
rect 180208 995132 195980 995160
rect 180208 995120 180214 995132
rect 195974 995120 195980 995132
rect 196032 995120 196038 995172
rect 235902 995120 235908 995172
rect 235960 995160 235966 995172
rect 247126 995160 247132 995172
rect 235960 995132 247132 995160
rect 235960 995120 235966 995132
rect 247126 995120 247132 995132
rect 247184 995120 247190 995172
rect 287146 995120 287152 995172
rect 287204 995160 287210 995172
rect 304442 995160 304448 995172
rect 287204 995132 304448 995160
rect 287204 995120 287210 995132
rect 304442 995120 304448 995132
rect 304500 995120 304506 995172
rect 504266 995120 504272 995172
rect 504324 995160 504330 995172
rect 509206 995160 509234 995200
rect 504324 995132 509234 995160
rect 504324 995120 504330 995132
rect 515214 995120 515220 995172
rect 515272 995160 515278 995172
rect 516686 995160 516692 995172
rect 515272 995132 516692 995160
rect 515272 995120 515278 995132
rect 516686 995120 516692 995132
rect 516744 995120 516750 995172
rect 518866 995160 518894 995200
rect 574738 995188 574744 995240
rect 574796 995228 574802 995240
rect 636148 995228 636154 995240
rect 574796 995200 636154 995228
rect 574796 995188 574802 995200
rect 636148 995188 636154 995200
rect 636206 995188 636212 995240
rect 533706 995160 533712 995172
rect 518866 995132 533712 995160
rect 533706 995120 533712 995132
rect 533764 995120 533770 995172
rect 620278 995120 620284 995172
rect 620336 995160 620342 995172
rect 638954 995160 638960 995172
rect 620336 995132 638960 995160
rect 620336 995120 620342 995132
rect 638954 995120 638960 995132
rect 639012 995120 639018 995172
rect 78306 995052 78312 995104
rect 78364 995092 78370 995104
rect 97258 995092 97264 995104
rect 78364 995064 97264 995092
rect 78364 995052 78370 995064
rect 97258 995052 97264 995064
rect 97316 995052 97322 995104
rect 128446 995052 128452 995104
rect 128504 995092 128510 995104
rect 154574 995092 154580 995104
rect 128504 995064 154580 995092
rect 128504 995052 128510 995064
rect 154574 995052 154580 995064
rect 154632 995052 154638 995104
rect 180610 995052 180616 995104
rect 180668 995092 180674 995104
rect 202138 995092 202144 995104
rect 180668 995064 202144 995092
rect 180668 995052 180674 995064
rect 202138 995052 202144 995064
rect 202196 995052 202202 995104
rect 217410 995052 217416 995104
rect 217468 995092 217474 995104
rect 218882 995092 218888 995104
rect 217468 995064 218888 995092
rect 217468 995052 217474 995064
rect 218882 995052 218888 995064
rect 218940 995052 218946 995104
rect 231578 995052 231584 995104
rect 231636 995092 231642 995104
rect 251542 995092 251548 995104
rect 231636 995064 251548 995092
rect 231636 995052 231642 995064
rect 251542 995052 251548 995064
rect 251600 995052 251606 995104
rect 286502 995052 286508 995104
rect 286560 995092 286566 995104
rect 305638 995092 305644 995104
rect 286560 995064 305644 995092
rect 286560 995052 286566 995064
rect 305638 995052 305644 995064
rect 305696 995052 305702 995104
rect 460198 995052 460204 995104
rect 460256 995092 460262 995104
rect 482278 995092 482284 995104
rect 460256 995064 482284 995092
rect 460256 995052 460262 995064
rect 482278 995052 482284 995064
rect 482336 995052 482342 995104
rect 504358 995052 504364 995104
rect 504416 995092 504422 995104
rect 534350 995092 534356 995104
rect 504416 995064 534356 995092
rect 504416 995052 504422 995064
rect 534350 995052 534356 995064
rect 534408 995052 534414 995104
rect 568666 995052 568672 995104
rect 568724 995092 568730 995104
rect 634814 995092 634820 995104
rect 568724 995064 634820 995092
rect 568724 995052 568730 995064
rect 634814 995052 634820 995064
rect 634872 995052 634878 995104
rect 77018 994984 77024 995036
rect 77076 995024 77082 995036
rect 106642 995024 106648 995036
rect 77076 994996 106648 995024
rect 77076 994984 77082 994996
rect 106642 994984 106648 994996
rect 106700 994984 106706 995036
rect 165982 994984 165988 995036
rect 166040 995024 166046 995036
rect 167546 995024 167552 995036
rect 166040 994996 167552 995024
rect 166040 994984 166046 994996
rect 167546 994984 167552 994996
rect 167604 994984 167610 995036
rect 183278 994984 183284 995036
rect 183336 995024 183342 995036
rect 208394 995024 208400 995036
rect 183336 994996 208400 995024
rect 183336 994984 183342 994996
rect 208394 994984 208400 994996
rect 208452 994984 208458 995036
rect 232866 994984 232872 995036
rect 232924 995024 232930 995036
rect 257338 995024 257344 995036
rect 232924 994996 257344 995024
rect 232924 994984 232930 994996
rect 257338 994984 257344 994996
rect 257396 994984 257402 995036
rect 282822 994984 282828 995036
rect 282880 995024 282886 995036
rect 311894 995024 311900 995036
rect 282880 994996 311900 995024
rect 282880 994984 282886 994996
rect 311894 994984 311900 994996
rect 311952 994984 311958 995036
rect 357066 994984 357072 995036
rect 357124 995024 357130 995036
rect 398834 995024 398840 995036
rect 357124 994996 398840 995024
rect 357124 994984 357130 994996
rect 398834 994984 398840 994996
rect 398892 994984 398898 995036
rect 457438 994984 457444 995036
rect 457496 995024 457502 995036
rect 485958 995024 485964 995036
rect 457496 994996 485964 995024
rect 457496 994984 457502 994996
rect 485958 994984 485964 994996
rect 486016 994984 486022 995036
rect 499206 994984 499212 995036
rect 499264 995024 499270 995036
rect 535546 995024 535552 995036
rect 499264 994996 535552 995024
rect 499264 994984 499270 994996
rect 535546 994984 535552 994996
rect 535604 994984 535610 995036
rect 556154 994984 556160 995036
rect 556212 995024 556218 995036
rect 637022 995024 637028 995036
rect 556212 994996 637028 995024
rect 556212 994984 556218 994996
rect 637022 994984 637028 994996
rect 637080 994984 637086 995036
rect 440234 994236 440240 994288
rect 440292 994276 440298 994288
rect 446122 994276 446128 994288
rect 440292 994248 446128 994276
rect 440292 994236 440298 994248
rect 446122 994236 446128 994248
rect 446180 994236 446186 994288
rect 562502 993012 562508 993064
rect 562560 993052 562566 993064
rect 660298 993052 660304 993064
rect 562560 993024 660304 993052
rect 562560 993012 562566 993024
rect 660298 993012 660304 993024
rect 660356 993012 660362 993064
rect 88334 992944 88340 992996
rect 88392 992984 88398 992996
rect 111794 992984 111800 992996
rect 88392 992956 111800 992984
rect 88392 992944 88398 992956
rect 111794 992944 111800 992956
rect 111852 992944 111858 992996
rect 498010 992944 498016 992996
rect 498068 992984 498074 992996
rect 666646 992984 666652 992996
rect 498068 992956 666652 992984
rect 498068 992944 498074 992956
rect 666646 992944 666652 992956
rect 666704 992944 666710 992996
rect 46198 992876 46204 992928
rect 46256 992916 46262 992928
rect 110506 992916 110512 992928
rect 46256 992888 110512 992916
rect 46256 992876 46262 992888
rect 110506 992876 110512 992888
rect 110564 992876 110570 992928
rect 245654 992876 245660 992928
rect 245712 992916 245718 992928
rect 251450 992916 251456 992928
rect 245712 992888 251456 992916
rect 245712 992876 245718 992888
rect 251450 992876 251456 992888
rect 251508 992876 251514 992928
rect 353110 992876 353116 992928
rect 353168 992916 353174 992928
rect 666830 992916 666836 992928
rect 353168 992888 666836 992916
rect 353168 992876 353174 992888
rect 666830 992876 666836 992888
rect 666888 992876 666894 992928
rect 560938 991652 560944 991704
rect 560996 991692 561002 991704
rect 658918 991692 658924 991704
rect 560996 991664 658924 991692
rect 560996 991652 561002 991664
rect 658918 991652 658924 991664
rect 658976 991652 658982 991704
rect 549162 991584 549168 991636
rect 549220 991624 549226 991636
rect 666554 991624 666560 991636
rect 549220 991596 666560 991624
rect 549220 991584 549226 991596
rect 666554 991584 666560 991596
rect 666612 991584 666618 991636
rect 367830 991516 367836 991568
rect 367888 991556 367894 991568
rect 381630 991556 381636 991568
rect 367888 991528 381636 991556
rect 367888 991516 367894 991528
rect 381630 991516 381636 991528
rect 381688 991516 381694 991568
rect 420730 991516 420736 991568
rect 420788 991556 420794 991568
rect 666738 991556 666744 991568
rect 420788 991528 666744 991556
rect 420788 991516 420794 991528
rect 666738 991516 666744 991528
rect 666796 991516 666802 991568
rect 44818 991448 44824 991500
rect 44876 991488 44882 991500
rect 107930 991488 107936 991500
rect 44876 991460 107936 991488
rect 44876 991448 44882 991460
rect 107930 991448 107936 991460
rect 107988 991448 107994 991500
rect 203150 991448 203156 991500
rect 203208 991488 203214 991500
rect 213914 991488 213920 991500
rect 203208 991460 213920 991488
rect 203208 991448 203214 991460
rect 213914 991448 213920 991460
rect 213972 991448 213978 991500
rect 215938 991448 215944 991500
rect 215996 991488 216002 991500
rect 235626 991488 235632 991500
rect 215996 991460 235632 991488
rect 215996 991448 216002 991460
rect 235626 991448 235632 991460
rect 235684 991448 235690 991500
rect 303522 991448 303528 991500
rect 303580 991488 303586 991500
rect 665450 991488 665456 991500
rect 303580 991460 665456 991488
rect 303580 991448 303586 991460
rect 665450 991448 665456 991460
rect 665508 991448 665514 991500
rect 47578 990088 47584 990140
rect 47636 990128 47642 990140
rect 109034 990128 109040 990140
rect 47636 990100 109040 990128
rect 47636 990088 47642 990100
rect 109034 990088 109040 990100
rect 109092 990088 109098 990140
rect 138290 990088 138296 990140
rect 138348 990128 138354 990140
rect 162854 990128 162860 990140
rect 138348 990100 162860 990128
rect 138348 990088 138354 990100
rect 162854 990088 162860 990100
rect 162912 990088 162918 990140
rect 269758 990088 269764 990140
rect 269816 990128 269822 990140
rect 300486 990128 300492 990140
rect 269816 990100 300492 990128
rect 269816 990088 269822 990100
rect 300486 990088 300492 990100
rect 300544 990088 300550 990140
rect 370498 990088 370504 990140
rect 370556 990128 370562 990140
rect 430298 990128 430304 990140
rect 370556 990100 430304 990128
rect 370556 990088 370562 990100
rect 430298 990088 430304 990100
rect 430356 990088 430362 990140
rect 435358 990088 435364 990140
rect 435416 990128 435422 990140
rect 478966 990128 478972 990140
rect 435416 990100 478972 990128
rect 435416 990088 435422 990100
rect 478966 990088 478972 990100
rect 479024 990088 479030 990140
rect 514018 990088 514024 990140
rect 514076 990128 514082 990140
rect 560110 990128 560116 990140
rect 514076 990100 560116 990128
rect 514076 990088 514082 990100
rect 560110 990088 560116 990100
rect 560168 990088 560174 990140
rect 562318 990088 562324 990140
rect 562376 990128 562382 990140
rect 663058 990128 663064 990140
rect 562376 990100 663064 990128
rect 562376 990088 562382 990100
rect 663058 990088 663064 990100
rect 663116 990088 663122 990140
rect 566458 988728 566464 988780
rect 566516 988768 566522 988780
rect 592494 988768 592500 988780
rect 566516 988740 592500 988768
rect 566516 988728 566522 988740
rect 592494 988728 592500 988740
rect 592552 988728 592558 988780
rect 330478 987368 330484 987420
rect 330536 987408 330542 987420
rect 365438 987408 365444 987420
rect 330536 987380 365444 987408
rect 330536 987368 330542 987380
rect 365438 987368 365444 987380
rect 365496 987368 365502 987420
rect 512638 987368 512644 987420
rect 512696 987408 512702 987420
rect 543826 987408 543832 987420
rect 512696 987380 543832 987408
rect 512696 987368 512702 987380
rect 543826 987368 543832 987380
rect 543884 987368 543890 987420
rect 565078 987368 565084 987420
rect 565136 987408 565142 987420
rect 624970 987408 624976 987420
rect 565136 987380 624976 987408
rect 565136 987368 565142 987380
rect 624970 987368 624976 987380
rect 625028 987368 625034 987420
rect 88334 986620 88340 986672
rect 88392 986660 88398 986672
rect 89622 986660 89628 986672
rect 88392 986632 89628 986660
rect 88392 986620 88398 986632
rect 89622 986620 89628 986632
rect 89680 986620 89686 986672
rect 265618 986620 265624 986672
rect 265676 986660 265682 986672
rect 268102 986660 268108 986672
rect 265676 986632 268108 986660
rect 265676 986620 265682 986632
rect 268102 986620 268108 986632
rect 268160 986620 268166 986672
rect 367738 986008 367744 986060
rect 367796 986048 367802 986060
rect 397822 986048 397828 986060
rect 367796 986020 397828 986048
rect 367796 986008 367802 986020
rect 397822 986008 397828 986020
rect 397880 986008 397886 986060
rect 73430 985940 73436 985992
rect 73488 985980 73494 985992
rect 102778 985980 102784 985992
rect 73488 985952 102784 985980
rect 73488 985940 73494 985952
rect 102778 985940 102784 985952
rect 102836 985940 102842 985992
rect 266998 985940 267004 985992
rect 267056 985980 267062 985992
rect 284294 985980 284300 985992
rect 267056 985952 284300 985980
rect 267056 985940 267062 985952
rect 284294 985940 284300 985952
rect 284352 985940 284358 985992
rect 318058 985940 318064 985992
rect 318116 985980 318122 985992
rect 349154 985980 349160 985992
rect 318116 985952 349160 985980
rect 318116 985940 318122 985952
rect 349154 985940 349160 985952
rect 349212 985940 349218 985992
rect 369118 985940 369124 985992
rect 369176 985980 369182 985992
rect 414106 985980 414112 985992
rect 369176 985952 414112 985980
rect 369176 985940 369182 985952
rect 414106 985940 414112 985952
rect 414164 985940 414170 985992
rect 467098 985940 467104 985992
rect 467156 985980 467162 985992
rect 495158 985980 495164 985992
rect 467156 985952 495164 985980
rect 467156 985940 467162 985952
rect 495158 985940 495164 985952
rect 495216 985940 495222 985992
rect 571978 985940 571984 985992
rect 572036 985980 572042 985992
rect 608778 985980 608784 985992
rect 572036 985952 608784 985980
rect 572036 985940 572042 985952
rect 608778 985940 608784 985952
rect 608836 985940 608842 985992
rect 163498 985872 163504 985924
rect 163556 985912 163562 985924
rect 170766 985912 170772 985924
rect 163556 985884 170772 985912
rect 163556 985872 163562 985884
rect 170766 985872 170772 985884
rect 170824 985872 170830 985924
rect 520918 985736 520924 985788
rect 520976 985776 520982 985788
rect 527634 985776 527640 985788
rect 520976 985748 527640 985776
rect 520976 985736 520982 985748
rect 527634 985736 527640 985748
rect 527692 985736 527698 985788
rect 280798 984784 280804 984836
rect 280856 984824 280862 984836
rect 649994 984824 650000 984836
rect 280856 984796 650000 984824
rect 280856 984784 280862 984796
rect 649994 984784 650000 984796
rect 650052 984784 650058 984836
rect 228358 984716 228364 984768
rect 228416 984756 228422 984768
rect 651374 984756 651380 984768
rect 228416 984728 651380 984756
rect 228416 984716 228422 984728
rect 651374 984716 651380 984728
rect 651432 984716 651438 984768
rect 177298 984648 177304 984700
rect 177356 984688 177362 984700
rect 650086 984688 650092 984700
rect 177356 984660 650092 984688
rect 177356 984648 177362 984660
rect 650086 984648 650092 984660
rect 650144 984648 650150 984700
rect 126238 984580 126244 984632
rect 126296 984620 126302 984632
rect 651466 984620 651472 984632
rect 126296 984592 651472 984620
rect 126296 984580 126302 984592
rect 651466 984580 651472 984592
rect 651524 984580 651530 984632
rect 42702 975672 42708 975724
rect 42760 975712 42766 975724
rect 62114 975712 62120 975724
rect 42760 975684 62120 975712
rect 42760 975672 42766 975684
rect 62114 975672 62120 975684
rect 62172 975672 62178 975724
rect 651650 975672 651656 975724
rect 651708 975712 651714 975724
rect 672718 975712 672724 975724
rect 651708 975684 672724 975712
rect 651708 975672 651714 975684
rect 672718 975672 672724 975684
rect 672776 975672 672782 975724
rect 42150 967240 42156 967292
rect 42208 967280 42214 967292
rect 42702 967280 42708 967292
rect 42208 967252 42708 967280
rect 42208 967240 42214 967252
rect 42702 967240 42708 967252
rect 42760 967240 42766 967292
rect 42150 963976 42156 964028
rect 42208 964016 42214 964028
rect 42794 964016 42800 964028
rect 42208 963988 42800 964016
rect 42208 963976 42214 963988
rect 42794 963976 42800 963988
rect 42852 963976 42858 964028
rect 42150 962820 42156 962872
rect 42208 962860 42214 962872
rect 42886 962860 42892 962872
rect 42208 962832 42892 962860
rect 42208 962820 42214 962832
rect 42886 962820 42892 962832
rect 42944 962820 42950 962872
rect 44910 961868 44916 961920
rect 44968 961908 44974 961920
rect 62114 961908 62120 961920
rect 44968 961880 62120 961908
rect 44968 961868 44974 961880
rect 62114 961868 62120 961880
rect 62172 961868 62178 961920
rect 669958 961868 669964 961920
rect 670016 961908 670022 961920
rect 674834 961908 674840 961920
rect 670016 961880 674840 961908
rect 670016 961868 670022 961880
rect 674834 961868 674840 961880
rect 674892 961868 674898 961920
rect 675018 961324 675024 961376
rect 675076 961364 675082 961376
rect 675386 961364 675392 961376
rect 675076 961336 675392 961364
rect 675076 961324 675082 961336
rect 675386 961324 675392 961336
rect 675444 961324 675450 961376
rect 42058 959692 42064 959744
rect 42116 959732 42122 959744
rect 44174 959732 44180 959744
rect 42116 959704 44180 959732
rect 42116 959692 42122 959704
rect 44174 959692 44180 959704
rect 44232 959692 44238 959744
rect 42150 959080 42156 959132
rect 42208 959120 42214 959132
rect 42978 959120 42984 959132
rect 42208 959092 42984 959120
rect 42208 959080 42214 959092
rect 42978 959080 42984 959092
rect 43036 959080 43042 959132
rect 674742 958196 674748 958248
rect 674800 958236 674806 958248
rect 675386 958236 675392 958248
rect 674800 958208 675392 958236
rect 674800 958196 674806 958208
rect 675386 958196 675392 958208
rect 675444 958196 675450 958248
rect 659010 957788 659016 957840
rect 659068 957828 659074 957840
rect 675018 957828 675024 957840
rect 659068 957800 675024 957828
rect 659068 957788 659074 957800
rect 675018 957788 675024 957800
rect 675076 957788 675082 957840
rect 673362 956972 673368 957024
rect 673420 957012 673426 957024
rect 675386 957012 675392 957024
rect 673420 956984 675392 957012
rect 673420 956972 673426 956984
rect 675386 956972 675392 956984
rect 675444 956972 675450 957024
rect 673178 956088 673184 956140
rect 673236 956128 673242 956140
rect 675478 956128 675484 956140
rect 673236 956100 675484 956128
rect 673236 956088 673242 956100
rect 675478 956088 675484 956100
rect 675536 956088 675542 956140
rect 675018 955476 675024 955528
rect 675076 955516 675082 955528
rect 675478 955516 675484 955528
rect 675076 955488 675484 955516
rect 675076 955476 675082 955488
rect 675478 955476 675484 955488
rect 675536 955476 675542 955528
rect 42150 955340 42156 955392
rect 42208 955380 42214 955392
rect 42334 955380 42340 955392
rect 42208 955352 42340 955380
rect 42208 955340 42214 955352
rect 42334 955340 42340 955352
rect 42392 955340 42398 955392
rect 41782 954592 41788 954644
rect 41840 954592 41846 954644
rect 41800 954440 41828 954592
rect 41782 954388 41788 954440
rect 41840 954388 41846 954440
rect 32398 952824 32404 952876
rect 32456 952864 32462 952876
rect 41782 952864 41788 952876
rect 32456 952836 41788 952864
rect 32456 952824 32462 952836
rect 41782 952824 41788 952836
rect 41840 952824 41846 952876
rect 37918 952212 37924 952264
rect 37976 952252 37982 952264
rect 42334 952252 42340 952264
rect 37976 952224 42340 952252
rect 37976 952212 37982 952224
rect 42334 952212 42340 952224
rect 42392 952212 42398 952264
rect 675754 952008 675760 952060
rect 675812 952008 675818 952060
rect 675772 951788 675800 952008
rect 675754 951736 675760 951788
rect 675812 951736 675818 951788
rect 675754 949424 675760 949476
rect 675812 949464 675818 949476
rect 678238 949464 678244 949476
rect 675812 949436 678244 949464
rect 675812 949424 675818 949436
rect 678238 949424 678244 949436
rect 678296 949424 678302 949476
rect 651558 948064 651564 948116
rect 651616 948104 651622 948116
rect 674190 948104 674196 948116
rect 651616 948076 674196 948104
rect 651616 948064 651622 948076
rect 674190 948064 674196 948076
rect 674248 948064 674254 948116
rect 27614 947316 27620 947368
rect 27672 947356 27678 947368
rect 62114 947356 62120 947368
rect 27672 947328 62120 947356
rect 27672 947316 27678 947328
rect 62114 947316 62120 947328
rect 62172 947316 62178 947368
rect 35802 943236 35808 943288
rect 35860 943276 35866 943288
rect 45738 943276 45744 943288
rect 35860 943248 45744 943276
rect 35860 943236 35866 943248
rect 45738 943236 45744 943248
rect 45796 943236 45802 943288
rect 35710 943168 35716 943220
rect 35768 943208 35774 943220
rect 44910 943208 44916 943220
rect 35768 943180 44916 943208
rect 35768 943168 35774 943180
rect 44910 943168 44916 943180
rect 44968 943168 44974 943220
rect 652018 939768 652024 939820
rect 652076 939808 652082 939820
rect 676030 939808 676036 939820
rect 652076 939780 676036 939808
rect 652076 939768 652082 939780
rect 676030 939768 676036 939780
rect 676088 939768 676094 939820
rect 674190 939156 674196 939208
rect 674248 939196 674254 939208
rect 676030 939196 676036 939208
rect 674248 939168 676036 939196
rect 674248 939156 674254 939168
rect 676030 939156 676036 939168
rect 676088 939156 676094 939208
rect 672718 938680 672724 938732
rect 672776 938720 672782 938732
rect 676214 938720 676220 938732
rect 672776 938692 676220 938720
rect 672776 938680 672782 938692
rect 676214 938680 676220 938692
rect 676272 938680 676278 938732
rect 660298 938544 660304 938596
rect 660356 938584 660362 938596
rect 676030 938584 676036 938596
rect 660356 938556 676036 938584
rect 660356 938544 660362 938556
rect 676030 938544 676036 938556
rect 676088 938544 676094 938596
rect 674650 938272 674656 938324
rect 674708 938312 674714 938324
rect 676030 938312 676036 938324
rect 674708 938284 676036 938312
rect 674708 938272 674714 938284
rect 676030 938272 676036 938284
rect 676088 938272 676094 938324
rect 673822 937456 673828 937508
rect 673880 937496 673886 937508
rect 676030 937496 676036 937508
rect 673880 937468 676036 937496
rect 673880 937456 673886 937468
rect 676030 937456 676036 937468
rect 676088 937456 676094 937508
rect 663058 937320 663064 937372
rect 663116 937360 663122 937372
rect 676214 937360 676220 937372
rect 663116 937332 676220 937360
rect 663116 937320 663122 937332
rect 676214 937320 676220 937332
rect 676272 937320 676278 937372
rect 658918 937184 658924 937236
rect 658976 937224 658982 937236
rect 676214 937224 676220 937236
rect 658976 937196 676220 937224
rect 658976 937184 658982 937196
rect 676214 937184 676220 937196
rect 676272 937184 676278 937236
rect 45738 936980 45744 937032
rect 45796 937020 45802 937032
rect 62114 937020 62120 937032
rect 45796 936992 62120 937020
rect 45796 936980 45802 936992
rect 62114 936980 62120 936992
rect 62172 936980 62178 937032
rect 651558 936980 651564 937032
rect 651616 937020 651622 937032
rect 659010 937020 659016 937032
rect 651616 936992 659016 937020
rect 651616 936980 651622 936992
rect 659010 936980 659016 936992
rect 659068 936980 659074 937032
rect 672350 935756 672356 935808
rect 672408 935796 672414 935808
rect 676030 935796 676036 935808
rect 672408 935768 676036 935796
rect 672408 935756 672414 935768
rect 676030 935756 676036 935768
rect 676088 935756 676094 935808
rect 672810 935688 672816 935740
rect 672868 935728 672874 935740
rect 676122 935728 676128 935740
rect 672868 935700 676128 935728
rect 672868 935688 672874 935700
rect 676122 935688 676128 935700
rect 676180 935688 676186 935740
rect 661678 935620 661684 935672
rect 661736 935660 661742 935672
rect 676214 935660 676220 935672
rect 661736 935632 676220 935660
rect 661736 935620 661742 935632
rect 676214 935620 676220 935632
rect 676272 935620 676278 935672
rect 39942 932356 39948 932408
rect 40000 932396 40006 932408
rect 41690 932396 41696 932408
rect 40000 932368 41696 932396
rect 40000 932356 40006 932368
rect 41690 932356 41696 932368
rect 41748 932356 41754 932408
rect 41690 932152 41696 932204
rect 41748 932192 41754 932204
rect 47578 932192 47584 932204
rect 41748 932164 47584 932192
rect 41748 932152 41754 932164
rect 47578 932152 47584 932164
rect 47636 932152 47642 932204
rect 673178 931608 673184 931660
rect 673236 931648 673242 931660
rect 676030 931648 676036 931660
rect 673236 931620 676036 931648
rect 673236 931608 673242 931620
rect 676030 931608 676036 931620
rect 676088 931608 676094 931660
rect 674742 930724 674748 930776
rect 674800 930764 674806 930776
rect 676214 930764 676220 930776
rect 674800 930736 676220 930764
rect 674800 930724 674806 930736
rect 676214 930724 676220 930736
rect 676272 930724 676278 930776
rect 673362 930248 673368 930300
rect 673420 930288 673426 930300
rect 676214 930288 676220 930300
rect 673420 930260 676220 930288
rect 673420 930248 673426 930260
rect 676214 930248 676220 930260
rect 676272 930248 676278 930300
rect 671338 927392 671344 927444
rect 671396 927432 671402 927444
rect 683114 927432 683120 927444
rect 671396 927404 683120 927432
rect 671396 927392 671402 927404
rect 683114 927392 683120 927404
rect 683172 927392 683178 927444
rect 47670 923244 47676 923296
rect 47728 923284 47734 923296
rect 62114 923284 62120 923296
rect 47728 923256 62120 923284
rect 47728 923244 47734 923256
rect 62114 923244 62120 923256
rect 62172 923244 62178 923296
rect 651558 921816 651564 921868
rect 651616 921856 651622 921868
rect 670050 921856 670056 921868
rect 651616 921828 670056 921856
rect 651616 921816 651622 921828
rect 670050 921816 670056 921828
rect 670108 921816 670114 921868
rect 54478 909440 54484 909492
rect 54536 909480 54542 909492
rect 62114 909480 62120 909492
rect 54536 909452 62120 909480
rect 54536 909440 54542 909452
rect 62114 909440 62120 909452
rect 62172 909440 62178 909492
rect 651558 909440 651564 909492
rect 651616 909480 651622 909492
rect 661678 909480 661684 909492
rect 651616 909452 661684 909480
rect 651616 909440 651622 909452
rect 661678 909440 661684 909452
rect 661736 909440 661742 909492
rect 51718 896996 51724 897048
rect 51776 897036 51782 897048
rect 62114 897036 62120 897048
rect 51776 897008 62120 897036
rect 51776 896996 51782 897008
rect 62114 896996 62120 897008
rect 62172 896996 62178 897048
rect 651558 895636 651564 895688
rect 651616 895676 651622 895688
rect 660298 895676 660304 895688
rect 651616 895648 660304 895676
rect 651616 895636 651622 895648
rect 660298 895636 660304 895648
rect 660356 895636 660362 895688
rect 48958 884620 48964 884672
rect 49016 884660 49022 884672
rect 62114 884660 62120 884672
rect 49016 884632 62120 884660
rect 49016 884620 49022 884632
rect 62114 884620 62120 884632
rect 62172 884620 62178 884672
rect 674466 873536 674472 873588
rect 674524 873576 674530 873588
rect 675386 873576 675392 873588
rect 674524 873548 675392 873576
rect 674524 873536 674530 873548
rect 675386 873536 675392 873548
rect 675444 873536 675450 873588
rect 673178 872652 673184 872704
rect 673236 872692 673242 872704
rect 675386 872692 675392 872704
rect 673236 872664 675392 872692
rect 673236 872652 673242 872664
rect 675386 872652 675392 872664
rect 675444 872652 675450 872704
rect 674558 872176 674564 872228
rect 674616 872216 674622 872228
rect 675386 872216 675392 872228
rect 674616 872188 675392 872216
rect 674616 872176 674622 872188
rect 675386 872176 675392 872188
rect 675444 872176 675450 872228
rect 44818 870816 44824 870868
rect 44876 870856 44882 870868
rect 62114 870856 62120 870868
rect 44876 870828 62120 870856
rect 44876 870816 44882 870828
rect 62114 870816 62120 870828
rect 62172 870816 62178 870868
rect 674282 869796 674288 869848
rect 674340 869836 674346 869848
rect 675386 869836 675392 869848
rect 674340 869808 675392 869836
rect 674340 869796 674346 869808
rect 675386 869796 675392 869808
rect 675444 869796 675450 869848
rect 672994 869660 673000 869712
rect 673052 869700 673058 869712
rect 675386 869700 675392 869712
rect 673052 869672 675392 869700
rect 673052 869660 673058 869672
rect 675386 869660 675392 869672
rect 675444 869660 675450 869712
rect 673086 869592 673092 869644
rect 673144 869632 673150 869644
rect 674926 869632 674932 869644
rect 673144 869604 674932 869632
rect 673144 869592 673150 869604
rect 674926 869592 674932 869604
rect 674984 869592 674990 869644
rect 651558 869388 651564 869440
rect 651616 869428 651622 869440
rect 671430 869428 671436 869440
rect 651616 869400 671436 869428
rect 651616 869388 651622 869400
rect 671430 869388 671436 869400
rect 671488 869388 671494 869440
rect 674926 868708 674932 868760
rect 674984 868748 674990 868760
rect 675386 868748 675392 868760
rect 674984 868720 675392 868748
rect 674984 868708 674990 868720
rect 675386 868708 675392 868720
rect 675444 868708 675450 868760
rect 652018 868640 652024 868692
rect 652076 868680 652082 868692
rect 652076 868652 663794 868680
rect 652076 868640 652082 868652
rect 663766 868612 663794 868652
rect 674926 868612 674932 868624
rect 663766 868584 674932 868612
rect 674926 868572 674932 868584
rect 674984 868572 674990 868624
rect 674374 868504 674380 868556
rect 674432 868544 674438 868556
rect 675478 868544 675484 868556
rect 674432 868516 675484 868544
rect 674432 868504 674438 868516
rect 675478 868504 675484 868516
rect 675536 868504 675542 868556
rect 674926 866192 674932 866244
rect 674984 866232 674990 866244
rect 675386 866232 675392 866244
rect 674984 866204 675392 866232
rect 674984 866192 674990 866204
rect 675386 866192 675392 866204
rect 675444 866192 675450 866244
rect 672902 862792 672908 862844
rect 672960 862832 672966 862844
rect 675478 862832 675484 862844
rect 672960 862804 675484 862832
rect 672960 862792 672966 862804
rect 675478 862792 675484 862804
rect 675536 862792 675542 862844
rect 43622 858372 43628 858424
rect 43680 858412 43686 858424
rect 62114 858412 62120 858424
rect 43680 858384 62120 858412
rect 43680 858372 43686 858384
rect 62114 858372 62120 858384
rect 62172 858372 62178 858424
rect 651558 855584 651564 855636
rect 651616 855624 651622 855636
rect 664438 855624 664444 855636
rect 651616 855596 664444 855624
rect 651616 855584 651622 855596
rect 664438 855584 664444 855596
rect 664496 855584 664502 855636
rect 53098 844568 53104 844620
rect 53156 844608 53162 844620
rect 62114 844608 62120 844620
rect 53156 844580 62120 844608
rect 53156 844568 53162 844580
rect 62114 844568 62120 844580
rect 62172 844568 62178 844620
rect 651558 841780 651564 841832
rect 651616 841820 651622 841832
rect 663058 841820 663064 841832
rect 651616 841792 663064 841820
rect 651616 841780 651622 841792
rect 663058 841780 663064 841792
rect 663116 841780 663122 841832
rect 50338 832124 50344 832176
rect 50396 832164 50402 832176
rect 62114 832164 62120 832176
rect 50396 832136 62120 832164
rect 50396 832124 50402 832136
rect 62114 832124 62120 832136
rect 62172 832124 62178 832176
rect 651558 829404 651564 829456
rect 651616 829444 651622 829456
rect 658918 829444 658924 829456
rect 651616 829416 658924 829444
rect 651616 829404 651622 829416
rect 658918 829404 658924 829416
rect 658976 829404 658982 829456
rect 43530 818320 43536 818372
rect 43588 818360 43594 818372
rect 62114 818360 62120 818372
rect 43588 818332 62120 818360
rect 43588 818320 43594 818332
rect 62114 818320 62120 818332
rect 62172 818320 62178 818372
rect 41322 817504 41328 817556
rect 41380 817544 41386 817556
rect 48958 817544 48964 817556
rect 41380 817516 48964 817544
rect 41380 817504 41386 817516
rect 48958 817504 48964 817516
rect 49016 817504 49022 817556
rect 41230 817368 41236 817420
rect 41288 817408 41294 817420
rect 51718 817408 51724 817420
rect 41288 817380 51724 817408
rect 41288 817368 41294 817380
rect 51718 817368 51724 817380
rect 51776 817368 51782 817420
rect 651558 815600 651564 815652
rect 651616 815640 651622 815652
rect 665818 815640 665824 815652
rect 651616 815612 665824 815640
rect 651616 815600 651622 815612
rect 665818 815600 665824 815612
rect 665876 815600 665882 815652
rect 40770 811520 40776 811572
rect 40828 811560 40834 811572
rect 41782 811560 41788 811572
rect 40828 811532 41788 811560
rect 40828 811520 40834 811532
rect 41782 811520 41788 811532
rect 41840 811520 41846 811572
rect 39850 807236 39856 807288
rect 39908 807276 39914 807288
rect 41782 807276 41788 807288
rect 39908 807248 41788 807276
rect 39908 807236 39914 807248
rect 41782 807236 41788 807248
rect 41840 807236 41846 807288
rect 49050 805944 49056 805996
rect 49108 805984 49114 805996
rect 62114 805984 62120 805996
rect 49108 805956 62120 805984
rect 49108 805944 49114 805956
rect 62114 805944 62120 805956
rect 62172 805944 62178 805996
rect 42150 803836 42156 803888
rect 42208 803876 42214 803888
rect 42610 803876 42616 803888
rect 42208 803848 42616 803876
rect 42208 803836 42214 803848
rect 42610 803836 42616 803848
rect 42668 803836 42674 803888
rect 42058 803768 42064 803820
rect 42116 803808 42122 803820
rect 42702 803808 42708 803820
rect 42116 803780 42708 803808
rect 42116 803768 42122 803780
rect 42702 803768 42708 803780
rect 42760 803768 42766 803820
rect 651558 803156 651564 803208
rect 651616 803196 651622 803208
rect 672718 803196 672724 803208
rect 651616 803168 672724 803196
rect 651616 803156 651622 803168
rect 672718 803156 672724 803168
rect 672776 803156 672782 803208
rect 35158 801116 35164 801168
rect 35216 801156 35222 801168
rect 43070 801156 43076 801168
rect 35216 801128 43076 801156
rect 35216 801116 35222 801128
rect 43070 801116 43076 801128
rect 43128 801116 43134 801168
rect 32398 801048 32404 801100
rect 32456 801088 32462 801100
rect 42886 801088 42892 801100
rect 32456 801060 42892 801088
rect 32456 801048 32462 801060
rect 42886 801048 42892 801060
rect 42944 801048 42950 801100
rect 40770 800504 40776 800556
rect 40828 800544 40834 800556
rect 42978 800544 42984 800556
rect 40828 800516 42984 800544
rect 40828 800504 40834 800516
rect 42978 800504 42984 800516
rect 43036 800504 43042 800556
rect 42150 799960 42156 800012
rect 42208 800000 42214 800012
rect 42334 800000 42340 800012
rect 42208 799972 42340 800000
rect 42208 799960 42214 799972
rect 42334 799960 42340 799972
rect 42392 799960 42398 800012
rect 43162 799008 43168 799060
rect 43220 799048 43226 799060
rect 47670 799048 47676 799060
rect 43220 799020 47676 799048
rect 43220 799008 43226 799020
rect 47670 799008 47676 799020
rect 47728 799008 47734 799060
rect 42150 798124 42156 798176
rect 42208 798164 42214 798176
rect 42610 798164 42616 798176
rect 42208 798136 42616 798164
rect 42208 798124 42214 798136
rect 42610 798124 42616 798136
rect 42668 798124 42674 798176
rect 42150 797240 42156 797292
rect 42208 797280 42214 797292
rect 43162 797280 43168 797292
rect 42208 797252 43168 797280
rect 42208 797240 42214 797252
rect 43162 797240 43168 797252
rect 43220 797240 43226 797292
rect 42150 796288 42156 796340
rect 42208 796328 42214 796340
rect 42702 796328 42708 796340
rect 42208 796300 42708 796328
rect 42208 796288 42214 796300
rect 42702 796288 42708 796300
rect 42760 796288 42766 796340
rect 42702 796152 42708 796204
rect 42760 796192 42766 796204
rect 42886 796192 42892 796204
rect 42760 796164 42892 796192
rect 42760 796152 42766 796164
rect 42886 796152 42892 796164
rect 42944 796152 42950 796204
rect 42150 794996 42156 795048
rect 42208 795036 42214 795048
rect 42426 795036 42432 795048
rect 42208 795008 42432 795036
rect 42208 794996 42214 795008
rect 42426 794996 42432 795008
rect 42484 794996 42490 795048
rect 42886 794928 42892 794980
rect 42944 794968 42950 794980
rect 44358 794968 44364 794980
rect 42944 794940 44364 794968
rect 42944 794928 42950 794940
rect 44358 794928 44364 794940
rect 44416 794928 44422 794980
rect 42426 794860 42432 794912
rect 42484 794900 42490 794912
rect 42978 794900 42984 794912
rect 42484 794872 42984 794900
rect 42484 794860 42490 794872
rect 42978 794860 42984 794872
rect 43036 794860 43042 794912
rect 42150 794248 42156 794300
rect 42208 794288 42214 794300
rect 42702 794288 42708 794300
rect 42208 794260 42708 794288
rect 42208 794248 42214 794260
rect 42702 794248 42708 794260
rect 42760 794248 42766 794300
rect 42702 794112 42708 794164
rect 42760 794152 42766 794164
rect 43070 794152 43076 794164
rect 42760 794124 43076 794152
rect 42760 794112 42766 794124
rect 43070 794112 43076 794124
rect 43128 794112 43134 794164
rect 42150 793772 42156 793824
rect 42208 793812 42214 793824
rect 42886 793812 42892 793824
rect 42208 793784 42892 793812
rect 42208 793772 42214 793784
rect 42886 793772 42892 793784
rect 42944 793772 42950 793824
rect 54478 793500 54484 793552
rect 54536 793540 54542 793552
rect 62114 793540 62120 793552
rect 54536 793512 62120 793540
rect 54536 793500 54542 793512
rect 62114 793500 62120 793512
rect 62172 793500 62178 793552
rect 42150 793160 42156 793212
rect 42208 793200 42214 793212
rect 42426 793200 42432 793212
rect 42208 793172 42432 793200
rect 42208 793160 42214 793172
rect 42426 793160 42432 793172
rect 42484 793160 42490 793212
rect 42426 793024 42432 793076
rect 42484 793064 42490 793076
rect 42794 793064 42800 793076
rect 42484 793036 42800 793064
rect 42484 793024 42490 793036
rect 42794 793024 42800 793036
rect 42852 793024 42858 793076
rect 42150 790644 42156 790696
rect 42208 790684 42214 790696
rect 42794 790684 42800 790696
rect 42208 790656 42800 790684
rect 42208 790644 42214 790656
rect 42794 790644 42800 790656
rect 42852 790644 42858 790696
rect 42150 790100 42156 790152
rect 42208 790140 42214 790152
rect 42426 790140 42432 790152
rect 42208 790112 42432 790140
rect 42208 790100 42214 790112
rect 42426 790100 42432 790112
rect 42484 790100 42490 790152
rect 42150 789420 42156 789472
rect 42208 789460 42214 789472
rect 42334 789460 42340 789472
rect 42208 789432 42340 789460
rect 42208 789420 42214 789432
rect 42334 789420 42340 789432
rect 42392 789420 42398 789472
rect 651650 789352 651656 789404
rect 651708 789392 651714 789404
rect 661770 789392 661776 789404
rect 651708 789364 661776 789392
rect 651708 789352 651714 789364
rect 661770 789352 661776 789364
rect 661828 789352 661834 789404
rect 42150 788808 42156 788860
rect 42208 788848 42214 788860
rect 42702 788848 42708 788860
rect 42208 788820 42708 788848
rect 42208 788808 42214 788820
rect 42702 788808 42708 788820
rect 42760 788808 42766 788860
rect 670602 787992 670608 788044
rect 670660 788032 670666 788044
rect 675386 788032 675392 788044
rect 670660 788004 675392 788032
rect 670660 787992 670666 788004
rect 675386 787992 675392 788004
rect 675444 787992 675450 788044
rect 674190 787312 674196 787364
rect 674248 787352 674254 787364
rect 675386 787352 675392 787364
rect 674248 787324 675392 787352
rect 674248 787312 674254 787324
rect 675386 787312 675392 787324
rect 675444 787312 675450 787364
rect 42150 786972 42156 787024
rect 42208 787012 42214 787024
rect 42426 787012 42432 787024
rect 42208 786984 42432 787012
rect 42208 786972 42214 786984
rect 42426 786972 42432 786984
rect 42484 786972 42490 787024
rect 672626 786700 672632 786752
rect 672684 786740 672690 786752
rect 675386 786740 675392 786752
rect 672684 786712 675392 786740
rect 672684 786700 672690 786712
rect 675386 786700 675392 786712
rect 675444 786700 675450 786752
rect 42150 785612 42156 785664
rect 42208 785652 42214 785664
rect 42702 785652 42708 785664
rect 42208 785624 42708 785652
rect 42208 785612 42214 785624
rect 42702 785612 42708 785624
rect 42760 785612 42766 785664
rect 674006 784252 674012 784304
rect 674064 784292 674070 784304
rect 675386 784292 675392 784304
rect 674064 784264 675392 784292
rect 674064 784252 674070 784264
rect 675386 784252 675392 784264
rect 675444 784252 675450 784304
rect 673270 782892 673276 782944
rect 673328 782932 673334 782944
rect 675478 782932 675484 782944
rect 673328 782904 675484 782932
rect 673328 782892 673334 782904
rect 675478 782892 675484 782904
rect 675536 782892 675542 782944
rect 672534 780716 672540 780768
rect 672592 780756 672598 780768
rect 675478 780756 675484 780768
rect 672592 780728 675484 780756
rect 672592 780716 672598 780728
rect 675478 780716 675484 780728
rect 675536 780716 675542 780768
rect 673638 779968 673644 780020
rect 673696 780008 673702 780020
rect 675478 780008 675484 780020
rect 673696 779980 675484 780008
rect 673696 779968 673702 779980
rect 675478 779968 675484 779980
rect 675536 779968 675542 780020
rect 51718 779696 51724 779748
rect 51776 779736 51782 779748
rect 62114 779736 62120 779748
rect 51776 779708 62120 779736
rect 51776 779696 51782 779708
rect 62114 779696 62120 779708
rect 62172 779696 62178 779748
rect 658918 778948 658924 779000
rect 658976 778988 658982 779000
rect 674742 778988 674748 779000
rect 658976 778960 674748 778988
rect 658976 778948 658982 778960
rect 674742 778948 674748 778960
rect 674800 778948 674806 779000
rect 673914 778608 673920 778660
rect 673972 778648 673978 778660
rect 675478 778648 675484 778660
rect 673972 778620 675484 778648
rect 673972 778608 673978 778620
rect 675478 778608 675484 778620
rect 675536 778608 675542 778660
rect 672442 777316 672448 777368
rect 672500 777356 672506 777368
rect 675386 777356 675392 777368
rect 672500 777328 675392 777356
rect 672500 777316 672506 777328
rect 675386 777316 675392 777328
rect 675444 777316 675450 777368
rect 674742 777044 674748 777096
rect 674800 777084 674806 777096
rect 675386 777084 675392 777096
rect 674800 777056 675392 777084
rect 674800 777044 674806 777056
rect 675386 777044 675392 777056
rect 675444 777044 675450 777096
rect 651558 775548 651564 775600
rect 651616 775588 651622 775600
rect 658918 775588 658924 775600
rect 651616 775560 658924 775588
rect 651616 775548 651622 775560
rect 658918 775548 658924 775560
rect 658976 775548 658982 775600
rect 35802 774188 35808 774240
rect 35860 774228 35866 774240
rect 53098 774228 53104 774240
rect 35860 774200 53104 774228
rect 35860 774188 35866 774200
rect 53098 774188 53104 774200
rect 53156 774188 53162 774240
rect 672166 773576 672172 773628
rect 672224 773616 672230 773628
rect 675478 773616 675484 773628
rect 672224 773588 675484 773616
rect 672224 773576 672230 773588
rect 675478 773576 675484 773588
rect 675536 773576 675542 773628
rect 46198 767320 46204 767372
rect 46256 767360 46262 767372
rect 62114 767360 62120 767372
rect 46256 767332 62120 767360
rect 46256 767320 46262 767332
rect 62114 767320 62120 767332
rect 62172 767320 62178 767372
rect 651558 763172 651564 763224
rect 651616 763212 651622 763224
rect 664530 763212 664536 763224
rect 651616 763184 664536 763212
rect 651616 763172 651622 763184
rect 664530 763172 664536 763184
rect 664588 763172 664594 763224
rect 41506 761744 41512 761796
rect 41564 761784 41570 761796
rect 48958 761784 48964 761796
rect 41564 761756 48964 761784
rect 41564 761744 41570 761756
rect 48958 761744 48964 761756
rect 49016 761744 49022 761796
rect 670050 760792 670056 760844
rect 670108 760832 670114 760844
rect 676214 760832 676220 760844
rect 670108 760804 676220 760832
rect 670108 760792 670114 760804
rect 676214 760792 676220 760804
rect 676272 760792 676278 760844
rect 661678 760656 661684 760708
rect 661736 760696 661742 760708
rect 676122 760696 676128 760708
rect 661736 760668 676128 760696
rect 661736 760656 661742 760668
rect 676122 760656 676128 760668
rect 676180 760656 676186 760708
rect 660298 760520 660304 760572
rect 660356 760560 660362 760572
rect 676030 760560 676036 760572
rect 660356 760532 676036 760560
rect 660356 760520 660362 760532
rect 676030 760520 676036 760532
rect 676088 760520 676094 760572
rect 674650 760316 674656 760368
rect 674708 760356 674714 760368
rect 676030 760356 676036 760368
rect 674708 760328 676036 760356
rect 674708 760316 674714 760328
rect 676030 760316 676036 760328
rect 676088 760316 676094 760368
rect 31018 759636 31024 759688
rect 31076 759676 31082 759688
rect 41874 759676 41880 759688
rect 31076 759648 41880 759676
rect 31076 759636 31082 759648
rect 41874 759636 41880 759648
rect 41932 759636 41938 759688
rect 673822 759500 673828 759552
rect 673880 759540 673886 759552
rect 676030 759540 676036 759552
rect 673880 759512 676036 759540
rect 673880 759500 673886 759512
rect 676030 759500 676036 759512
rect 676088 759500 676094 759552
rect 673362 759092 673368 759144
rect 673420 759132 673426 759144
rect 676214 759132 676220 759144
rect 673420 759104 676220 759132
rect 673420 759092 673426 759104
rect 676214 759092 676220 759104
rect 676272 759092 676278 759144
rect 672258 759024 672264 759076
rect 672316 759064 672322 759076
rect 676030 759064 676036 759076
rect 672316 759036 676036 759064
rect 672316 759024 672322 759036
rect 676030 759024 676036 759036
rect 676088 759024 676094 759076
rect 33778 758480 33784 758532
rect 33836 758520 33842 758532
rect 42426 758520 42432 758532
rect 33836 758492 42432 758520
rect 33836 758480 33842 758492
rect 42426 758480 42432 758492
rect 42484 758480 42490 758532
rect 32490 758344 32496 758396
rect 32548 758384 32554 758396
rect 42702 758384 42708 758396
rect 32548 758356 42708 758384
rect 32548 758344 32554 758356
rect 42702 758344 42708 758356
rect 42760 758344 42766 758396
rect 32398 758276 32404 758328
rect 32456 758316 32462 758328
rect 43162 758316 43168 758328
rect 32456 758288 43168 758316
rect 32456 758276 32462 758288
rect 43162 758276 43168 758288
rect 43220 758276 43226 758328
rect 674650 758208 674656 758260
rect 674708 758248 674714 758260
rect 676030 758248 676036 758260
rect 674708 758220 676036 758248
rect 674708 758208 674714 758220
rect 676030 758208 676036 758220
rect 676088 758208 676094 758260
rect 41874 756984 41880 757036
rect 41932 756984 41938 757036
rect 41892 756764 41920 756984
rect 41874 756712 41880 756764
rect 41932 756712 41938 756764
rect 43254 756236 43260 756288
rect 43312 756276 43318 756288
rect 44818 756276 44824 756288
rect 43312 756248 44824 756276
rect 43312 756236 43318 756248
rect 44818 756236 44824 756248
rect 44876 756236 44882 756288
rect 674282 755556 674288 755608
rect 674340 755596 674346 755608
rect 676214 755596 676220 755608
rect 674340 755568 676220 755596
rect 674340 755556 674346 755568
rect 676214 755556 676220 755568
rect 676272 755556 676278 755608
rect 42426 755528 42432 755540
rect 42168 755500 42432 755528
rect 42168 755472 42196 755500
rect 42426 755488 42432 755500
rect 42484 755488 42490 755540
rect 42150 755420 42156 755472
rect 42208 755420 42214 755472
rect 42610 755216 42616 755268
rect 42668 755256 42674 755268
rect 43162 755256 43168 755268
rect 42668 755228 43168 755256
rect 42668 755216 42674 755228
rect 43162 755216 43168 755228
rect 43220 755216 43226 755268
rect 42150 755148 42156 755200
rect 42208 755148 42214 755200
rect 42168 754928 42196 755148
rect 672902 754944 672908 754996
rect 672960 754984 672966 754996
rect 676030 754984 676036 754996
rect 672960 754956 676036 754984
rect 672960 754944 672966 754956
rect 676030 754944 676036 754956
rect 676088 754944 676094 754996
rect 42150 754876 42156 754928
rect 42208 754876 42214 754928
rect 674466 754332 674472 754384
rect 674524 754372 674530 754384
rect 676214 754372 676220 754384
rect 674524 754344 676220 754372
rect 674524 754332 674530 754344
rect 676214 754332 676220 754344
rect 676272 754332 676278 754384
rect 42058 754060 42064 754112
rect 42116 754100 42122 754112
rect 43254 754100 43260 754112
rect 42116 754072 43260 754100
rect 42116 754060 42122 754072
rect 43254 754060 43260 754072
rect 43312 754060 43318 754112
rect 673178 753584 673184 753636
rect 673236 753624 673242 753636
rect 676030 753624 676036 753636
rect 673236 753596 676036 753624
rect 673236 753584 673242 753596
rect 676030 753584 676036 753596
rect 676088 753584 676094 753636
rect 44910 753516 44916 753568
rect 44968 753556 44974 753568
rect 62114 753556 62120 753568
rect 44968 753528 62120 753556
rect 44968 753516 44974 753528
rect 62114 753516 62120 753528
rect 62172 753516 62178 753568
rect 674374 753108 674380 753160
rect 674432 753148 674438 753160
rect 676214 753148 676220 753160
rect 674432 753120 676220 753148
rect 674432 753108 674438 753120
rect 676214 753108 676220 753120
rect 676272 753108 676278 753160
rect 674558 752700 674564 752752
rect 674616 752740 674622 752752
rect 676214 752740 676220 752752
rect 674616 752712 676220 752740
rect 674616 752700 674622 752712
rect 676214 752700 676220 752712
rect 676272 752700 676278 752752
rect 672994 752224 673000 752276
rect 673052 752264 673058 752276
rect 676214 752264 676220 752276
rect 673052 752236 676220 752264
rect 673052 752224 673058 752236
rect 676214 752224 676220 752236
rect 676272 752224 676278 752276
rect 43070 752088 43076 752140
rect 43128 752128 43134 752140
rect 44450 752128 44456 752140
rect 43128 752100 44456 752128
rect 43128 752088 43134 752100
rect 44450 752088 44456 752100
rect 44508 752088 44514 752140
rect 42150 751068 42156 751120
rect 42208 751108 42214 751120
rect 42978 751108 42984 751120
rect 42208 751080 42984 751108
rect 42208 751068 42214 751080
rect 42978 751068 42984 751080
rect 43036 751068 43042 751120
rect 673086 750864 673092 750916
rect 673144 750904 673150 750916
rect 676214 750904 676220 750916
rect 673144 750876 676220 750904
rect 673144 750864 673150 750876
rect 676214 750864 676220 750876
rect 676272 750864 676278 750916
rect 42150 749776 42156 749828
rect 42208 749816 42214 749828
rect 43070 749816 43076 749828
rect 42208 749788 43076 749816
rect 42208 749776 42214 749788
rect 43070 749776 43076 749788
rect 43128 749776 43134 749828
rect 651558 749436 651564 749488
rect 651616 749476 651622 749488
rect 672810 749476 672816 749488
rect 651616 749448 672816 749476
rect 651616 749436 651622 749448
rect 672810 749436 672816 749448
rect 672868 749436 672874 749488
rect 42978 749368 42984 749420
rect 43036 749408 43042 749420
rect 44542 749408 44548 749420
rect 43036 749380 44548 749408
rect 43036 749368 43042 749380
rect 44542 749368 44548 749380
rect 44600 749368 44606 749420
rect 670050 749368 670056 749420
rect 670108 749408 670114 749420
rect 683114 749408 683120 749420
rect 670108 749380 683120 749408
rect 670108 749368 670114 749380
rect 683114 749368 683120 749380
rect 683172 749368 683178 749420
rect 42978 747028 42984 747040
rect 42076 747000 42984 747028
rect 42076 746972 42104 747000
rect 42978 746988 42984 747000
rect 43036 746988 43042 747040
rect 42058 746920 42064 746972
rect 42116 746920 42122 746972
rect 42150 746920 42156 746972
rect 42208 746960 42214 746972
rect 42702 746960 42708 746972
rect 42208 746932 42708 746960
rect 42208 746920 42214 746932
rect 42702 746920 42708 746932
rect 42760 746920 42766 746972
rect 42702 746784 42708 746836
rect 42760 746824 42766 746836
rect 42886 746824 42892 746836
rect 42760 746796 42892 746824
rect 42760 746784 42766 746796
rect 42886 746784 42892 746796
rect 42944 746784 42950 746836
rect 42610 746648 42616 746700
rect 42668 746688 42674 746700
rect 43070 746688 43076 746700
rect 42668 746660 43076 746688
rect 42668 746648 42674 746660
rect 43070 746648 43076 746660
rect 43128 746648 43134 746700
rect 42150 746036 42156 746088
rect 42208 746076 42214 746088
rect 42702 746076 42708 746088
rect 42208 746048 42708 746076
rect 42208 746036 42214 746048
rect 42702 746036 42708 746048
rect 42760 746036 42766 746088
rect 42702 745900 42708 745952
rect 42760 745940 42766 745952
rect 44358 745940 44364 745952
rect 42760 745912 44364 745940
rect 42760 745900 42766 745912
rect 44358 745900 44364 745912
rect 44416 745900 44422 745952
rect 42150 745424 42156 745476
rect 42208 745464 42214 745476
rect 43070 745464 43076 745476
rect 42208 745436 43076 745464
rect 42208 745424 42214 745436
rect 43070 745424 43076 745436
rect 43128 745424 43134 745476
rect 42150 743724 42156 743776
rect 42208 743764 42214 743776
rect 42702 743764 42708 743776
rect 42208 743736 42708 743764
rect 42208 743724 42214 743736
rect 42702 743724 42708 743736
rect 42760 743724 42766 743776
rect 42150 743248 42156 743300
rect 42208 743288 42214 743300
rect 42610 743288 42616 743300
rect 42208 743260 42616 743288
rect 42208 743248 42214 743260
rect 42610 743248 42616 743260
rect 42668 743248 42674 743300
rect 671982 743180 671988 743232
rect 672040 743220 672046 743232
rect 675386 743220 675392 743232
rect 672040 743192 675392 743220
rect 672040 743180 672046 743192
rect 675386 743180 675392 743192
rect 675444 743180 675450 743232
rect 672350 742500 672356 742552
rect 672408 742540 672414 742552
rect 675386 742540 675392 742552
rect 672408 742512 675392 742540
rect 672408 742500 672414 742512
rect 675386 742500 675392 742512
rect 675444 742500 675450 742552
rect 50430 741072 50436 741124
rect 50488 741112 50494 741124
rect 62114 741112 62120 741124
rect 50488 741084 62120 741112
rect 50488 741072 50494 741084
rect 62114 741072 62120 741084
rect 62172 741072 62178 741124
rect 673178 739100 673184 739152
rect 673236 739140 673242 739152
rect 675386 739140 675392 739152
rect 673236 739112 675392 739140
rect 673236 739100 673242 739112
rect 675386 739100 675392 739112
rect 675444 739100 675450 739152
rect 673730 738216 673736 738268
rect 673788 738256 673794 738268
rect 675386 738256 675392 738268
rect 673788 738228 675392 738256
rect 673788 738216 673794 738228
rect 675386 738216 675392 738228
rect 675444 738216 675450 738268
rect 674282 735632 674288 735684
rect 674340 735672 674346 735684
rect 675386 735672 675392 735684
rect 674340 735644 675392 735672
rect 674340 735632 674346 735644
rect 675386 735632 675392 735644
rect 675444 735632 675450 735684
rect 651558 735564 651564 735616
rect 651616 735604 651622 735616
rect 660298 735604 660304 735616
rect 651616 735576 660304 735604
rect 651616 735564 651622 735576
rect 660298 735564 660304 735576
rect 660356 735564 660362 735616
rect 673086 734952 673092 735004
rect 673144 734992 673150 735004
rect 675386 734992 675392 735004
rect 673144 734964 675392 734992
rect 673144 734952 673150 734964
rect 675386 734952 675392 734964
rect 675444 734952 675450 735004
rect 658918 734816 658924 734868
rect 658976 734856 658982 734868
rect 658976 734828 663794 734856
rect 658976 734816 658982 734828
rect 663766 734380 663794 734828
rect 674558 734380 674564 734392
rect 663766 734352 674564 734380
rect 674558 734340 674564 734352
rect 674616 734340 674622 734392
rect 674466 733592 674472 733644
rect 674524 733632 674530 733644
rect 675386 733632 675392 733644
rect 674524 733604 675392 733632
rect 674524 733592 674530 733604
rect 675386 733592 675392 733604
rect 675444 733592 675450 733644
rect 674558 732028 674564 732080
rect 674616 732068 674622 732080
rect 675386 732068 675392 732080
rect 674616 732040 675392 732068
rect 674616 732028 674622 732040
rect 675386 732028 675392 732040
rect 675444 732028 675450 732080
rect 31386 731348 31392 731400
rect 31444 731388 31450 731400
rect 44726 731388 44732 731400
rect 31444 731360 44732 731388
rect 31444 731348 31450 731360
rect 44726 731348 44732 731360
rect 44784 731348 44790 731400
rect 31570 731280 31576 731332
rect 31628 731320 31634 731332
rect 31628 731292 35894 731320
rect 31628 731280 31634 731292
rect 35866 731252 35894 731292
rect 49050 731252 49056 731264
rect 35866 731224 49056 731252
rect 49050 731212 49056 731224
rect 49108 731212 49114 731264
rect 31662 731144 31668 731196
rect 31720 731184 31726 731196
rect 31720 731156 35894 731184
rect 31720 731144 31726 731156
rect 35866 731116 35894 731156
rect 51718 731116 51724 731128
rect 35866 731088 51724 731116
rect 51718 731076 51724 731088
rect 51776 731076 51782 731128
rect 31478 731008 31484 731060
rect 31536 731048 31542 731060
rect 31536 731020 35894 731048
rect 31536 731008 31542 731020
rect 35866 730980 35894 731020
rect 54478 730980 54484 730992
rect 35866 730952 54484 730980
rect 54478 730940 54484 730952
rect 54536 730940 54542 730992
rect 674466 730464 674472 730516
rect 674524 730504 674530 730516
rect 675386 730504 675392 730516
rect 674524 730476 675392 730504
rect 674524 730464 674530 730476
rect 675386 730464 675392 730476
rect 675444 730464 675450 730516
rect 673822 728628 673828 728680
rect 673880 728668 673886 728680
rect 675478 728668 675484 728680
rect 673880 728640 675484 728668
rect 673880 728628 673886 728640
rect 675478 728628 675484 728640
rect 675536 728628 675542 728680
rect 47670 727268 47676 727320
rect 47728 727308 47734 727320
rect 62114 727308 62120 727320
rect 47728 727280 62120 727308
rect 47728 727268 47734 727280
rect 62114 727268 62120 727280
rect 62172 727268 62178 727320
rect 652018 723120 652024 723172
rect 652076 723160 652082 723172
rect 658918 723160 658924 723172
rect 652076 723132 658924 723160
rect 652076 723120 652082 723132
rect 658918 723120 658924 723132
rect 658976 723120 658982 723172
rect 41506 719652 41512 719704
rect 41564 719692 41570 719704
rect 50338 719692 50344 719704
rect 41564 719664 50344 719692
rect 41564 719652 41570 719664
rect 50338 719652 50344 719664
rect 50396 719652 50402 719704
rect 42150 716864 42156 716916
rect 42208 716904 42214 716916
rect 42518 716904 42524 716916
rect 42208 716876 42524 716904
rect 42208 716864 42214 716876
rect 42518 716864 42524 716876
rect 42576 716864 42582 716916
rect 664438 716252 664444 716304
rect 664496 716292 664502 716304
rect 676030 716292 676036 716304
rect 664496 716264 676036 716292
rect 664496 716252 664502 716264
rect 676030 716252 676036 716264
rect 676088 716252 676094 716304
rect 40862 716184 40868 716236
rect 40920 716224 40926 716236
rect 41874 716224 41880 716236
rect 40920 716196 41880 716224
rect 40920 716184 40926 716196
rect 41874 716184 41880 716196
rect 41932 716184 41938 716236
rect 671430 716116 671436 716168
rect 671488 716156 671494 716168
rect 676030 716156 676036 716168
rect 671488 716128 676036 716156
rect 671488 716116 671494 716128
rect 676030 716116 676036 716128
rect 676088 716116 676094 716168
rect 34422 715504 34428 715556
rect 34480 715544 34486 715556
rect 42150 715544 42156 715556
rect 34480 715516 42156 715544
rect 34480 715504 34486 715516
rect 42150 715504 42156 715516
rect 42208 715504 42214 715556
rect 673362 715300 673368 715352
rect 673420 715340 673426 715352
rect 675938 715340 675944 715352
rect 673420 715312 675944 715340
rect 673420 715300 673426 715312
rect 675938 715300 675944 715312
rect 675996 715300 676002 715352
rect 663058 714960 663064 715012
rect 663116 715000 663122 715012
rect 676030 715000 676036 715012
rect 663116 714972 676036 715000
rect 663116 714960 663122 714972
rect 676030 714960 676036 714972
rect 676088 714960 676094 715012
rect 44818 714824 44824 714876
rect 44876 714864 44882 714876
rect 62114 714864 62120 714876
rect 44876 714836 62120 714864
rect 44876 714824 44882 714836
rect 62114 714824 62120 714836
rect 62172 714824 62178 714876
rect 672902 714824 672908 714876
rect 672960 714864 672966 714876
rect 676030 714864 676036 714876
rect 672960 714836 676036 714864
rect 672960 714824 672966 714836
rect 676030 714824 676036 714836
rect 676088 714824 676094 714876
rect 40678 714756 40684 714808
rect 40736 714796 40742 714808
rect 42426 714796 42432 714808
rect 40736 714768 42432 714796
rect 40736 714756 40742 714768
rect 42426 714756 42432 714768
rect 42484 714756 42490 714808
rect 672258 714484 672264 714536
rect 672316 714524 672322 714536
rect 676030 714524 676036 714536
rect 672316 714496 676036 714524
rect 672316 714484 672322 714496
rect 676030 714484 676036 714496
rect 676088 714484 676094 714536
rect 672258 714008 672264 714060
rect 672316 714048 672322 714060
rect 676030 714048 676036 714060
rect 672316 714020 676036 714048
rect 672316 714008 672322 714020
rect 676030 714008 676036 714020
rect 676088 714008 676094 714060
rect 41874 713804 41880 713856
rect 41932 713804 41938 713856
rect 42150 713804 42156 713856
rect 42208 713844 42214 713856
rect 42208 713816 42564 713844
rect 42208 713804 42214 713816
rect 41892 713584 41920 713804
rect 41874 713532 41880 713584
rect 41932 713532 41938 713584
rect 42536 712156 42564 713816
rect 674650 713668 674656 713720
rect 674708 713708 674714 713720
rect 676030 713708 676036 713720
rect 674708 713680 676036 713708
rect 674708 713668 674714 713680
rect 676030 713668 676036 713680
rect 676088 713668 676094 713720
rect 673454 713192 673460 713244
rect 673512 713232 673518 713244
rect 676030 713232 676036 713244
rect 673512 713204 676036 713232
rect 673512 713192 673518 713204
rect 676030 713192 676036 713204
rect 676088 713192 676094 713244
rect 673546 712376 673552 712428
rect 673604 712416 673610 712428
rect 676030 712416 676036 712428
rect 673604 712388 676036 712416
rect 673604 712376 673610 712388
rect 676030 712376 676036 712388
rect 676088 712376 676094 712428
rect 42518 712104 42524 712156
rect 42576 712104 42582 712156
rect 672626 712036 672632 712088
rect 672684 712076 672690 712088
rect 676030 712076 676036 712088
rect 672684 712048 676036 712076
rect 672684 712036 672690 712048
rect 676030 712036 676036 712048
rect 676088 712036 676094 712088
rect 670602 711220 670608 711272
rect 670660 711260 670666 711272
rect 676030 711260 676036 711272
rect 670660 711232 676036 711260
rect 670660 711220 670666 711232
rect 676030 711220 676036 711232
rect 676088 711220 676094 711272
rect 42518 710948 42524 711000
rect 42576 710988 42582 711000
rect 42978 710988 42984 711000
rect 42576 710960 42984 710988
rect 42576 710948 42582 710960
rect 42978 710948 42984 710960
rect 43036 710948 43042 711000
rect 42150 710880 42156 710932
rect 42208 710920 42214 710932
rect 43530 710920 43536 710932
rect 42208 710892 43536 710920
rect 42208 710880 42214 710892
rect 43530 710880 43536 710892
rect 43588 710880 43594 710932
rect 672534 710404 672540 710456
rect 672592 710444 672598 710456
rect 676030 710444 676036 710456
rect 672592 710416 676036 710444
rect 672592 710404 672598 710416
rect 676030 710404 676036 710416
rect 676088 710404 676094 710456
rect 672166 709996 672172 710048
rect 672224 710036 672230 710048
rect 676030 710036 676036 710048
rect 672224 710008 676036 710036
rect 672224 709996 672230 710008
rect 676030 709996 676036 710008
rect 676088 709996 676094 710048
rect 674190 709588 674196 709640
rect 674248 709628 674254 709640
rect 676030 709628 676036 709640
rect 674248 709600 676036 709628
rect 674248 709588 674254 709600
rect 676030 709588 676036 709600
rect 676088 709588 676094 709640
rect 43162 709316 43168 709368
rect 43220 709356 43226 709368
rect 44542 709356 44548 709368
rect 43220 709328 44548 709356
rect 43220 709316 43226 709328
rect 44542 709316 44548 709328
rect 44600 709316 44606 709368
rect 651558 709316 651564 709368
rect 651616 709356 651622 709368
rect 671430 709356 671436 709368
rect 651616 709328 671436 709356
rect 651616 709316 651622 709328
rect 671430 709316 671436 709328
rect 671488 709316 671494 709368
rect 674006 709180 674012 709232
rect 674064 709220 674070 709232
rect 676030 709220 676036 709232
rect 674064 709192 676036 709220
rect 674064 709180 674070 709192
rect 676030 709180 676036 709192
rect 676088 709180 676094 709232
rect 42150 708568 42156 708620
rect 42208 708608 42214 708620
rect 42518 708608 42524 708620
rect 42208 708580 42524 708608
rect 42208 708568 42214 708580
rect 42518 708568 42524 708580
rect 42576 708568 42582 708620
rect 672442 708364 672448 708416
rect 672500 708404 672506 708416
rect 676030 708404 676036 708416
rect 672500 708376 676036 708404
rect 672500 708364 672506 708376
rect 676030 708364 676036 708376
rect 676088 708364 676094 708416
rect 676030 708228 676036 708280
rect 676088 708268 676094 708280
rect 677318 708268 677324 708280
rect 676088 708240 677324 708268
rect 676088 708228 676094 708240
rect 677318 708228 677324 708240
rect 677376 708228 677382 708280
rect 42150 708024 42156 708076
rect 42208 708064 42214 708076
rect 43162 708064 43168 708076
rect 42208 708036 43168 708064
rect 42208 708024 42214 708036
rect 43162 708024 43168 708036
rect 43220 708024 43226 708076
rect 673270 707548 673276 707600
rect 673328 707588 673334 707600
rect 676030 707588 676036 707600
rect 673328 707560 676036 707588
rect 673328 707548 673334 707560
rect 676030 707548 676036 707560
rect 676088 707548 676094 707600
rect 42150 707208 42156 707260
rect 42208 707248 42214 707260
rect 44358 707248 44364 707260
rect 42208 707220 44364 707248
rect 42208 707208 42214 707220
rect 44358 707208 44364 707220
rect 44416 707208 44422 707260
rect 673638 707140 673644 707192
rect 673696 707180 673702 707192
rect 676030 707180 676036 707192
rect 673696 707152 676036 707180
rect 673696 707140 673702 707152
rect 676030 707140 676036 707152
rect 676088 707140 676094 707192
rect 42150 706732 42156 706784
rect 42208 706772 42214 706784
rect 42518 706772 42524 706784
rect 42208 706744 42524 706772
rect 42208 706732 42214 706744
rect 42518 706732 42524 706744
rect 42576 706732 42582 706784
rect 673914 706732 673920 706784
rect 673972 706772 673978 706784
rect 676030 706772 676036 706784
rect 673972 706744 676036 706772
rect 673972 706732 673978 706744
rect 676030 706732 676036 706744
rect 676088 706732 676094 706784
rect 42058 704216 42064 704268
rect 42116 704256 42122 704268
rect 43070 704256 43076 704268
rect 42116 704228 43076 704256
rect 42116 704216 42122 704228
rect 43070 704216 43076 704228
rect 43128 704216 43134 704268
rect 670142 703808 670148 703860
rect 670200 703848 670206 703860
rect 676030 703848 676036 703860
rect 670200 703820 676036 703848
rect 670200 703808 670206 703820
rect 676030 703808 676036 703820
rect 676088 703808 676094 703860
rect 42150 703536 42156 703588
rect 42208 703576 42214 703588
rect 42978 703576 42984 703588
rect 42208 703548 42984 703576
rect 42208 703536 42214 703548
rect 42978 703536 42984 703548
rect 43036 703536 43042 703588
rect 42426 702992 42432 703044
rect 42484 702992 42490 703044
rect 42058 702856 42064 702908
rect 42116 702896 42122 702908
rect 42444 702896 42472 702992
rect 42116 702868 42472 702896
rect 42116 702856 42122 702868
rect 42242 702516 42248 702568
rect 42300 702516 42306 702568
rect 42058 702244 42064 702296
rect 42116 702284 42122 702296
rect 42260 702284 42288 702516
rect 42116 702256 42288 702284
rect 42116 702244 42122 702256
rect 42150 700408 42156 700460
rect 42208 700448 42214 700460
rect 42426 700448 42432 700460
rect 42208 700420 42432 700448
rect 42208 700408 42214 700420
rect 42426 700408 42432 700420
rect 42484 700408 42490 700460
rect 42150 699864 42156 699916
rect 42208 699904 42214 699916
rect 42886 699904 42892 699916
rect 42208 699876 42892 699904
rect 42208 699864 42214 699876
rect 42886 699864 42892 699876
rect 42944 699864 42950 699916
rect 671890 698164 671896 698216
rect 671948 698204 671954 698216
rect 675386 698204 675392 698216
rect 671948 698176 675392 698204
rect 671948 698164 671954 698176
rect 675386 698164 675392 698176
rect 675444 698164 675450 698216
rect 674650 694152 674656 694204
rect 674708 694192 674714 694204
rect 675478 694192 675484 694204
rect 674708 694164 675484 694192
rect 674708 694152 674714 694164
rect 675478 694152 675484 694164
rect 675536 694152 675542 694204
rect 673270 692928 673276 692980
rect 673328 692968 673334 692980
rect 675478 692968 675484 692980
rect 673328 692940 675484 692968
rect 673328 692928 673334 692940
rect 675478 692928 675484 692940
rect 675536 692928 675542 692980
rect 35710 692044 35716 692096
rect 35768 692084 35774 692096
rect 44910 692084 44916 692096
rect 35768 692056 44916 692084
rect 35768 692044 35774 692056
rect 44910 692044 44916 692056
rect 44968 692044 44974 692096
rect 672626 690412 672632 690464
rect 672684 690452 672690 690464
rect 675386 690452 675392 690464
rect 672684 690424 675392 690452
rect 672684 690412 672690 690424
rect 675386 690412 675392 690424
rect 675444 690412 675450 690464
rect 673914 690004 673920 690056
rect 673972 690044 673978 690056
rect 675386 690044 675392 690056
rect 673972 690016 675392 690044
rect 673972 690004 673978 690016
rect 675386 690004 675392 690016
rect 675444 690004 675450 690056
rect 674374 689324 674380 689376
rect 674432 689364 674438 689376
rect 675478 689364 675484 689376
rect 674432 689336 675484 689364
rect 674432 689324 674438 689336
rect 675478 689324 675484 689336
rect 675536 689324 675542 689376
rect 658918 689256 658924 689308
rect 658976 689296 658982 689308
rect 674742 689296 674748 689308
rect 658976 689268 674748 689296
rect 658976 689256 658982 689268
rect 674742 689256 674748 689268
rect 674800 689256 674806 689308
rect 49050 688644 49056 688696
rect 49108 688684 49114 688696
rect 62114 688684 62120 688696
rect 49108 688656 62120 688684
rect 49108 688644 49114 688656
rect 62114 688644 62120 688656
rect 62172 688644 62178 688696
rect 672994 688644 673000 688696
rect 673052 688684 673058 688696
rect 675386 688684 675392 688696
rect 673052 688656 675392 688684
rect 673052 688644 673058 688656
rect 675386 688644 675392 688656
rect 675444 688644 675450 688696
rect 35802 687896 35808 687948
rect 35860 687936 35866 687948
rect 47670 687936 47676 687948
rect 35860 687908 47676 687936
rect 35860 687896 35866 687908
rect 47670 687896 47676 687908
rect 47728 687896 47734 687948
rect 35618 687760 35624 687812
rect 35676 687800 35682 687812
rect 50430 687800 50436 687812
rect 35676 687772 50436 687800
rect 35676 687760 35682 687772
rect 50430 687760 50436 687772
rect 50488 687760 50494 687812
rect 673362 687284 673368 687336
rect 673420 687324 673426 687336
rect 675386 687324 675392 687336
rect 673420 687296 675392 687324
rect 673420 687284 673426 687296
rect 675386 687284 675392 687296
rect 675444 687284 675450 687336
rect 674742 687012 674748 687064
rect 674800 687052 674806 687064
rect 675478 687052 675484 687064
rect 674800 687024 675484 687052
rect 674800 687012 674806 687024
rect 675478 687012 675484 687024
rect 675536 687012 675542 687064
rect 670602 686060 670608 686112
rect 670660 686100 670666 686112
rect 675386 686100 675392 686112
rect 670660 686072 675392 686100
rect 670660 686060 670666 686072
rect 675386 686060 675392 686072
rect 675444 686060 675450 686112
rect 672534 684224 672540 684276
rect 672592 684264 672598 684276
rect 675386 684264 675392 684276
rect 672592 684236 675392 684264
rect 672592 684224 672598 684236
rect 675386 684224 675392 684236
rect 675444 684224 675450 684276
rect 651834 683136 651840 683188
rect 651892 683176 651898 683188
rect 658918 683176 658924 683188
rect 651892 683148 658924 683176
rect 651892 683136 651898 683148
rect 658918 683136 658924 683148
rect 658976 683136 658982 683188
rect 40678 683000 40684 683052
rect 40736 683040 40742 683052
rect 41690 683040 41696 683052
rect 40736 683012 41696 683040
rect 40736 683000 40742 683012
rect 41690 683000 41696 683012
rect 41748 683000 41754 683052
rect 40770 681776 40776 681828
rect 40828 681816 40834 681828
rect 41690 681816 41696 681828
rect 40828 681788 41696 681816
rect 40828 681776 40834 681788
rect 41690 681776 41696 681788
rect 41748 681776 41754 681828
rect 30466 676812 30472 676864
rect 30524 676852 30530 676864
rect 51718 676852 51724 676864
rect 30524 676824 51724 676852
rect 30524 676812 30530 676824
rect 51718 676812 51724 676824
rect 51776 676812 51782 676864
rect 47670 674840 47676 674892
rect 47728 674880 47734 674892
rect 62114 674880 62120 674892
rect 47728 674852 62120 674880
rect 47728 674840 47734 674852
rect 62114 674840 62120 674852
rect 62172 674840 62178 674892
rect 35158 672800 35164 672852
rect 35216 672840 35222 672852
rect 42426 672840 42432 672852
rect 35216 672812 42432 672840
rect 35216 672800 35222 672812
rect 42426 672800 42432 672812
rect 42484 672800 42490 672852
rect 31018 672732 31024 672784
rect 31076 672772 31082 672784
rect 41874 672772 41880 672784
rect 31076 672744 41880 672772
rect 31076 672732 31082 672744
rect 41874 672732 41880 672744
rect 41932 672732 41938 672784
rect 40770 670964 40776 671016
rect 40828 671004 40834 671016
rect 42058 671004 42064 671016
rect 40828 670976 42064 671004
rect 40828 670964 40834 670976
rect 42058 670964 42064 670976
rect 42116 670964 42122 671016
rect 40678 670896 40684 670948
rect 40736 670936 40742 670948
rect 42702 670936 42708 670948
rect 40736 670908 42708 670936
rect 40736 670896 40742 670908
rect 42702 670896 42708 670908
rect 42760 670896 42766 670948
rect 672718 670896 672724 670948
rect 672776 670936 672782 670948
rect 676214 670936 676220 670948
rect 672776 670908 676220 670936
rect 672776 670896 672782 670908
rect 676214 670896 676220 670908
rect 676272 670896 676278 670948
rect 665818 670760 665824 670812
rect 665876 670800 665882 670812
rect 676030 670800 676036 670812
rect 665876 670772 676036 670800
rect 665876 670760 665882 670772
rect 676030 670760 676036 670772
rect 676088 670760 676094 670812
rect 41874 670556 41880 670608
rect 41932 670556 41938 670608
rect 41966 670556 41972 670608
rect 42024 670596 42030 670608
rect 42978 670596 42984 670608
rect 42024 670568 42984 670596
rect 42024 670556 42030 670568
rect 42978 670556 42984 670568
rect 43036 670556 43042 670608
rect 41892 670404 41920 670556
rect 41874 670352 41880 670404
rect 41932 670352 41938 670404
rect 672258 669672 672264 669724
rect 672316 669712 672322 669724
rect 676214 669712 676220 669724
rect 672316 669684 676220 669712
rect 672316 669672 672322 669684
rect 676214 669672 676220 669684
rect 676272 669672 676278 669724
rect 672902 669536 672908 669588
rect 672960 669576 672966 669588
rect 676122 669576 676128 669588
rect 672960 669548 676128 669576
rect 672960 669536 672966 669548
rect 676122 669536 676128 669548
rect 676180 669536 676186 669588
rect 661770 669400 661776 669452
rect 661828 669440 661834 669452
rect 676306 669440 676312 669452
rect 661828 669412 676312 669440
rect 661828 669400 661834 669412
rect 676306 669400 676312 669412
rect 676364 669400 676370 669452
rect 42702 669332 42708 669384
rect 42760 669372 42766 669384
rect 46198 669372 46204 669384
rect 42760 669344 46204 669372
rect 42760 669332 42766 669344
rect 46198 669332 46204 669344
rect 46256 669332 46262 669384
rect 651558 669332 651564 669384
rect 651616 669372 651622 669384
rect 659010 669372 659016 669384
rect 651616 669344 659016 669372
rect 651616 669332 651622 669344
rect 659010 669332 659016 669344
rect 659068 669332 659074 669384
rect 674190 668856 674196 668908
rect 674248 668896 674254 668908
rect 676030 668896 676036 668908
rect 674248 668868 676036 668896
rect 674248 668856 674254 668868
rect 676030 668856 676036 668868
rect 676088 668856 676094 668908
rect 42978 668720 42984 668772
rect 43036 668720 43042 668772
rect 42886 668516 42892 668568
rect 42944 668556 42950 668568
rect 42996 668556 43024 668720
rect 673454 668652 673460 668704
rect 673512 668692 673518 668704
rect 676214 668692 676220 668704
rect 673512 668664 676220 668692
rect 673512 668652 673518 668664
rect 676214 668652 676220 668664
rect 676272 668652 676278 668704
rect 42944 668528 43024 668556
rect 42944 668516 42950 668528
rect 44450 667944 44456 667956
rect 42812 667916 44456 667944
rect 42150 667836 42156 667888
rect 42208 667876 42214 667888
rect 42702 667876 42708 667888
rect 42208 667848 42708 667876
rect 42208 667836 42214 667848
rect 42702 667836 42708 667848
rect 42760 667836 42766 667888
rect 42702 667700 42708 667752
rect 42760 667740 42766 667752
rect 42812 667740 42840 667916
rect 44450 667904 44456 667916
rect 44508 667904 44514 667956
rect 672718 667904 672724 667956
rect 672776 667944 672782 667956
rect 676030 667944 676036 667956
rect 672776 667916 676036 667944
rect 672776 667904 672782 667916
rect 676030 667904 676036 667916
rect 676088 667904 676094 667956
rect 673546 667836 673552 667888
rect 673604 667876 673610 667888
rect 676214 667876 676220 667888
rect 673604 667848 676220 667876
rect 673604 667836 673610 667848
rect 676214 667836 676220 667848
rect 676272 667836 676278 667888
rect 42760 667712 42840 667740
rect 42760 667700 42766 667712
rect 42150 666680 42156 666732
rect 42208 666720 42214 666732
rect 42702 666720 42708 666732
rect 42208 666692 42708 666720
rect 42208 666680 42214 666692
rect 42702 666680 42708 666692
rect 42760 666680 42766 666732
rect 672258 666544 672264 666596
rect 672316 666584 672322 666596
rect 676214 666584 676220 666596
rect 672316 666556 676220 666584
rect 672316 666544 672322 666556
rect 676214 666544 676220 666556
rect 676272 666544 676278 666596
rect 42702 666476 42708 666528
rect 42760 666516 42766 666528
rect 43070 666516 43076 666528
rect 42760 666488 43076 666516
rect 42760 666476 42766 666488
rect 43070 666476 43076 666488
rect 43128 666476 43134 666528
rect 674466 666476 674472 666528
rect 674524 666516 674530 666528
rect 676030 666516 676036 666528
rect 674524 666488 676036 666516
rect 674524 666476 674530 666488
rect 676030 666476 676036 666488
rect 676088 666476 676094 666528
rect 671982 665320 671988 665372
rect 672040 665360 672046 665372
rect 676214 665360 676220 665372
rect 672040 665332 676220 665360
rect 672040 665320 672046 665332
rect 676214 665320 676220 665332
rect 676272 665320 676278 665372
rect 674282 665252 674288 665304
rect 674340 665292 674346 665304
rect 676030 665292 676036 665304
rect 674340 665264 676036 665292
rect 674340 665252 674346 665264
rect 676030 665252 676036 665264
rect 676088 665252 676094 665304
rect 673822 664980 673828 665032
rect 673880 665020 673886 665032
rect 676214 665020 676220 665032
rect 673880 664992 676220 665020
rect 673880 664980 673886 664992
rect 676214 664980 676220 664992
rect 676272 664980 676278 665032
rect 42150 664164 42156 664216
rect 42208 664204 42214 664216
rect 42702 664204 42708 664216
rect 42208 664176 42708 664204
rect 42208 664164 42214 664176
rect 42702 664164 42708 664176
rect 42760 664164 42766 664216
rect 672350 663960 672356 664012
rect 672408 664000 672414 664012
rect 676214 664000 676220 664012
rect 672408 663972 676220 664000
rect 672408 663960 672414 663972
rect 676214 663960 676220 663972
rect 676272 663960 676278 664012
rect 673178 663756 673184 663808
rect 673236 663796 673242 663808
rect 676214 663796 676220 663808
rect 673236 663768 676220 663796
rect 673236 663756 673242 663768
rect 676214 663756 676220 663768
rect 676272 663756 676278 663808
rect 43530 662396 43536 662448
rect 43588 662436 43594 662448
rect 62114 662436 62120 662448
rect 43588 662408 62120 662436
rect 43588 662396 43594 662408
rect 62114 662396 62120 662408
rect 62172 662396 62178 662448
rect 673730 662328 673736 662380
rect 673788 662368 673794 662380
rect 676030 662368 676036 662380
rect 673788 662340 676036 662368
rect 673788 662328 673794 662340
rect 676030 662328 676036 662340
rect 676088 662328 676094 662380
rect 674558 661580 674564 661632
rect 674616 661620 674622 661632
rect 676030 661620 676036 661632
rect 674616 661592 676036 661620
rect 674616 661580 674622 661592
rect 676030 661580 676036 661592
rect 676088 661580 676094 661632
rect 673086 661104 673092 661156
rect 673144 661144 673150 661156
rect 676214 661144 676220 661156
rect 673144 661116 676220 661144
rect 673144 661104 673150 661116
rect 676214 661104 676220 661116
rect 676272 661104 676278 661156
rect 42150 661036 42156 661088
rect 42208 661076 42214 661088
rect 43070 661076 43076 661088
rect 42208 661048 43076 661076
rect 42208 661036 42214 661048
rect 43070 661036 43076 661048
rect 43128 661036 43134 661088
rect 42150 659676 42156 659728
rect 42208 659716 42214 659728
rect 42886 659716 42892 659728
rect 42208 659688 42892 659716
rect 42208 659676 42214 659688
rect 42886 659676 42892 659688
rect 42944 659676 42950 659728
rect 42150 658996 42156 659048
rect 42208 659036 42214 659048
rect 42702 659036 42708 659048
rect 42208 659008 42708 659036
rect 42208 658996 42214 659008
rect 42702 658996 42708 659008
rect 42760 658996 42766 659048
rect 42886 658248 42892 658300
rect 42944 658288 42950 658300
rect 44358 658288 44364 658300
rect 42944 658260 44364 658288
rect 42944 658248 42950 658260
rect 44358 658248 44364 658260
rect 44416 658248 44422 658300
rect 42150 657228 42156 657280
rect 42208 657268 42214 657280
rect 42518 657268 42524 657280
rect 42208 657240 42524 657268
rect 42208 657228 42214 657240
rect 42518 657228 42524 657240
rect 42576 657228 42582 657280
rect 651558 656888 651564 656940
rect 651616 656928 651622 656940
rect 663058 656928 663064 656940
rect 651616 656900 663064 656928
rect 651616 656888 651622 656900
rect 663058 656888 663064 656900
rect 663116 656888 663122 656940
rect 42150 656820 42156 656872
rect 42208 656860 42214 656872
rect 42886 656860 42892 656872
rect 42208 656832 42892 656860
rect 42208 656820 42214 656832
rect 42886 656820 42892 656832
rect 42944 656820 42950 656872
rect 42150 656140 42156 656192
rect 42208 656180 42214 656192
rect 42334 656180 42340 656192
rect 42208 656152 42340 656180
rect 42208 656140 42214 656152
rect 42334 656140 42340 656152
rect 42392 656140 42398 656192
rect 671982 652740 671988 652792
rect 672040 652780 672046 652792
rect 675386 652780 675392 652792
rect 672040 652752 675392 652780
rect 672040 652740 672046 652752
rect 675386 652740 675392 652752
rect 675444 652740 675450 652792
rect 54478 650020 54484 650072
rect 54536 650060 54542 650072
rect 62114 650060 62120 650072
rect 54536 650032 62120 650060
rect 54536 650020 54542 650032
rect 62114 650020 62120 650032
rect 62172 650020 62178 650072
rect 674558 649816 674564 649868
rect 674616 649856 674622 649868
rect 675386 649856 675392 649868
rect 674616 649828 675392 649856
rect 674616 649816 674622 649828
rect 675386 649816 675392 649828
rect 675444 649816 675450 649868
rect 673178 647708 673184 647760
rect 673236 647748 673242 647760
rect 675478 647748 675484 647760
rect 673236 647720 675484 647748
rect 673236 647708 673242 647720
rect 675478 647708 675484 647720
rect 675536 647708 675542 647760
rect 672902 645532 672908 645584
rect 672960 645572 672966 645584
rect 675386 645572 675392 645584
rect 672960 645544 675392 645572
rect 672960 645532 672966 645544
rect 675386 645532 675392 645544
rect 675444 645532 675450 645584
rect 674282 644784 674288 644836
rect 674340 644824 674346 644836
rect 675386 644824 675392 644836
rect 674340 644796 675392 644824
rect 674340 644784 674346 644796
rect 675386 644784 675392 644796
rect 675444 644784 675450 644836
rect 35802 644580 35808 644632
rect 35860 644620 35866 644632
rect 47670 644620 47676 644632
rect 35860 644592 47676 644620
rect 35860 644580 35866 644592
rect 47670 644580 47676 644592
rect 47728 644580 47734 644632
rect 35618 644512 35624 644564
rect 35676 644552 35682 644564
rect 49050 644552 49056 644564
rect 35676 644524 49056 644552
rect 35676 644512 35682 644524
rect 49050 644512 49056 644524
rect 49108 644512 49114 644564
rect 659010 643696 659016 643748
rect 659068 643736 659074 643748
rect 674466 643736 674472 643748
rect 659068 643708 674472 643736
rect 659068 643696 659074 643708
rect 674466 643696 674472 643708
rect 674524 643696 674530 643748
rect 673086 643356 673092 643408
rect 673144 643396 673150 643408
rect 675386 643396 675392 643408
rect 673144 643368 675392 643396
rect 673144 643356 673150 643368
rect 675386 643356 675392 643368
rect 675444 643356 675450 643408
rect 651558 643084 651564 643136
rect 651616 643124 651622 643136
rect 668670 643124 668676 643136
rect 651616 643096 668676 643124
rect 651616 643084 651622 643096
rect 668670 643084 668676 643096
rect 668728 643084 668734 643136
rect 674466 641860 674472 641912
rect 674524 641900 674530 641912
rect 675386 641900 675392 641912
rect 674524 641872 675392 641900
rect 674524 641860 674530 641872
rect 675386 641860 675392 641872
rect 675444 641860 675450 641912
rect 674006 639072 674012 639124
rect 674064 639112 674070 639124
rect 675386 639112 675392 639124
rect 674064 639084 675392 639112
rect 674064 639072 674070 639084
rect 675386 639072 675392 639084
rect 675444 639072 675450 639124
rect 47670 636216 47676 636268
rect 47728 636256 47734 636268
rect 62114 636256 62120 636268
rect 47728 636228 62120 636256
rect 47728 636216 47734 636228
rect 62114 636216 62120 636228
rect 62172 636216 62178 636268
rect 32398 629892 32404 629944
rect 32456 629932 32462 629944
rect 41782 629932 41788 629944
rect 32456 629904 41788 629932
rect 32456 629892 32462 629904
rect 41782 629892 41788 629904
rect 41840 629892 41846 629944
rect 651558 629280 651564 629332
rect 651616 629320 651622 629332
rect 661770 629320 661776 629332
rect 651616 629292 661776 629320
rect 651616 629280 651622 629292
rect 661770 629280 661776 629292
rect 661828 629280 661834 629332
rect 33778 628532 33784 628584
rect 33836 628572 33842 628584
rect 42518 628572 42524 628584
rect 33836 628544 42524 628572
rect 33836 628532 33842 628544
rect 42518 628532 42524 628544
rect 42576 628532 42582 628584
rect 41782 627376 41788 627428
rect 41840 627376 41846 627428
rect 41800 627088 41828 627376
rect 41782 627036 41788 627088
rect 41840 627036 41846 627088
rect 42978 626560 42984 626612
rect 43036 626600 43042 626612
rect 44818 626600 44824 626612
rect 43036 626572 44824 626600
rect 43036 626560 43042 626572
rect 44818 626560 44824 626572
rect 44876 626560 44882 626612
rect 672810 625472 672816 625524
rect 672868 625512 672874 625524
rect 676122 625512 676128 625524
rect 672868 625484 676128 625512
rect 672868 625472 672874 625484
rect 676122 625472 676128 625484
rect 676180 625472 676186 625524
rect 664530 625336 664536 625388
rect 664588 625376 664594 625388
rect 676214 625376 676220 625388
rect 664588 625348 676220 625376
rect 664588 625336 664594 625348
rect 676214 625336 676220 625348
rect 676272 625336 676278 625388
rect 42150 625268 42156 625320
rect 42208 625308 42214 625320
rect 42518 625308 42524 625320
rect 42208 625280 42524 625308
rect 42208 625268 42214 625280
rect 42518 625268 42524 625280
rect 42576 625268 42582 625320
rect 660298 625132 660304 625184
rect 660356 625172 660362 625184
rect 676214 625172 676220 625184
rect 660356 625144 676220 625172
rect 660356 625132 660362 625144
rect 676214 625132 676220 625144
rect 676272 625132 676278 625184
rect 42150 624656 42156 624708
rect 42208 624696 42214 624708
rect 42978 624696 42984 624708
rect 42208 624668 42984 624696
rect 42208 624656 42214 624668
rect 42978 624656 42984 624668
rect 43036 624656 43042 624708
rect 674190 624316 674196 624368
rect 674248 624356 674254 624368
rect 676030 624356 676036 624368
rect 674248 624328 676036 624356
rect 674248 624316 674254 624328
rect 676030 624316 676036 624328
rect 676088 624316 676094 624368
rect 42518 623840 42524 623892
rect 42576 623840 42582 623892
rect 672350 623840 672356 623892
rect 672408 623880 672414 623892
rect 676030 623880 676036 623892
rect 672408 623852 676036 623880
rect 672408 623840 672414 623852
rect 676030 623840 676036 623852
rect 676088 623840 676094 623892
rect 42150 623432 42156 623484
rect 42208 623472 42214 623484
rect 42536 623472 42564 623840
rect 43622 623772 43628 623824
rect 43680 623812 43686 623824
rect 62114 623812 62120 623824
rect 43680 623784 62120 623812
rect 43680 623772 43686 623784
rect 62114 623772 62120 623784
rect 62172 623772 62178 623824
rect 672442 623772 672448 623824
rect 672500 623812 672506 623824
rect 676214 623812 676220 623824
rect 672500 623784 676220 623812
rect 672500 623772 672506 623784
rect 676214 623772 676220 623784
rect 676272 623772 676278 623824
rect 42208 623444 42564 623472
rect 42208 623432 42214 623444
rect 672258 622684 672264 622736
rect 672316 622724 672322 622736
rect 676030 622724 676036 622736
rect 672316 622696 676036 622724
rect 672316 622684 672322 622696
rect 676030 622684 676036 622696
rect 676088 622684 676094 622736
rect 672718 622548 672724 622600
rect 672776 622588 672782 622600
rect 676122 622588 676128 622600
rect 672776 622560 676128 622588
rect 672776 622548 672782 622560
rect 676122 622548 676128 622560
rect 676180 622548 676186 622600
rect 672258 622412 672264 622464
rect 672316 622452 672322 622464
rect 676214 622452 676220 622464
rect 672316 622424 676220 622452
rect 672316 622412 672322 622424
rect 676214 622412 676220 622424
rect 676272 622412 676278 622464
rect 673638 622208 673644 622260
rect 673696 622248 673702 622260
rect 676030 622248 676036 622260
rect 673696 622220 676036 622248
rect 673696 622208 673702 622220
rect 676030 622208 676036 622220
rect 676088 622208 676094 622260
rect 42058 622140 42064 622192
rect 42116 622180 42122 622192
rect 42518 622180 42524 622192
rect 42116 622152 42524 622180
rect 42116 622140 42122 622152
rect 42518 622140 42524 622152
rect 42576 622140 42582 622192
rect 42518 622004 42524 622056
rect 42576 622044 42582 622056
rect 42794 622044 42800 622056
rect 42576 622016 42800 622044
rect 42576 622004 42582 622016
rect 42794 622004 42800 622016
rect 42852 622004 42858 622056
rect 671890 621256 671896 621308
rect 671948 621296 671954 621308
rect 676214 621296 676220 621308
rect 671948 621268 676220 621296
rect 671948 621256 671954 621268
rect 676214 621256 676220 621268
rect 676272 621256 676278 621308
rect 670602 621120 670608 621172
rect 670660 621160 670666 621172
rect 676030 621160 676036 621172
rect 670660 621132 676036 621160
rect 670660 621120 670666 621132
rect 676030 621120 676036 621132
rect 676088 621120 676094 621172
rect 42058 620780 42064 620832
rect 42116 620820 42122 620832
rect 43070 620820 43076 620832
rect 42116 620792 43076 620820
rect 42116 620780 42122 620792
rect 43070 620780 43076 620792
rect 43128 620780 43134 620832
rect 42058 620304 42064 620356
rect 42116 620344 42122 620356
rect 42518 620344 42524 620356
rect 42116 620316 42524 620344
rect 42116 620304 42122 620316
rect 42518 620304 42524 620316
rect 42576 620304 42582 620356
rect 42518 620168 42524 620220
rect 42576 620208 42582 620220
rect 42886 620208 42892 620220
rect 42576 620180 42892 620208
rect 42576 620168 42582 620180
rect 42886 620168 42892 620180
rect 42944 620168 42950 620220
rect 672626 619896 672632 619948
rect 672684 619936 672690 619948
rect 676214 619936 676220 619948
rect 672684 619908 676220 619936
rect 672684 619896 672690 619908
rect 676214 619896 676220 619908
rect 676272 619896 676278 619948
rect 672534 619760 672540 619812
rect 672592 619800 672598 619812
rect 676030 619800 676036 619812
rect 672592 619772 676036 619800
rect 672592 619760 672598 619772
rect 676030 619760 676036 619772
rect 676088 619760 676094 619812
rect 674650 619148 674656 619200
rect 674708 619188 674714 619200
rect 676214 619188 676220 619200
rect 674708 619160 676220 619188
rect 674708 619148 674714 619160
rect 676214 619148 676220 619160
rect 676272 619148 676278 619200
rect 44450 618304 44456 618316
rect 42628 618276 44456 618304
rect 42150 617856 42156 617908
rect 42208 617896 42214 617908
rect 42518 617896 42524 617908
rect 42208 617868 42524 617896
rect 42208 617856 42214 617868
rect 42518 617856 42524 617868
rect 42576 617856 42582 617908
rect 42518 617720 42524 617772
rect 42576 617760 42582 617772
rect 42628 617760 42656 618276
rect 44450 618264 44456 618276
rect 44508 618264 44514 618316
rect 674374 617788 674380 617840
rect 674432 617828 674438 617840
rect 676030 617828 676036 617840
rect 674432 617800 676036 617828
rect 674432 617788 674438 617800
rect 676030 617788 676036 617800
rect 676088 617788 676094 617840
rect 42576 617732 42656 617760
rect 42576 617720 42582 617732
rect 42058 617108 42064 617160
rect 42116 617148 42122 617160
rect 42518 617148 42524 617160
rect 42116 617120 42524 617148
rect 42116 617108 42122 617120
rect 42518 617108 42524 617120
rect 42576 617108 42582 617160
rect 673362 617040 673368 617092
rect 673420 617080 673426 617092
rect 676122 617080 676128 617092
rect 673420 617052 676128 617080
rect 673420 617040 673426 617052
rect 676122 617040 676128 617052
rect 676180 617040 676186 617092
rect 673914 616972 673920 617024
rect 673972 617012 673978 617024
rect 676030 617012 676036 617024
rect 673972 616984 676036 617012
rect 673972 616972 673978 616984
rect 676030 616972 676036 616984
rect 676088 616972 676094 617024
rect 652386 616836 652392 616888
rect 652444 616876 652450 616888
rect 659010 616876 659016 616888
rect 652444 616848 659016 616876
rect 652444 616836 652450 616848
rect 659010 616836 659016 616848
rect 659068 616836 659074 616888
rect 673270 616836 673276 616888
rect 673328 616876 673334 616888
rect 676214 616876 676220 616888
rect 673328 616848 676220 616876
rect 673328 616836 673334 616848
rect 676214 616836 676220 616848
rect 676272 616836 676278 616888
rect 672994 615476 673000 615528
rect 673052 615516 673058 615528
rect 676214 615516 676220 615528
rect 673052 615488 676220 615516
rect 673052 615476 673058 615488
rect 676214 615476 676220 615488
rect 676272 615476 676278 615528
rect 672718 614116 672724 614168
rect 672776 614156 672782 614168
rect 683114 614156 683120 614168
rect 672776 614128 683120 614156
rect 672776 614116 672782 614128
rect 683114 614116 683120 614128
rect 683172 614116 683178 614168
rect 42150 613436 42156 613488
rect 42208 613476 42214 613488
rect 42518 613476 42524 613488
rect 42208 613448 42524 613476
rect 42208 613436 42214 613448
rect 42518 613436 42524 613448
rect 42576 613436 42582 613488
rect 675202 610648 675208 610700
rect 675260 610688 675266 610700
rect 675662 610688 675668 610700
rect 675260 610660 675668 610688
rect 675260 610648 675266 610660
rect 675662 610648 675668 610660
rect 675720 610648 675726 610700
rect 44818 609968 44824 610020
rect 44876 610008 44882 610020
rect 62114 610008 62120 610020
rect 44876 609980 62120 610008
rect 44876 609968 44882 609980
rect 62114 609968 62120 609980
rect 62172 609968 62178 610020
rect 673362 607588 673368 607640
rect 673420 607628 673426 607640
rect 675386 607628 675392 607640
rect 673420 607600 675392 607628
rect 673420 607588 673426 607600
rect 675386 607588 675392 607600
rect 675444 607588 675450 607640
rect 674466 604732 674472 604784
rect 674524 604772 674530 604784
rect 675386 604772 675392 604784
rect 674524 604744 675392 604772
rect 674524 604732 674530 604744
rect 675386 604732 675392 604744
rect 675444 604732 675450 604784
rect 674650 604324 674656 604376
rect 674708 604364 674714 604376
rect 675386 604364 675392 604376
rect 674708 604336 675392 604364
rect 674708 604324 674714 604336
rect 675386 604324 675392 604336
rect 675444 604324 675450 604376
rect 673822 603440 673828 603492
rect 673880 603480 673886 603492
rect 675478 603480 675484 603492
rect 673880 603452 675484 603480
rect 673880 603440 673886 603452
rect 675478 603440 675484 603452
rect 675536 603440 675542 603492
rect 651558 603100 651564 603152
rect 651616 603140 651622 603152
rect 660298 603140 660304 603152
rect 651616 603112 660304 603140
rect 651616 603100 651622 603112
rect 660298 603100 660304 603112
rect 660356 603100 660362 603152
rect 673270 603032 673276 603084
rect 673328 603072 673334 603084
rect 675386 603072 675392 603084
rect 673328 603044 675392 603072
rect 673328 603032 673334 603044
rect 675386 603032 675392 603044
rect 675444 603032 675450 603084
rect 35802 601672 35808 601724
rect 35860 601712 35866 601724
rect 47670 601712 47676 601724
rect 35860 601684 47676 601712
rect 35860 601672 35866 601684
rect 47670 601672 47676 601684
rect 47728 601672 47734 601724
rect 43622 601644 43628 601656
rect 35866 601616 43628 601644
rect 35866 601588 35894 601616
rect 43622 601604 43628 601616
rect 43680 601604 43686 601656
rect 35802 601536 35808 601588
rect 35860 601548 35894 601588
rect 35860 601536 35866 601548
rect 35710 601468 35716 601520
rect 35768 601508 35774 601520
rect 44358 601508 44364 601520
rect 35768 601480 44364 601508
rect 35768 601468 35774 601480
rect 44358 601468 44364 601480
rect 44416 601468 44422 601520
rect 35802 601332 35808 601384
rect 35860 601372 35866 601384
rect 54478 601372 54484 601384
rect 35860 601344 54484 601372
rect 35860 601332 35866 601344
rect 54478 601332 54484 601344
rect 54536 601332 54542 601384
rect 674374 599768 674380 599820
rect 674432 599808 674438 599820
rect 675478 599808 675484 599820
rect 674432 599780 675484 599808
rect 674432 599768 674438 599780
rect 675478 599768 675484 599780
rect 675536 599768 675542 599820
rect 659010 599564 659016 599616
rect 659068 599604 659074 599616
rect 659068 599576 663794 599604
rect 659068 599564 659074 599576
rect 663766 599196 663794 599576
rect 674742 599196 674748 599208
rect 663766 599168 674748 599196
rect 674742 599156 674748 599168
rect 674800 599156 674806 599208
rect 674190 598408 674196 598460
rect 674248 598448 674254 598460
rect 675478 598448 675484 598460
rect 674248 598420 675484 598448
rect 674248 598408 674254 598420
rect 675478 598408 675484 598420
rect 675536 598408 675542 598460
rect 46198 597524 46204 597576
rect 46256 597564 46262 597576
rect 62114 597564 62120 597576
rect 46256 597536 62120 597564
rect 46256 597524 46262 597536
rect 62114 597524 62120 597536
rect 62172 597524 62178 597576
rect 674742 596844 674748 596896
rect 674800 596884 674806 596896
rect 675386 596884 675392 596896
rect 674800 596856 675392 596884
rect 674800 596844 674806 596856
rect 675386 596844 675392 596856
rect 675444 596844 675450 596896
rect 672626 595280 672632 595332
rect 672684 595320 672690 595332
rect 675386 595320 675392 595332
rect 672684 595292 675392 595320
rect 672684 595280 672690 595292
rect 675386 595280 675392 595292
rect 675444 595280 675450 595332
rect 672810 593376 672816 593428
rect 672868 593416 672874 593428
rect 675478 593416 675484 593428
rect 672868 593388 675484 593416
rect 672868 593376 672874 593388
rect 675478 593376 675484 593388
rect 675536 593376 675542 593428
rect 651558 590656 651564 590708
rect 651616 590696 651622 590708
rect 664438 590696 664444 590708
rect 651616 590668 664444 590696
rect 651616 590656 651622 590668
rect 664438 590656 664444 590668
rect 664496 590656 664502 590708
rect 41506 589908 41512 589960
rect 41564 589948 41570 589960
rect 54478 589948 54484 589960
rect 41564 589920 54484 589948
rect 41564 589908 41570 589920
rect 54478 589908 54484 589920
rect 54536 589908 54542 589960
rect 33778 585828 33784 585880
rect 33836 585868 33842 585880
rect 41874 585868 41880 585880
rect 33836 585840 41880 585868
rect 33836 585828 33842 585840
rect 41874 585828 41880 585840
rect 41932 585828 41938 585880
rect 32398 585760 32404 585812
rect 32456 585800 32462 585812
rect 41782 585800 41788 585812
rect 32456 585772 41788 585800
rect 32456 585760 32462 585772
rect 41782 585760 41788 585772
rect 41840 585760 41846 585812
rect 40770 584604 40776 584656
rect 40828 584644 40834 584656
rect 42426 584644 42432 584656
rect 40828 584616 42432 584644
rect 40828 584604 40834 584616
rect 42426 584604 42432 584616
rect 42484 584604 42490 584656
rect 40678 584536 40684 584588
rect 40736 584576 40742 584588
rect 41966 584576 41972 584588
rect 40736 584548 41972 584576
rect 40736 584536 40742 584548
rect 41966 584536 41972 584548
rect 42024 584536 42030 584588
rect 41874 584196 41880 584248
rect 41932 584196 41938 584248
rect 42058 584196 42064 584248
rect 42116 584236 42122 584248
rect 42702 584236 42708 584248
rect 42116 584208 42708 584236
rect 42116 584196 42122 584208
rect 42702 584196 42708 584208
rect 42760 584196 42766 584248
rect 41892 583976 41920 584196
rect 41874 583924 41880 583976
rect 41932 583924 41938 583976
rect 47762 583720 47768 583772
rect 47820 583760 47826 583772
rect 62114 583760 62120 583772
rect 47820 583732 62120 583760
rect 47820 583720 47826 583732
rect 62114 583720 62120 583732
rect 62172 583720 62178 583772
rect 42886 581612 42892 581664
rect 42944 581652 42950 581664
rect 43070 581652 43076 581664
rect 42944 581624 43076 581652
rect 42944 581612 42950 581624
rect 43070 581612 43076 581624
rect 43128 581612 43134 581664
rect 42150 581272 42156 581324
rect 42208 581312 42214 581324
rect 43530 581312 43536 581324
rect 42208 581284 43536 581312
rect 42208 581272 42214 581284
rect 43530 581272 43536 581284
rect 43588 581272 43594 581324
rect 652018 581000 652024 581052
rect 652076 581040 652082 581052
rect 676030 581040 676036 581052
rect 652076 581012 676036 581040
rect 652076 581000 652082 581012
rect 676030 581000 676036 581012
rect 676088 581000 676094 581052
rect 672442 580048 672448 580100
rect 672500 580088 672506 580100
rect 676214 580088 676220 580100
rect 672500 580060 676220 580088
rect 672500 580048 672506 580060
rect 676214 580048 676220 580060
rect 676272 580048 676278 580100
rect 671430 579912 671436 579964
rect 671488 579952 671494 579964
rect 676122 579952 676128 579964
rect 671488 579924 676128 579952
rect 671488 579912 671494 579924
rect 676122 579912 676128 579924
rect 676180 579912 676186 579964
rect 658918 579776 658924 579828
rect 658976 579816 658982 579828
rect 676030 579816 676036 579828
rect 658976 579788 676036 579816
rect 658976 579776 658982 579788
rect 676030 579776 676036 579788
rect 676088 579776 676094 579828
rect 42886 579640 42892 579692
rect 42944 579680 42950 579692
rect 44450 579680 44456 579692
rect 42944 579652 44456 579680
rect 42944 579640 42950 579652
rect 44450 579640 44456 579652
rect 44508 579640 44514 579692
rect 673730 579232 673736 579284
rect 673788 579272 673794 579284
rect 676214 579272 676220 579284
rect 673788 579244 676220 579272
rect 673788 579232 673794 579244
rect 676214 579232 676220 579244
rect 676272 579232 676278 579284
rect 673914 578552 673920 578604
rect 673972 578592 673978 578604
rect 676030 578592 676036 578604
rect 673972 578564 676036 578592
rect 673972 578552 673978 578564
rect 676030 578552 676036 578564
rect 676088 578552 676094 578604
rect 42150 578416 42156 578468
rect 42208 578456 42214 578468
rect 42886 578456 42892 578468
rect 42208 578428 42892 578456
rect 42208 578416 42214 578428
rect 42886 578416 42892 578428
rect 42944 578416 42950 578468
rect 43162 578212 43168 578264
rect 43220 578252 43226 578264
rect 44358 578252 44364 578264
rect 43220 578224 44364 578252
rect 43220 578212 43226 578224
rect 44358 578212 44364 578224
rect 44416 578212 44422 578264
rect 672350 578212 672356 578264
rect 672408 578252 672414 578264
rect 676214 578252 676220 578264
rect 672408 578224 676220 578252
rect 672408 578212 672414 578224
rect 676214 578212 676220 578224
rect 676272 578212 676278 578264
rect 673638 577396 673644 577448
rect 673696 577436 673702 577448
rect 676030 577436 676036 577448
rect 673696 577408 676036 577436
rect 673696 577396 673702 577408
rect 676030 577396 676036 577408
rect 676088 577396 676094 577448
rect 672258 576988 672264 577040
rect 672316 577028 672322 577040
rect 676214 577028 676220 577040
rect 672316 577000 676220 577028
rect 672316 576988 672322 577000
rect 676214 576988 676220 577000
rect 676272 576988 676278 577040
rect 42150 576920 42156 576972
rect 42208 576960 42214 576972
rect 43162 576960 43168 576972
rect 42208 576932 43168 576960
rect 42208 576920 42214 576932
rect 43162 576920 43168 576932
rect 43220 576920 43226 576972
rect 672534 576920 672540 576972
rect 672592 576960 672598 576972
rect 676030 576960 676036 576972
rect 672592 576932 676036 576960
rect 672592 576920 672598 576932
rect 676030 576920 676036 576932
rect 676088 576920 676094 576972
rect 651558 576852 651564 576904
rect 651616 576892 651622 576904
rect 659010 576892 659016 576904
rect 651616 576864 659016 576892
rect 651616 576852 651622 576864
rect 659010 576852 659016 576864
rect 659068 576852 659074 576904
rect 672442 576852 672448 576904
rect 672500 576892 672506 576904
rect 676122 576892 676128 576904
rect 672500 576864 676128 576892
rect 672500 576852 672506 576864
rect 676122 576852 676128 576864
rect 676180 576852 676186 576904
rect 42426 576308 42432 576360
rect 42484 576348 42490 576360
rect 42978 576348 42984 576360
rect 42484 576320 42984 576348
rect 42484 576308 42490 576320
rect 42978 576308 42984 576320
rect 43036 576308 43042 576360
rect 671982 575560 671988 575612
rect 672040 575600 672046 575612
rect 676214 575600 676220 575612
rect 672040 575572 676220 575600
rect 672040 575560 672046 575572
rect 676214 575560 676220 575572
rect 676272 575560 676278 575612
rect 674558 575356 674564 575408
rect 674616 575396 674622 575408
rect 676030 575396 676036 575408
rect 674616 575368 676036 575396
rect 674616 575356 674622 575368
rect 676030 575356 676036 575368
rect 676088 575356 676094 575408
rect 42150 574540 42156 574592
rect 42208 574580 42214 574592
rect 42426 574580 42432 574592
rect 42208 574552 42432 574580
rect 42208 574540 42214 574552
rect 42426 574540 42432 574552
rect 42484 574540 42490 574592
rect 674006 574540 674012 574592
rect 674064 574580 674070 574592
rect 676030 574580 676036 574592
rect 674064 574552 676036 574580
rect 674064 574540 674070 574552
rect 676030 574540 676036 574552
rect 676088 574540 676094 574592
rect 672902 574200 672908 574252
rect 672960 574240 672966 574252
rect 676214 574240 676220 574252
rect 672960 574212 676220 574240
rect 672960 574200 672966 574212
rect 676214 574200 676220 574212
rect 676272 574200 676278 574252
rect 42150 574064 42156 574116
rect 42208 574104 42214 574116
rect 42334 574104 42340 574116
rect 42208 574076 42340 574104
rect 42208 574064 42214 574076
rect 42334 574064 42340 574076
rect 42392 574064 42398 574116
rect 42150 573452 42156 573504
rect 42208 573492 42214 573504
rect 43070 573492 43076 573504
rect 42208 573464 43076 573492
rect 42208 573452 42214 573464
rect 43070 573452 43076 573464
rect 43128 573452 43134 573504
rect 674282 571684 674288 571736
rect 674340 571724 674346 571736
rect 676030 571724 676036 571736
rect 674340 571696 676036 571724
rect 674340 571684 674346 571696
rect 676030 571684 676036 571696
rect 676088 571684 676094 571736
rect 42334 571480 42340 571532
rect 42392 571480 42398 571532
rect 673178 571480 673184 571532
rect 673236 571520 673242 571532
rect 676214 571520 676220 571532
rect 673236 571492 676220 571520
rect 673236 571480 673242 571492
rect 676214 571480 676220 571492
rect 676272 571480 676278 571532
rect 42058 570868 42064 570920
rect 42116 570908 42122 570920
rect 42352 570908 42380 571480
rect 43530 571344 43536 571396
rect 43588 571384 43594 571396
rect 62114 571384 62120 571396
rect 43588 571356 62120 571384
rect 43588 571344 43594 571356
rect 62114 571344 62120 571356
rect 62172 571344 62178 571396
rect 42116 570880 42380 570908
rect 42116 570868 42122 570880
rect 673086 569916 673092 569968
rect 673144 569956 673150 569968
rect 676214 569956 676220 569968
rect 673144 569928 676220 569956
rect 673144 569916 673150 569928
rect 676214 569916 676220 569928
rect 676272 569916 676278 569968
rect 42058 569576 42064 569628
rect 42116 569616 42122 569628
rect 42702 569616 42708 569628
rect 42116 569588 42708 569616
rect 42116 569576 42122 569588
rect 42702 569576 42708 569588
rect 42760 569576 42766 569628
rect 668578 568556 668584 568608
rect 668636 568596 668642 568608
rect 683114 568596 683120 568608
rect 668636 568568 683120 568596
rect 668636 568556 668642 568568
rect 683114 568556 683120 568568
rect 683172 568556 683178 568608
rect 652110 563048 652116 563100
rect 652168 563088 652174 563100
rect 658918 563088 658924 563100
rect 652168 563060 658924 563088
rect 652168 563048 652174 563060
rect 658918 563048 658924 563060
rect 658976 563048 658982 563100
rect 35618 562300 35624 562352
rect 35676 562340 35682 562352
rect 43530 562340 43536 562352
rect 35676 562312 43536 562340
rect 35676 562300 35682 562312
rect 43530 562300 43536 562312
rect 43588 562300 43594 562352
rect 671982 561892 671988 561944
rect 672040 561932 672046 561944
rect 675386 561932 675392 561944
rect 672040 561904 675392 561932
rect 672040 561892 672046 561904
rect 675386 561892 675392 561904
rect 675444 561892 675450 561944
rect 673086 560192 673092 560244
rect 673144 560232 673150 560244
rect 675202 560232 675208 560244
rect 673144 560204 675208 560232
rect 673144 560192 673150 560204
rect 675202 560192 675208 560204
rect 675260 560192 675266 560244
rect 675202 559648 675208 559700
rect 675260 559688 675266 559700
rect 675386 559688 675392 559700
rect 675260 559660 675392 559688
rect 675260 559648 675266 559660
rect 675386 559648 675392 559660
rect 675444 559648 675450 559700
rect 35710 558288 35716 558340
rect 35768 558328 35774 558340
rect 46198 558328 46204 558340
rect 35768 558300 46204 558328
rect 35768 558288 35774 558300
rect 46198 558288 46204 558300
rect 46256 558288 46262 558340
rect 35802 558152 35808 558204
rect 35860 558192 35866 558204
rect 47762 558192 47768 558204
rect 35860 558164 47768 558192
rect 35860 558152 35866 558164
rect 47762 558152 47768 558164
rect 47820 558152 47826 558204
rect 47670 557540 47676 557592
rect 47728 557580 47734 557592
rect 62114 557580 62120 557592
rect 47728 557552 62120 557580
rect 47728 557540 47734 557552
rect 62114 557540 62120 557552
rect 62172 557540 62178 557592
rect 673178 557540 673184 557592
rect 673236 557580 673242 557592
rect 675478 557580 675484 557592
rect 673236 557552 675484 557580
rect 673236 557540 673242 557552
rect 675478 557540 675484 557552
rect 675536 557540 675542 557592
rect 674282 555228 674288 555280
rect 674340 555268 674346 555280
rect 675386 555268 675392 555280
rect 674340 555240 675392 555268
rect 674340 555228 674346 555240
rect 675386 555228 675392 555240
rect 675444 555228 675450 555280
rect 672994 554752 673000 554804
rect 673052 554792 673058 554804
rect 675294 554792 675300 554804
rect 673052 554764 675300 554792
rect 673052 554752 673058 554764
rect 675294 554752 675300 554764
rect 675352 554752 675358 554804
rect 674558 554140 674564 554192
rect 674616 554180 674622 554192
rect 675294 554180 675300 554192
rect 674616 554152 675300 554180
rect 674616 554140 674622 554152
rect 675294 554140 675300 554152
rect 675352 554140 675358 554192
rect 658918 554004 658924 554056
rect 658976 554044 658982 554056
rect 675294 554044 675300 554056
rect 658976 554016 675300 554044
rect 658976 554004 658982 554016
rect 675294 554004 675300 554016
rect 675352 554004 675358 554056
rect 672902 553460 672908 553512
rect 672960 553500 672966 553512
rect 675386 553500 675392 553512
rect 672960 553472 675392 553500
rect 672960 553460 672966 553472
rect 675386 553460 675392 553472
rect 675444 553460 675450 553512
rect 651558 550604 651564 550656
rect 651616 550644 651622 550656
rect 661678 550644 661684 550656
rect 651616 550616 661684 550644
rect 651616 550604 651622 550616
rect 661678 550604 661684 550616
rect 661736 550604 661742 550656
rect 674926 549176 674932 549228
rect 674984 549216 674990 549228
rect 675294 549216 675300 549228
rect 674984 549188 675300 549216
rect 674984 549176 674990 549188
rect 675294 549176 675300 549188
rect 675352 549176 675358 549228
rect 674742 548292 674748 548344
rect 674800 548332 674806 548344
rect 675294 548332 675300 548344
rect 674800 548304 675300 548332
rect 674800 548292 674806 548304
rect 675294 548292 675300 548304
rect 675352 548292 675358 548344
rect 31662 547136 31668 547188
rect 31720 547176 31726 547188
rect 35802 547176 35808 547188
rect 31720 547148 35808 547176
rect 31720 547136 31726 547148
rect 35802 547136 35808 547148
rect 35860 547176 35866 547188
rect 55858 547176 55864 547188
rect 35860 547148 55864 547176
rect 35860 547136 35866 547148
rect 55858 547136 55864 547148
rect 55916 547136 55922 547188
rect 31018 542988 31024 543040
rect 31076 543028 31082 543040
rect 41782 543028 41788 543040
rect 31076 543000 41788 543028
rect 31076 542988 31082 543000
rect 41782 542988 41788 543000
rect 41840 542988 41846 543040
rect 40678 542308 40684 542360
rect 40736 542348 40742 542360
rect 42702 542348 42708 542360
rect 40736 542320 42708 542348
rect 40736 542308 40742 542320
rect 42702 542308 42708 542320
rect 42760 542308 42766 542360
rect 41782 541016 41788 541068
rect 41840 541016 41846 541068
rect 41800 540796 41828 541016
rect 41782 540744 41788 540796
rect 41840 540744 41846 540796
rect 43162 539588 43168 539640
rect 43220 539628 43226 539640
rect 44818 539628 44824 539640
rect 43220 539600 44824 539628
rect 43220 539588 43226 539600
rect 44818 539588 44824 539600
rect 44876 539588 44882 539640
rect 42058 538908 42064 538960
rect 42116 538948 42122 538960
rect 42702 538948 42708 538960
rect 42116 538920 42708 538948
rect 42116 538908 42122 538920
rect 42702 538908 42708 538920
rect 42760 538908 42766 538960
rect 44542 538268 44548 538280
rect 42076 538240 44548 538268
rect 42076 537124 42104 538240
rect 44542 538228 44548 538240
rect 44600 538228 44606 538280
rect 42150 538160 42156 538212
rect 42208 538200 42214 538212
rect 43162 538200 43168 538212
rect 42208 538172 43168 538200
rect 42208 538160 42214 538172
rect 43162 538160 43168 538172
rect 43220 538160 43226 538212
rect 42058 537072 42064 537124
rect 42116 537072 42122 537124
rect 42610 536800 42616 536852
rect 42668 536840 42674 536852
rect 44450 536840 44456 536852
rect 42668 536812 44456 536840
rect 42668 536800 42674 536812
rect 44450 536800 44456 536812
rect 44508 536800 44514 536852
rect 651558 536800 651564 536852
rect 651616 536840 651622 536852
rect 664530 536840 664536 536852
rect 651616 536812 664536 536840
rect 651616 536800 651622 536812
rect 664530 536800 664536 536812
rect 664588 536800 664594 536852
rect 42610 535984 42616 536036
rect 42668 535984 42674 536036
rect 42150 535780 42156 535832
rect 42208 535820 42214 535832
rect 42628 535820 42656 535984
rect 42208 535792 42656 535820
rect 42208 535780 42214 535792
rect 668670 535712 668676 535764
rect 668728 535752 668734 535764
rect 676214 535752 676220 535764
rect 668728 535724 676220 535752
rect 668728 535712 668734 535724
rect 676214 535712 676220 535724
rect 676272 535712 676278 535764
rect 663058 535576 663064 535628
rect 663116 535616 663122 535628
rect 676030 535616 676036 535628
rect 663116 535588 676036 535616
rect 663116 535576 663122 535588
rect 676030 535576 676036 535588
rect 676088 535576 676094 535628
rect 42058 535236 42064 535288
rect 42116 535276 42122 535288
rect 43070 535276 43076 535288
rect 42116 535248 43076 535276
rect 42116 535236 42122 535248
rect 43070 535236 43076 535248
rect 43128 535236 43134 535288
rect 673730 534896 673736 534948
rect 673788 534936 673794 534948
rect 676030 534936 676036 534948
rect 673788 534908 676036 534936
rect 673788 534896 673794 534908
rect 676030 534896 676036 534908
rect 676088 534896 676094 534948
rect 661770 534216 661776 534268
rect 661828 534256 661834 534268
rect 676214 534256 676220 534268
rect 661828 534228 676220 534256
rect 661828 534216 661834 534228
rect 676214 534216 676220 534228
rect 676272 534216 676278 534268
rect 673914 534080 673920 534132
rect 673972 534120 673978 534132
rect 676030 534120 676036 534132
rect 673972 534092 676036 534120
rect 673972 534080 673978 534092
rect 676030 534080 676036 534092
rect 676088 534080 676094 534132
rect 42150 533944 42156 533996
rect 42208 533984 42214 533996
rect 42610 533984 42616 533996
rect 42208 533956 42616 533984
rect 42208 533944 42214 533956
rect 42610 533944 42616 533956
rect 42668 533944 42674 533996
rect 672442 532856 672448 532908
rect 672500 532896 672506 532908
rect 676214 532896 676220 532908
rect 672500 532868 676220 532896
rect 672500 532856 672506 532868
rect 676214 532856 676220 532868
rect 676272 532856 676278 532908
rect 51810 532720 51816 532772
rect 51868 532760 51874 532772
rect 62114 532760 62120 532772
rect 51868 532732 62120 532760
rect 51868 532720 51874 532732
rect 62114 532720 62120 532732
rect 62172 532720 62178 532772
rect 42150 531428 42156 531480
rect 42208 531468 42214 531480
rect 42610 531468 42616 531480
rect 42208 531440 42616 531468
rect 42208 531428 42214 531440
rect 42610 531428 42616 531440
rect 42668 531428 42674 531480
rect 42610 531292 42616 531344
rect 42668 531332 42674 531344
rect 42978 531332 42984 531344
rect 42668 531304 42984 531332
rect 42668 531292 42674 531304
rect 42978 531292 42984 531304
rect 43036 531292 43042 531344
rect 672534 531292 672540 531344
rect 672592 531332 672598 531344
rect 676214 531332 676220 531344
rect 672592 531304 676220 531332
rect 672592 531292 672598 531304
rect 676214 531292 676220 531304
rect 676272 531292 676278 531344
rect 674466 530408 674472 530460
rect 674524 530448 674530 530460
rect 676030 530448 676036 530460
rect 674524 530420 676036 530448
rect 674524 530408 674530 530420
rect 676030 530408 676036 530420
rect 676088 530408 676094 530460
rect 42150 530068 42156 530120
rect 42208 530108 42214 530120
rect 42610 530108 42616 530120
rect 42208 530080 42616 530108
rect 42208 530068 42214 530080
rect 42610 530068 42616 530080
rect 42668 530068 42674 530120
rect 672626 530000 672632 530052
rect 672684 530040 672690 530052
rect 676214 530040 676220 530052
rect 672684 530012 676220 530040
rect 672684 530000 672690 530012
rect 676214 530000 676220 530012
rect 676272 530000 676278 530052
rect 42334 529632 42340 529644
rect 42260 529604 42340 529632
rect 42150 529456 42156 529508
rect 42208 529496 42214 529508
rect 42260 529496 42288 529604
rect 42334 529592 42340 529604
rect 42392 529592 42398 529644
rect 42208 529468 42288 529496
rect 42208 529456 42214 529468
rect 674650 528844 674656 528896
rect 674708 528884 674714 528896
rect 676030 528884 676036 528896
rect 674708 528856 676036 528884
rect 674708 528844 674714 528856
rect 676030 528844 676036 528856
rect 676088 528844 676094 528896
rect 673362 528776 673368 528828
rect 673420 528816 673426 528828
rect 676214 528816 676220 528828
rect 673420 528788 676220 528816
rect 673420 528776 673426 528788
rect 676214 528776 676220 528788
rect 676272 528776 676278 528828
rect 672810 528640 672816 528692
rect 672868 528680 672874 528692
rect 676122 528680 676128 528692
rect 672868 528652 676128 528680
rect 672868 528640 672874 528652
rect 676122 528640 676128 528652
rect 676180 528640 676186 528692
rect 42978 528572 42984 528624
rect 43036 528612 43042 528624
rect 44358 528612 44364 528624
rect 43036 528584 44364 528612
rect 43036 528572 43042 528584
rect 44358 528572 44364 528584
rect 44416 528572 44422 528624
rect 673822 528368 673828 528420
rect 673880 528408 673886 528420
rect 676030 528408 676036 528420
rect 673880 528380 676036 528408
rect 673880 528368 673886 528380
rect 676030 528368 676036 528380
rect 676088 528368 676094 528420
rect 42058 527212 42064 527264
rect 42116 527252 42122 527264
rect 42334 527252 42340 527264
rect 42116 527224 42340 527252
rect 42116 527212 42122 527224
rect 42334 527212 42340 527224
rect 42392 527212 42398 527264
rect 42150 527144 42156 527196
rect 42208 527184 42214 527196
rect 42978 527184 42984 527196
rect 42208 527156 42984 527184
rect 42208 527144 42214 527156
rect 42978 527144 42984 527156
rect 43036 527144 43042 527196
rect 674374 526736 674380 526788
rect 674432 526776 674438 526788
rect 676030 526776 676036 526788
rect 674432 526748 676036 526776
rect 674432 526736 674438 526748
rect 676030 526736 676036 526748
rect 676088 526736 676094 526788
rect 42150 526600 42156 526652
rect 42208 526640 42214 526652
rect 42610 526640 42616 526652
rect 42208 526612 42616 526640
rect 42208 526600 42214 526612
rect 42610 526600 42616 526612
rect 42668 526600 42674 526652
rect 674190 526328 674196 526380
rect 674248 526368 674254 526380
rect 676030 526368 676036 526380
rect 674248 526340 676036 526368
rect 674248 526328 674254 526340
rect 676030 526328 676036 526340
rect 676088 526328 676094 526380
rect 673270 525920 673276 525972
rect 673328 525960 673334 525972
rect 676214 525960 676220 525972
rect 673328 525932 676220 525960
rect 673328 525920 673334 525932
rect 676214 525920 676220 525932
rect 676272 525920 676278 525972
rect 668670 524424 668676 524476
rect 668728 524464 668734 524476
rect 683114 524464 683120 524476
rect 668728 524436 683120 524464
rect 668728 524424 668734 524436
rect 683114 524424 683120 524436
rect 683172 524424 683178 524476
rect 651558 522996 651564 523048
rect 651616 523036 651622 523048
rect 663150 523036 663156 523048
rect 651616 523008 663156 523036
rect 651616 522996 651622 523008
rect 663150 522996 663156 523008
rect 663208 522996 663214 523048
rect 676122 520956 676128 521008
rect 676180 520996 676186 521008
rect 683298 520996 683304 521008
rect 676180 520968 683304 520996
rect 676180 520956 676186 520968
rect 683298 520956 683304 520968
rect 683356 520956 683362 521008
rect 676030 520888 676036 520940
rect 676088 520928 676094 520940
rect 683666 520928 683672 520940
rect 676088 520900 683672 520928
rect 676088 520888 676094 520900
rect 683666 520888 683672 520900
rect 683724 520888 683730 520940
rect 40678 518916 40684 518968
rect 40736 518956 40742 518968
rect 62114 518956 62120 518968
rect 40736 518928 62120 518956
rect 40736 518916 40742 518928
rect 62114 518916 62120 518928
rect 62172 518916 62178 518968
rect 651558 510620 651564 510672
rect 651616 510660 651622 510672
rect 665818 510660 665824 510672
rect 651616 510632 665824 510660
rect 651616 510620 651622 510632
rect 665818 510620 665824 510632
rect 665876 510620 665882 510672
rect 49050 506472 49056 506524
rect 49108 506512 49114 506524
rect 62114 506512 62120 506524
rect 49108 506484 62120 506512
rect 49108 506472 49114 506484
rect 62114 506472 62120 506484
rect 62172 506472 62178 506524
rect 40862 497428 40868 497480
rect 40920 497468 40926 497480
rect 62758 497468 62764 497480
rect 40920 497440 62764 497468
rect 40920 497428 40926 497440
rect 62758 497428 62764 497440
rect 62816 497428 62822 497480
rect 651558 496816 651564 496868
rect 651616 496856 651622 496868
rect 658918 496856 658924 496868
rect 651616 496828 658924 496856
rect 651616 496816 651622 496828
rect 658918 496816 658924 496828
rect 658976 496816 658982 496868
rect 53190 492668 53196 492720
rect 53248 492708 53254 492720
rect 62114 492708 62120 492720
rect 53248 492680 62120 492708
rect 53248 492668 53254 492680
rect 62114 492668 62120 492680
rect 62172 492668 62178 492720
rect 664438 491648 664444 491700
rect 664496 491688 664502 491700
rect 675938 491688 675944 491700
rect 664496 491660 675944 491688
rect 664496 491648 664502 491660
rect 675938 491648 675944 491660
rect 675996 491648 676002 491700
rect 660298 491512 660304 491564
rect 660356 491552 660362 491564
rect 676030 491552 676036 491564
rect 660356 491524 676036 491552
rect 660356 491512 660362 491524
rect 676030 491512 676036 491524
rect 676088 491512 676094 491564
rect 659010 491376 659016 491428
rect 659068 491416 659074 491428
rect 676030 491416 676036 491428
rect 659068 491388 676036 491416
rect 659068 491376 659074 491388
rect 676030 491376 676036 491388
rect 676088 491376 676094 491428
rect 675938 489268 675944 489320
rect 675996 489308 676002 489320
rect 677318 489308 677324 489320
rect 675996 489280 677324 489308
rect 675996 489268 676002 489280
rect 677318 489268 677324 489280
rect 677376 489268 677382 489320
rect 675938 488588 675944 488640
rect 675996 488628 676002 488640
rect 676122 488628 676128 488640
rect 675996 488600 676128 488628
rect 675996 488588 676002 488600
rect 676122 488588 676128 488600
rect 676180 488588 676186 488640
rect 675938 488452 675944 488504
rect 675996 488492 676002 488504
rect 677502 488492 677508 488504
rect 675996 488464 677508 488492
rect 675996 488452 676002 488464
rect 677502 488452 677508 488464
rect 677560 488452 677566 488504
rect 674926 488316 674932 488368
rect 674984 488356 674990 488368
rect 675938 488356 675944 488368
rect 674984 488328 675944 488356
rect 674984 488316 674990 488328
rect 675938 488316 675944 488328
rect 675996 488316 676002 488368
rect 675846 487976 675852 488028
rect 675904 488016 675910 488028
rect 677226 488016 677232 488028
rect 675904 487988 677232 488016
rect 675904 487976 675910 487988
rect 677226 487976 677232 487988
rect 677284 487976 677290 488028
rect 674282 486004 674288 486056
rect 674340 486044 674346 486056
rect 675938 486044 675944 486056
rect 674340 486016 675944 486044
rect 674340 486004 674346 486016
rect 675938 486004 675944 486016
rect 675996 486004 676002 486056
rect 673086 484576 673092 484628
rect 673144 484616 673150 484628
rect 675938 484616 675944 484628
rect 673144 484588 675944 484616
rect 673144 484576 673150 484588
rect 675938 484576 675944 484588
rect 675996 484576 676002 484628
rect 651558 484372 651564 484424
rect 651616 484412 651622 484424
rect 660390 484412 660396 484424
rect 651616 484384 660396 484412
rect 651616 484372 651622 484384
rect 660390 484372 660396 484384
rect 660448 484372 660454 484424
rect 671982 484372 671988 484424
rect 672040 484412 672046 484424
rect 675846 484412 675852 484424
rect 672040 484384 675852 484412
rect 672040 484372 672046 484384
rect 675846 484372 675852 484384
rect 675904 484372 675910 484424
rect 674558 483556 674564 483608
rect 674616 483596 674622 483608
rect 675938 483596 675944 483608
rect 674616 483568 675944 483596
rect 674616 483556 674622 483568
rect 675938 483556 675944 483568
rect 675996 483556 676002 483608
rect 673178 483080 673184 483132
rect 673236 483120 673242 483132
rect 675938 483120 675944 483132
rect 673236 483092 675944 483120
rect 673236 483080 673242 483092
rect 675938 483080 675944 483092
rect 675996 483080 676002 483132
rect 672994 481856 673000 481908
rect 673052 481896 673058 481908
rect 675846 481896 675852 481908
rect 673052 481868 675852 481896
rect 673052 481856 673058 481868
rect 675846 481856 675852 481868
rect 675904 481856 675910 481908
rect 672902 481720 672908 481772
rect 672960 481760 672966 481772
rect 675938 481760 675944 481772
rect 672960 481732 675944 481760
rect 672960 481720 672966 481732
rect 675938 481720 675944 481732
rect 675996 481720 676002 481772
rect 50522 480224 50528 480276
rect 50580 480264 50586 480276
rect 62114 480264 62120 480276
rect 50580 480236 62120 480264
rect 50580 480224 50586 480236
rect 62114 480224 62120 480236
rect 62172 480224 62178 480276
rect 674190 480224 674196 480276
rect 674248 480264 674254 480276
rect 678974 480264 678980 480276
rect 674248 480236 678980 480264
rect 674248 480224 674254 480236
rect 678974 480224 678980 480236
rect 679032 480224 679038 480276
rect 651650 470568 651656 470620
rect 651708 470608 651714 470620
rect 664438 470608 664444 470620
rect 651708 470580 664444 470608
rect 651708 470568 651714 470580
rect 664438 470568 664444 470580
rect 664496 470568 664502 470620
rect 55950 466420 55956 466472
rect 56008 466460 56014 466472
rect 62114 466460 62120 466472
rect 56008 466432 62120 466460
rect 56008 466420 56014 466432
rect 62114 466420 62120 466432
rect 62172 466420 62178 466472
rect 651558 456764 651564 456816
rect 651616 456804 651622 456816
rect 671522 456804 671528 456816
rect 651616 456776 671528 456804
rect 651616 456764 651622 456776
rect 671522 456764 671528 456776
rect 671580 456764 671586 456816
rect 50430 454044 50436 454096
rect 50488 454084 50494 454096
rect 62114 454084 62120 454096
rect 50488 454056 62120 454084
rect 50488 454044 50494 454056
rect 62114 454044 62120 454056
rect 62172 454044 62178 454096
rect 651558 444388 651564 444440
rect 651616 444428 651622 444440
rect 659010 444428 659016 444440
rect 651616 444400 659016 444428
rect 651616 444388 651622 444400
rect 659010 444388 659016 444400
rect 659068 444388 659074 444440
rect 44910 440240 44916 440292
rect 44968 440280 44974 440292
rect 62114 440280 62120 440292
rect 44968 440252 62120 440280
rect 44968 440240 44974 440252
rect 62114 440240 62120 440252
rect 62172 440240 62178 440292
rect 40678 432556 40684 432608
rect 40736 432596 40742 432608
rect 41782 432596 41788 432608
rect 40736 432568 41788 432596
rect 40736 432556 40742 432568
rect 41782 432556 41788 432568
rect 41840 432556 41846 432608
rect 43346 430584 43352 430636
rect 43404 430624 43410 430636
rect 51810 430624 51816 430636
rect 43404 430596 51816 430624
rect 43404 430584 43410 430596
rect 51810 430584 51816 430596
rect 51868 430584 51874 430636
rect 651558 430584 651564 430636
rect 651616 430624 651622 430636
rect 660298 430624 660304 430636
rect 651616 430596 660304 430624
rect 651616 430584 651622 430596
rect 660298 430584 660304 430596
rect 660356 430584 660362 430636
rect 40862 430108 40868 430160
rect 40920 430148 40926 430160
rect 41782 430148 41788 430160
rect 40920 430120 41788 430148
rect 40920 430108 40926 430120
rect 41782 430108 41788 430120
rect 41840 430108 41846 430160
rect 54570 427796 54576 427848
rect 54628 427836 54634 427848
rect 62114 427836 62120 427848
rect 54628 427808 62120 427836
rect 54628 427796 54634 427808
rect 62114 427796 62120 427808
rect 62172 427796 62178 427848
rect 40770 425688 40776 425740
rect 40828 425728 40834 425740
rect 41782 425728 41788 425740
rect 40828 425700 41788 425728
rect 40828 425688 40834 425700
rect 41782 425688 41788 425700
rect 41840 425688 41846 425740
rect 41782 419432 41788 419484
rect 41840 419472 41846 419484
rect 44818 419472 44824 419484
rect 41840 419444 44824 419472
rect 41840 419432 41846 419444
rect 44818 419432 44824 419444
rect 44876 419432 44882 419484
rect 651558 416780 651564 416832
rect 651616 416820 651622 416832
rect 663058 416820 663064 416832
rect 651616 416792 663064 416820
rect 651616 416780 651622 416792
rect 663058 416780 663064 416792
rect 663116 416780 663122 416832
rect 51810 415420 51816 415472
rect 51868 415460 51874 415472
rect 62114 415460 62120 415472
rect 51868 415432 62120 415460
rect 51868 415420 51874 415432
rect 62114 415420 62120 415432
rect 62172 415420 62178 415472
rect 32398 414808 32404 414860
rect 32456 414848 32462 414860
rect 41874 414848 41880 414860
rect 32456 414820 41880 414848
rect 32456 414808 32462 414820
rect 41874 414808 41880 414820
rect 41932 414808 41938 414860
rect 31018 414672 31024 414724
rect 31076 414712 31082 414724
rect 42518 414712 42524 414724
rect 31076 414684 42524 414712
rect 31076 414672 31082 414684
rect 42518 414672 42524 414684
rect 42576 414672 42582 414724
rect 41874 413380 41880 413432
rect 41932 413380 41938 413432
rect 41892 413160 41920 413380
rect 41874 413108 41880 413160
rect 41932 413108 41938 413160
rect 42150 410660 42156 410712
rect 42208 410700 42214 410712
rect 47670 410700 47676 410712
rect 42208 410672 47676 410700
rect 42208 410660 42214 410672
rect 47670 410660 47676 410672
rect 47728 410660 47734 410712
rect 42058 408144 42064 408196
rect 42116 408184 42122 408196
rect 43070 408184 43076 408196
rect 42116 408156 43076 408184
rect 42116 408144 42122 408156
rect 43070 408144 43076 408156
rect 43128 408144 43134 408196
rect 42150 407600 42156 407652
rect 42208 407640 42214 407652
rect 42518 407640 42524 407652
rect 42208 407612 42524 407640
rect 42208 407600 42214 407612
rect 42518 407600 42524 407612
rect 42576 407600 42582 407652
rect 42058 406784 42064 406836
rect 42116 406824 42122 406836
rect 44450 406824 44456 406836
rect 42116 406796 44456 406824
rect 42116 406784 42122 406796
rect 44450 406784 44456 406796
rect 44508 406784 44514 406836
rect 652018 404336 652024 404388
rect 652076 404376 652082 404388
rect 661770 404376 661776 404388
rect 652076 404348 661776 404376
rect 652076 404336 652082 404348
rect 661770 404336 661776 404348
rect 661828 404336 661834 404388
rect 42150 403860 42156 403912
rect 42208 403900 42214 403912
rect 42794 403900 42800 403912
rect 42208 403872 42800 403900
rect 42208 403860 42214 403872
rect 42794 403860 42800 403872
rect 42852 403860 42858 403912
rect 664530 403384 664536 403436
rect 664588 403424 664594 403436
rect 676214 403424 676220 403436
rect 664588 403396 676220 403424
rect 664588 403384 664594 403396
rect 676214 403384 676220 403396
rect 676272 403384 676278 403436
rect 663150 403248 663156 403300
rect 663208 403288 663214 403300
rect 676214 403288 676220 403300
rect 663208 403260 676220 403288
rect 663208 403248 663214 403260
rect 676214 403248 676220 403260
rect 676272 403248 676278 403300
rect 661678 403112 661684 403164
rect 661736 403152 661742 403164
rect 676398 403152 676404 403164
rect 661736 403124 676404 403152
rect 661736 403112 661742 403124
rect 676398 403112 676404 403124
rect 676456 403112 676462 403164
rect 42150 402908 42156 402960
rect 42208 402948 42214 402960
rect 44358 402948 44364 402960
rect 42208 402920 44364 402948
rect 42208 402908 42214 402920
rect 44358 402908 44364 402920
rect 44416 402908 44422 402960
rect 43530 401616 43536 401668
rect 43588 401656 43594 401668
rect 62114 401656 62120 401668
rect 43588 401628 62120 401656
rect 43588 401616 43594 401628
rect 62114 401616 62120 401628
rect 62172 401616 62178 401668
rect 673178 401616 673184 401668
rect 673236 401656 673242 401668
rect 676214 401656 676220 401668
rect 673236 401628 676220 401656
rect 673236 401616 673242 401628
rect 676214 401616 676220 401628
rect 676272 401616 676278 401668
rect 673362 400256 673368 400308
rect 673420 400296 673426 400308
rect 676214 400296 676220 400308
rect 673420 400268 676220 400296
rect 673420 400256 673426 400268
rect 676214 400256 676220 400268
rect 676272 400256 676278 400308
rect 673270 400188 673276 400240
rect 673328 400228 673334 400240
rect 676122 400228 676128 400240
rect 673328 400200 676128 400228
rect 673328 400188 673334 400200
rect 676122 400188 676128 400200
rect 676180 400188 676186 400240
rect 674742 399576 674748 399628
rect 674800 399616 674806 399628
rect 676214 399616 676220 399628
rect 674800 399588 676220 399616
rect 674800 399576 674806 399588
rect 676214 399576 676220 399588
rect 676272 399576 676278 399628
rect 675018 398216 675024 398268
rect 675076 398256 675082 398268
rect 676030 398256 676036 398268
rect 675076 398228 676036 398256
rect 675076 398216 675082 398228
rect 676030 398216 676036 398228
rect 676088 398216 676094 398268
rect 674926 397468 674932 397520
rect 674984 397508 674990 397520
rect 676030 397508 676036 397520
rect 674984 397480 676036 397508
rect 674984 397468 674990 397480
rect 676030 397468 676036 397480
rect 676088 397468 676094 397520
rect 674650 394000 674656 394052
rect 674708 394040 674714 394052
rect 676030 394040 676036 394052
rect 674708 394012 676036 394040
rect 674708 394000 674714 394012
rect 676030 394000 676036 394012
rect 676088 394000 676094 394052
rect 673086 393320 673092 393372
rect 673144 393360 673150 393372
rect 676214 393360 676220 393372
rect 673144 393332 676220 393360
rect 673144 393320 673150 393332
rect 676214 393320 676220 393332
rect 676272 393320 676278 393372
rect 670234 391960 670240 392012
rect 670292 392000 670298 392012
rect 683114 392000 683120 392012
rect 670292 391972 683120 392000
rect 670292 391960 670298 391972
rect 683114 391960 683120 391972
rect 683172 391960 683178 392012
rect 651558 390532 651564 390584
rect 651616 390572 651622 390584
rect 671430 390572 671436 390584
rect 651616 390544 671436 390572
rect 651616 390532 651622 390544
rect 671430 390532 671436 390544
rect 671488 390532 671494 390584
rect 43622 389172 43628 389224
rect 43680 389212 43686 389224
rect 62114 389212 62120 389224
rect 43680 389184 62120 389212
rect 43680 389172 43686 389184
rect 62114 389172 62120 389184
rect 62172 389172 62178 389224
rect 35710 387744 35716 387796
rect 35768 387784 35774 387796
rect 44266 387784 44272 387796
rect 35768 387756 44272 387784
rect 35768 387744 35774 387756
rect 44266 387744 44272 387756
rect 44324 387744 44330 387796
rect 675202 387744 675208 387796
rect 675260 387784 675266 387796
rect 676950 387784 676956 387796
rect 675260 387756 676956 387784
rect 675260 387744 675266 387756
rect 676950 387744 676956 387756
rect 677008 387744 677014 387796
rect 675110 387676 675116 387728
rect 675168 387716 675174 387728
rect 676490 387716 676496 387728
rect 675168 387688 676496 387716
rect 675168 387676 675174 387688
rect 676490 387676 676496 387688
rect 676548 387676 676554 387728
rect 35802 387608 35808 387660
rect 35860 387648 35866 387660
rect 50522 387648 50528 387660
rect 35860 387620 50528 387648
rect 35860 387608 35866 387620
rect 50522 387608 50528 387620
rect 50580 387608 50586 387660
rect 675294 387608 675300 387660
rect 675352 387648 675358 387660
rect 678238 387648 678244 387660
rect 675352 387620 678244 387648
rect 675352 387608 675358 387620
rect 678238 387608 678244 387620
rect 678296 387608 678302 387660
rect 35618 387472 35624 387524
rect 35676 387512 35682 387524
rect 53190 387512 53196 387524
rect 35676 387484 53196 387512
rect 35676 387472 35682 387484
rect 53190 387472 53196 387484
rect 53248 387472 53254 387524
rect 35802 387336 35808 387388
rect 35860 387376 35866 387388
rect 55950 387376 55956 387388
rect 35860 387348 55956 387376
rect 35860 387336 35866 387348
rect 55950 387336 55956 387348
rect 56008 387336 56014 387388
rect 675018 386112 675024 386164
rect 675076 386152 675082 386164
rect 675386 386152 675392 386164
rect 675076 386124 675392 386152
rect 675076 386112 675082 386124
rect 675386 386112 675392 386124
rect 675444 386112 675450 386164
rect 675018 385976 675024 386028
rect 675076 386016 675082 386028
rect 675294 386016 675300 386028
rect 675076 385988 675300 386016
rect 675076 385976 675082 385988
rect 675294 385976 675300 385988
rect 675352 385976 675358 386028
rect 675202 385772 675208 385824
rect 675260 385812 675266 385824
rect 675260 385784 675432 385812
rect 675260 385772 675266 385784
rect 675404 385620 675432 385784
rect 675386 385568 675392 385620
rect 675444 385568 675450 385620
rect 675018 383868 675024 383920
rect 675076 383908 675082 383920
rect 675294 383908 675300 383920
rect 675076 383880 675300 383908
rect 675076 383868 675082 383880
rect 675294 383868 675300 383880
rect 675352 383868 675358 383920
rect 674926 383052 674932 383104
rect 674984 383092 674990 383104
rect 675386 383092 675392 383104
rect 674984 383064 675392 383092
rect 674984 383052 674990 383064
rect 675386 383052 675392 383064
rect 675444 383052 675450 383104
rect 675110 381080 675116 381132
rect 675168 381120 675174 381132
rect 675386 381120 675392 381132
rect 675168 381092 675392 381120
rect 675168 381080 675174 381092
rect 675386 381080 675392 381092
rect 675444 381080 675450 381132
rect 651558 378156 651564 378208
rect 651616 378196 651622 378208
rect 664530 378196 664536 378208
rect 651616 378168 664536 378196
rect 651616 378156 651622 378168
rect 664530 378156 664536 378168
rect 664588 378156 664594 378208
rect 673086 376728 673092 376780
rect 673144 376768 673150 376780
rect 675294 376768 675300 376780
rect 673144 376740 675300 376768
rect 673144 376728 673150 376740
rect 675294 376728 675300 376740
rect 675352 376728 675358 376780
rect 674650 376660 674656 376712
rect 674708 376700 674714 376712
rect 675478 376700 675484 376712
rect 674708 376672 675484 376700
rect 674708 376660 674714 376672
rect 675478 376660 675484 376672
rect 675536 376660 675542 376712
rect 35802 375980 35808 376032
rect 35860 376020 35866 376032
rect 41506 376020 41512 376032
rect 35860 375992 41512 376020
rect 35860 375980 35866 375992
rect 41506 375980 41512 375992
rect 41564 376020 41570 376032
rect 53190 376020 53196 376032
rect 41564 375992 53196 376020
rect 41564 375980 41570 375992
rect 53190 375980 53196 375992
rect 53248 375980 53254 376032
rect 47670 375368 47676 375420
rect 47728 375408 47734 375420
rect 62114 375408 62120 375420
rect 47728 375380 62120 375408
rect 47728 375368 47734 375380
rect 62114 375368 62120 375380
rect 62172 375368 62178 375420
rect 31018 371832 31024 371884
rect 31076 371872 31082 371884
rect 42334 371872 42340 371884
rect 31076 371844 42340 371872
rect 31076 371832 31082 371844
rect 42334 371832 42340 371844
rect 42392 371832 42398 371884
rect 40862 371220 40868 371272
rect 40920 371260 40926 371272
rect 42702 371260 42708 371272
rect 40920 371232 42708 371260
rect 40920 371220 40926 371232
rect 42702 371220 42708 371232
rect 42760 371220 42766 371272
rect 40678 370540 40684 370592
rect 40736 370580 40742 370592
rect 41782 370580 41788 370592
rect 40736 370552 41788 370580
rect 40736 370540 40742 370552
rect 41782 370540 41788 370552
rect 41840 370540 41846 370592
rect 42150 369656 42156 369708
rect 42208 369696 42214 369708
rect 42334 369696 42340 369708
rect 42208 369668 42340 369696
rect 42208 369656 42214 369668
rect 42334 369656 42340 369668
rect 42392 369656 42398 369708
rect 42150 368092 42156 368144
rect 42208 368132 42214 368144
rect 42702 368132 42708 368144
rect 42208 368104 42708 368132
rect 42208 368092 42214 368104
rect 42702 368092 42708 368104
rect 42760 368092 42766 368144
rect 42150 366800 42156 366852
rect 42208 366840 42214 366852
rect 42702 366840 42708 366852
rect 42208 366812 42708 366840
rect 42208 366800 42214 366812
rect 42702 366800 42708 366812
rect 42760 366800 42766 366852
rect 42150 364964 42156 365016
rect 42208 365004 42214 365016
rect 43070 365004 43076 365016
rect 42208 364976 43076 365004
rect 42208 364964 42214 364976
rect 43070 364964 43076 364976
rect 43128 364964 43134 365016
rect 652018 364352 652024 364404
rect 652076 364392 652082 364404
rect 674374 364392 674380 364404
rect 652076 364364 674380 364392
rect 652076 364352 652082 364364
rect 674374 364352 674380 364364
rect 674432 364352 674438 364404
rect 42150 364284 42156 364336
rect 42208 364324 42214 364336
rect 44542 364324 44548 364336
rect 42208 364296 44548 364324
rect 42208 364284 42214 364296
rect 44542 364284 44548 364296
rect 44600 364284 44606 364336
rect 42702 364216 42708 364268
rect 42760 364256 42766 364268
rect 49050 364256 49056 364268
rect 42760 364228 49056 364256
rect 42760 364216 42766 364228
rect 49050 364216 49056 364228
rect 49108 364216 49114 364268
rect 51902 362924 51908 362976
rect 51960 362964 51966 362976
rect 62114 362964 62120 362976
rect 51960 362936 62120 362964
rect 51960 362924 51966 362936
rect 62114 362924 62120 362936
rect 62172 362924 62178 362976
rect 42058 360680 42064 360732
rect 42116 360720 42122 360732
rect 42978 360720 42984 360732
rect 42116 360692 42984 360720
rect 42116 360680 42122 360692
rect 42978 360680 42984 360692
rect 43036 360680 43042 360732
rect 42150 359456 42156 359508
rect 42208 359496 42214 359508
rect 42886 359496 42892 359508
rect 42208 359468 42892 359496
rect 42208 359456 42214 359468
rect 42886 359456 42892 359468
rect 42944 359456 42950 359508
rect 665818 357824 665824 357876
rect 665876 357864 665882 357876
rect 675938 357864 675944 357876
rect 665876 357836 675944 357864
rect 665876 357824 665882 357836
rect 675938 357824 675944 357836
rect 675996 357824 676002 357876
rect 660390 357688 660396 357740
rect 660448 357728 660454 357740
rect 676030 357728 676036 357740
rect 660448 357700 676036 357728
rect 660448 357688 660454 357700
rect 676030 357688 676036 357700
rect 676088 357688 676094 357740
rect 658918 357552 658924 357604
rect 658976 357592 658982 357604
rect 675846 357592 675852 357604
rect 658976 357564 675852 357592
rect 658976 357552 658982 357564
rect 675846 357552 675852 357564
rect 675904 357552 675910 357604
rect 673178 357484 673184 357536
rect 673236 357524 673242 357536
rect 676030 357524 676036 357536
rect 673236 357496 676036 357524
rect 673236 357484 673242 357496
rect 676030 357484 676036 357496
rect 676088 357484 676094 357536
rect 674650 357008 674656 357060
rect 674708 357048 674714 357060
rect 676030 357048 676036 357060
rect 674708 357020 676036 357048
rect 674708 357008 674714 357020
rect 676030 357008 676036 357020
rect 676088 357008 676094 357060
rect 673270 356668 673276 356720
rect 673328 356708 673334 356720
rect 676030 356708 676036 356720
rect 673328 356680 676036 356708
rect 673328 356668 673334 356680
rect 676030 356668 676036 356680
rect 676088 356668 676094 356720
rect 674466 356192 674472 356244
rect 674524 356232 674530 356244
rect 676030 356232 676036 356244
rect 674524 356204 676036 356232
rect 674524 356192 674530 356204
rect 676030 356192 676036 356204
rect 676088 356192 676094 356244
rect 42150 355988 42156 356040
rect 42208 356028 42214 356040
rect 44450 356028 44456 356040
rect 42208 356000 44456 356028
rect 42208 355988 42214 356000
rect 44450 355988 44456 356000
rect 44508 355988 44514 356040
rect 673362 355852 673368 355904
rect 673420 355892 673426 355904
rect 676030 355892 676036 355904
rect 673420 355864 676036 355892
rect 673420 355852 673426 355864
rect 676030 355852 676036 355864
rect 676088 355852 676094 355904
rect 672902 355376 672908 355428
rect 672960 355416 672966 355428
rect 676030 355416 676036 355428
rect 672960 355388 676036 355416
rect 672960 355376 672966 355388
rect 676030 355376 676036 355388
rect 676088 355376 676094 355428
rect 673270 354560 673276 354612
rect 673328 354600 673334 354612
rect 676030 354600 676036 354612
rect 673328 354572 676036 354600
rect 673328 354560 673334 354572
rect 676030 354560 676036 354572
rect 676088 354560 676094 354612
rect 676030 351024 676036 351076
rect 676088 351064 676094 351076
rect 676766 351064 676772 351076
rect 676088 351036 676772 351064
rect 676088 351024 676094 351036
rect 676766 351024 676772 351036
rect 676824 351024 676830 351076
rect 673362 350888 673368 350940
rect 673420 350928 673426 350940
rect 676030 350928 676036 350940
rect 673420 350900 676036 350928
rect 673420 350888 673426 350900
rect 676030 350888 676036 350900
rect 676088 350888 676094 350940
rect 651558 350548 651564 350600
rect 651616 350588 651622 350600
rect 674098 350588 674104 350600
rect 651616 350560 674104 350588
rect 651616 350548 651622 350560
rect 674098 350548 674104 350560
rect 674156 350548 674162 350600
rect 674558 350548 674564 350600
rect 674616 350588 674622 350600
rect 676030 350588 676036 350600
rect 674616 350560 676036 350588
rect 674616 350548 674622 350560
rect 676030 350548 676036 350560
rect 676088 350548 676094 350600
rect 673178 349256 673184 349308
rect 673236 349296 673242 349308
rect 676030 349296 676036 349308
rect 673236 349268 676036 349296
rect 673236 349256 673242 349268
rect 676030 349256 676036 349268
rect 676088 349256 676094 349308
rect 46198 349120 46204 349172
rect 46256 349160 46262 349172
rect 62114 349160 62120 349172
rect 46256 349132 62120 349160
rect 46256 349120 46262 349132
rect 62114 349120 62120 349132
rect 62172 349120 62178 349172
rect 673086 348848 673092 348900
rect 673144 348888 673150 348900
rect 676030 348888 676036 348900
rect 673144 348860 676036 348888
rect 673144 348848 673150 348860
rect 676030 348848 676036 348860
rect 676088 348848 676094 348900
rect 672810 346400 672816 346452
rect 672868 346440 672874 346452
rect 676030 346440 676036 346452
rect 672868 346412 676036 346440
rect 672868 346400 672874 346412
rect 676030 346400 676036 346412
rect 676088 346400 676094 346452
rect 35710 344428 35716 344480
rect 35768 344468 35774 344480
rect 44910 344468 44916 344480
rect 35768 344440 44916 344468
rect 35768 344428 35774 344440
rect 44910 344428 44916 344440
rect 44968 344428 44974 344480
rect 35802 344292 35808 344344
rect 35860 344332 35866 344344
rect 51810 344332 51816 344344
rect 35860 344304 51816 344332
rect 35860 344292 35866 344304
rect 51810 344292 51816 344304
rect 51868 344292 51874 344344
rect 35618 344156 35624 344208
rect 35676 344196 35682 344208
rect 54570 344196 54576 344208
rect 35676 344168 54576 344196
rect 35676 344156 35682 344168
rect 54570 344156 54576 344168
rect 54628 344156 54634 344208
rect 651650 338104 651656 338156
rect 651708 338144 651714 338156
rect 672994 338144 673000 338156
rect 651708 338116 673000 338144
rect 651708 338104 651714 338116
rect 672994 338104 673000 338116
rect 673052 338104 673058 338156
rect 44910 336744 44916 336796
rect 44968 336784 44974 336796
rect 62114 336784 62120 336796
rect 44968 336756 62120 336784
rect 44968 336744 44974 336756
rect 62114 336744 62120 336756
rect 62172 336744 62178 336796
rect 674834 336676 674840 336728
rect 674892 336716 674898 336728
rect 675386 336716 675392 336728
rect 674892 336688 675392 336716
rect 674892 336676 674898 336688
rect 675386 336676 675392 336688
rect 675444 336676 675450 336728
rect 673362 336540 673368 336592
rect 673420 336580 673426 336592
rect 675386 336580 675392 336592
rect 673420 336552 675392 336580
rect 673420 336540 673426 336552
rect 675386 336540 675392 336552
rect 675444 336540 675450 336592
rect 30374 333208 30380 333260
rect 30432 333248 30438 333260
rect 49050 333248 49056 333260
rect 30432 333220 49056 333248
rect 30432 333208 30438 333220
rect 49050 333208 49056 333220
rect 49108 333208 49114 333260
rect 673178 332596 673184 332648
rect 673236 332636 673242 332648
rect 675386 332636 675392 332648
rect 673236 332608 675392 332636
rect 673236 332596 673242 332608
rect 675386 332596 675392 332608
rect 675444 332596 675450 332648
rect 673086 331576 673092 331628
rect 673144 331616 673150 331628
rect 675386 331616 675392 331628
rect 673144 331588 675392 331616
rect 673144 331576 673150 331588
rect 675386 331576 675392 331588
rect 675444 331576 675450 331628
rect 674558 330556 674564 330608
rect 674616 330596 674622 330608
rect 675386 330596 675392 330608
rect 674616 330568 675392 330596
rect 674616 330556 674622 330568
rect 675386 330556 675392 330568
rect 675444 330556 675450 330608
rect 675110 327632 675116 327684
rect 675168 327672 675174 327684
rect 675478 327672 675484 327684
rect 675168 327644 675484 327672
rect 675168 327632 675174 327644
rect 675478 327632 675484 327644
rect 675536 327632 675542 327684
rect 42058 326748 42064 326800
rect 42116 326788 42122 326800
rect 43070 326788 43076 326800
rect 42116 326760 43076 326788
rect 42116 326748 42122 326760
rect 43070 326748 43076 326760
rect 43128 326748 43134 326800
rect 675754 325796 675760 325848
rect 675812 325796 675818 325848
rect 675772 325644 675800 325796
rect 675754 325592 675760 325644
rect 675812 325592 675818 325644
rect 651558 324300 651564 324352
rect 651616 324340 651622 324352
rect 671614 324340 671620 324352
rect 651616 324312 671620 324340
rect 651616 324300 651622 324312
rect 671614 324300 671620 324312
rect 671672 324300 671678 324352
rect 42150 323280 42156 323332
rect 42208 323320 42214 323332
rect 42610 323320 42616 323332
rect 42208 323292 42616 323320
rect 42208 323280 42214 323292
rect 42610 323280 42616 323292
rect 42668 323280 42674 323332
rect 43714 322940 43720 322992
rect 43772 322980 43778 322992
rect 62114 322980 62120 322992
rect 43772 322952 62120 322980
rect 43772 322940 43778 322952
rect 62114 322940 62120 322952
rect 62172 322940 62178 322992
rect 42058 322872 42064 322924
rect 42116 322912 42122 322924
rect 42978 322912 42984 322924
rect 42116 322884 42984 322912
rect 42116 322872 42122 322884
rect 42978 322872 42984 322884
rect 43036 322872 43042 322924
rect 42610 321512 42616 321564
rect 42668 321552 42674 321564
rect 50430 321552 50436 321564
rect 42668 321524 50436 321552
rect 42668 321512 42674 321524
rect 50430 321512 50436 321524
rect 50488 321512 50494 321564
rect 42150 321444 42156 321496
rect 42208 321484 42214 321496
rect 42886 321484 42892 321496
rect 42208 321456 42892 321484
rect 42208 321444 42214 321456
rect 42886 321444 42892 321456
rect 42944 321444 42950 321496
rect 42150 319948 42156 320000
rect 42208 319988 42214 320000
rect 44542 319988 44548 320000
rect 42208 319960 44548 319988
rect 42208 319948 42214 319960
rect 44542 319948 44548 319960
rect 44600 319948 44606 320000
rect 42150 316684 42156 316736
rect 42208 316724 42214 316736
rect 44450 316724 44456 316736
rect 42208 316696 44456 316724
rect 42208 316684 42214 316696
rect 44450 316684 44456 316696
rect 44508 316684 44514 316736
rect 671522 313488 671528 313540
rect 671580 313528 671586 313540
rect 676214 313528 676220 313540
rect 671580 313500 676220 313528
rect 671580 313488 671586 313500
rect 676214 313488 676220 313500
rect 676272 313488 676278 313540
rect 664438 313352 664444 313404
rect 664496 313392 664502 313404
rect 676030 313392 676036 313404
rect 664496 313364 676036 313392
rect 664496 313352 664502 313364
rect 676030 313352 676036 313364
rect 676088 313352 676094 313404
rect 674650 312468 674656 312520
rect 674708 312508 674714 312520
rect 676030 312508 676036 312520
rect 674708 312480 676036 312508
rect 674708 312468 674714 312480
rect 676030 312468 676036 312480
rect 676088 312468 676094 312520
rect 659010 311992 659016 312044
rect 659068 312032 659074 312044
rect 676214 312032 676220 312044
rect 659068 312004 676220 312032
rect 659068 311992 659074 312004
rect 676214 311992 676220 312004
rect 676272 311992 676278 312044
rect 674742 311856 674748 311908
rect 674800 311896 674806 311908
rect 676214 311896 676220 311908
rect 674800 311868 676220 311896
rect 674800 311856 674806 311868
rect 676214 311856 676220 311868
rect 676272 311856 676278 311908
rect 674466 311652 674472 311704
rect 674524 311692 674530 311704
rect 676030 311692 676036 311704
rect 674524 311664 676036 311692
rect 674524 311652 674530 311664
rect 676030 311652 676036 311664
rect 676088 311652 676094 311704
rect 674650 311040 674656 311092
rect 674708 311080 674714 311092
rect 676214 311080 676220 311092
rect 674708 311052 676220 311080
rect 674708 311040 674714 311052
rect 676214 311040 676220 311052
rect 676272 311040 676278 311092
rect 672902 310632 672908 310684
rect 672960 310672 672966 310684
rect 676214 310672 676220 310684
rect 672960 310644 676220 310672
rect 672960 310632 672966 310644
rect 676214 310632 676220 310644
rect 676272 310632 676278 310684
rect 55950 310496 55956 310548
rect 56008 310536 56014 310548
rect 62114 310536 62120 310548
rect 56008 310508 62120 310536
rect 56008 310496 56014 310508
rect 62114 310496 62120 310508
rect 62172 310496 62178 310548
rect 652386 310496 652392 310548
rect 652444 310536 652450 310548
rect 672902 310536 672908 310548
rect 652444 310508 672908 310536
rect 652444 310496 652450 310508
rect 672902 310496 672908 310508
rect 672960 310496 672966 310548
rect 673270 309408 673276 309460
rect 673328 309448 673334 309460
rect 676214 309448 676220 309460
rect 673328 309420 676220 309448
rect 673328 309408 673334 309420
rect 676214 309408 676220 309420
rect 676272 309408 676278 309460
rect 673362 309340 673368 309392
rect 673420 309380 673426 309392
rect 676122 309380 676128 309392
rect 673420 309352 676128 309380
rect 673420 309340 673426 309352
rect 676122 309340 676128 309352
rect 676180 309340 676186 309392
rect 673362 309204 673368 309256
rect 673420 309244 673426 309256
rect 676306 309244 676312 309256
rect 673420 309216 676312 309244
rect 673420 309204 673426 309216
rect 676306 309204 676312 309216
rect 676364 309204 676370 309256
rect 41966 307028 41972 307080
rect 42024 307068 42030 307080
rect 51902 307068 51908 307080
rect 42024 307040 51908 307068
rect 42024 307028 42030 307040
rect 51902 307028 51908 307040
rect 51960 307028 51966 307080
rect 674558 304512 674564 304564
rect 674616 304552 674622 304564
rect 676214 304552 676220 304564
rect 674616 304524 676220 304552
rect 674616 304512 674622 304524
rect 676214 304512 676220 304524
rect 676272 304512 676278 304564
rect 673178 303696 673184 303748
rect 673236 303736 673242 303748
rect 676214 303736 676220 303748
rect 673236 303708 676220 303736
rect 673236 303696 673242 303708
rect 676214 303696 676220 303708
rect 676272 303696 676278 303748
rect 673086 303628 673092 303680
rect 673144 303668 673150 303680
rect 676122 303668 676128 303680
rect 673144 303640 676128 303668
rect 673144 303628 673150 303640
rect 676122 303628 676128 303640
rect 676180 303628 676186 303680
rect 674282 302200 674288 302252
rect 674340 302240 674346 302252
rect 683114 302240 683120 302252
rect 674340 302212 683120 302240
rect 674340 302200 674346 302212
rect 683114 302200 683120 302212
rect 683172 302200 683178 302252
rect 42058 300908 42064 300960
rect 42116 300948 42122 300960
rect 47670 300948 47676 300960
rect 42116 300920 47676 300948
rect 42116 300908 42122 300920
rect 47670 300908 47676 300920
rect 47728 300908 47734 300960
rect 43622 298120 43628 298172
rect 43680 298160 43686 298172
rect 62114 298160 62120 298172
rect 43680 298132 62120 298160
rect 43680 298120 43686 298132
rect 62114 298120 62120 298132
rect 62172 298120 62178 298172
rect 675110 298120 675116 298172
rect 675168 298160 675174 298172
rect 676398 298160 676404 298172
rect 675168 298132 676404 298160
rect 675168 298120 675174 298132
rect 676398 298120 676404 298132
rect 676456 298120 676462 298172
rect 675754 298052 675760 298104
rect 675812 298092 675818 298104
rect 679710 298092 679716 298104
rect 675812 298064 679716 298092
rect 675812 298052 675818 298064
rect 679710 298052 679716 298064
rect 679768 298052 679774 298104
rect 675202 297984 675208 298036
rect 675260 298024 675266 298036
rect 676858 298024 676864 298036
rect 675260 297996 676864 298024
rect 675260 297984 675266 297996
rect 676858 297984 676864 297996
rect 676916 297984 676922 298036
rect 675754 296148 675760 296200
rect 675812 296148 675818 296200
rect 675772 295996 675800 296148
rect 675754 295944 675760 295996
rect 675812 295944 675818 295996
rect 675202 295196 675208 295248
rect 675260 295236 675266 295248
rect 675386 295236 675392 295248
rect 675260 295208 675392 295236
rect 675260 295196 675266 295208
rect 675386 295196 675392 295208
rect 675444 295196 675450 295248
rect 675110 294040 675116 294092
rect 675168 294040 675174 294092
rect 675018 293972 675024 294024
rect 675076 294012 675082 294024
rect 675128 294012 675156 294040
rect 675076 293984 675156 294012
rect 675076 293972 675082 293984
rect 675018 291728 675024 291780
rect 675076 291768 675082 291780
rect 675386 291768 675392 291780
rect 675076 291740 675392 291768
rect 675076 291728 675082 291740
rect 675386 291728 675392 291740
rect 675444 291728 675450 291780
rect 674558 291048 674564 291100
rect 674616 291088 674622 291100
rect 675386 291088 675392 291100
rect 674616 291060 675392 291088
rect 674616 291048 674622 291060
rect 675386 291048 675392 291060
rect 675444 291048 675450 291100
rect 673086 287920 673092 287972
rect 673144 287960 673150 287972
rect 675386 287960 675392 287972
rect 673144 287932 675392 287960
rect 673144 287920 673150 287932
rect 675386 287920 675392 287932
rect 675444 287920 675450 287972
rect 673178 286560 673184 286612
rect 673236 286600 673242 286612
rect 675386 286600 675392 286612
rect 673236 286572 675392 286600
rect 673236 286560 673242 286572
rect 675386 286560 675392 286572
rect 675444 286560 675450 286612
rect 46290 284316 46296 284368
rect 46348 284356 46354 284368
rect 62114 284356 62120 284368
rect 46348 284328 62120 284356
rect 46348 284316 46354 284328
rect 62114 284316 62120 284328
rect 62172 284316 62178 284368
rect 651558 284316 651564 284368
rect 651616 284356 651622 284368
rect 671522 284356 671528 284368
rect 651616 284328 671528 284356
rect 651616 284316 651622 284328
rect 671522 284316 671528 284328
rect 671580 284316 671586 284368
rect 42150 283568 42156 283620
rect 42208 283608 42214 283620
rect 42426 283608 42432 283620
rect 42208 283580 42432 283608
rect 42208 283568 42214 283580
rect 42426 283568 42432 283580
rect 42484 283568 42490 283620
rect 42150 281052 42156 281104
rect 42208 281092 42214 281104
rect 43530 281092 43536 281104
rect 42208 281064 43536 281092
rect 42208 281052 42214 281064
rect 43530 281052 43536 281064
rect 43588 281052 43594 281104
rect 42150 279828 42156 279880
rect 42208 279868 42214 279880
rect 42978 279868 42984 279880
rect 42208 279840 42984 279868
rect 42208 279828 42214 279840
rect 42978 279828 42984 279840
rect 43036 279828 43042 279880
rect 42058 278604 42064 278656
rect 42116 278644 42122 278656
rect 44174 278644 44180 278656
rect 42116 278616 44180 278644
rect 42116 278604 42122 278616
rect 44174 278604 44180 278616
rect 44232 278604 44238 278656
rect 43438 278128 43444 278180
rect 43496 278168 43502 278180
rect 647326 278168 647332 278180
rect 43496 278140 647332 278168
rect 43496 278128 43502 278140
rect 647326 278128 647332 278140
rect 647384 278128 647390 278180
rect 53190 278060 53196 278112
rect 53248 278100 53254 278112
rect 659654 278100 659660 278112
rect 53248 278072 659660 278100
rect 53248 278060 53254 278072
rect 659654 278060 659660 278072
rect 659712 278060 659718 278112
rect 44818 277992 44824 278044
rect 44876 278032 44882 278044
rect 658274 278032 658280 278044
rect 44876 278004 658280 278032
rect 44876 277992 44882 278004
rect 658274 277992 658280 278004
rect 658332 277992 658338 278044
rect 339402 277584 339408 277636
rect 339460 277624 339466 277636
rect 454770 277624 454776 277636
rect 339460 277596 454776 277624
rect 339460 277584 339466 277596
rect 454770 277584 454776 277596
rect 454828 277584 454834 277636
rect 389082 277516 389088 277568
rect 389140 277556 389146 277568
rect 587158 277556 587164 277568
rect 389140 277528 587164 277556
rect 389140 277516 389146 277528
rect 587158 277516 587164 277528
rect 587216 277516 587222 277568
rect 394418 277448 394424 277500
rect 394476 277488 394482 277500
rect 601418 277488 601424 277500
rect 394476 277460 601424 277488
rect 394476 277448 394482 277460
rect 601418 277448 601424 277460
rect 601476 277448 601482 277500
rect 398374 277380 398380 277432
rect 398432 277420 398438 277432
rect 611998 277420 612004 277432
rect 398432 277392 612004 277420
rect 398432 277380 398438 277392
rect 611998 277380 612004 277392
rect 612056 277380 612062 277432
rect 351822 277312 351828 277364
rect 351880 277352 351886 277364
rect 489086 277352 489092 277364
rect 351880 277324 489092 277352
rect 351880 277312 351886 277324
rect 489086 277312 489092 277324
rect 489144 277312 489150 277364
rect 354582 277244 354588 277296
rect 354640 277284 354646 277296
rect 496170 277284 496176 277296
rect 354640 277256 496176 277284
rect 354640 277244 354646 277256
rect 496170 277244 496176 277256
rect 496228 277244 496234 277296
rect 357342 277176 357348 277228
rect 357400 277216 357406 277228
rect 503254 277216 503260 277228
rect 357400 277188 503260 277216
rect 357400 277176 357406 277188
rect 503254 277176 503260 277188
rect 503312 277176 503318 277228
rect 42150 277108 42156 277160
rect 42208 277148 42214 277160
rect 42886 277148 42892 277160
rect 42208 277120 42892 277148
rect 42208 277108 42214 277120
rect 42886 277108 42892 277120
rect 42944 277108 42950 277160
rect 360102 277108 360108 277160
rect 360160 277148 360166 277160
rect 510338 277148 510344 277160
rect 360160 277120 510344 277148
rect 360160 277108 360166 277120
rect 510338 277108 510344 277120
rect 510396 277108 510402 277160
rect 384942 277040 384948 277092
rect 385000 277080 385006 277092
rect 574186 277080 574192 277092
rect 385000 277052 574192 277080
rect 385000 277040 385006 277052
rect 574186 277040 574192 277052
rect 574244 277040 574250 277092
rect 381998 276972 382004 277024
rect 382056 277012 382062 277024
rect 567102 277012 567108 277024
rect 382056 276984 567108 277012
rect 382056 276972 382062 276984
rect 567102 276972 567108 276984
rect 567160 276972 567166 277024
rect 384574 276904 384580 276956
rect 384632 276944 384638 276956
rect 575382 276944 575388 276956
rect 384632 276916 575388 276944
rect 384632 276904 384638 276916
rect 575382 276904 575388 276916
rect 575440 276904 575446 276956
rect 387242 276836 387248 276888
rect 387300 276876 387306 276888
rect 582466 276876 582472 276888
rect 387300 276848 582472 276876
rect 387300 276836 387306 276848
rect 582466 276836 582472 276848
rect 582524 276836 582530 276888
rect 391750 276768 391756 276820
rect 391808 276808 391814 276820
rect 593138 276808 593144 276820
rect 391808 276780 593144 276808
rect 391808 276768 391814 276780
rect 593138 276768 593144 276780
rect 593196 276768 593202 276820
rect 394602 276700 394608 276752
rect 394660 276740 394666 276752
rect 600222 276740 600228 276752
rect 394660 276712 600228 276740
rect 394660 276700 394666 276712
rect 600222 276700 600228 276712
rect 600280 276700 600286 276752
rect 408402 276632 408408 276684
rect 408460 276672 408466 276684
rect 638034 276672 638040 276684
rect 408460 276644 638040 276672
rect 408460 276632 408466 276644
rect 638034 276632 638040 276644
rect 638092 276632 638098 276684
rect 335262 276564 335268 276616
rect 335320 276604 335326 276616
rect 444190 276604 444196 276616
rect 335320 276576 444196 276604
rect 335320 276564 335326 276576
rect 444190 276564 444196 276576
rect 444248 276564 444254 276616
rect 333882 276496 333888 276548
rect 333940 276536 333946 276548
rect 439406 276536 439412 276548
rect 333940 276508 439412 276536
rect 333940 276496 333946 276508
rect 439406 276496 439412 276508
rect 439464 276496 439470 276548
rect 330754 276428 330760 276480
rect 330812 276468 330818 276480
rect 432322 276468 432328 276480
rect 330812 276440 432328 276468
rect 330812 276428 330818 276440
rect 432322 276428 432328 276440
rect 432380 276428 432386 276480
rect 329742 276360 329748 276412
rect 329800 276400 329806 276412
rect 428826 276400 428832 276412
rect 329800 276372 428832 276400
rect 329800 276360 329806 276372
rect 428826 276360 428832 276372
rect 428884 276360 428890 276412
rect 326982 276292 326988 276344
rect 327040 276332 327046 276344
rect 421650 276332 421656 276344
rect 327040 276304 421656 276332
rect 327040 276292 327046 276304
rect 421650 276292 421656 276304
rect 421708 276292 421714 276344
rect 405642 276020 405648 276072
rect 405700 276060 405706 276072
rect 405700 276032 474688 276060
rect 405700 276020 405706 276032
rect 142706 275952 142712 276004
rect 142764 275992 142770 276004
rect 181162 275992 181168 276004
rect 142764 275964 181168 275992
rect 142764 275952 142770 275964
rect 181162 275952 181168 275964
rect 181220 275952 181226 276004
rect 185210 275952 185216 276004
rect 185268 275992 185274 276004
rect 217318 275992 217324 276004
rect 185268 275964 217324 275992
rect 185268 275952 185274 275964
rect 217318 275952 217324 275964
rect 217376 275952 217382 276004
rect 346118 275952 346124 276004
rect 346176 275992 346182 276004
rect 473722 275992 473728 276004
rect 346176 275964 473728 275992
rect 346176 275952 346182 275964
rect 473722 275952 473728 275964
rect 473780 275952 473786 276004
rect 474660 275992 474688 276032
rect 629754 275992 629760 276004
rect 474660 275964 629760 275992
rect 629754 275952 629760 275964
rect 629812 275952 629818 276004
rect 153286 275884 153292 275936
rect 153344 275924 153350 275936
rect 204898 275924 204904 275936
rect 153344 275896 204904 275924
rect 153344 275884 153350 275896
rect 204898 275884 204904 275896
rect 204956 275884 204962 275936
rect 348786 275884 348792 275936
rect 348844 275924 348850 275936
rect 480806 275924 480812 275936
rect 348844 275896 480812 275924
rect 348844 275884 348850 275896
rect 480806 275884 480812 275896
rect 480864 275884 480870 275936
rect 481174 275884 481180 275936
rect 481232 275924 481238 275936
rect 581270 275924 581276 275936
rect 481232 275896 581276 275924
rect 481232 275884 481238 275896
rect 581270 275884 581276 275896
rect 581328 275884 581334 275936
rect 167546 275816 167552 275868
rect 167604 275856 167610 275868
rect 223206 275856 223212 275868
rect 167604 275828 223212 275856
rect 167604 275816 167610 275828
rect 223206 275816 223212 275828
rect 223264 275816 223270 275868
rect 343358 275816 343364 275868
rect 343416 275856 343422 275868
rect 466638 275856 466644 275868
rect 343416 275828 466644 275856
rect 343416 275816 343422 275828
rect 466638 275816 466644 275828
rect 466696 275816 466702 275868
rect 466730 275816 466736 275868
rect 466788 275856 466794 275868
rect 603718 275856 603724 275868
rect 466788 275828 603724 275856
rect 466788 275816 466794 275828
rect 603718 275816 603724 275828
rect 603776 275816 603782 275868
rect 160462 275748 160468 275800
rect 160520 275788 160526 275800
rect 220630 275788 220636 275800
rect 160520 275760 220636 275788
rect 160520 275748 160526 275760
rect 220630 275748 220636 275760
rect 220688 275748 220694 275800
rect 250254 275748 250260 275800
rect 250312 275788 250318 275800
rect 251174 275788 251180 275800
rect 250312 275760 251180 275788
rect 250312 275748 250318 275760
rect 251174 275748 251180 275760
rect 251232 275748 251238 275800
rect 258534 275748 258540 275800
rect 258592 275788 258598 275800
rect 264606 275788 264612 275800
rect 258592 275760 264612 275788
rect 258592 275748 258598 275760
rect 264606 275748 264612 275760
rect 264664 275748 264670 275800
rect 354490 275748 354496 275800
rect 354548 275788 354554 275800
rect 494974 275788 494980 275800
rect 354548 275760 494980 275788
rect 354548 275748 354554 275760
rect 494974 275748 494980 275760
rect 495032 275748 495038 275800
rect 495066 275748 495072 275800
rect 495124 275788 495130 275800
rect 588354 275788 588360 275800
rect 495124 275760 588360 275788
rect 495124 275748 495130 275760
rect 588354 275748 588360 275760
rect 588412 275748 588418 275800
rect 107194 275680 107200 275732
rect 107252 275720 107258 275732
rect 208394 275720 208400 275732
rect 107252 275692 208400 275720
rect 107252 275680 107258 275692
rect 208394 275680 208400 275692
rect 208452 275680 208458 275732
rect 213638 275680 213644 275732
rect 213696 275720 213702 275732
rect 223022 275720 223028 275732
rect 213696 275692 223028 275720
rect 213696 275680 213702 275692
rect 223022 275680 223028 275692
rect 223080 275680 223086 275732
rect 251450 275680 251456 275732
rect 251508 275720 251514 275732
rect 252370 275720 252376 275732
rect 251508 275692 252376 275720
rect 251508 275680 251514 275692
rect 252370 275680 252376 275692
rect 252428 275680 252434 275732
rect 357250 275680 357256 275732
rect 357308 275720 357314 275732
rect 502058 275720 502064 275732
rect 357308 275692 502064 275720
rect 357308 275680 357314 275692
rect 502058 275680 502064 275692
rect 502116 275680 502122 275732
rect 507854 275680 507860 275732
rect 507912 275720 507918 275732
rect 507912 275692 518894 275720
rect 507912 275680 507918 275692
rect 100110 275612 100116 275664
rect 100168 275652 100174 275664
rect 205818 275652 205824 275664
rect 100168 275624 205824 275652
rect 100168 275612 100174 275624
rect 205818 275612 205824 275624
rect 205876 275612 205882 275664
rect 212442 275612 212448 275664
rect 212500 275652 212506 275664
rect 224954 275652 224960 275664
rect 212500 275624 224960 275652
rect 212500 275612 212506 275624
rect 224954 275612 224960 275624
rect 225012 275612 225018 275664
rect 360010 275612 360016 275664
rect 360068 275652 360074 275664
rect 509142 275652 509148 275664
rect 360068 275624 509148 275652
rect 360068 275612 360074 275624
rect 509142 275612 509148 275624
rect 509200 275612 509206 275664
rect 518866 275652 518894 275692
rect 577682 275680 577688 275732
rect 577740 275720 577746 275732
rect 599026 275720 599032 275732
rect 577740 275692 599032 275720
rect 577740 275680 577746 275692
rect 599026 275680 599032 275692
rect 599084 275680 599090 275732
rect 591942 275652 591948 275664
rect 518866 275624 591948 275652
rect 591942 275612 591948 275624
rect 592000 275612 592006 275664
rect 592034 275612 592040 275664
rect 592092 275652 592098 275664
rect 614390 275652 614396 275664
rect 592092 275624 614396 275652
rect 592092 275612 592098 275624
rect 614390 275612 614396 275624
rect 614448 275612 614454 275664
rect 93026 275544 93032 275596
rect 93084 275584 93090 275596
rect 201402 275584 201408 275596
rect 93084 275556 201408 275584
rect 93084 275544 93090 275556
rect 201402 275544 201408 275556
rect 201460 275544 201466 275596
rect 210050 275544 210056 275596
rect 210108 275584 210114 275596
rect 231762 275584 231768 275596
rect 210108 275556 231768 275584
rect 210108 275544 210114 275556
rect 231762 275544 231768 275556
rect 231820 275544 231826 275596
rect 234890 275544 234896 275596
rect 234948 275584 234954 275596
rect 245654 275584 245660 275596
rect 234948 275556 245660 275584
rect 234948 275544 234954 275556
rect 245654 275544 245660 275556
rect 245712 275544 245718 275596
rect 362310 275544 362316 275596
rect 362368 275584 362374 275596
rect 516226 275584 516232 275596
rect 362368 275556 516232 275584
rect 362368 275544 362374 275556
rect 516226 275544 516232 275556
rect 516284 275544 516290 275596
rect 581638 275544 581644 275596
rect 581696 275584 581702 275596
rect 607306 275584 607312 275596
rect 581696 275556 607312 275584
rect 581696 275544 581702 275556
rect 607306 275544 607312 275556
rect 607364 275544 607370 275596
rect 90634 275476 90640 275528
rect 90692 275516 90698 275528
rect 201678 275516 201684 275528
rect 90692 275488 201684 275516
rect 90692 275476 90698 275488
rect 201678 275476 201684 275488
rect 201736 275476 201742 275528
rect 223114 275476 223120 275528
rect 223172 275516 223178 275528
rect 244274 275516 244280 275528
rect 223172 275488 244280 275516
rect 223172 275476 223178 275488
rect 244274 275476 244280 275488
rect 244332 275476 244338 275528
rect 365438 275476 365444 275528
rect 365496 275516 365502 275528
rect 523402 275516 523408 275528
rect 365496 275488 523408 275516
rect 365496 275476 365502 275488
rect 523402 275476 523408 275488
rect 523460 275476 523466 275528
rect 523586 275476 523592 275528
rect 523644 275516 523650 275528
rect 594702 275516 594708 275528
rect 523644 275488 594708 275516
rect 523644 275476 523650 275488
rect 594702 275476 594708 275488
rect 594760 275476 594766 275528
rect 594794 275476 594800 275528
rect 594852 275516 594858 275528
rect 617978 275516 617984 275528
rect 594852 275488 617984 275516
rect 594852 275476 594858 275488
rect 617978 275476 617984 275488
rect 618036 275476 618042 275528
rect 81250 275408 81256 275460
rect 81308 275448 81314 275460
rect 197814 275448 197820 275460
rect 81308 275420 197820 275448
rect 81308 275408 81314 275420
rect 197814 275408 197820 275420
rect 197872 275408 197878 275460
rect 215938 275408 215944 275460
rect 215996 275448 216002 275460
rect 240042 275448 240048 275460
rect 215996 275420 240048 275448
rect 215996 275408 216002 275420
rect 240042 275408 240048 275420
rect 240100 275408 240106 275460
rect 333790 275408 333796 275460
rect 333848 275448 333854 275460
rect 438210 275448 438216 275460
rect 333848 275420 438216 275448
rect 333848 275408 333854 275420
rect 438210 275408 438216 275420
rect 438268 275408 438274 275460
rect 438854 275408 438860 275460
rect 438912 275448 438918 275460
rect 622670 275448 622676 275460
rect 438912 275420 622676 275448
rect 438912 275408 438918 275420
rect 622670 275408 622676 275420
rect 622728 275408 622734 275460
rect 66990 275340 66996 275392
rect 67048 275380 67054 275392
rect 185578 275380 185584 275392
rect 67048 275352 185584 275380
rect 67048 275340 67054 275352
rect 185578 275340 185584 275352
rect 185636 275340 185642 275392
rect 188798 275340 188804 275392
rect 188856 275380 188862 275392
rect 215846 275380 215852 275392
rect 188856 275352 215852 275380
rect 188856 275340 188862 275352
rect 215846 275340 215852 275352
rect 215904 275340 215910 275392
rect 220722 275340 220728 275392
rect 220780 275380 220786 275392
rect 243354 275380 243360 275392
rect 220780 275352 243360 275380
rect 220780 275340 220786 275352
rect 243354 275340 243360 275352
rect 243412 275340 243418 275392
rect 244366 275340 244372 275392
rect 244424 275380 244430 275392
rect 259362 275380 259368 275392
rect 244424 275352 259368 275380
rect 244424 275340 244430 275352
rect 259362 275340 259368 275352
rect 259420 275340 259426 275392
rect 398834 275340 398840 275392
rect 398892 275380 398898 275392
rect 413370 275380 413376 275392
rect 398892 275352 413376 275380
rect 398892 275340 398898 275352
rect 413370 275340 413376 275352
rect 413428 275340 413434 275392
rect 419534 275340 419540 275392
rect 419592 275380 419598 275392
rect 643922 275380 643928 275392
rect 419592 275352 643928 275380
rect 419592 275340 419598 275352
rect 643922 275340 643928 275352
rect 643980 275340 643986 275392
rect 71774 275272 71780 275324
rect 71832 275312 71838 275324
rect 193858 275312 193864 275324
rect 71832 275284 193864 275312
rect 71832 275272 71838 275284
rect 193858 275272 193864 275284
rect 193916 275272 193922 275324
rect 208854 275272 208860 275324
rect 208912 275312 208918 275324
rect 234614 275312 234620 275324
rect 208912 275284 234620 275312
rect 208912 275272 208918 275284
rect 234614 275272 234620 275284
rect 234672 275272 234678 275324
rect 239582 275272 239588 275324
rect 239640 275312 239646 275324
rect 252922 275312 252928 275324
rect 239640 275284 252928 275312
rect 239640 275272 239646 275284
rect 252922 275272 252928 275284
rect 252980 275272 252986 275324
rect 259730 275272 259736 275324
rect 259788 275312 259794 275324
rect 265066 275312 265072 275324
rect 259788 275284 265072 275312
rect 259788 275272 259794 275284
rect 265066 275272 265072 275284
rect 265124 275272 265130 275324
rect 389266 275272 389272 275324
rect 389324 275312 389330 275324
rect 409874 275312 409880 275324
rect 389324 275284 409880 275312
rect 389324 275272 389330 275284
rect 409874 275272 409880 275284
rect 409932 275272 409938 275324
rect 411162 275272 411168 275324
rect 411220 275312 411226 275324
rect 646314 275312 646320 275324
rect 411220 275284 646320 275312
rect 411220 275272 411226 275284
rect 646314 275272 646320 275284
rect 646372 275272 646378 275324
rect 174630 275204 174636 275256
rect 174688 275244 174694 275256
rect 207014 275244 207020 275256
rect 174688 275216 207020 275244
rect 174688 275204 174694 275216
rect 207014 275204 207020 275216
rect 207072 275204 207078 275256
rect 340598 275204 340604 275256
rect 340656 275244 340662 275256
rect 459554 275244 459560 275256
rect 340656 275216 459560 275244
rect 340656 275204 340662 275216
rect 459554 275204 459560 275216
rect 459612 275204 459618 275256
rect 459738 275204 459744 275256
rect 459796 275244 459802 275256
rect 577774 275244 577780 275256
rect 459796 275216 577780 275244
rect 459796 275204 459802 275216
rect 577774 275204 577780 275216
rect 577832 275204 577838 275256
rect 181714 275136 181720 275188
rect 181772 275176 181778 275188
rect 213178 275176 213184 275188
rect 181772 275148 213184 275176
rect 181772 275136 181778 275148
rect 213178 275136 213184 275148
rect 213236 275136 213242 275188
rect 337838 275136 337844 275188
rect 337896 275176 337902 275188
rect 452470 275176 452476 275188
rect 337896 275148 452476 275176
rect 337896 275136 337902 275148
rect 452470 275136 452476 275148
rect 452528 275136 452534 275188
rect 178126 275068 178132 275120
rect 178184 275108 178190 275120
rect 195974 275108 195980 275120
rect 178184 275080 195980 275108
rect 178184 275068 178190 275080
rect 195974 275068 195980 275080
rect 196032 275068 196038 275120
rect 375926 275068 375932 275120
rect 375984 275108 375990 275120
rect 487890 275108 487896 275120
rect 375984 275080 487896 275108
rect 375984 275068 375990 275080
rect 487890 275068 487896 275080
rect 487948 275068 487954 275120
rect 335170 275000 335176 275052
rect 335228 275040 335234 275052
rect 445294 275040 445300 275052
rect 335228 275012 445300 275040
rect 335228 275000 335234 275012
rect 445294 275000 445300 275012
rect 445352 275000 445358 275052
rect 88334 274932 88340 274984
rect 88392 274972 88398 274984
rect 90358 274972 90364 274984
rect 88392 274944 90364 274972
rect 88392 274932 88398 274944
rect 90358 274932 90364 274944
rect 90416 274932 90422 274984
rect 262122 274932 262128 274984
rect 262180 274972 262186 274984
rect 264974 274972 264980 274984
rect 262180 274944 264980 274972
rect 262180 274932 262186 274944
rect 264974 274932 264980 274944
rect 265032 274932 265038 274984
rect 330662 274932 330668 274984
rect 330720 274972 330726 274984
rect 431126 274972 431132 274984
rect 330720 274944 431132 274972
rect 330720 274932 330726 274944
rect 431126 274932 431132 274944
rect 431184 274932 431190 274984
rect 74074 274864 74080 274916
rect 74132 274904 74138 274916
rect 77202 274904 77208 274916
rect 74132 274876 77208 274904
rect 74132 274864 74138 274876
rect 77202 274864 77208 274876
rect 77260 274864 77266 274916
rect 252646 274864 252652 274916
rect 252704 274904 252710 274916
rect 252704 274876 260236 274904
rect 252704 274864 252710 274876
rect 96614 274796 96620 274848
rect 96672 274836 96678 274848
rect 100018 274836 100024 274848
rect 96672 274808 100024 274836
rect 96672 274796 96678 274808
rect 100018 274796 100024 274808
rect 100076 274796 100082 274848
rect 70578 274660 70584 274712
rect 70636 274700 70642 274712
rect 73798 274700 73804 274712
rect 70636 274672 73804 274700
rect 70636 274660 70642 274672
rect 73798 274660 73804 274672
rect 73856 274660 73862 274712
rect 103698 274660 103704 274712
rect 103756 274700 103762 274712
rect 106918 274700 106924 274712
rect 103756 274672 106924 274700
rect 103756 274660 103762 274672
rect 106918 274660 106924 274672
rect 106976 274660 106982 274712
rect 207750 274660 207756 274712
rect 207808 274700 207814 274712
rect 210602 274700 210608 274712
rect 207808 274672 210608 274700
rect 207808 274660 207814 274672
rect 210602 274660 210608 274672
rect 210660 274660 210666 274712
rect 227806 274660 227812 274712
rect 227864 274700 227870 274712
rect 229922 274700 229928 274712
rect 227864 274672 229928 274700
rect 227864 274660 227870 274672
rect 229922 274660 229928 274672
rect 229980 274660 229986 274712
rect 159266 274592 159272 274644
rect 159324 274632 159330 274644
rect 226886 274632 226892 274644
rect 159324 274604 226892 274632
rect 159324 274592 159330 274604
rect 226886 274592 226892 274604
rect 226944 274592 226950 274644
rect 260208 274632 260236 274876
rect 260926 274864 260932 274916
rect 260984 274904 260990 274916
rect 265434 274904 265440 274916
rect 260984 274876 265440 274904
rect 260984 274864 260990 274876
rect 265434 274864 265440 274876
rect 265492 274864 265498 274916
rect 403434 274864 403440 274916
rect 403492 274904 403498 274916
rect 424042 274904 424048 274916
rect 403492 274876 424048 274904
rect 403492 274864 403498 274876
rect 424042 274864 424048 274876
rect 424100 274864 424106 274916
rect 409138 274796 409144 274848
rect 409196 274836 409202 274848
rect 420546 274836 420552 274848
rect 409196 274808 420552 274836
rect 409196 274796 409202 274808
rect 420546 274796 420552 274808
rect 420604 274796 420610 274848
rect 264422 274728 264428 274780
rect 264480 274768 264486 274780
rect 266722 274768 266728 274780
rect 264480 274740 266728 274768
rect 264480 274728 264486 274740
rect 266722 274728 266728 274740
rect 266780 274728 266786 274780
rect 263226 274660 263232 274712
rect 263284 274700 263290 274712
rect 266446 274700 266452 274712
rect 263284 274672 266452 274700
rect 263284 274660 263290 274672
rect 266446 274660 266452 274672
rect 266504 274660 266510 274712
rect 266814 274660 266820 274712
rect 266872 274700 266878 274712
rect 267734 274700 267740 274712
rect 266872 274672 267740 274700
rect 266872 274660 266878 274672
rect 267734 274660 267740 274672
rect 267792 274660 267798 274712
rect 262398 274632 262404 274644
rect 260208 274604 262404 274632
rect 262398 274592 262404 274604
rect 262456 274592 262462 274644
rect 311158 274592 311164 274644
rect 311216 274632 311222 274644
rect 333054 274632 333060 274644
rect 311216 274604 333060 274632
rect 311216 274592 311222 274604
rect 333054 274592 333060 274604
rect 333112 274592 333118 274644
rect 350442 274592 350448 274644
rect 350500 274632 350506 274644
rect 483198 274632 483204 274644
rect 350500 274604 483204 274632
rect 350500 274592 350506 274604
rect 483198 274592 483204 274604
rect 483256 274592 483262 274644
rect 128538 274524 128544 274576
rect 128596 274564 128602 274576
rect 196710 274564 196716 274576
rect 128596 274536 196716 274564
rect 128596 274524 128602 274536
rect 196710 274524 196716 274536
rect 196768 274524 196774 274576
rect 199470 274524 199476 274576
rect 199528 274564 199534 274576
rect 242066 274564 242072 274576
rect 199528 274536 242072 274564
rect 199528 274524 199534 274536
rect 242066 274524 242072 274536
rect 242124 274524 242130 274576
rect 312446 274524 312452 274576
rect 312504 274564 312510 274576
rect 336550 274564 336556 274576
rect 312504 274536 336556 274564
rect 312504 274524 312510 274536
rect 336550 274524 336556 274536
rect 336608 274524 336614 274576
rect 351730 274524 351736 274576
rect 351788 274564 351794 274576
rect 486694 274564 486700 274576
rect 351788 274536 486700 274564
rect 351788 274524 351794 274536
rect 486694 274524 486700 274536
rect 486752 274524 486758 274576
rect 150986 274456 150992 274508
rect 151044 274496 151050 274508
rect 223758 274496 223764 274508
rect 151044 274468 223764 274496
rect 151044 274456 151050 274468
rect 223758 274456 223764 274468
rect 223816 274456 223822 274508
rect 320818 274456 320824 274508
rect 320876 274496 320882 274508
rect 349614 274496 349620 274508
rect 320876 274468 349620 274496
rect 320876 274456 320882 274468
rect 349614 274456 349620 274468
rect 349672 274456 349678 274508
rect 353202 274456 353208 274508
rect 353260 274496 353266 274508
rect 490282 274496 490288 274508
rect 353260 274468 490288 274496
rect 353260 274456 353266 274468
rect 490282 274456 490288 274468
rect 490340 274456 490346 274508
rect 493318 274456 493324 274508
rect 493376 274496 493382 274508
rect 505646 274496 505652 274508
rect 493376 274468 505652 274496
rect 493376 274456 493382 274468
rect 505646 274456 505652 274468
rect 505704 274456 505710 274508
rect 148594 274388 148600 274440
rect 148652 274428 148658 274440
rect 222746 274428 222752 274440
rect 148652 274400 222752 274428
rect 148652 274388 148658 274400
rect 222746 274388 222752 274400
rect 222804 274388 222810 274440
rect 295978 274388 295984 274440
rect 296036 274428 296042 274440
rect 329466 274428 329472 274440
rect 296036 274400 329472 274428
rect 296036 274388 296042 274400
rect 329466 274388 329472 274400
rect 329524 274388 329530 274440
rect 354398 274388 354404 274440
rect 354456 274428 354462 274440
rect 493778 274428 493784 274440
rect 354456 274400 493784 274428
rect 354456 274388 354462 274400
rect 493778 274388 493784 274400
rect 493836 274388 493842 274440
rect 121362 274320 121368 274372
rect 121420 274360 121426 274372
rect 196618 274360 196624 274372
rect 121420 274332 196624 274360
rect 121420 274320 121426 274332
rect 196618 274320 196624 274332
rect 196676 274320 196682 274372
rect 198274 274320 198280 274372
rect 198332 274360 198338 274372
rect 241606 274360 241612 274372
rect 198332 274332 241612 274360
rect 198332 274320 198338 274332
rect 241606 274320 241612 274332
rect 241664 274320 241670 274372
rect 291010 274320 291016 274372
rect 291068 274360 291074 274372
rect 324774 274360 324780 274372
rect 291068 274332 324780 274360
rect 291068 274320 291074 274332
rect 324774 274320 324780 274332
rect 324832 274320 324838 274372
rect 355962 274320 355968 274372
rect 356020 274360 356026 274372
rect 497366 274360 497372 274372
rect 356020 274332 497372 274360
rect 356020 274320 356026 274332
rect 497366 274320 497372 274332
rect 497424 274320 497430 274372
rect 42150 274252 42156 274304
rect 42208 274292 42214 274304
rect 44542 274292 44548 274304
rect 42208 274264 44548 274292
rect 42208 274252 42214 274264
rect 44542 274252 44548 274264
rect 44600 274252 44606 274304
rect 137922 274252 137928 274304
rect 137980 274292 137986 274304
rect 219618 274292 219624 274304
rect 137980 274264 219624 274292
rect 137980 274252 137986 274264
rect 219618 274252 219624 274264
rect 219676 274252 219682 274304
rect 289078 274252 289084 274304
rect 289136 274292 289142 274304
rect 318794 274292 318800 274304
rect 289136 274264 318800 274292
rect 289136 274252 289142 274264
rect 318794 274252 318800 274264
rect 318852 274252 318858 274304
rect 322198 274252 322204 274304
rect 322256 274292 322262 274304
rect 356698 274292 356704 274304
rect 322256 274264 356704 274292
rect 322256 274252 322262 274264
rect 356698 274252 356704 274264
rect 356756 274252 356762 274304
rect 357158 274252 357164 274304
rect 357216 274292 357222 274304
rect 500862 274292 500868 274304
rect 357216 274264 500868 274292
rect 357216 274252 357222 274264
rect 500862 274252 500868 274264
rect 500920 274252 500926 274304
rect 123754 274184 123760 274236
rect 123812 274224 123818 274236
rect 214098 274224 214104 274236
rect 123812 274196 214104 274224
rect 123812 274184 123818 274196
rect 214098 274184 214104 274196
rect 214156 274184 214162 274236
rect 291102 274184 291108 274236
rect 291160 274224 291166 274236
rect 325970 274224 325976 274236
rect 291160 274196 325976 274224
rect 291160 274184 291166 274196
rect 325970 274184 325976 274196
rect 326028 274184 326034 274236
rect 362770 274184 362776 274236
rect 362828 274224 362834 274236
rect 518618 274224 518624 274236
rect 362828 274196 518624 274224
rect 362828 274184 362834 274196
rect 518618 274184 518624 274196
rect 518676 274184 518682 274236
rect 523678 274184 523684 274236
rect 523736 274224 523742 274236
rect 533982 274224 533988 274236
rect 523736 274196 533988 274224
rect 523736 274184 523742 274196
rect 533982 274184 533988 274196
rect 534040 274184 534046 274236
rect 113174 274116 113180 274168
rect 113232 274156 113238 274168
rect 209958 274156 209964 274168
rect 113232 274128 209964 274156
rect 113232 274116 113238 274128
rect 209958 274116 209964 274128
rect 210016 274116 210022 274168
rect 243170 274116 243176 274168
rect 243228 274156 243234 274168
rect 258626 274156 258632 274168
rect 243228 274128 258632 274156
rect 243228 274116 243234 274128
rect 258626 274116 258632 274128
rect 258684 274116 258690 274168
rect 273162 274116 273168 274168
rect 273220 274156 273226 274168
rect 279786 274156 279792 274168
rect 273220 274128 279792 274156
rect 273220 274116 273226 274128
rect 279786 274116 279792 274128
rect 279844 274116 279850 274168
rect 292482 274116 292488 274168
rect 292540 274156 292546 274168
rect 328270 274156 328276 274168
rect 292540 274128 328276 274156
rect 292540 274116 292546 274128
rect 328270 274116 328276 274128
rect 328328 274116 328334 274168
rect 348970 274116 348976 274168
rect 349028 274156 349034 274168
rect 479334 274156 479340 274168
rect 349028 274128 479340 274156
rect 349028 274116 349034 274128
rect 479334 274116 479340 274128
rect 479392 274116 479398 274168
rect 479518 274116 479524 274168
rect 479576 274156 479582 274168
rect 640426 274156 640432 274168
rect 479576 274128 640432 274156
rect 479576 274116 479582 274128
rect 640426 274116 640432 274128
rect 640484 274116 640490 274168
rect 111978 274048 111984 274100
rect 112036 274088 112042 274100
rect 208946 274088 208952 274100
rect 112036 274060 208952 274088
rect 112036 274048 112042 274060
rect 208946 274048 208952 274060
rect 209004 274048 209010 274100
rect 231394 274048 231400 274100
rect 231452 274088 231458 274100
rect 254302 274088 254308 274100
rect 231452 274060 254308 274088
rect 231452 274048 231458 274060
rect 254302 274048 254308 274060
rect 254360 274048 254366 274100
rect 296438 274048 296444 274100
rect 296496 274088 296502 274100
rect 342438 274088 342444 274100
rect 296496 274060 342444 274088
rect 296496 274048 296502 274060
rect 342438 274048 342444 274060
rect 342496 274048 342502 274100
rect 371050 274048 371056 274100
rect 371108 274088 371114 274100
rect 539870 274088 539876 274100
rect 371108 274060 539876 274088
rect 371108 274048 371114 274060
rect 539870 274048 539876 274060
rect 539928 274048 539934 274100
rect 97718 273980 97724 274032
rect 97776 274020 97782 274032
rect 203610 274020 203616 274032
rect 97776 273992 203616 274020
rect 97776 273980 97782 273992
rect 203610 273980 203616 273992
rect 203668 273980 203674 274032
rect 223022 273980 223028 274032
rect 223080 274020 223086 274032
rect 247218 274020 247224 274032
rect 223080 273992 247224 274020
rect 223080 273980 223086 273992
rect 247218 273980 247224 273992
rect 247276 273980 247282 274032
rect 277302 273980 277308 274032
rect 277360 274020 277366 274032
rect 289262 274020 289268 274032
rect 277360 273992 289268 274020
rect 277360 273980 277366 273992
rect 289262 273980 289268 273992
rect 289320 273980 289326 274032
rect 300762 273980 300768 274032
rect 300820 274020 300826 274032
rect 353110 274020 353116 274032
rect 300820 273992 353116 274020
rect 300820 273980 300826 273992
rect 353110 273980 353116 273992
rect 353168 273980 353174 274032
rect 375650 273980 375656 274032
rect 375708 274020 375714 274032
rect 551738 274020 551744 274032
rect 375708 273992 551744 274020
rect 375708 273980 375714 273992
rect 551738 273980 551744 273992
rect 551796 273980 551802 274032
rect 89530 273912 89536 273964
rect 89588 273952 89594 273964
rect 200482 273952 200488 273964
rect 89588 273924 200488 273952
rect 89588 273912 89594 273924
rect 200482 273912 200488 273924
rect 200540 273912 200546 273964
rect 205358 273912 205364 273964
rect 205416 273952 205422 273964
rect 244550 273952 244556 273964
rect 205416 273924 244556 273952
rect 205416 273912 205422 273924
rect 244550 273912 244556 273924
rect 244608 273912 244614 273964
rect 251174 273912 251180 273964
rect 251232 273952 251238 273964
rect 261478 273952 261484 273964
rect 251232 273924 261484 273952
rect 251232 273912 251238 273924
rect 261478 273912 261484 273924
rect 261536 273912 261542 273964
rect 287698 273912 287704 273964
rect 287756 273952 287762 273964
rect 304626 273952 304632 273964
rect 287756 273924 304632 273952
rect 287756 273912 287762 273924
rect 304626 273912 304632 273924
rect 304684 273912 304690 273964
rect 304718 273912 304724 273964
rect 304776 273952 304782 273964
rect 363782 273952 363788 273964
rect 304776 273924 363788 273952
rect 304776 273912 304782 273924
rect 363782 273912 363788 273924
rect 363840 273912 363846 273964
rect 379422 273912 379428 273964
rect 379480 273952 379486 273964
rect 562410 273952 562416 273964
rect 379480 273924 562416 273952
rect 379480 273912 379486 273924
rect 562410 273912 562416 273924
rect 562468 273912 562474 273964
rect 172238 273844 172244 273896
rect 172296 273884 172302 273896
rect 232038 273884 232044 273896
rect 172296 273856 232044 273884
rect 172296 273844 172302 273856
rect 232038 273844 232044 273856
rect 232096 273844 232102 273896
rect 244274 273844 244280 273896
rect 244332 273884 244338 273896
rect 251358 273884 251364 273896
rect 244332 273856 251364 273884
rect 244332 273844 244338 273856
rect 251358 273844 251364 273856
rect 251416 273844 251422 273896
rect 304258 273844 304264 273896
rect 304316 273884 304322 273896
rect 323578 273884 323584 273896
rect 304316 273856 323584 273884
rect 304316 273844 304322 273856
rect 323578 273844 323584 273856
rect 323636 273844 323642 273896
rect 347682 273844 347688 273896
rect 347740 273884 347746 273896
rect 476114 273884 476120 273896
rect 347740 273856 476120 273884
rect 347740 273844 347746 273856
rect 476114 273844 476120 273856
rect 476172 273844 476178 273896
rect 169846 273776 169852 273828
rect 169904 273816 169910 273828
rect 231026 273816 231032 273828
rect 169904 273788 231032 273816
rect 169904 273776 169910 273788
rect 231026 273776 231032 273788
rect 231084 273776 231090 273828
rect 319438 273776 319444 273828
rect 319496 273816 319502 273828
rect 338942 273816 338948 273828
rect 319496 273788 338948 273816
rect 319496 273776 319502 273788
rect 338942 273776 338948 273788
rect 339000 273776 339006 273828
rect 346210 273776 346216 273828
rect 346268 273816 346274 273828
rect 472526 273816 472532 273828
rect 346268 273788 472532 273816
rect 346268 273776 346274 273788
rect 472526 273776 472532 273788
rect 472584 273776 472590 273828
rect 194686 273708 194692 273760
rect 194744 273748 194750 273760
rect 240134 273748 240140 273760
rect 194744 273720 240140 273748
rect 194744 273708 194750 273720
rect 240134 273708 240140 273720
rect 240192 273708 240198 273760
rect 316678 273708 316684 273760
rect 316736 273748 316742 273760
rect 331858 273748 331864 273760
rect 316736 273720 331864 273748
rect 316736 273708 316742 273720
rect 331858 273708 331864 273720
rect 331916 273708 331922 273760
rect 344554 273708 344560 273760
rect 344612 273748 344618 273760
rect 468938 273748 468944 273760
rect 344612 273720 468944 273748
rect 344612 273708 344618 273720
rect 468938 273708 468944 273720
rect 468996 273708 469002 273760
rect 197078 273640 197084 273692
rect 197136 273680 197142 273692
rect 238018 273680 238024 273692
rect 197136 273652 238024 273680
rect 197136 273640 197142 273652
rect 238018 273640 238024 273652
rect 238076 273640 238082 273692
rect 309778 273640 309784 273692
rect 309836 273680 309842 273692
rect 322382 273680 322388 273692
rect 309836 273652 322388 273680
rect 309836 273640 309842 273652
rect 322382 273640 322388 273652
rect 322440 273640 322446 273692
rect 343450 273640 343456 273692
rect 343508 273680 343514 273692
rect 465442 273680 465448 273692
rect 343508 273652 465448 273680
rect 343508 273640 343514 273652
rect 465442 273640 465448 273652
rect 465500 273640 465506 273692
rect 341886 273572 341892 273624
rect 341944 273612 341950 273624
rect 461854 273612 461860 273624
rect 341944 273584 461860 273612
rect 341944 273572 341950 273584
rect 461854 273572 461860 273584
rect 461912 273572 461918 273624
rect 185578 273504 185584 273556
rect 185636 273544 185642 273556
rect 192478 273544 192484 273556
rect 185636 273516 192484 273544
rect 185636 273504 185642 273516
rect 192478 273504 192484 273516
rect 192536 273504 192542 273556
rect 340690 273504 340696 273556
rect 340748 273544 340754 273556
rect 458358 273544 458364 273556
rect 340748 273516 458364 273544
rect 340748 273504 340754 273516
rect 458358 273504 458364 273516
rect 458416 273504 458422 273556
rect 324958 273436 324964 273488
rect 325016 273476 325022 273488
rect 402790 273476 402796 273488
rect 325016 273448 402796 273476
rect 325016 273436 325022 273448
rect 402790 273436 402796 273448
rect 402848 273436 402854 273488
rect 402882 273436 402888 273488
rect 402940 273476 402946 273488
rect 438854 273476 438860 273488
rect 402940 273448 438860 273476
rect 402940 273436 402946 273448
rect 438854 273436 438860 273448
rect 438912 273436 438918 273488
rect 42058 273300 42064 273352
rect 42116 273340 42122 273352
rect 44450 273340 44456 273352
rect 42116 273312 44456 273340
rect 42116 273300 42122 273312
rect 44450 273300 44456 273312
rect 44508 273300 44514 273352
rect 279418 273232 279424 273284
rect 279476 273272 279482 273284
rect 285766 273272 285772 273284
rect 279476 273244 285772 273272
rect 279476 273232 279482 273244
rect 285766 273232 285772 273244
rect 285824 273232 285830 273284
rect 307018 273232 307024 273284
rect 307076 273272 307082 273284
rect 315298 273272 315304 273284
rect 307076 273244 315304 273272
rect 307076 273232 307082 273244
rect 315298 273232 315304 273244
rect 315356 273232 315362 273284
rect 158070 273164 158076 273216
rect 158128 273204 158134 273216
rect 226334 273204 226340 273216
rect 158128 273176 226340 273204
rect 158128 273164 158134 273176
rect 226334 273164 226340 273176
rect 226392 273164 226398 273216
rect 300118 273164 300124 273216
rect 300176 273204 300182 273216
rect 319990 273204 319996 273216
rect 300176 273176 319996 273204
rect 300176 273164 300182 273176
rect 319990 273164 319996 273176
rect 320048 273164 320054 273216
rect 364242 273164 364248 273216
rect 364300 273204 364306 273216
rect 522206 273204 522212 273216
rect 364300 273176 522212 273204
rect 364300 273164 364306 273176
rect 522206 273164 522212 273176
rect 522264 273164 522270 273216
rect 152182 273096 152188 273148
rect 152240 273136 152246 273148
rect 223666 273136 223672 273148
rect 152240 273108 223672 273136
rect 152240 273096 152246 273108
rect 223666 273096 223672 273108
rect 223724 273096 223730 273148
rect 301498 273096 301504 273148
rect 301556 273136 301562 273148
rect 321186 273136 321192 273148
rect 301556 273108 321192 273136
rect 301556 273096 301562 273108
rect 321186 273096 321192 273108
rect 321244 273096 321250 273148
rect 369762 273096 369768 273148
rect 369820 273136 369826 273148
rect 536374 273136 536380 273148
rect 369820 273108 536380 273136
rect 369820 273096 369826 273108
rect 536374 273096 536380 273108
rect 536432 273096 536438 273148
rect 42150 273028 42156 273080
rect 42208 273068 42214 273080
rect 42702 273068 42708 273080
rect 42208 273040 42708 273068
rect 42208 273028 42214 273040
rect 42702 273028 42708 273040
rect 42760 273028 42766 273080
rect 141510 273028 141516 273080
rect 141568 273068 141574 273080
rect 220814 273068 220820 273080
rect 141568 273040 220820 273068
rect 141568 273028 141574 273040
rect 220814 273028 220820 273040
rect 220872 273028 220878 273080
rect 314470 273028 314476 273080
rect 314528 273068 314534 273080
rect 387426 273068 387432 273080
rect 314528 273040 387432 273068
rect 314528 273028 314534 273040
rect 387426 273028 387432 273040
rect 387484 273028 387490 273080
rect 388438 273028 388444 273080
rect 388496 273068 388502 273080
rect 565906 273068 565912 273080
rect 388496 273040 565912 273068
rect 388496 273028 388502 273040
rect 565906 273028 565912 273040
rect 565964 273028 565970 273080
rect 120258 272960 120264 273012
rect 120316 273000 120322 273012
rect 212718 273000 212724 273012
rect 120316 272972 212724 273000
rect 120316 272960 120322 272972
rect 212718 272960 212724 272972
rect 212776 272960 212782 273012
rect 219526 272960 219532 273012
rect 219584 273000 219590 273012
rect 219584 272972 238754 273000
rect 219584 272960 219590 272972
rect 117866 272892 117872 272944
rect 117924 272932 117930 272944
rect 211982 272932 211988 272944
rect 117924 272904 211988 272932
rect 117924 272892 117930 272904
rect 211982 272892 211988 272904
rect 212040 272892 212046 272944
rect 236730 272932 236736 272944
rect 224926 272904 236736 272932
rect 101306 272824 101312 272876
rect 101364 272864 101370 272876
rect 204806 272864 204812 272876
rect 101364 272836 204812 272864
rect 101364 272824 101370 272836
rect 204806 272824 204812 272836
rect 204864 272824 204870 272876
rect 94222 272756 94228 272808
rect 94280 272796 94286 272808
rect 201586 272796 201592 272808
rect 94280 272768 201592 272796
rect 94280 272756 94286 272768
rect 201586 272756 201592 272768
rect 201644 272756 201650 272808
rect 204162 272756 204168 272808
rect 204220 272796 204226 272808
rect 224926 272796 224954 272904
rect 236730 272892 236736 272904
rect 236788 272892 236794 272944
rect 238726 272864 238754 272972
rect 314286 272960 314292 273012
rect 314344 273000 314350 273012
rect 388622 273000 388628 273012
rect 314344 272972 388628 273000
rect 314344 272960 314350 272972
rect 388622 272960 388628 272972
rect 388680 272960 388686 273012
rect 397270 272960 397276 273012
rect 397328 273000 397334 273012
rect 581638 273000 581644 273012
rect 397328 272972 581644 273000
rect 397328 272960 397334 272972
rect 581638 272960 581644 272972
rect 581696 272960 581702 273012
rect 315850 272892 315856 272944
rect 315908 272932 315914 272944
rect 390922 272932 390928 272944
rect 315908 272904 390928 272932
rect 315908 272892 315914 272904
rect 390922 272892 390928 272904
rect 390980 272892 390986 272944
rect 398926 272892 398932 272944
rect 398984 272932 398990 272944
rect 591942 272932 591948 272944
rect 398984 272904 591948 272932
rect 398984 272892 398990 272904
rect 591942 272892 591948 272904
rect 592000 272892 592006 272944
rect 249978 272864 249984 272876
rect 238726 272836 249984 272864
rect 249978 272824 249984 272836
rect 250036 272824 250042 272876
rect 289170 272824 289176 272876
rect 289228 272864 289234 272876
rect 301130 272864 301136 272876
rect 289228 272836 301136 272864
rect 289228 272824 289234 272836
rect 301130 272824 301136 272836
rect 301188 272824 301194 272876
rect 317230 272824 317236 272876
rect 317288 272864 317294 272876
rect 394510 272864 394516 272876
rect 317288 272836 394516 272864
rect 317288 272824 317294 272836
rect 394510 272824 394516 272836
rect 394568 272824 394574 272876
rect 400306 272824 400312 272876
rect 400364 272864 400370 272876
rect 594794 272864 594800 272876
rect 400364 272836 594800 272864
rect 400364 272824 400370 272836
rect 594794 272824 594800 272836
rect 594852 272824 594858 272876
rect 239214 272796 239220 272808
rect 204220 272768 224954 272796
rect 234586 272768 239220 272796
rect 204220 272756 204226 272768
rect 78858 272688 78864 272740
rect 78916 272728 78922 272740
rect 191098 272728 191104 272740
rect 78916 272700 191104 272728
rect 78916 272688 78922 272700
rect 191098 272688 191104 272700
rect 191156 272688 191162 272740
rect 191190 272688 191196 272740
rect 191248 272728 191254 272740
rect 234586 272728 234614 272768
rect 239214 272756 239220 272768
rect 239272 272756 239278 272808
rect 291838 272756 291844 272808
rect 291896 272796 291902 272808
rect 311710 272796 311716 272808
rect 291896 272768 311716 272796
rect 291896 272756 291902 272768
rect 311710 272756 311716 272768
rect 311768 272756 311774 272808
rect 322658 272756 322664 272808
rect 322716 272796 322722 272808
rect 411806 272796 411812 272808
rect 322716 272768 411812 272796
rect 322716 272756 322722 272768
rect 411806 272756 411812 272768
rect 411864 272756 411870 272808
rect 411898 272756 411904 272808
rect 411956 272796 411962 272808
rect 610802 272796 610808 272808
rect 411956 272768 610808 272796
rect 411956 272756 411962 272768
rect 610802 272756 610808 272768
rect 610860 272756 610866 272808
rect 191248 272700 234614 272728
rect 191248 272688 191254 272700
rect 240042 272688 240048 272740
rect 240100 272728 240106 272740
rect 248598 272728 248604 272740
rect 240100 272700 248604 272728
rect 240100 272688 240106 272700
rect 248598 272688 248604 272700
rect 248656 272688 248662 272740
rect 282822 272688 282828 272740
rect 282880 272728 282886 272740
rect 305822 272728 305828 272740
rect 282880 272700 305828 272728
rect 282880 272688 282886 272700
rect 305822 272688 305828 272700
rect 305880 272688 305886 272740
rect 318610 272688 318616 272740
rect 318668 272728 318674 272740
rect 398006 272728 398012 272740
rect 318668 272700 398012 272728
rect 318668 272688 318674 272700
rect 398006 272688 398012 272700
rect 398064 272688 398070 272740
rect 401962 272688 401968 272740
rect 402020 272728 402026 272740
rect 621474 272728 621480 272740
rect 402020 272700 621480 272728
rect 402020 272688 402026 272700
rect 621474 272688 621480 272700
rect 621532 272688 621538 272740
rect 84746 272620 84752 272672
rect 84804 272660 84810 272672
rect 198918 272660 198924 272672
rect 84804 272632 198924 272660
rect 84804 272620 84810 272632
rect 198918 272620 198924 272632
rect 198976 272620 198982 272672
rect 206554 272620 206560 272672
rect 206612 272660 206618 272672
rect 244366 272660 244372 272672
rect 206612 272632 244372 272660
rect 206612 272620 206618 272632
rect 244366 272620 244372 272632
rect 244424 272620 244430 272672
rect 285582 272620 285588 272672
rect 285640 272660 285646 272672
rect 312906 272660 312912 272672
rect 285640 272632 312912 272660
rect 285640 272620 285646 272632
rect 312906 272620 312912 272632
rect 312964 272620 312970 272672
rect 319990 272620 319996 272672
rect 320048 272660 320054 272672
rect 401594 272660 401600 272672
rect 320048 272632 401600 272660
rect 320048 272620 320054 272632
rect 401594 272620 401600 272632
rect 401652 272620 401658 272672
rect 403250 272620 403256 272672
rect 403308 272660 403314 272672
rect 625062 272660 625068 272672
rect 403308 272632 625068 272660
rect 403308 272620 403314 272632
rect 625062 272620 625068 272632
rect 625120 272620 625126 272672
rect 77202 272552 77208 272604
rect 77260 272592 77266 272604
rect 194686 272592 194692 272604
rect 77260 272564 194692 272592
rect 77260 272552 77266 272564
rect 194686 272552 194692 272564
rect 194744 272552 194750 272604
rect 201770 272552 201776 272604
rect 201828 272592 201834 272604
rect 243170 272592 243176 272604
rect 201828 272564 243176 272592
rect 201828 272552 201834 272564
rect 243170 272552 243176 272564
rect 243228 272552 243234 272604
rect 246758 272552 246764 272604
rect 246816 272592 246822 272604
rect 259638 272592 259644 272604
rect 246816 272564 259644 272592
rect 246816 272552 246822 272564
rect 259638 272552 259644 272564
rect 259696 272552 259702 272604
rect 288342 272552 288348 272604
rect 288400 272592 288406 272604
rect 317690 272592 317696 272604
rect 288400 272564 317696 272592
rect 288400 272552 288406 272564
rect 317690 272552 317696 272564
rect 317748 272552 317754 272604
rect 321370 272552 321376 272604
rect 321428 272592 321434 272604
rect 405182 272592 405188 272604
rect 321428 272564 405188 272592
rect 321428 272552 321434 272564
rect 405182 272552 405188 272564
rect 405240 272552 405246 272604
rect 405550 272552 405556 272604
rect 405608 272592 405614 272604
rect 632146 272592 632152 272604
rect 405608 272564 632152 272592
rect 405608 272552 405614 272564
rect 632146 272552 632152 272564
rect 632204 272552 632210 272604
rect 72970 272484 72976 272536
rect 73028 272524 73034 272536
rect 194778 272524 194784 272536
rect 73028 272496 194784 272524
rect 73028 272484 73034 272496
rect 194778 272484 194784 272496
rect 194836 272484 194842 272536
rect 195882 272484 195888 272536
rect 195940 272524 195946 272536
rect 240962 272524 240968 272536
rect 195940 272496 240968 272524
rect 195940 272484 195946 272496
rect 240962 272484 240968 272496
rect 241020 272484 241026 272536
rect 245562 272484 245568 272536
rect 245620 272524 245626 272536
rect 259730 272524 259736 272536
rect 245620 272496 259736 272524
rect 245620 272484 245626 272496
rect 259730 272484 259736 272496
rect 259788 272484 259794 272536
rect 274174 272484 274180 272536
rect 274232 272524 274238 272536
rect 282178 272524 282184 272536
rect 274232 272496 282184 272524
rect 274232 272484 274238 272496
rect 282178 272484 282184 272496
rect 282236 272484 282242 272536
rect 286870 272484 286876 272536
rect 286928 272524 286934 272536
rect 316494 272524 316500 272536
rect 286928 272496 316500 272524
rect 286928 272484 286934 272496
rect 316494 272484 316500 272496
rect 316552 272484 316558 272536
rect 321462 272484 321468 272536
rect 321520 272524 321526 272536
rect 408678 272524 408684 272536
rect 321520 272496 408684 272524
rect 321520 272484 321526 272496
rect 408678 272484 408684 272496
rect 408736 272484 408742 272536
rect 409782 272484 409788 272536
rect 409840 272524 409846 272536
rect 642726 272524 642732 272536
rect 409840 272496 642732 272524
rect 409840 272484 409846 272496
rect 642726 272484 642732 272496
rect 642784 272484 642790 272536
rect 162762 272416 162768 272468
rect 162820 272456 162826 272468
rect 228818 272456 228824 272468
rect 162820 272428 228824 272456
rect 162820 272416 162826 272428
rect 228818 272416 228824 272428
rect 228876 272416 228882 272468
rect 362678 272416 362684 272468
rect 362736 272456 362742 272468
rect 515122 272456 515128 272468
rect 362736 272428 515128 272456
rect 362736 272416 362742 272428
rect 515122 272416 515128 272428
rect 515180 272416 515186 272468
rect 187602 272348 187608 272400
rect 187660 272388 187666 272400
rect 235258 272388 235264 272400
rect 187660 272360 235264 272388
rect 187660 272348 187666 272360
rect 235258 272348 235264 272360
rect 235316 272348 235322 272400
rect 359918 272348 359924 272400
rect 359976 272388 359982 272400
rect 507946 272388 507952 272400
rect 359976 272360 507952 272388
rect 359976 272348 359982 272360
rect 507946 272348 507952 272360
rect 508004 272348 508010 272400
rect 193490 272280 193496 272332
rect 193548 272320 193554 272332
rect 240226 272320 240232 272332
rect 193548 272292 240232 272320
rect 193548 272280 193554 272292
rect 240226 272280 240232 272292
rect 240284 272280 240290 272332
rect 332502 272280 332508 272332
rect 332560 272320 332566 272332
rect 332560 272292 431954 272320
rect 332560 272280 332566 272292
rect 182910 272212 182916 272264
rect 182968 272252 182974 272264
rect 225598 272252 225604 272264
rect 182968 272224 225604 272252
rect 182968 272212 182974 272224
rect 225598 272212 225604 272224
rect 225656 272212 225662 272264
rect 329098 272212 329104 272264
rect 329156 272252 329162 272264
rect 426434 272252 426440 272264
rect 329156 272224 426440 272252
rect 329156 272212 329162 272224
rect 426434 272212 426440 272224
rect 426492 272212 426498 272264
rect 431926 272252 431954 272292
rect 435358 272280 435364 272332
rect 435416 272320 435422 272332
rect 441798 272320 441804 272332
rect 435416 272292 441804 272320
rect 435416 272280 435422 272292
rect 441798 272280 441804 272292
rect 441856 272280 441862 272332
rect 491294 272280 491300 272332
rect 491352 272320 491358 272332
rect 492214 272320 492220 272332
rect 491352 272292 492220 272320
rect 491352 272280 491358 272292
rect 492214 272280 492220 272292
rect 492272 272280 492278 272332
rect 437014 272252 437020 272264
rect 431926 272224 437020 272252
rect 437014 272212 437020 272224
rect 437072 272212 437078 272264
rect 325602 272144 325608 272196
rect 325660 272184 325666 272196
rect 419350 272184 419356 272196
rect 325660 272156 419356 272184
rect 325660 272144 325666 272156
rect 419350 272144 419356 272156
rect 419408 272144 419414 272196
rect 420178 272144 420184 272196
rect 420236 272184 420242 272196
rect 434714 272184 434720 272196
rect 420236 272156 434720 272184
rect 420236 272144 420242 272156
rect 434714 272144 434720 272156
rect 434772 272144 434778 272196
rect 324130 272076 324136 272128
rect 324188 272116 324194 272128
rect 415762 272116 415768 272128
rect 324188 272088 415768 272116
rect 324188 272076 324194 272088
rect 415762 272076 415768 272088
rect 415820 272076 415826 272128
rect 328362 272008 328368 272060
rect 328420 272048 328426 272060
rect 403434 272048 403440 272060
rect 328420 272020 403440 272048
rect 328420 272008 328426 272020
rect 403434 272008 403440 272020
rect 403492 272008 403498 272060
rect 395798 271940 395804 271992
rect 395856 271980 395862 271992
rect 466730 271980 466736 271992
rect 395856 271952 466736 271980
rect 395856 271940 395862 271952
rect 466730 271940 466736 271952
rect 466788 271940 466794 271992
rect 387058 271872 387064 271924
rect 387116 271912 387122 271924
rect 399202 271912 399208 271924
rect 387116 271884 399208 271912
rect 387116 271872 387122 271884
rect 399202 271872 399208 271884
rect 399260 271872 399266 271924
rect 161566 271804 161572 271856
rect 161624 271844 161630 271856
rect 227990 271844 227996 271856
rect 161624 271816 227996 271844
rect 161624 271804 161630 271816
rect 227990 271804 227996 271816
rect 228048 271804 228054 271856
rect 296530 271804 296536 271856
rect 296588 271844 296594 271856
rect 340138 271844 340144 271856
rect 296588 271816 340144 271844
rect 296588 271804 296594 271816
rect 340138 271804 340144 271816
rect 340196 271804 340202 271856
rect 368106 271804 368112 271856
rect 368164 271844 368170 271856
rect 531590 271844 531596 271856
rect 368164 271816 531596 271844
rect 368164 271804 368170 271816
rect 531590 271804 531596 271816
rect 531648 271804 531654 271856
rect 155678 271736 155684 271788
rect 155736 271776 155742 271788
rect 226150 271776 226156 271788
rect 155736 271748 226156 271776
rect 155736 271736 155742 271748
rect 226150 271736 226156 271748
rect 226208 271736 226214 271788
rect 287790 271736 287796 271788
rect 287848 271776 287854 271788
rect 294046 271776 294052 271788
rect 287848 271748 294052 271776
rect 287848 271736 287854 271748
rect 294046 271736 294052 271748
rect 294104 271736 294110 271788
rect 297818 271736 297824 271788
rect 297876 271776 297882 271788
rect 343634 271776 343640 271788
rect 297876 271748 343640 271776
rect 297876 271736 297882 271748
rect 343634 271736 343640 271748
rect 343692 271736 343698 271788
rect 369486 271736 369492 271788
rect 369544 271776 369550 271788
rect 535178 271776 535184 271788
rect 369544 271748 535184 271776
rect 369544 271736 369550 271748
rect 535178 271736 535184 271748
rect 535236 271736 535242 271788
rect 145006 271668 145012 271720
rect 145064 271708 145070 271720
rect 222286 271708 222292 271720
rect 145064 271680 222292 271708
rect 145064 271668 145070 271680
rect 222286 271668 222292 271680
rect 222344 271668 222350 271720
rect 302142 271668 302148 271720
rect 302200 271708 302206 271720
rect 354306 271708 354312 271720
rect 302200 271680 354312 271708
rect 302200 271668 302206 271680
rect 354306 271668 354312 271680
rect 354364 271668 354370 271720
rect 370774 271668 370780 271720
rect 370832 271708 370838 271720
rect 538766 271708 538772 271720
rect 370832 271680 538772 271708
rect 370832 271668 370838 271680
rect 538766 271668 538772 271680
rect 538824 271668 538830 271720
rect 136818 271600 136824 271652
rect 136876 271640 136882 271652
rect 218238 271640 218244 271652
rect 136876 271612 218244 271640
rect 136876 271600 136882 271612
rect 218238 271600 218244 271612
rect 218296 271600 218302 271652
rect 252922 271600 252928 271652
rect 252980 271640 252986 271652
rect 257430 271640 257436 271652
rect 252980 271612 257436 271640
rect 252980 271600 252986 271612
rect 257430 271600 257436 271612
rect 257488 271600 257494 271652
rect 304810 271600 304816 271652
rect 304868 271640 304874 271652
rect 362586 271640 362592 271652
rect 304868 271612 362592 271640
rect 304868 271600 304874 271612
rect 362586 271600 362592 271612
rect 362644 271600 362650 271652
rect 372154 271600 372160 271652
rect 372212 271640 372218 271652
rect 542262 271640 542268 271652
rect 372212 271612 542268 271640
rect 372212 271600 372218 271612
rect 542262 271600 542268 271612
rect 542320 271600 542326 271652
rect 83550 271532 83556 271584
rect 83608 271572 83614 271584
rect 164878 271572 164884 271584
rect 83608 271544 164884 271572
rect 83608 271532 83614 271544
rect 164878 271532 164884 271544
rect 164936 271532 164942 271584
rect 165154 271532 165160 271584
rect 165212 271572 165218 271584
rect 229278 271572 229284 271584
rect 165212 271544 229284 271572
rect 165212 271532 165218 271544
rect 229278 271532 229284 271544
rect 229336 271532 229342 271584
rect 306282 271532 306288 271584
rect 306340 271572 306346 271584
rect 366082 271572 366088 271584
rect 306340 271544 366088 271572
rect 306340 271532 306346 271544
rect 366082 271532 366088 271544
rect 366140 271532 366146 271584
rect 373810 271532 373816 271584
rect 373868 271572 373874 271584
rect 547046 271572 547052 271584
rect 373868 271544 547052 271572
rect 373868 271532 373874 271544
rect 547046 271532 547052 271544
rect 547104 271532 547110 271584
rect 135622 271464 135628 271516
rect 135680 271504 135686 271516
rect 218698 271504 218704 271516
rect 135680 271476 218704 271504
rect 135680 271464 135686 271476
rect 218698 271464 218704 271476
rect 218756 271464 218762 271516
rect 224954 271464 224960 271516
rect 225012 271504 225018 271516
rect 247310 271504 247316 271516
rect 225012 271476 247316 271504
rect 225012 271464 225018 271476
rect 247310 271464 247316 271476
rect 247368 271464 247374 271516
rect 307570 271464 307576 271516
rect 307628 271504 307634 271516
rect 369302 271504 369308 271516
rect 307628 271476 369308 271504
rect 307628 271464 307634 271476
rect 369302 271464 369308 271476
rect 369360 271464 369366 271516
rect 375282 271464 375288 271516
rect 375340 271504 375346 271516
rect 550542 271504 550548 271516
rect 375340 271476 550548 271504
rect 375340 271464 375346 271476
rect 550542 271464 550548 271476
rect 550600 271464 550606 271516
rect 114278 271396 114284 271448
rect 114336 271436 114342 271448
rect 200850 271436 200856 271448
rect 114336 271408 200856 271436
rect 114336 271396 114342 271408
rect 200850 271396 200856 271408
rect 200908 271396 200914 271448
rect 202966 271396 202972 271448
rect 203024 271436 203030 271448
rect 242986 271436 242992 271448
rect 203024 271408 242992 271436
rect 203024 271396 203030 271408
rect 242986 271396 242992 271408
rect 243044 271396 243050 271448
rect 307478 271396 307484 271448
rect 307536 271436 307542 271448
rect 370866 271436 370872 271448
rect 307536 271408 370872 271436
rect 307536 271396 307542 271408
rect 370866 271396 370872 271408
rect 370924 271396 370930 271448
rect 376570 271396 376576 271448
rect 376628 271436 376634 271448
rect 554130 271436 554136 271448
rect 376628 271408 554136 271436
rect 376628 271396 376634 271408
rect 554130 271396 554136 271408
rect 554188 271396 554194 271448
rect 127342 271328 127348 271380
rect 127400 271368 127406 271380
rect 215478 271368 215484 271380
rect 127400 271340 215484 271368
rect 127400 271328 127406 271340
rect 215478 271328 215484 271340
rect 215536 271328 215542 271380
rect 230198 271328 230204 271380
rect 230256 271368 230262 271380
rect 254026 271368 254032 271380
rect 230256 271340 254032 271368
rect 230256 271328 230262 271340
rect 254026 271328 254032 271340
rect 254084 271328 254090 271380
rect 308950 271328 308956 271380
rect 309008 271368 309014 271380
rect 373258 271368 373264 271380
rect 309008 271340 373264 271368
rect 309008 271328 309014 271340
rect 373258 271328 373264 271340
rect 373316 271328 373322 271380
rect 376478 271328 376484 271380
rect 376536 271368 376542 271380
rect 555234 271368 555240 271380
rect 376536 271340 555240 271368
rect 376536 271328 376542 271340
rect 555234 271328 555240 271340
rect 555292 271328 555298 271380
rect 116670 271260 116676 271312
rect 116728 271300 116734 271312
rect 211246 271300 211252 271312
rect 116728 271272 211252 271300
rect 116728 271260 116734 271272
rect 211246 271260 211252 271272
rect 211304 271260 211310 271312
rect 226610 271260 226616 271312
rect 226668 271300 226674 271312
rect 252738 271300 252744 271312
rect 226668 271272 252744 271300
rect 226668 271260 226674 271272
rect 252738 271260 252744 271272
rect 252796 271260 252802 271312
rect 279970 271260 279976 271312
rect 280028 271300 280034 271312
rect 297542 271300 297548 271312
rect 280028 271272 297548 271300
rect 280028 271260 280034 271272
rect 297542 271260 297548 271272
rect 297600 271260 297606 271312
rect 310330 271260 310336 271312
rect 310388 271300 310394 271312
rect 376754 271300 376760 271312
rect 310388 271272 376760 271300
rect 310388 271260 310394 271272
rect 376754 271260 376760 271272
rect 376812 271260 376818 271312
rect 377950 271260 377956 271312
rect 378008 271300 378014 271312
rect 557626 271300 557632 271312
rect 378008 271272 557632 271300
rect 378008 271260 378014 271272
rect 557626 271260 557632 271272
rect 557684 271260 557690 271312
rect 104894 271192 104900 271244
rect 104952 271232 104958 271244
rect 206278 271232 206284 271244
rect 104952 271204 206284 271232
rect 104952 271192 104958 271204
rect 206278 271192 206284 271204
rect 206336 271192 206342 271244
rect 224218 271192 224224 271244
rect 224276 271232 224282 271244
rect 251266 271232 251272 271244
rect 224276 271204 251272 271232
rect 224276 271192 224282 271204
rect 251266 271192 251272 271204
rect 251324 271192 251330 271244
rect 253842 271192 253848 271244
rect 253900 271232 253906 271244
rect 262306 271232 262312 271244
rect 253900 271204 262312 271232
rect 253900 271192 253906 271204
rect 262306 271192 262312 271204
rect 262364 271192 262370 271244
rect 281350 271192 281356 271244
rect 281408 271232 281414 271244
rect 299934 271232 299940 271244
rect 281408 271204 299940 271232
rect 281408 271192 281414 271204
rect 299934 271192 299940 271204
rect 299992 271192 299998 271244
rect 311710 271192 311716 271244
rect 311768 271232 311774 271244
rect 380342 271232 380348 271244
rect 311768 271204 380348 271232
rect 311768 271192 311774 271204
rect 380342 271192 380348 271204
rect 380400 271192 380406 271244
rect 380618 271192 380624 271244
rect 380676 271232 380682 271244
rect 564710 271232 564716 271244
rect 380676 271204 564716 271232
rect 380676 271192 380682 271204
rect 564710 271192 564716 271204
rect 564768 271192 564774 271244
rect 68186 271124 68192 271176
rect 68244 271164 68250 271176
rect 193214 271164 193220 271176
rect 68244 271136 193220 271164
rect 68244 271124 68250 271136
rect 193214 271124 193220 271136
rect 193272 271124 193278 271176
rect 200574 271124 200580 271176
rect 200632 271164 200638 271176
rect 242158 271164 242164 271176
rect 200632 271136 242164 271164
rect 200632 271124 200638 271136
rect 242158 271124 242164 271136
rect 242216 271124 242222 271176
rect 242250 271124 242256 271176
rect 242308 271164 242314 271176
rect 258258 271164 258264 271176
rect 242308 271136 258264 271164
rect 242308 271124 242314 271136
rect 258258 271124 258264 271136
rect 258316 271124 258322 271176
rect 284018 271124 284024 271176
rect 284076 271164 284082 271176
rect 308214 271164 308220 271176
rect 284076 271136 308220 271164
rect 284076 271124 284082 271136
rect 308214 271124 308220 271136
rect 308272 271124 308278 271176
rect 315298 271124 315304 271176
rect 315356 271164 315362 271176
rect 383838 271164 383844 271176
rect 315356 271136 383844 271164
rect 315356 271124 315362 271136
rect 383838 271124 383844 271136
rect 383896 271124 383902 271176
rect 392578 271124 392584 271176
rect 392636 271164 392642 271176
rect 594334 271164 594340 271176
rect 392636 271136 594340 271164
rect 392636 271124 392642 271136
rect 594334 271124 594340 271136
rect 594392 271124 594398 271176
rect 166350 271056 166356 271108
rect 166408 271096 166414 271108
rect 230198 271096 230204 271108
rect 166408 271068 230204 271096
rect 166408 271056 166414 271068
rect 230198 271056 230204 271068
rect 230256 271056 230262 271108
rect 335998 271056 336004 271108
rect 336056 271096 336062 271108
rect 364978 271096 364984 271108
rect 336056 271068 364984 271096
rect 336056 271056 336062 271068
rect 364978 271056 364984 271068
rect 365036 271056 365042 271108
rect 366818 271056 366824 271108
rect 366876 271096 366882 271108
rect 528094 271096 528100 271108
rect 366876 271068 528100 271096
rect 366876 271056 366882 271068
rect 528094 271056 528100 271068
rect 528152 271056 528158 271108
rect 168650 270988 168656 271040
rect 168708 271028 168714 271040
rect 230658 271028 230664 271040
rect 168708 271000 230664 271028
rect 168708 270988 168714 271000
rect 230658 270988 230664 271000
rect 230716 270988 230722 271040
rect 326338 270988 326344 271040
rect 326396 271028 326402 271040
rect 350718 271028 350724 271040
rect 326396 271000 350724 271028
rect 326396 270988 326402 271000
rect 350718 270988 350724 271000
rect 350776 270988 350782 271040
rect 365530 270988 365536 271040
rect 365588 271028 365594 271040
rect 524506 271028 524512 271040
rect 365588 271000 524512 271028
rect 365588 270988 365594 271000
rect 524506 270988 524512 271000
rect 524564 270988 524570 271040
rect 175826 270920 175832 270972
rect 175884 270960 175890 270972
rect 233326 270960 233332 270972
rect 175884 270932 233332 270960
rect 175884 270920 175890 270932
rect 233326 270920 233332 270932
rect 233384 270920 233390 270972
rect 322290 270920 322296 270972
rect 322348 270960 322354 270972
rect 347222 270960 347228 270972
rect 322348 270932 347228 270960
rect 322348 270920 322354 270932
rect 347222 270920 347228 270932
rect 347280 270920 347286 270972
rect 364150 270920 364156 270972
rect 364208 270960 364214 270972
rect 521010 270960 521016 270972
rect 364208 270932 521016 270960
rect 364208 270920 364214 270932
rect 521010 270920 521016 270932
rect 521068 270920 521074 270972
rect 192294 270852 192300 270904
rect 192352 270892 192358 270904
rect 238846 270892 238852 270904
rect 192352 270864 238852 270892
rect 192352 270852 192358 270864
rect 238846 270852 238852 270864
rect 238904 270852 238910 270904
rect 362862 270852 362868 270904
rect 362920 270892 362926 270904
rect 517422 270892 517428 270904
rect 362920 270864 517428 270892
rect 362920 270852 362926 270864
rect 517422 270852 517428 270864
rect 517480 270852 517486 270904
rect 186406 270784 186412 270836
rect 186464 270824 186470 270836
rect 227622 270824 227628 270836
rect 186464 270796 227628 270824
rect 186464 270784 186470 270796
rect 227622 270784 227628 270796
rect 227680 270784 227686 270836
rect 337930 270784 337936 270836
rect 337988 270824 337994 270836
rect 451274 270824 451280 270836
rect 337988 270796 451280 270824
rect 337988 270784 337994 270796
rect 451274 270784 451280 270796
rect 451332 270784 451338 270836
rect 329650 270716 329656 270768
rect 329708 270756 329714 270768
rect 429930 270756 429936 270768
rect 329708 270728 429936 270756
rect 329708 270716 329714 270728
rect 429930 270716 429936 270728
rect 429988 270716 429994 270768
rect 326890 270648 326896 270700
rect 326948 270688 326954 270700
rect 422846 270688 422852 270700
rect 326948 270660 422852 270688
rect 326948 270648 326954 270660
rect 422846 270648 422852 270660
rect 422904 270648 422910 270700
rect 344278 270580 344284 270632
rect 344336 270620 344342 270632
rect 374362 270620 374368 270632
rect 344336 270592 374368 270620
rect 344336 270580 344342 270592
rect 374362 270580 374368 270592
rect 374420 270580 374426 270632
rect 351638 270512 351644 270564
rect 351696 270552 351702 270564
rect 375926 270552 375932 270564
rect 351696 270524 375932 270552
rect 351696 270512 351702 270524
rect 375926 270512 375932 270524
rect 375984 270512 375990 270564
rect 154482 270444 154488 270496
rect 154540 270484 154546 270496
rect 225322 270484 225328 270496
rect 154540 270456 225328 270484
rect 154540 270444 154546 270456
rect 225322 270444 225328 270456
rect 225380 270444 225386 270496
rect 293862 270444 293868 270496
rect 293920 270484 293926 270496
rect 335354 270484 335360 270496
rect 293920 270456 335360 270484
rect 293920 270444 293926 270456
rect 335354 270444 335360 270456
rect 335412 270444 335418 270496
rect 346762 270444 346768 270496
rect 346820 270484 346826 270496
rect 474734 270484 474740 270496
rect 346820 270456 474740 270484
rect 346820 270444 346826 270456
rect 474734 270444 474740 270456
rect 474792 270444 474798 270496
rect 147582 270376 147588 270428
rect 147640 270416 147646 270428
rect 222654 270416 222660 270428
rect 147640 270388 222660 270416
rect 147640 270376 147646 270388
rect 222654 270376 222660 270388
rect 222712 270376 222718 270428
rect 296070 270376 296076 270428
rect 296128 270416 296134 270428
rect 340874 270416 340880 270428
rect 296128 270388 340880 270416
rect 296128 270376 296134 270388
rect 340874 270376 340880 270388
rect 340932 270376 340938 270428
rect 348050 270376 348056 270428
rect 348108 270416 348114 270428
rect 477494 270416 477500 270428
rect 348108 270388 477500 270416
rect 348108 270376 348114 270388
rect 477494 270376 477500 270388
rect 477552 270376 477558 270428
rect 110782 270308 110788 270360
rect 110840 270348 110846 270360
rect 140774 270348 140780 270360
rect 110840 270320 140780 270348
rect 110840 270308 110846 270320
rect 140774 270308 140780 270320
rect 140832 270308 140838 270360
rect 143902 270308 143908 270360
rect 143960 270348 143966 270360
rect 221274 270348 221280 270360
rect 143960 270320 221280 270348
rect 143960 270308 143966 270320
rect 221274 270308 221280 270320
rect 221332 270308 221338 270360
rect 297910 270308 297916 270360
rect 297968 270348 297974 270360
rect 345014 270348 345020 270360
rect 297968 270320 345020 270348
rect 297968 270308 297974 270320
rect 345014 270308 345020 270320
rect 345072 270308 345078 270360
rect 349062 270308 349068 270360
rect 349120 270348 349126 270360
rect 481634 270348 481640 270360
rect 349120 270320 481640 270348
rect 349120 270308 349126 270320
rect 481634 270308 481640 270320
rect 481692 270308 481698 270360
rect 140682 270240 140688 270292
rect 140740 270280 140746 270292
rect 219986 270280 219992 270292
rect 140740 270252 219992 270280
rect 140740 270240 140746 270252
rect 219986 270240 219992 270252
rect 220044 270240 220050 270292
rect 220630 270240 220636 270292
rect 220688 270280 220694 270292
rect 228450 270280 228456 270292
rect 220688 270252 228456 270280
rect 220688 270240 220694 270252
rect 228450 270240 228456 270252
rect 228508 270240 228514 270292
rect 298738 270240 298744 270292
rect 298796 270280 298802 270292
rect 347774 270280 347780 270292
rect 298796 270252 347780 270280
rect 298796 270240 298802 270252
rect 347774 270240 347780 270252
rect 347832 270240 347838 270292
rect 357526 270240 357532 270292
rect 357584 270280 357590 270292
rect 503714 270280 503720 270292
rect 357584 270252 503720 270280
rect 357584 270240 357590 270252
rect 503714 270240 503720 270252
rect 503772 270240 503778 270292
rect 133782 270172 133788 270224
rect 133840 270212 133846 270224
rect 216950 270212 216956 270224
rect 133840 270184 216956 270212
rect 133840 270172 133846 270184
rect 216950 270172 216956 270184
rect 217008 270172 217014 270224
rect 234614 270172 234620 270224
rect 234672 270212 234678 270224
rect 246206 270212 246212 270224
rect 234672 270184 246212 270212
rect 234672 270172 234678 270184
rect 246206 270172 246212 270184
rect 246264 270172 246270 270224
rect 300394 270172 300400 270224
rect 300452 270212 300458 270224
rect 351914 270212 351920 270224
rect 300452 270184 351920 270212
rect 300452 270172 300458 270184
rect 351914 270172 351920 270184
rect 351972 270172 351978 270224
rect 360194 270172 360200 270224
rect 360252 270212 360258 270224
rect 510614 270212 510620 270224
rect 360252 270184 510620 270212
rect 360252 270172 360258 270184
rect 510614 270172 510620 270184
rect 510672 270172 510678 270224
rect 129550 270104 129556 270156
rect 129608 270144 129614 270156
rect 215662 270144 215668 270156
rect 129608 270116 215668 270144
rect 129608 270104 129614 270116
rect 215662 270104 215668 270116
rect 215720 270104 215726 270156
rect 231762 270104 231768 270156
rect 231820 270144 231826 270156
rect 246666 270144 246672 270156
rect 231820 270116 246672 270144
rect 231820 270104 231826 270116
rect 246666 270104 246672 270116
rect 246724 270104 246730 270156
rect 297450 270104 297456 270156
rect 297508 270144 297514 270156
rect 343818 270144 343824 270156
rect 297508 270116 343824 270144
rect 297508 270104 297514 270116
rect 343818 270104 343824 270116
rect 343876 270104 343882 270156
rect 344002 270104 344008 270156
rect 344060 270144 344066 270156
rect 467834 270144 467840 270156
rect 344060 270116 467840 270144
rect 344060 270104 344066 270116
rect 467834 270104 467840 270116
rect 467892 270104 467898 270156
rect 469306 270104 469312 270156
rect 469364 270144 469370 270156
rect 625154 270144 625160 270156
rect 469364 270116 625160 270144
rect 469364 270104 469370 270116
rect 625154 270104 625160 270116
rect 625212 270104 625218 270156
rect 126882 270036 126888 270088
rect 126940 270076 126946 270088
rect 214650 270076 214656 270088
rect 126940 270048 214656 270076
rect 126940 270036 126946 270048
rect 214650 270036 214656 270048
rect 214708 270036 214714 270088
rect 241422 270036 241428 270088
rect 241480 270076 241486 270088
rect 258074 270076 258080 270088
rect 241480 270048 258080 270076
rect 241480 270036 241486 270048
rect 258074 270036 258080 270048
rect 258132 270036 258138 270088
rect 273346 270036 273352 270088
rect 273404 270076 273410 270088
rect 280154 270076 280160 270088
rect 273404 270048 280160 270076
rect 273404 270036 273410 270048
rect 280154 270036 280160 270048
rect 280212 270036 280218 270088
rect 282730 270036 282736 270088
rect 282788 270076 282794 270088
rect 289814 270076 289820 270088
rect 282788 270048 289820 270076
rect 282788 270036 282794 270048
rect 289814 270036 289820 270048
rect 289872 270036 289878 270088
rect 301406 270036 301412 270088
rect 301464 270076 301470 270088
rect 354674 270076 354680 270088
rect 301464 270048 354680 270076
rect 301464 270036 301470 270048
rect 354674 270036 354680 270048
rect 354732 270036 354738 270088
rect 365622 270036 365628 270088
rect 365680 270076 365686 270088
rect 524598 270076 524604 270088
rect 365680 270048 524604 270076
rect 365680 270036 365686 270048
rect 524598 270036 524604 270048
rect 524656 270036 524662 270088
rect 77110 269968 77116 270020
rect 77168 270008 77174 270020
rect 124214 270008 124220 270020
rect 77168 269980 124220 270008
rect 77168 269968 77174 269980
rect 124214 269968 124220 269980
rect 124272 269968 124278 270020
rect 125502 269968 125508 270020
rect 125560 270008 125566 270020
rect 215018 270008 215024 270020
rect 125560 269980 215024 270008
rect 125560 269968 125566 269980
rect 215018 269968 215024 269980
rect 215076 269968 215082 270020
rect 236086 269968 236092 270020
rect 236144 270008 236150 270020
rect 256418 270008 256424 270020
rect 236144 269980 256424 270008
rect 236144 269968 236150 269980
rect 256418 269968 256424 269980
rect 256476 269968 256482 270020
rect 274726 269968 274732 270020
rect 274784 270008 274790 270020
rect 284294 270008 284300 270020
rect 274784 269980 284300 270008
rect 274784 269968 274790 269980
rect 284294 269968 284300 269980
rect 284352 269968 284358 270020
rect 306006 269968 306012 270020
rect 306064 270008 306070 270020
rect 358814 270008 358820 270020
rect 306064 269980 358820 270008
rect 306064 269968 306070 269980
rect 358814 269968 358820 269980
rect 358872 269968 358878 270020
rect 372246 269968 372252 270020
rect 372304 270008 372310 270020
rect 542354 270008 542360 270020
rect 372304 269980 542360 270008
rect 372304 269968 372310 269980
rect 542354 269968 542360 269980
rect 542412 269968 542418 270020
rect 122742 269900 122748 269952
rect 122800 269940 122806 269952
rect 213270 269940 213276 269952
rect 122800 269912 213276 269940
rect 122800 269900 122806 269912
rect 213270 269900 213276 269912
rect 213328 269900 213334 269952
rect 237190 269900 237196 269952
rect 237248 269940 237254 269952
rect 256878 269940 256884 269952
rect 237248 269912 256884 269940
rect 237248 269900 237254 269912
rect 256878 269900 256884 269912
rect 256936 269900 256942 269952
rect 276014 269900 276020 269952
rect 276072 269940 276078 269952
rect 287054 269940 287060 269952
rect 276072 269912 287060 269940
rect 276072 269900 276078 269912
rect 287054 269900 287060 269912
rect 287112 269900 287118 269952
rect 303246 269900 303252 269952
rect 303304 269940 303310 269952
rect 360286 269940 360292 269952
rect 303304 269912 360292 269940
rect 303304 269900 303310 269912
rect 360286 269900 360292 269912
rect 360344 269900 360350 269952
rect 374362 269900 374368 269952
rect 374420 269940 374426 269952
rect 547874 269940 547880 269952
rect 374420 269912 547880 269940
rect 374420 269900 374426 269912
rect 547874 269900 547880 269912
rect 547932 269900 547938 269952
rect 85942 269832 85948 269884
rect 86000 269872 86006 269884
rect 116486 269872 116492 269884
rect 86000 269844 116492 269872
rect 86000 269832 86006 269844
rect 116486 269832 116492 269844
rect 116544 269832 116550 269884
rect 119062 269832 119068 269884
rect 119120 269872 119126 269884
rect 211890 269872 211896 269884
rect 119120 269844 211896 269872
rect 119120 269832 119126 269844
rect 211890 269832 211896 269844
rect 211948 269832 211954 269884
rect 233694 269832 233700 269884
rect 233752 269872 233758 269884
rect 255590 269872 255596 269884
rect 233752 269844 255596 269872
rect 233752 269832 233758 269844
rect 255590 269832 255596 269844
rect 255648 269832 255654 269884
rect 277854 269832 277860 269884
rect 277912 269872 277918 269884
rect 292574 269872 292580 269884
rect 277912 269844 292580 269872
rect 277912 269832 277918 269844
rect 292574 269832 292580 269844
rect 292632 269832 292638 269884
rect 305914 269832 305920 269884
rect 305972 269872 305978 269884
rect 367094 269872 367100 269884
rect 305972 269844 367100 269872
rect 305972 269832 305978 269844
rect 367094 269832 367100 269844
rect 367152 269832 367158 269884
rect 378042 269832 378048 269884
rect 378100 269872 378106 269884
rect 557718 269872 557724 269884
rect 378100 269844 557724 269872
rect 378100 269832 378106 269844
rect 557718 269832 557724 269844
rect 557776 269832 557782 269884
rect 108942 269764 108948 269816
rect 109000 269804 109006 269816
rect 207934 269804 207940 269816
rect 109000 269776 207940 269804
rect 109000 269764 109006 269776
rect 207934 269764 207940 269776
rect 207992 269764 207998 269816
rect 229922 269764 229928 269816
rect 229980 269804 229986 269816
rect 253382 269804 253388 269816
rect 229980 269776 253388 269804
rect 229980 269764 229986 269776
rect 253382 269764 253388 269776
rect 253440 269764 253446 269816
rect 279142 269764 279148 269816
rect 279200 269804 279206 269816
rect 295334 269804 295340 269816
rect 279200 269776 295340 269804
rect 279200 269764 279206 269776
rect 295334 269764 295340 269776
rect 295392 269764 295398 269816
rect 321922 269764 321928 269816
rect 321980 269804 321986 269816
rect 389266 269804 389272 269816
rect 321980 269776 389272 269804
rect 321980 269764 321986 269776
rect 389266 269764 389272 269776
rect 389324 269764 389330 269816
rect 390002 269764 390008 269816
rect 390060 269804 390066 269816
rect 590654 269804 590660 269816
rect 390060 269776 590660 269804
rect 390060 269764 390066 269776
rect 590654 269764 590660 269776
rect 590712 269764 590718 269816
rect 232866 269736 232872 269748
rect 177776 269708 232872 269736
rect 146202 269628 146208 269680
rect 146260 269668 146266 269680
rect 177574 269668 177580 269680
rect 146260 269640 177580 269668
rect 146260 269628 146266 269640
rect 177574 269628 177580 269640
rect 177632 269628 177638 269680
rect 173802 269560 173808 269612
rect 173860 269600 173866 269612
rect 177776 269600 177804 269708
rect 232866 269696 232872 269708
rect 232924 269696 232930 269748
rect 294782 269696 294788 269748
rect 294840 269736 294846 269748
rect 336734 269736 336740 269748
rect 294840 269708 336740 269736
rect 294840 269696 294846 269708
rect 336734 269696 336740 269708
rect 336792 269696 336798 269748
rect 345106 269696 345112 269748
rect 345164 269736 345170 269748
rect 470594 269736 470600 269748
rect 345164 269708 470600 269736
rect 345164 269696 345170 269708
rect 470594 269696 470600 269708
rect 470652 269696 470658 269748
rect 234154 269668 234160 269680
rect 173860 269572 177804 269600
rect 177868 269640 234160 269668
rect 173860 269560 173866 269572
rect 176930 269492 176936 269544
rect 176988 269532 176994 269544
rect 177868 269532 177896 269640
rect 234154 269628 234160 269640
rect 234212 269628 234218 269680
rect 293402 269628 293408 269680
rect 293460 269668 293466 269680
rect 333974 269668 333980 269680
rect 293460 269640 333980 269668
rect 293460 269628 293466 269640
rect 333974 269628 333980 269640
rect 334032 269628 334038 269680
rect 342438 269628 342444 269680
rect 342496 269668 342502 269680
rect 463694 269668 463700 269680
rect 342496 269640 463700 269668
rect 342496 269628 342502 269640
rect 463694 269628 463700 269640
rect 463752 269628 463758 269680
rect 179322 269560 179328 269612
rect 179380 269600 179386 269612
rect 234614 269600 234620 269612
rect 179380 269572 234620 269600
rect 179380 269560 179386 269572
rect 234614 269560 234620 269572
rect 234672 269560 234678 269612
rect 292114 269560 292120 269612
rect 292172 269600 292178 269612
rect 329834 269600 329840 269612
rect 292172 269572 329840 269600
rect 292172 269560 292178 269572
rect 329834 269560 329840 269572
rect 329892 269560 329898 269612
rect 341058 269560 341064 269612
rect 341116 269600 341122 269612
rect 459646 269600 459652 269612
rect 341116 269572 459652 269600
rect 341116 269560 341122 269572
rect 459646 269560 459652 269572
rect 459704 269560 459710 269612
rect 464706 269560 464712 269612
rect 464764 269600 464770 269612
rect 469214 269600 469220 269612
rect 464764 269572 469220 269600
rect 464764 269560 464770 269572
rect 469214 269560 469220 269572
rect 469272 269560 469278 269612
rect 176988 269504 177896 269532
rect 176988 269492 176994 269504
rect 180702 269492 180708 269544
rect 180760 269532 180766 269544
rect 235534 269532 235540 269544
rect 180760 269504 235540 269532
rect 180760 269492 180766 269504
rect 235534 269492 235540 269504
rect 235592 269492 235598 269544
rect 307754 269492 307760 269544
rect 307812 269532 307818 269544
rect 327074 269532 327080 269544
rect 307812 269504 327080 269532
rect 307812 269492 307818 269504
rect 327074 269492 327080 269504
rect 327132 269492 327138 269544
rect 339770 269492 339776 269544
rect 339828 269532 339834 269544
rect 456794 269532 456800 269544
rect 339828 269504 456800 269532
rect 339828 269492 339834 269504
rect 456794 269492 456800 269504
rect 456852 269492 456858 269544
rect 184842 269424 184848 269476
rect 184900 269464 184906 269476
rect 236914 269464 236920 269476
rect 184900 269436 236920 269464
rect 184900 269424 184906 269436
rect 236914 269424 236920 269436
rect 236972 269424 236978 269476
rect 338390 269424 338396 269476
rect 338448 269464 338454 269476
rect 452654 269464 452660 269476
rect 338448 269436 452660 269464
rect 338448 269424 338454 269436
rect 452654 269424 452660 269436
rect 452712 269424 452718 269476
rect 337102 269356 337108 269408
rect 337160 269396 337166 269408
rect 449894 269396 449900 269408
rect 337160 269368 449900 269396
rect 337160 269356 337166 269368
rect 449894 269356 449900 269368
rect 449952 269356 449958 269408
rect 335722 269288 335728 269340
rect 335780 269328 335786 269340
rect 445754 269328 445760 269340
rect 335780 269300 445760 269328
rect 335780 269288 335786 269300
rect 445754 269288 445760 269300
rect 445812 269288 445818 269340
rect 518986 269288 518992 269340
rect 519044 269328 519050 269340
rect 525794 269328 525800 269340
rect 519044 269300 525800 269328
rect 519044 269288 519050 269300
rect 525794 269288 525800 269300
rect 525852 269288 525858 269340
rect 323578 269220 323584 269272
rect 323636 269260 323642 269272
rect 376938 269260 376944 269272
rect 323636 269232 376944 269260
rect 323636 269220 323642 269232
rect 376938 269220 376944 269232
rect 376996 269220 377002 269272
rect 223206 269084 223212 269136
rect 223264 269124 223270 269136
rect 231118 269124 231124 269136
rect 223264 269096 231124 269124
rect 223264 269084 223270 269096
rect 231118 269084 231124 269096
rect 231176 269084 231182 269136
rect 516134 269084 516140 269136
rect 516192 269124 516198 269136
rect 518894 269124 518900 269136
rect 516192 269096 518900 269124
rect 516192 269084 516198 269096
rect 518894 269084 518900 269096
rect 518952 269084 518958 269136
rect 102502 269016 102508 269068
rect 102560 269056 102566 269068
rect 206186 269056 206192 269068
rect 102560 269028 206192 269056
rect 102560 269016 102566 269028
rect 206186 269016 206192 269028
rect 206244 269016 206250 269068
rect 323210 269016 323216 269068
rect 323268 269056 323274 269068
rect 398834 269056 398840 269068
rect 323268 269028 398840 269056
rect 323268 269016 323274 269028
rect 398834 269016 398840 269028
rect 398892 269016 398898 269068
rect 408678 269016 408684 269068
rect 408736 269056 408742 269068
rect 583754 269056 583760 269068
rect 408736 269028 583760 269056
rect 408736 269016 408742 269028
rect 583754 269016 583760 269028
rect 583812 269016 583818 269068
rect 99282 268948 99288 269000
rect 99340 268988 99346 269000
rect 204438 268988 204444 269000
rect 99340 268960 204444 268988
rect 99340 268948 99346 268960
rect 204438 268948 204444 268960
rect 204496 268948 204502 269000
rect 222102 268948 222108 269000
rect 222160 268988 222166 269000
rect 236638 268988 236644 269000
rect 222160 268960 236644 268988
rect 222160 268948 222166 268960
rect 236638 268948 236644 268960
rect 236696 268948 236702 269000
rect 309042 268948 309048 269000
rect 309100 268988 309106 269000
rect 375374 268988 375380 269000
rect 309100 268960 375380 268988
rect 309100 268948 309106 268960
rect 375374 268948 375380 268960
rect 375432 268948 375438 269000
rect 393130 268948 393136 269000
rect 393188 268988 393194 269000
rect 577682 268988 577688 269000
rect 393188 268960 577688 268988
rect 393188 268948 393194 268960
rect 577682 268948 577688 268960
rect 577740 268948 577746 269000
rect 95418 268880 95424 268932
rect 95476 268920 95482 268932
rect 203518 268920 203524 268932
rect 95476 268892 203524 268920
rect 95476 268880 95482 268892
rect 203518 268880 203524 268892
rect 203576 268880 203582 268932
rect 225414 268880 225420 268932
rect 225472 268920 225478 268932
rect 245286 268920 245292 268932
rect 225472 268892 245292 268920
rect 225472 268880 225478 268892
rect 245286 268880 245292 268892
rect 245344 268880 245350 268932
rect 310422 268880 310428 268932
rect 310480 268920 310486 268932
rect 378134 268920 378140 268932
rect 310480 268892 378140 268920
rect 310480 268880 310486 268892
rect 378134 268880 378140 268892
rect 378192 268880 378198 268932
rect 382182 268880 382188 268932
rect 382240 268920 382246 268932
rect 568574 268920 568580 268932
rect 382240 268892 568580 268920
rect 382240 268880 382246 268892
rect 568574 268880 568580 268892
rect 568632 268880 568638 268932
rect 92382 268812 92388 268864
rect 92440 268852 92446 268864
rect 202138 268852 202144 268864
rect 92440 268824 202144 268852
rect 92440 268812 92446 268824
rect 202138 268812 202144 268824
rect 202196 268812 202202 268864
rect 218330 268812 218336 268864
rect 218388 268852 218394 268864
rect 239306 268852 239312 268864
rect 218388 268824 239312 268852
rect 218388 268812 218394 268824
rect 239306 268812 239312 268824
rect 239364 268812 239370 268864
rect 284846 268812 284852 268864
rect 284904 268852 284910 268864
rect 298094 268852 298100 268864
rect 284904 268824 298100 268852
rect 284904 268812 284910 268824
rect 298094 268812 298100 268824
rect 298152 268812 298158 268864
rect 311802 268812 311808 268864
rect 311860 268852 311866 268864
rect 382274 268852 382280 268864
rect 311860 268824 382280 268852
rect 311860 268812 311866 268824
rect 382274 268812 382280 268824
rect 382332 268812 382338 268864
rect 394602 268812 394608 268864
rect 394660 268852 394666 268864
rect 601694 268852 601700 268864
rect 394660 268824 601700 268852
rect 394660 268812 394666 268824
rect 601694 268812 601700 268824
rect 601752 268812 601758 268864
rect 87138 268744 87144 268796
rect 87196 268784 87202 268796
rect 200390 268784 200396 268796
rect 87196 268756 200396 268784
rect 87196 268744 87202 268756
rect 200390 268744 200396 268756
rect 200448 268744 200454 268796
rect 201402 268744 201408 268796
rect 201460 268784 201466 268796
rect 203058 268784 203064 268796
rect 201460 268756 203064 268784
rect 201460 268744 201466 268756
rect 203058 268744 203064 268756
rect 203116 268744 203122 268796
rect 204898 268744 204904 268796
rect 204956 268784 204962 268796
rect 225782 268784 225788 268796
rect 204956 268756 225788 268784
rect 204956 268744 204962 268756
rect 225782 268744 225788 268756
rect 225840 268744 225846 268796
rect 229002 268744 229008 268796
rect 229060 268784 229066 268796
rect 253750 268784 253756 268796
rect 229060 268756 253756 268784
rect 229060 268744 229066 268756
rect 253750 268744 253756 268756
rect 253808 268744 253814 268796
rect 278682 268744 278688 268796
rect 278740 268784 278746 268796
rect 294138 268784 294144 268796
rect 278740 268756 294144 268784
rect 278740 268744 278746 268756
rect 294138 268744 294144 268756
rect 294196 268744 294202 268796
rect 312998 268744 313004 268796
rect 313056 268784 313062 268796
rect 385218 268784 385224 268796
rect 313056 268756 385224 268784
rect 313056 268744 313062 268756
rect 385218 268744 385224 268756
rect 385276 268744 385282 268796
rect 395430 268744 395436 268796
rect 395488 268784 395494 268796
rect 604454 268784 604460 268796
rect 395488 268756 604460 268784
rect 395488 268744 395494 268756
rect 604454 268744 604460 268756
rect 604512 268744 604518 268796
rect 82722 268676 82728 268728
rect 82780 268716 82786 268728
rect 198550 268716 198556 268728
rect 82780 268688 198556 268716
rect 82780 268676 82786 268688
rect 198550 268676 198556 268688
rect 198608 268676 198614 268728
rect 207014 268676 207020 268728
rect 207072 268716 207078 268728
rect 233786 268716 233792 268728
rect 207072 268688 233792 268716
rect 207072 268676 207078 268688
rect 233786 268676 233792 268688
rect 233844 268676 233850 268728
rect 290918 268676 290924 268728
rect 290976 268716 290982 268728
rect 306374 268716 306380 268728
rect 290976 268688 306380 268716
rect 290976 268676 290982 268688
rect 306374 268676 306380 268688
rect 306432 268676 306438 268728
rect 314378 268676 314384 268728
rect 314436 268716 314442 268728
rect 389174 268716 389180 268728
rect 314436 268688 389180 268716
rect 314436 268676 314442 268688
rect 389174 268676 389180 268688
rect 389232 268676 389238 268728
rect 395890 268676 395896 268728
rect 395948 268716 395954 268728
rect 605834 268716 605840 268728
rect 395948 268688 605840 268716
rect 395948 268676 395954 268688
rect 605834 268676 605840 268688
rect 605892 268676 605898 268728
rect 80054 268608 80060 268660
rect 80112 268648 80118 268660
rect 197262 268648 197268 268660
rect 80112 268620 197268 268648
rect 80112 268608 80118 268620
rect 197262 268608 197268 268620
rect 197320 268608 197326 268660
rect 215202 268608 215208 268660
rect 215260 268648 215266 268660
rect 244182 268648 244188 268660
rect 215260 268620 244188 268648
rect 215260 268608 215266 268620
rect 244182 268608 244188 268620
rect 244240 268608 244246 268660
rect 245654 268608 245660 268660
rect 245712 268648 245718 268660
rect 256050 268648 256056 268660
rect 245712 268620 256056 268648
rect 245712 268608 245718 268620
rect 256050 268608 256056 268620
rect 256108 268608 256114 268660
rect 280522 268608 280528 268660
rect 280580 268648 280586 268660
rect 291194 268648 291200 268660
rect 280580 268620 291200 268648
rect 280580 268608 280586 268620
rect 291194 268608 291200 268620
rect 291252 268608 291258 268660
rect 291470 268608 291476 268660
rect 291528 268648 291534 268660
rect 310514 268648 310520 268660
rect 291528 268620 310520 268648
rect 291528 268608 291534 268620
rect 310514 268608 310520 268620
rect 310572 268608 310578 268660
rect 315666 268608 315672 268660
rect 315724 268648 315730 268660
rect 393314 268648 393320 268660
rect 315724 268620 393320 268648
rect 315724 268608 315730 268620
rect 393314 268608 393320 268620
rect 393372 268608 393378 268660
rect 397178 268608 397184 268660
rect 397236 268648 397242 268660
rect 608594 268648 608600 268660
rect 397236 268620 608600 268648
rect 397236 268608 397242 268620
rect 608594 268608 608600 268620
rect 608652 268608 608658 268660
rect 77662 268540 77668 268592
rect 77720 268580 77726 268592
rect 196526 268580 196532 268592
rect 77720 268552 196532 268580
rect 77720 268540 77726 268552
rect 196526 268540 196532 268552
rect 196584 268540 196590 268592
rect 217134 268540 217140 268592
rect 217192 268580 217198 268592
rect 249334 268580 249340 268592
rect 217192 268552 249340 268580
rect 217192 268540 217198 268552
rect 249334 268540 249340 268552
rect 249392 268540 249398 268592
rect 283006 268540 283012 268592
rect 283064 268580 283070 268592
rect 302418 268580 302424 268592
rect 283064 268552 302424 268580
rect 283064 268540 283070 268552
rect 302418 268540 302424 268552
rect 302476 268540 302482 268592
rect 317046 268540 317052 268592
rect 317104 268580 317110 268592
rect 396074 268580 396080 268592
rect 317104 268552 396080 268580
rect 317104 268540 317110 268552
rect 396074 268540 396080 268552
rect 396132 268540 396138 268592
rect 399846 268540 399852 268592
rect 399904 268580 399910 268592
rect 615678 268580 615684 268592
rect 399904 268552 615684 268580
rect 399904 268540 399910 268552
rect 615678 268540 615684 268552
rect 615736 268540 615742 268592
rect 75822 268472 75828 268524
rect 75880 268512 75886 268524
rect 195422 268512 195428 268524
rect 75880 268484 195428 268512
rect 75880 268472 75886 268484
rect 195422 268472 195428 268484
rect 195480 268472 195486 268524
rect 211338 268472 211344 268524
rect 211396 268512 211402 268524
rect 247126 268512 247132 268524
rect 211396 268484 247132 268512
rect 211396 268472 211402 268484
rect 247126 268472 247132 268484
rect 247184 268472 247190 268524
rect 281442 268472 281448 268524
rect 281500 268512 281506 268524
rect 302234 268512 302240 268524
rect 281500 268484 302240 268512
rect 281500 268472 281506 268484
rect 302234 268472 302240 268484
rect 302292 268472 302298 268524
rect 318334 268472 318340 268524
rect 318392 268512 318398 268524
rect 400214 268512 400220 268524
rect 318392 268484 400220 268512
rect 318392 268472 318398 268484
rect 400214 268472 400220 268484
rect 400272 268472 400278 268524
rect 401134 268472 401140 268524
rect 401192 268512 401198 268524
rect 619634 268512 619640 268524
rect 401192 268484 619640 268512
rect 401192 268472 401198 268484
rect 619634 268472 619640 268484
rect 619692 268472 619698 268524
rect 69382 268404 69388 268456
rect 69440 268444 69446 268456
rect 193674 268444 193680 268456
rect 69440 268416 193680 268444
rect 69440 268404 69446 268416
rect 193674 268404 193680 268416
rect 193732 268404 193738 268456
rect 210602 268404 210608 268456
rect 210660 268444 210666 268456
rect 245746 268444 245752 268456
rect 210660 268416 245752 268444
rect 210660 268404 210666 268416
rect 245746 268404 245752 268416
rect 245804 268404 245810 268456
rect 249702 268404 249708 268456
rect 249760 268444 249766 268456
rect 261386 268444 261392 268456
rect 249760 268416 261392 268444
rect 249760 268404 249766 268416
rect 261386 268404 261392 268416
rect 261444 268404 261450 268456
rect 274266 268404 274272 268456
rect 274324 268444 274330 268456
rect 282914 268444 282920 268456
rect 274324 268416 282920 268444
rect 274324 268404 274330 268416
rect 282914 268404 282920 268416
rect 282972 268404 282978 268456
rect 286778 268404 286784 268456
rect 286836 268444 286842 268456
rect 309134 268444 309140 268456
rect 286836 268416 309140 268444
rect 286836 268404 286842 268416
rect 309134 268404 309140 268416
rect 309192 268404 309198 268456
rect 319714 268404 319720 268456
rect 319772 268444 319778 268456
rect 402974 268444 402980 268456
rect 319772 268416 402980 268444
rect 319772 268404 319778 268416
rect 402974 268404 402980 268416
rect 403032 268404 403038 268456
rect 403894 268404 403900 268456
rect 403952 268444 403958 268456
rect 626534 268444 626540 268456
rect 403952 268416 626540 268444
rect 403952 268404 403958 268416
rect 626534 268404 626540 268416
rect 626592 268404 626598 268456
rect 66162 268336 66168 268388
rect 66220 268376 66226 268388
rect 192386 268376 192392 268388
rect 66220 268348 192392 268376
rect 66220 268336 66226 268348
rect 192386 268336 192392 268348
rect 192444 268336 192450 268388
rect 195974 268336 195980 268388
rect 196032 268376 196038 268388
rect 235074 268376 235080 268388
rect 196032 268348 235080 268376
rect 196032 268336 196038 268348
rect 235074 268336 235080 268348
rect 235132 268336 235138 268388
rect 248322 268336 248328 268388
rect 248380 268376 248386 268388
rect 260926 268376 260932 268388
rect 248380 268348 260932 268376
rect 248380 268336 248386 268348
rect 260926 268336 260932 268348
rect 260984 268336 260990 268388
rect 275646 268336 275652 268388
rect 275704 268376 275710 268388
rect 285858 268376 285864 268388
rect 275704 268348 285864 268376
rect 275704 268336 275710 268348
rect 285858 268336 285864 268348
rect 285916 268336 285922 268388
rect 286226 268336 286232 268388
rect 286284 268376 286290 268388
rect 313274 268376 313280 268388
rect 286284 268348 313280 268376
rect 286284 268336 286290 268348
rect 313274 268336 313280 268348
rect 313332 268336 313338 268388
rect 322382 268336 322388 268388
rect 322440 268376 322446 268388
rect 409966 268376 409972 268388
rect 322440 268348 409972 268376
rect 322440 268336 322446 268348
rect 409966 268336 409972 268348
rect 410024 268336 410030 268388
rect 410426 268336 410432 268388
rect 410484 268376 410490 268388
rect 636194 268376 636200 268388
rect 410484 268348 636200 268376
rect 410484 268336 410490 268348
rect 636194 268336 636200 268348
rect 636252 268336 636258 268388
rect 106182 268268 106188 268320
rect 106240 268308 106246 268320
rect 207474 268308 207480 268320
rect 106240 268280 207480 268308
rect 106240 268268 106246 268280
rect 207474 268268 207480 268280
rect 207532 268268 207538 268320
rect 307662 268268 307668 268320
rect 307720 268308 307726 268320
rect 371234 268308 371240 268320
rect 307720 268280 371240 268308
rect 307720 268268 307726 268280
rect 371234 268268 371240 268280
rect 371292 268268 371298 268320
rect 371878 268268 371884 268320
rect 371936 268308 371942 268320
rect 394694 268308 394700 268320
rect 371936 268280 394700 268308
rect 371936 268268 371942 268280
rect 394694 268268 394700 268280
rect 394752 268268 394758 268320
rect 110322 268200 110328 268252
rect 110380 268240 110386 268252
rect 208854 268240 208860 268252
rect 110380 268212 208860 268240
rect 110380 268200 110386 268212
rect 208854 268200 208860 268212
rect 208912 268200 208918 268252
rect 303706 268200 303712 268252
rect 303764 268240 303770 268252
rect 360378 268240 360384 268252
rect 303764 268212 360384 268240
rect 303764 268200 303770 268212
rect 360378 268200 360384 268212
rect 360436 268200 360442 268252
rect 362954 268200 362960 268252
rect 363012 268240 363018 268252
rect 385126 268240 385132 268252
rect 363012 268212 385132 268240
rect 363012 268200 363018 268212
rect 385126 268200 385132 268212
rect 385184 268200 385190 268252
rect 390462 268200 390468 268252
rect 390520 268240 390526 268252
rect 507854 268240 507860 268252
rect 390520 268212 507860 268240
rect 390520 268200 390526 268212
rect 507854 268200 507860 268212
rect 507912 268200 507918 268252
rect 115842 268132 115848 268184
rect 115900 268172 115906 268184
rect 210602 268172 210608 268184
rect 115900 268144 210608 268172
rect 115900 268132 115906 268144
rect 210602 268132 210608 268144
rect 210660 268132 210666 268184
rect 302326 268132 302332 268184
rect 302384 268172 302390 268184
rect 357434 268172 357440 268184
rect 302384 268144 357440 268172
rect 302384 268132 302390 268144
rect 357434 268132 357440 268144
rect 357492 268132 357498 268184
rect 361482 268132 361488 268184
rect 361540 268172 361546 268184
rect 380894 268172 380900 268184
rect 361540 268144 380900 268172
rect 361540 268132 361546 268144
rect 380894 268132 380900 268144
rect 380952 268132 380958 268184
rect 389174 268132 389180 268184
rect 389232 268172 389238 268184
rect 495066 268172 495072 268184
rect 389232 268144 495072 268172
rect 389232 268132 389238 268144
rect 495066 268132 495072 268144
rect 495124 268132 495130 268184
rect 131022 268064 131028 268116
rect 131080 268104 131086 268116
rect 216858 268104 216864 268116
rect 131080 268076 216864 268104
rect 131080 268064 131086 268076
rect 216858 268064 216864 268076
rect 216916 268064 216922 268116
rect 335354 268064 335360 268116
rect 335412 268104 335418 268116
rect 368474 268104 368480 268116
rect 335412 268076 368480 268104
rect 335412 268064 335418 268076
rect 368474 268064 368480 268076
rect 368532 268064 368538 268116
rect 386506 268064 386512 268116
rect 386564 268104 386570 268116
rect 481174 268104 481180 268116
rect 386564 268076 481180 268104
rect 386564 268064 386570 268076
rect 481174 268064 481180 268076
rect 481232 268064 481238 268116
rect 663058 268064 663064 268116
rect 663116 268104 663122 268116
rect 676214 268104 676220 268116
rect 663116 268076 676220 268104
rect 663116 268064 663122 268076
rect 676214 268064 676220 268076
rect 676272 268064 676278 268116
rect 135162 267996 135168 268048
rect 135220 268036 135226 268048
rect 218146 268036 218152 268048
rect 135220 268008 218152 268036
rect 135220 267996 135226 268008
rect 218146 267996 218152 268008
rect 218204 267996 218210 268048
rect 331122 267996 331128 268048
rect 331180 268036 331186 268048
rect 413922 268036 413928 268048
rect 331180 268008 413928 268036
rect 331180 267996 331186 268008
rect 413922 267996 413928 268008
rect 413980 267996 413986 268048
rect 414014 267996 414020 268048
rect 414072 268036 414078 268048
rect 426618 268036 426624 268048
rect 414072 268008 426624 268036
rect 414072 267996 414078 268008
rect 426618 267996 426624 268008
rect 426676 267996 426682 268048
rect 190362 267928 190368 267980
rect 190420 267968 190426 267980
rect 230474 267968 230480 267980
rect 190420 267940 230480 267968
rect 190420 267928 190426 267940
rect 230474 267928 230480 267940
rect 230532 267928 230538 267980
rect 385126 267928 385132 267980
rect 385184 267968 385190 267980
rect 459738 267968 459744 267980
rect 385184 267940 459744 267968
rect 385184 267928 385190 267940
rect 459738 267928 459744 267940
rect 459796 267928 459802 267980
rect 661770 267928 661776 267980
rect 661828 267968 661834 267980
rect 676214 267968 676220 267980
rect 661828 267940 676220 267968
rect 661828 267928 661834 267940
rect 676214 267928 676220 267940
rect 676272 267928 676278 267980
rect 181162 267860 181168 267912
rect 181220 267900 181226 267912
rect 221734 267900 221740 267912
rect 181220 267872 221740 267900
rect 181220 267860 181226 267872
rect 221734 267860 221740 267872
rect 221792 267860 221798 267912
rect 342162 267860 342168 267912
rect 342220 267900 342226 267912
rect 407114 267900 407120 267912
rect 342220 267872 407120 267900
rect 342220 267860 342226 267872
rect 407114 267860 407120 267872
rect 407172 267860 407178 267912
rect 354674 267792 354680 267844
rect 354732 267832 354738 267844
rect 416774 267832 416780 267844
rect 354732 267804 416780 267832
rect 354732 267792 354738 267804
rect 416774 267792 416780 267804
rect 416832 267792 416838 267844
rect 243354 267724 243360 267776
rect 243412 267764 243418 267776
rect 250714 267764 250720 267776
rect 243412 267736 250720 267764
rect 243412 267724 243418 267736
rect 250714 267724 250720 267736
rect 250772 267724 250778 267776
rect 369670 267724 369676 267776
rect 369728 267764 369734 267776
rect 391934 267764 391940 267776
rect 369728 267736 391940 267764
rect 369728 267724 369734 267736
rect 391934 267724 391940 267736
rect 391992 267724 391998 267776
rect 392026 267724 392032 267776
rect 392084 267764 392090 267776
rect 523586 267764 523592 267776
rect 392084 267736 523592 267764
rect 392084 267724 392090 267736
rect 523586 267724 523592 267736
rect 523644 267724 523650 267776
rect 660298 267724 660304 267776
rect 660356 267764 660362 267776
rect 676122 267764 676128 267776
rect 660356 267736 676128 267764
rect 660356 267724 660362 267736
rect 676122 267724 676128 267736
rect 676180 267724 676186 267776
rect 140774 267656 140780 267708
rect 140832 267696 140838 267708
rect 209682 267696 209688 267708
rect 140832 267668 209688 267696
rect 140832 267656 140838 267668
rect 209682 267656 209688 267668
rect 209740 267656 209746 267708
rect 284938 267656 284944 267708
rect 284996 267696 285002 267708
rect 291838 267696 291844 267708
rect 284996 267668 291844 267696
rect 284996 267656 285002 267668
rect 291838 267656 291844 267668
rect 291896 267656 291902 267708
rect 299198 267656 299204 267708
rect 299256 267696 299262 267708
rect 320818 267696 320824 267708
rect 299256 267668 320824 267696
rect 299256 267656 299262 267668
rect 320818 267656 320824 267668
rect 320876 267656 320882 267708
rect 341978 267656 341984 267708
rect 342036 267696 342042 267708
rect 462314 267696 462320 267708
rect 342036 267668 462320 267696
rect 342036 267656 342042 267668
rect 462314 267656 462320 267668
rect 462372 267656 462378 267708
rect 157242 267588 157248 267640
rect 157300 267628 157306 267640
rect 227070 267628 227076 267640
rect 157300 267600 227076 267628
rect 157300 267588 157306 267600
rect 227070 267588 227076 267600
rect 227128 267588 227134 267640
rect 283190 267588 283196 267640
rect 283248 267628 283254 267640
rect 290918 267628 290924 267640
rect 283248 267600 290924 267628
rect 283248 267588 283254 267600
rect 290918 267588 290924 267600
rect 290976 267588 290982 267640
rect 298278 267588 298284 267640
rect 298336 267628 298342 267640
rect 322290 267628 322296 267640
rect 298336 267600 322296 267628
rect 298336 267588 298342 267600
rect 322290 267588 322296 267600
rect 322348 267588 322354 267640
rect 323670 267588 323676 267640
rect 323728 267628 323734 267640
rect 331122 267628 331128 267640
rect 323728 267600 331128 267628
rect 323728 267588 323734 267600
rect 331122 267588 331128 267600
rect 331180 267588 331186 267640
rect 347314 267588 347320 267640
rect 347372 267628 347378 267640
rect 476298 267628 476304 267640
rect 347372 267600 476304 267628
rect 347372 267588 347378 267600
rect 476298 267588 476304 267600
rect 476356 267588 476362 267640
rect 124214 267520 124220 267572
rect 124272 267560 124278 267572
rect 196342 267560 196348 267572
rect 124272 267532 196348 267560
rect 124272 267520 124278 267532
rect 196342 267520 196348 267532
rect 196400 267520 196406 267572
rect 196710 267520 196716 267572
rect 196768 267560 196774 267572
rect 216398 267560 216404 267572
rect 196768 267532 216404 267560
rect 196768 267520 196774 267532
rect 216398 267520 216404 267532
rect 216456 267520 216462 267572
rect 284478 267520 284484 267572
rect 284536 267560 284542 267572
rect 291470 267560 291476 267572
rect 284536 267532 291476 267560
rect 284536 267520 284542 267532
rect 291470 267520 291476 267532
rect 291528 267520 291534 267572
rect 299658 267520 299664 267572
rect 299716 267560 299722 267572
rect 326338 267560 326344 267572
rect 299716 267532 326344 267560
rect 299716 267520 299722 267532
rect 326338 267520 326344 267532
rect 326396 267520 326402 267572
rect 330846 267520 330852 267572
rect 330904 267560 330910 267572
rect 350350 267560 350356 267572
rect 330904 267532 350356 267560
rect 330904 267520 330910 267532
rect 350350 267520 350356 267532
rect 350408 267520 350414 267572
rect 483382 267560 483388 267572
rect 350460 267532 483388 267560
rect 150342 267452 150348 267504
rect 150400 267492 150406 267504
rect 224402 267492 224408 267504
rect 150400 267464 224408 267492
rect 150400 267452 150406 267464
rect 224402 267452 224408 267464
rect 224460 267452 224466 267504
rect 236730 267452 236736 267504
rect 236788 267492 236794 267504
rect 244458 267492 244464 267504
rect 236788 267464 244464 267492
rect 236788 267452 236794 267464
rect 244458 267452 244464 267464
rect 244516 267452 244522 267504
rect 272058 267452 272064 267504
rect 272116 267492 272122 267504
rect 277394 267492 277400 267504
rect 272116 267464 277400 267492
rect 272116 267452 272122 267464
rect 277394 267452 277400 267464
rect 277452 267452 277458 267504
rect 288526 267452 288532 267504
rect 288584 267492 288590 267504
rect 301498 267492 301504 267504
rect 288584 267464 301504 267492
rect 288584 267452 288590 267464
rect 301498 267452 301504 267464
rect 301556 267452 301562 267504
rect 306374 267452 306380 267504
rect 306432 267492 306438 267504
rect 335354 267492 335360 267504
rect 306432 267464 335360 267492
rect 306432 267452 306438 267464
rect 335354 267452 335360 267464
rect 335412 267452 335418 267504
rect 349982 267452 349988 267504
rect 350040 267492 350046 267504
rect 350460 267492 350488 267532
rect 483382 267520 483388 267532
rect 483440 267520 483446 267572
rect 350040 267464 350488 267492
rect 350040 267452 350046 267464
rect 352650 267452 352656 267504
rect 352708 267492 352714 267504
rect 491386 267492 491392 267504
rect 352708 267464 491392 267492
rect 352708 267452 352714 267464
rect 491386 267452 491392 267464
rect 491444 267452 491450 267504
rect 139302 267384 139308 267436
rect 139360 267424 139366 267436
rect 220354 267424 220360 267436
rect 139360 267396 220360 267424
rect 139360 267384 139366 267396
rect 220354 267384 220360 267396
rect 220412 267384 220418 267436
rect 288066 267384 288072 267436
rect 288124 267424 288130 267436
rect 300118 267424 300124 267436
rect 288124 267396 300124 267424
rect 288124 267384 288130 267396
rect 300118 267384 300124 267396
rect 300176 267384 300182 267436
rect 304994 267384 305000 267436
rect 305052 267424 305058 267436
rect 335998 267424 336004 267436
rect 305052 267396 336004 267424
rect 305052 267384 305058 267396
rect 335998 267384 336004 267396
rect 336056 267384 336062 267436
rect 339310 267384 339316 267436
rect 339368 267424 339374 267436
rect 339368 267396 345014 267424
rect 339368 267384 339374 267396
rect 116486 267316 116492 267368
rect 116544 267356 116550 267368
rect 199930 267356 199936 267368
rect 116544 267328 199936 267356
rect 116544 267316 116550 267328
rect 199930 267316 199936 267328
rect 199988 267316 199994 267368
rect 200086 267328 200896 267356
rect 132402 267248 132408 267300
rect 132460 267288 132466 267300
rect 200086 267288 200114 267328
rect 132460 267260 200114 267288
rect 200868 267288 200896 267328
rect 227622 267316 227628 267368
rect 227680 267356 227686 267368
rect 237282 267356 237288 267368
rect 227680 267328 237288 267356
rect 227680 267316 227686 267328
rect 237282 267316 237288 267328
rect 237340 267316 237346 267368
rect 289446 267316 289452 267368
rect 289504 267356 289510 267368
rect 304258 267356 304264 267368
rect 289504 267328 304264 267356
rect 289504 267316 289510 267328
rect 304258 267316 304264 267328
rect 304316 267316 304322 267368
rect 308582 267316 308588 267368
rect 308640 267356 308646 267368
rect 344278 267356 344284 267368
rect 308640 267328 344284 267356
rect 308640 267316 308646 267328
rect 344278 267316 344284 267328
rect 344336 267316 344342 267368
rect 344986 267356 345014 267396
rect 355318 267384 355324 267436
rect 355376 267424 355382 267436
rect 498194 267424 498200 267436
rect 355376 267396 498200 267424
rect 355376 267384 355382 267396
rect 498194 267384 498200 267396
rect 498252 267384 498258 267436
rect 346394 267356 346400 267368
rect 344986 267328 346400 267356
rect 346394 267316 346400 267328
rect 346452 267316 346458 267368
rect 346854 267316 346860 267368
rect 346912 267356 346918 267368
rect 347682 267356 347688 267368
rect 346912 267328 347688 267356
rect 346912 267316 346918 267328
rect 347682 267316 347688 267328
rect 347740 267316 347746 267368
rect 348234 267316 348240 267368
rect 348292 267356 348298 267368
rect 348970 267356 348976 267368
rect 348292 267328 348976 267356
rect 348292 267316 348298 267328
rect 348970 267316 348976 267328
rect 349028 267316 349034 267368
rect 349522 267316 349528 267368
rect 349580 267356 349586 267368
rect 350442 267356 350448 267368
rect 349580 267328 350448 267356
rect 349580 267316 349586 267328
rect 350442 267316 350448 267328
rect 350500 267316 350506 267368
rect 350902 267316 350908 267368
rect 350960 267356 350966 267368
rect 351730 267356 351736 267368
rect 350960 267328 351736 267356
rect 350960 267316 350966 267328
rect 351730 267316 351736 267328
rect 351788 267316 351794 267368
rect 352190 267316 352196 267368
rect 352248 267356 352254 267368
rect 353202 267356 353208 267368
rect 352248 267328 353208 267356
rect 352248 267316 352254 267328
rect 353202 267316 353208 267328
rect 353260 267316 353266 267368
rect 353570 267316 353576 267368
rect 353628 267356 353634 267368
rect 354398 267356 354404 267368
rect 353628 267328 354404 267356
rect 353628 267316 353634 267328
rect 354398 267316 354404 267328
rect 354456 267316 354462 267368
rect 360654 267316 360660 267368
rect 360712 267356 360718 267368
rect 511994 267356 512000 267368
rect 360712 267328 512000 267356
rect 360712 267316 360718 267328
rect 511994 267316 512000 267328
rect 512052 267316 512058 267368
rect 217686 267288 217692 267300
rect 200868 267260 217692 267288
rect 132460 267248 132466 267260
rect 217686 267248 217692 267260
rect 217744 267248 217750 267300
rect 225598 267248 225604 267300
rect 225656 267288 225662 267300
rect 235994 267288 236000 267300
rect 225656 267260 236000 267288
rect 225656 267248 225662 267260
rect 235994 267248 236000 267260
rect 236052 267248 236058 267300
rect 236638 267248 236644 267300
rect 236696 267288 236702 267300
rect 251082 267288 251088 267300
rect 236696 267260 251088 267288
rect 236696 267248 236702 267260
rect 251082 267248 251088 267260
rect 251140 267248 251146 267300
rect 276934 267248 276940 267300
rect 276992 267288 276998 267300
rect 282730 267288 282736 267300
rect 276992 267260 282736 267288
rect 276992 267248 276998 267260
rect 282730 267248 282736 267260
rect 282788 267248 282794 267300
rect 290734 267248 290740 267300
rect 290792 267288 290798 267300
rect 307754 267288 307760 267300
rect 290792 267260 307760 267288
rect 290792 267248 290798 267260
rect 307754 267248 307760 267260
rect 307812 267248 307818 267300
rect 311250 267248 311256 267300
rect 311308 267288 311314 267300
rect 361482 267288 361488 267300
rect 311308 267260 361488 267288
rect 311308 267248 311314 267260
rect 361482 267248 361488 267260
rect 361540 267248 361546 267300
rect 362954 267288 362960 267300
rect 361592 267260 362960 267288
rect 106918 267180 106924 267232
rect 106976 267220 106982 267232
rect 200758 267220 200764 267232
rect 106976 267192 200764 267220
rect 106976 267180 106982 267192
rect 200758 267180 200764 267192
rect 200816 267180 200822 267232
rect 200850 267180 200856 267232
rect 200908 267220 200914 267232
rect 200908 267192 209774 267220
rect 200908 267180 200914 267192
rect 100018 267112 100024 267164
rect 100076 267152 100082 267164
rect 204346 267152 204352 267164
rect 100076 267124 204352 267152
rect 100076 267112 100082 267124
rect 204346 267112 204352 267124
rect 204404 267112 204410 267164
rect 90358 267044 90364 267096
rect 90416 267084 90422 267096
rect 201218 267084 201224 267096
rect 90416 267056 201224 267084
rect 90416 267044 90422 267056
rect 201218 267044 201224 267056
rect 201276 267044 201282 267096
rect 209746 267084 209774 267192
rect 217318 267180 217324 267232
rect 217376 267220 217382 267232
rect 237742 267220 237748 267232
rect 217376 267192 237748 267220
rect 217376 267180 217382 267192
rect 237742 267180 237748 267192
rect 237800 267180 237806 267232
rect 238018 267180 238024 267232
rect 238076 267220 238082 267232
rect 241790 267220 241796 267232
rect 238076 267192 241796 267220
rect 238076 267180 238082 267192
rect 241790 267180 241796 267192
rect 241848 267180 241854 267232
rect 245286 267180 245292 267232
rect 245344 267220 245350 267232
rect 252462 267220 252468 267232
rect 245344 267192 252468 267220
rect 245344 267180 245350 267192
rect 252462 267180 252468 267192
rect 252520 267180 252526 267232
rect 256602 267180 256608 267232
rect 256660 267220 256666 267232
rect 264054 267220 264060 267232
rect 256660 267192 264060 267220
rect 256660 267180 256666 267192
rect 264054 267180 264060 267192
rect 264112 267180 264118 267232
rect 288986 267180 288992 267232
rect 289044 267220 289050 267232
rect 309778 267220 309784 267232
rect 289044 267192 309784 267220
rect 289044 267180 289050 267192
rect 309778 267180 309784 267192
rect 309836 267180 309842 267232
rect 312538 267180 312544 267232
rect 312596 267220 312602 267232
rect 361592 267220 361620 267260
rect 362954 267248 362960 267260
rect 363012 267248 363018 267300
rect 363322 267248 363328 267300
rect 363380 267288 363386 267300
rect 516134 267288 516140 267300
rect 363380 267260 516140 267288
rect 363380 267248 363386 267260
rect 516134 267248 516140 267260
rect 516192 267248 516198 267300
rect 312596 267192 361620 267220
rect 312596 267180 312602 267192
rect 361850 267180 361856 267232
rect 361908 267220 361914 267232
rect 362678 267220 362684 267232
rect 361908 267192 362684 267220
rect 361908 267180 361914 267192
rect 362678 267180 362684 267192
rect 362736 267180 362742 267232
rect 368014 267180 368020 267232
rect 368072 267220 368078 267232
rect 368072 267192 369808 267220
rect 368072 267180 368078 267192
rect 233142 267112 233148 267164
rect 233200 267152 233206 267164
rect 255130 267152 255136 267164
rect 233200 267124 255136 267152
rect 233200 267112 233206 267124
rect 255130 267112 255136 267124
rect 255188 267112 255194 267164
rect 255222 267112 255228 267164
rect 255280 267152 255286 267164
rect 263594 267152 263600 267164
rect 255280 267124 263600 267152
rect 255280 267112 255286 267124
rect 263594 267112 263600 267124
rect 263652 267112 263658 267164
rect 286318 267112 286324 267164
rect 286376 267152 286382 267164
rect 307018 267152 307024 267164
rect 286376 267124 307024 267152
rect 286376 267112 286382 267124
rect 307018 267112 307024 267124
rect 307076 267112 307082 267164
rect 315206 267112 315212 267164
rect 315264 267152 315270 267164
rect 369670 267152 369676 267164
rect 315264 267124 369676 267152
rect 315264 267112 315270 267124
rect 369670 267112 369676 267124
rect 369728 267112 369734 267164
rect 369780 267152 369808 267192
rect 371326 267180 371332 267232
rect 371384 267220 371390 267232
rect 371384 267192 373994 267220
rect 371384 267180 371390 267192
rect 371878 267152 371884 267164
rect 369780 267124 371884 267152
rect 371878 267112 371884 267124
rect 371936 267112 371942 267164
rect 373966 267152 373994 267192
rect 378778 267180 378784 267232
rect 378836 267220 378842 267232
rect 523678 267220 523684 267232
rect 378836 267192 523684 267220
rect 378836 267180 378842 267192
rect 523678 267180 523684 267192
rect 523736 267180 523742 267232
rect 540974 267152 540980 267164
rect 373966 267124 540980 267152
rect 540974 267112 540980 267124
rect 541032 267112 541038 267164
rect 211062 267084 211068 267096
rect 209746 267056 211068 267084
rect 211062 267044 211068 267056
rect 211120 267044 211126 267096
rect 213178 267044 213184 267096
rect 213236 267084 213242 267096
rect 213236 267056 213868 267084
rect 213236 267044 213242 267056
rect 73798 266976 73804 267028
rect 73856 267016 73862 267028
rect 194134 267016 194140 267028
rect 73856 266988 194140 267016
rect 73856 266976 73862 266988
rect 194134 266976 194140 266988
rect 194192 266976 194198 267028
rect 202414 266976 202420 267028
rect 202472 267016 202478 267028
rect 213730 267016 213736 267028
rect 202472 266988 213736 267016
rect 202472 266976 202478 266988
rect 213730 266976 213736 266988
rect 213788 266976 213794 267028
rect 213840 267016 213868 267056
rect 215846 267044 215852 267096
rect 215904 267084 215910 267096
rect 239122 267084 239128 267096
rect 215904 267056 239128 267084
rect 215904 267044 215910 267056
rect 239122 267044 239128 267056
rect 239180 267044 239186 267096
rect 239306 267044 239312 267096
rect 239364 267084 239370 267096
rect 249794 267084 249800 267096
rect 239364 267056 249800 267084
rect 239364 267044 239370 267056
rect 249794 267044 249800 267056
rect 249852 267044 249858 267096
rect 252370 267044 252376 267096
rect 252428 267084 252434 267096
rect 262214 267084 262220 267096
rect 252428 267056 262220 267084
rect 252428 267044 252434 267056
rect 262214 267044 262220 267056
rect 262272 267044 262278 267096
rect 292574 267044 292580 267096
rect 292632 267084 292638 267096
rect 316678 267084 316684 267096
rect 292632 267056 316684 267084
rect 292632 267044 292638 267056
rect 316678 267044 316684 267056
rect 316736 267044 316742 267096
rect 317874 267044 317880 267096
rect 317932 267084 317938 267096
rect 387058 267084 387064 267096
rect 317932 267056 387064 267084
rect 317932 267044 317938 267056
rect 387058 267044 387064 267056
rect 387116 267044 387122 267096
rect 398806 267056 401640 267084
rect 236454 267016 236460 267028
rect 213840 266988 236460 267016
rect 236454 266976 236460 266988
rect 236512 266976 236518 267028
rect 238662 266976 238668 267028
rect 238720 267016 238726 267028
rect 257338 267016 257344 267028
rect 238720 266988 257344 267016
rect 238720 266976 238726 266988
rect 257338 266976 257344 266988
rect 257396 266976 257402 267028
rect 257982 266976 257988 267028
rect 258040 267016 258046 267028
rect 264514 267016 264520 267028
rect 258040 266988 264520 267016
rect 258040 266976 258046 266988
rect 264514 266976 264520 266988
rect 264572 266976 264578 267028
rect 278314 266976 278320 267028
rect 278372 267016 278378 267028
rect 287790 267016 287796 267028
rect 278372 266988 287796 267016
rect 278372 266976 278378 266988
rect 287790 266976 287796 266988
rect 287848 266976 287854 267028
rect 295242 266976 295248 267028
rect 295300 267016 295306 267028
rect 319438 267016 319444 267028
rect 295300 266988 319444 267016
rect 295300 266976 295306 266988
rect 319438 266976 319444 266988
rect 319496 266976 319502 267028
rect 320542 266976 320548 267028
rect 320600 267016 320606 267028
rect 398806 267016 398834 267056
rect 320600 266988 398834 267016
rect 320600 266976 320606 266988
rect 400766 266976 400772 267028
rect 400824 267016 400830 267028
rect 401502 267016 401508 267028
rect 400824 266988 401508 267016
rect 400824 266976 400830 266988
rect 401502 266976 401508 266988
rect 401560 266976 401566 267028
rect 401612 267016 401640 267056
rect 402054 267044 402060 267096
rect 402112 267084 402118 267096
rect 402882 267084 402888 267096
rect 402112 267056 402888 267084
rect 402112 267044 402118 267056
rect 402882 267044 402888 267056
rect 402940 267044 402946 267096
rect 404722 267044 404728 267096
rect 404780 267084 404786 267096
rect 405642 267084 405648 267096
rect 404780 267056 405648 267084
rect 404780 267044 404786 267056
rect 405642 267044 405648 267056
rect 405700 267044 405706 267096
rect 410518 267044 410524 267096
rect 410576 267084 410582 267096
rect 414750 267084 414756 267096
rect 410576 267056 414756 267084
rect 410576 267044 410582 267056
rect 414750 267044 414756 267056
rect 414808 267044 414814 267096
rect 632238 267084 632244 267096
rect 414860 267056 632244 267084
rect 405918 267016 405924 267028
rect 401612 266988 405924 267016
rect 405918 266976 405924 266988
rect 405976 266976 405982 267028
rect 406102 266976 406108 267028
rect 406160 267016 406166 267028
rect 414860 267016 414888 267056
rect 632238 267044 632244 267056
rect 632296 267044 632302 267096
rect 406160 266988 414888 267016
rect 406160 266976 406166 266988
rect 414934 266976 414940 267028
rect 414992 267016 414998 267028
rect 644474 267016 644480 267028
rect 414992 266988 644480 267016
rect 414992 266976 414998 266988
rect 644474 266976 644480 266988
rect 644532 266976 644538 267028
rect 164142 266908 164148 266960
rect 164200 266948 164206 266960
rect 312446 266948 312452 266960
rect 164200 266920 224356 266948
rect 164200 266908 164206 266920
rect 170950 266840 170956 266892
rect 171008 266880 171014 266892
rect 171008 266852 224172 266880
rect 171008 266840 171014 266852
rect 177574 266772 177580 266824
rect 177632 266812 177638 266824
rect 223022 266812 223028 266824
rect 177632 266784 223028 266812
rect 177632 266772 177638 266784
rect 223022 266772 223028 266784
rect 223080 266772 223086 266824
rect 164878 266704 164884 266756
rect 164936 266744 164942 266756
rect 199470 266744 199476 266756
rect 164936 266716 199476 266744
rect 164936 266704 164942 266716
rect 199470 266704 199476 266716
rect 199528 266704 199534 266756
rect 200758 266704 200764 266756
rect 200816 266744 200822 266756
rect 207014 266744 207020 266756
rect 200816 266716 207020 266744
rect 200816 266704 200822 266716
rect 207014 266704 207020 266716
rect 207072 266704 207078 266756
rect 224144 266744 224172 266852
rect 224328 266812 224356 266920
rect 296686 266920 312452 266948
rect 272518 266840 272524 266892
rect 272576 266880 272582 266892
rect 277762 266880 277768 266892
rect 272576 266852 277768 266880
rect 272576 266840 272582 266852
rect 277762 266840 277768 266852
rect 277820 266840 277826 266892
rect 294322 266840 294328 266892
rect 294380 266880 294386 266892
rect 296686 266880 296714 266920
rect 312446 266908 312452 266920
rect 312504 266908 312510 266960
rect 321002 266908 321008 266960
rect 321060 266948 321066 266960
rect 342162 266948 342168 266960
rect 321060 266920 342168 266948
rect 321060 266908 321066 266920
rect 342162 266908 342168 266920
rect 342220 266908 342226 266960
rect 345474 266908 345480 266960
rect 345532 266948 345538 266960
rect 346210 266948 346216 266960
rect 345532 266920 346216 266948
rect 345532 266908 345538 266920
rect 346210 266908 346216 266920
rect 346268 266908 346274 266960
rect 464706 266948 464712 266960
rect 346320 266920 464712 266948
rect 311158 266880 311164 266892
rect 294380 266852 296714 266880
rect 308784 266852 311164 266880
rect 294380 266840 294386 266852
rect 229738 266812 229744 266824
rect 224328 266784 229744 266812
rect 229738 266772 229744 266784
rect 229796 266772 229802 266824
rect 308784 266812 308812 266852
rect 311158 266840 311164 266852
rect 311216 266840 311222 266892
rect 331306 266840 331312 266892
rect 331364 266880 331370 266892
rect 331364 266852 334204 266880
rect 331364 266840 331370 266852
rect 322198 266812 322204 266824
rect 296686 266784 308812 266812
rect 311176 266784 322204 266812
rect 232406 266744 232412 266756
rect 224144 266716 232412 266744
rect 232406 266704 232412 266716
rect 232464 266704 232470 266756
rect 292942 266704 292948 266756
rect 293000 266744 293006 266756
rect 296686 266744 296714 266784
rect 293000 266716 296714 266744
rect 293000 266704 293006 266716
rect 301866 266704 301872 266756
rect 301924 266744 301930 266756
rect 311176 266744 311204 266784
rect 322198 266772 322204 266784
rect 322256 266772 322262 266824
rect 325970 266772 325976 266824
rect 326028 266812 326034 266824
rect 334066 266812 334072 266824
rect 326028 266784 334072 266812
rect 326028 266772 326034 266784
rect 334066 266772 334072 266784
rect 334124 266772 334130 266824
rect 301924 266716 311204 266744
rect 301924 266704 301930 266716
rect 328638 266704 328644 266756
rect 328696 266744 328702 266756
rect 328696 266716 333928 266744
rect 328696 266704 328702 266716
rect 282270 266636 282276 266688
rect 282328 266676 282334 266688
rect 287698 266676 287704 266688
rect 282328 266648 287704 266676
rect 282328 266636 282334 266648
rect 287698 266636 287704 266648
rect 287756 266636 287762 266688
rect 309870 266636 309876 266688
rect 309928 266676 309934 266688
rect 323578 266676 323584 266688
rect 309928 266648 323584 266676
rect 309928 266636 309934 266648
rect 323578 266636 323584 266648
rect 323636 266636 323642 266688
rect 196618 266568 196624 266620
rect 196676 266608 196682 266620
rect 202414 266608 202420 266620
rect 196676 266580 202420 266608
rect 196676 266568 196682 266580
rect 202414 266568 202420 266580
rect 202472 266568 202478 266620
rect 271598 266568 271604 266620
rect 271656 266608 271662 266620
rect 276290 266608 276296 266620
rect 271656 266580 276296 266608
rect 271656 266568 271662 266580
rect 276290 266568 276296 266580
rect 276348 266568 276354 266620
rect 277394 266568 277400 266620
rect 277452 266608 277458 266620
rect 280522 266608 280528 266620
rect 277452 266580 280528 266608
rect 277452 266568 277458 266580
rect 280522 266568 280528 266580
rect 280580 266568 280586 266620
rect 280982 266568 280988 266620
rect 281040 266608 281046 266620
rect 289170 266608 289176 266620
rect 281040 266580 289176 266608
rect 281040 266568 281046 266580
rect 289170 266568 289176 266580
rect 289228 266568 289234 266620
rect 328178 266568 328184 266620
rect 328236 266608 328242 266620
rect 329098 266608 329104 266620
rect 328236 266580 329104 266608
rect 328236 266568 328242 266580
rect 329098 266568 329104 266580
rect 329156 266568 329162 266620
rect 332594 266568 332600 266620
rect 332652 266608 332658 266620
rect 333790 266608 333796 266620
rect 332652 266580 333796 266608
rect 332652 266568 332658 266580
rect 333790 266568 333796 266580
rect 333848 266568 333854 266620
rect 333900 266608 333928 266716
rect 334176 266676 334204 266852
rect 336642 266840 336648 266892
rect 336700 266880 336706 266892
rect 336700 266852 343588 266880
rect 336700 266840 336706 266852
rect 334802 266772 334808 266824
rect 334860 266812 334866 266824
rect 335262 266812 335268 266824
rect 334860 266784 335268 266812
rect 334860 266772 334866 266784
rect 335262 266772 335268 266784
rect 335320 266772 335326 266824
rect 337470 266772 337476 266824
rect 337528 266812 337534 266824
rect 337930 266812 337936 266824
rect 337528 266784 337936 266812
rect 337528 266772 337534 266784
rect 337930 266772 337936 266784
rect 337988 266772 337994 266824
rect 340138 266772 340144 266824
rect 340196 266812 340202 266824
rect 340690 266812 340696 266824
rect 340196 266784 340696 266812
rect 340196 266772 340202 266784
rect 340690 266772 340696 266784
rect 340748 266772 340754 266824
rect 342806 266772 342812 266824
rect 342864 266812 342870 266824
rect 343450 266812 343456 266824
rect 342864 266784 343456 266812
rect 342864 266772 342870 266784
rect 343450 266772 343456 266784
rect 343508 266772 343514 266824
rect 343560 266812 343588 266852
rect 344646 266840 344652 266892
rect 344704 266880 344710 266892
rect 346320 266880 346348 266920
rect 464706 266908 464712 266920
rect 464764 266908 464770 266960
rect 344704 266852 346348 266880
rect 344704 266840 344710 266852
rect 346394 266840 346400 266892
rect 346452 266880 346458 266892
rect 455414 266880 455420 266892
rect 346452 266852 455420 266880
rect 346452 266840 346458 266852
rect 455414 266840 455420 266852
rect 455472 266840 455478 266892
rect 674742 266840 674748 266892
rect 674800 266880 674806 266892
rect 676214 266880 676220 266892
rect 674800 266852 676220 266880
rect 674800 266840 674806 266852
rect 676214 266840 676220 266852
rect 676272 266840 676278 266892
rect 448514 266812 448520 266824
rect 343560 266784 448520 266812
rect 448514 266772 448520 266784
rect 448572 266772 448578 266824
rect 334250 266704 334256 266756
rect 334308 266744 334314 266756
rect 435358 266744 435364 266756
rect 334308 266716 435364 266744
rect 334308 266704 334314 266716
rect 435358 266704 435364 266716
rect 435416 266704 435422 266756
rect 420178 266676 420184 266688
rect 334176 266648 420184 266676
rect 420178 266636 420184 266648
rect 420236 266636 420242 266688
rect 674650 266636 674656 266688
rect 674708 266676 674714 266688
rect 676030 266676 676036 266688
rect 674708 266648 676036 266676
rect 674708 266636 674714 266648
rect 676030 266636 676036 266648
rect 676088 266636 676094 266688
rect 414014 266608 414020 266620
rect 333900 266580 414020 266608
rect 414014 266568 414020 266580
rect 414072 266568 414078 266620
rect 271138 266500 271144 266552
rect 271196 266540 271202 266552
rect 274634 266540 274640 266552
rect 271196 266512 274640 266540
rect 271196 266500 271202 266512
rect 274634 266500 274640 266512
rect 274692 266500 274698 266552
rect 275186 266500 275192 266552
rect 275244 266540 275250 266552
rect 279418 266540 279424 266552
rect 275244 266512 279424 266540
rect 275244 266500 275250 266512
rect 279418 266500 279424 266512
rect 279476 266500 279482 266552
rect 319254 266500 319260 266552
rect 319312 266540 319318 266552
rect 324958 266540 324964 266552
rect 319312 266512 324964 266540
rect 319312 266500 319318 266512
rect 324958 266500 324964 266512
rect 325016 266500 325022 266552
rect 326338 266500 326344 266552
rect 326396 266540 326402 266552
rect 326982 266540 326988 266552
rect 326396 266512 326988 266540
rect 326396 266500 326402 266512
rect 326982 266500 326988 266512
rect 327040 266500 327046 266552
rect 327258 266500 327264 266552
rect 327316 266540 327322 266552
rect 328362 266540 328368 266552
rect 327316 266512 328368 266540
rect 327316 266500 327322 266512
rect 328362 266500 328368 266512
rect 328420 266500 328426 266552
rect 329006 266500 329012 266552
rect 329064 266540 329070 266552
rect 329742 266540 329748 266552
rect 329064 266512 329748 266540
rect 329064 266500 329070 266512
rect 329742 266500 329748 266512
rect 329800 266500 329806 266552
rect 329926 266500 329932 266552
rect 329984 266540 329990 266552
rect 330662 266540 330668 266552
rect 329984 266512 330668 266540
rect 329984 266500 329990 266512
rect 330662 266500 330668 266512
rect 330720 266500 330726 266552
rect 333054 266500 333060 266552
rect 333112 266540 333118 266552
rect 333882 266540 333888 266552
rect 333112 266512 333888 266540
rect 333112 266500 333118 266512
rect 333882 266500 333888 266512
rect 333940 266500 333946 266552
rect 334066 266500 334072 266552
rect 334124 266540 334130 266552
rect 409138 266540 409144 266552
rect 334124 266512 409144 266540
rect 334124 266500 334130 266512
rect 409138 266500 409144 266512
rect 409196 266500 409202 266552
rect 191098 266432 191104 266484
rect 191156 266472 191162 266484
rect 197722 266472 197728 266484
rect 191156 266444 197728 266472
rect 191156 266432 191162 266444
rect 197722 266432 197728 266444
rect 197780 266432 197786 266484
rect 230474 266432 230480 266484
rect 230532 266472 230538 266484
rect 238662 266472 238668 266484
rect 230532 266444 238668 266472
rect 230532 266432 230538 266444
rect 238662 266432 238668 266444
rect 238720 266432 238726 266484
rect 270678 266432 270684 266484
rect 270736 266472 270742 266484
rect 273254 266472 273260 266484
rect 270736 266444 273260 266472
rect 270736 266432 270742 266444
rect 273254 266432 273260 266444
rect 273312 266432 273318 266484
rect 280062 266432 280068 266484
rect 280120 266472 280126 266484
rect 284846 266472 284852 266484
rect 280120 266444 284852 266472
rect 280120 266432 280126 266444
rect 284846 266432 284852 266444
rect 284904 266432 284910 266484
rect 287606 266432 287612 266484
rect 287664 266472 287670 266484
rect 289078 266472 289084 266484
rect 287664 266444 289084 266472
rect 287664 266432 287670 266444
rect 289078 266432 289084 266444
rect 289136 266432 289142 266484
rect 289814 266432 289820 266484
rect 289872 266472 289878 266484
rect 291010 266472 291016 266484
rect 289872 266444 291016 266472
rect 289872 266432 289878 266444
rect 291010 266432 291016 266444
rect 291068 266432 291074 266484
rect 291654 266432 291660 266484
rect 291712 266472 291718 266484
rect 295978 266472 295984 266484
rect 291712 266444 295984 266472
rect 291712 266432 291718 266444
rect 295978 266432 295984 266444
rect 296036 266432 296042 266484
rect 302786 266432 302792 266484
rect 302844 266472 302850 266484
rect 306006 266472 306012 266484
rect 302844 266444 306012 266472
rect 302844 266432 302850 266444
rect 306006 266432 306012 266444
rect 306064 266432 306070 266484
rect 312078 266432 312084 266484
rect 312136 266472 312142 266484
rect 315298 266472 315304 266484
rect 312136 266444 315304 266472
rect 312136 266432 312142 266444
rect 315298 266432 315304 266444
rect 315356 266432 315362 266484
rect 316586 266432 316592 266484
rect 316644 266472 316650 266484
rect 368014 266472 368020 266484
rect 316644 266444 368020 266472
rect 316644 266432 316650 266444
rect 368014 266432 368020 266444
rect 368072 266432 368078 266484
rect 368658 266432 368664 266484
rect 368716 266472 368722 266484
rect 378778 266472 378784 266484
rect 368716 266444 378784 266472
rect 368716 266432 368722 266444
rect 378778 266432 378784 266444
rect 378836 266432 378842 266484
rect 387794 266432 387800 266484
rect 387852 266472 387858 266484
rect 387852 266444 393314 266472
rect 387852 266432 387858 266444
rect 193858 266364 193864 266416
rect 193916 266404 193922 266416
rect 194594 266404 194600 266416
rect 193916 266376 194600 266404
rect 193916 266364 193922 266376
rect 194594 266364 194600 266376
rect 194652 266364 194658 266416
rect 235258 266364 235264 266416
rect 235316 266404 235322 266416
rect 238202 266404 238208 266416
rect 235316 266376 238208 266404
rect 235316 266364 235322 266376
rect 238202 266364 238208 266376
rect 238260 266364 238266 266416
rect 242158 266364 242164 266416
rect 242216 266404 242222 266416
rect 243078 266404 243084 266416
rect 242216 266376 243084 266404
rect 242216 266364 242222 266376
rect 243078 266364 243084 266376
rect 243136 266364 243142 266416
rect 244182 266364 244188 266416
rect 244240 266404 244246 266416
rect 248414 266404 248420 266416
rect 244240 266376 248420 266404
rect 244240 266364 244246 266376
rect 248414 266364 248420 266376
rect 248472 266364 248478 266416
rect 270310 266364 270316 266416
rect 270368 266404 270374 266416
rect 272150 266404 272156 266416
rect 270368 266376 272156 266404
rect 270368 266364 270374 266376
rect 272150 266364 272156 266376
rect 272208 266364 272214 266416
rect 276474 266364 276480 266416
rect 276532 266404 276538 266416
rect 277302 266404 277308 266416
rect 276532 266376 277308 266404
rect 276532 266364 276538 266376
rect 277302 266364 277308 266376
rect 277360 266364 277366 266416
rect 280522 266364 280528 266416
rect 280580 266404 280586 266416
rect 281350 266404 281356 266416
rect 280580 266376 281356 266404
rect 280580 266364 280586 266376
rect 281350 266364 281356 266376
rect 281408 266364 281414 266416
rect 281810 266364 281816 266416
rect 281868 266404 281874 266416
rect 283006 266404 283012 266416
rect 281868 266376 283012 266404
rect 281868 266364 281874 266376
rect 283006 266364 283012 266376
rect 283064 266364 283070 266416
rect 284110 266364 284116 266416
rect 284168 266404 284174 266416
rect 286778 266404 286784 266416
rect 284168 266376 286784 266404
rect 284168 266364 284174 266376
rect 286778 266364 286784 266376
rect 286836 266364 286842 266416
rect 287146 266364 287152 266416
rect 287204 266404 287210 266416
rect 288342 266404 288348 266416
rect 287204 266376 288348 266404
rect 287204 266364 287210 266376
rect 288342 266364 288348 266376
rect 288400 266364 288406 266416
rect 290274 266364 290280 266416
rect 290332 266404 290338 266416
rect 291102 266404 291108 266416
rect 290332 266376 291108 266404
rect 290332 266364 290338 266376
rect 291102 266364 291108 266376
rect 291160 266364 291166 266416
rect 291194 266364 291200 266416
rect 291252 266404 291258 266416
rect 292482 266404 292488 266416
rect 291252 266376 292488 266404
rect 291252 266364 291258 266376
rect 292482 266364 292488 266376
rect 292540 266364 292546 266416
rect 295610 266364 295616 266416
rect 295668 266404 295674 266416
rect 296530 266404 296536 266416
rect 295668 266376 296536 266404
rect 295668 266364 295674 266376
rect 296530 266364 296536 266376
rect 296588 266364 296594 266416
rect 296990 266364 296996 266416
rect 297048 266404 297054 266416
rect 297818 266404 297824 266416
rect 297048 266376 297824 266404
rect 297048 266364 297054 266376
rect 297818 266364 297824 266376
rect 297876 266364 297882 266416
rect 300946 266364 300952 266416
rect 301004 266404 301010 266416
rect 302142 266404 302148 266416
rect 301004 266376 302148 266404
rect 301004 266364 301010 266376
rect 302142 266364 302148 266376
rect 302200 266364 302206 266416
rect 304074 266364 304080 266416
rect 304132 266404 304138 266416
rect 304810 266404 304816 266416
rect 304132 266376 304816 266404
rect 304132 266364 304138 266376
rect 304810 266364 304816 266376
rect 304868 266364 304874 266416
rect 305454 266364 305460 266416
rect 305512 266404 305518 266416
rect 306282 266404 306288 266416
rect 305512 266376 306288 266404
rect 305512 266364 305518 266376
rect 306282 266364 306288 266376
rect 306340 266364 306346 266416
rect 306742 266364 306748 266416
rect 306800 266404 306806 266416
rect 307570 266404 307576 266416
rect 306800 266376 307576 266404
rect 306800 266364 306806 266376
rect 307570 266364 307576 266376
rect 307628 266364 307634 266416
rect 308122 266364 308128 266416
rect 308180 266404 308186 266416
rect 308950 266404 308956 266416
rect 308180 266376 308956 266404
rect 308180 266364 308186 266376
rect 308950 266364 308956 266376
rect 309008 266364 309014 266416
rect 309410 266364 309416 266416
rect 309468 266404 309474 266416
rect 310330 266404 310336 266416
rect 309468 266376 310336 266404
rect 309468 266364 309474 266376
rect 310330 266364 310336 266376
rect 310388 266364 310394 266416
rect 310790 266364 310796 266416
rect 310848 266404 310854 266416
rect 311710 266404 311716 266416
rect 310848 266376 311716 266404
rect 310848 266364 310854 266376
rect 311710 266364 311716 266376
rect 311768 266364 311774 266416
rect 313458 266364 313464 266416
rect 313516 266404 313522 266416
rect 314470 266404 314476 266416
rect 313516 266376 314476 266404
rect 313516 266364 313522 266376
rect 314470 266364 314476 266376
rect 314528 266364 314534 266416
rect 314838 266364 314844 266416
rect 314896 266404 314902 266416
rect 315850 266404 315856 266416
rect 314896 266376 315856 266404
rect 314896 266364 314902 266376
rect 315850 266364 315856 266376
rect 315908 266364 315914 266416
rect 316126 266364 316132 266416
rect 316184 266404 316190 266416
rect 317230 266404 317236 266416
rect 316184 266376 317236 266404
rect 316184 266364 316190 266376
rect 317230 266364 317236 266376
rect 317288 266364 317294 266416
rect 317506 266364 317512 266416
rect 317564 266404 317570 266416
rect 318610 266404 318616 266416
rect 317564 266376 318616 266404
rect 317564 266364 317570 266376
rect 318610 266364 318616 266376
rect 318668 266364 318674 266416
rect 318794 266364 318800 266416
rect 318852 266404 318858 266416
rect 319990 266404 319996 266416
rect 318852 266376 319996 266404
rect 318852 266364 318858 266376
rect 319990 266364 319996 266376
rect 320048 266364 320054 266416
rect 320174 266364 320180 266416
rect 320232 266404 320238 266416
rect 321370 266404 321376 266416
rect 320232 266376 321376 266404
rect 320232 266364 320238 266376
rect 321370 266364 321376 266376
rect 321428 266364 321434 266416
rect 324590 266364 324596 266416
rect 324648 266404 324654 266416
rect 354674 266404 354680 266416
rect 324648 266376 354680 266404
rect 324648 266364 324654 266376
rect 354674 266364 354680 266376
rect 354732 266364 354738 266416
rect 354858 266364 354864 266416
rect 354916 266404 354922 266416
rect 355962 266404 355968 266416
rect 354916 266376 355968 266404
rect 354916 266364 354922 266376
rect 355962 266364 355968 266376
rect 356020 266364 356026 266416
rect 356238 266364 356244 266416
rect 356296 266404 356302 266416
rect 357158 266404 357164 266416
rect 356296 266376 357164 266404
rect 356296 266364 356302 266376
rect 357158 266364 357164 266376
rect 357216 266364 357222 266416
rect 358906 266364 358912 266416
rect 358964 266404 358970 266416
rect 359918 266404 359924 266416
rect 358964 266376 359924 266404
rect 358964 266364 358970 266376
rect 359918 266364 359924 266376
rect 359976 266364 359982 266416
rect 362402 266364 362408 266416
rect 362460 266404 362466 266416
rect 362862 266404 362868 266416
rect 362460 266376 362868 266404
rect 362460 266364 362466 266376
rect 362862 266364 362868 266376
rect 362920 266364 362926 266416
rect 364702 266364 364708 266416
rect 364760 266404 364766 266416
rect 365438 266404 365444 266416
rect 364760 266376 365444 266404
rect 364760 266364 364766 266376
rect 365438 266364 365444 266376
rect 365496 266364 365502 266416
rect 367370 266364 367376 266416
rect 367428 266404 367434 266416
rect 368382 266404 368388 266416
rect 367428 266376 368388 266404
rect 367428 266364 367434 266376
rect 368382 266364 368388 266376
rect 368440 266364 368446 266416
rect 370038 266364 370044 266416
rect 370096 266404 370102 266416
rect 371142 266404 371148 266416
rect 370096 266376 371148 266404
rect 370096 266364 370102 266376
rect 371142 266364 371148 266376
rect 371200 266364 371206 266416
rect 372706 266364 372712 266416
rect 372764 266404 372770 266416
rect 373902 266404 373908 266416
rect 372764 266376 373908 266404
rect 372764 266364 372770 266376
rect 373902 266364 373908 266376
rect 373960 266364 373966 266416
rect 376202 266364 376208 266416
rect 376260 266404 376266 266416
rect 376570 266404 376576 266416
rect 376260 266376 376576 266404
rect 376260 266364 376266 266376
rect 376570 266364 376576 266376
rect 376628 266364 376634 266416
rect 381170 266364 381176 266416
rect 381228 266404 381234 266416
rect 381998 266404 382004 266416
rect 381228 266376 382004 266404
rect 381228 266364 381234 266376
rect 381998 266364 382004 266376
rect 382056 266364 382062 266416
rect 383838 266364 383844 266416
rect 383896 266404 383902 266416
rect 384942 266404 384948 266416
rect 383896 266376 384948 266404
rect 383896 266364 383902 266376
rect 384942 266364 384948 266376
rect 385000 266364 385006 266416
rect 390922 266364 390928 266416
rect 390980 266404 390986 266416
rect 391750 266404 391756 266416
rect 390980 266376 391756 266404
rect 390980 266364 390986 266376
rect 391750 266364 391756 266376
rect 391808 266364 391814 266416
rect 393286 266404 393314 266444
rect 393590 266432 393596 266484
rect 393648 266472 393654 266484
rect 394510 266472 394516 266484
rect 393648 266444 394516 266472
rect 393648 266432 393654 266444
rect 394510 266432 394516 266444
rect 394568 266432 394574 266484
rect 394970 266432 394976 266484
rect 395028 266472 395034 266484
rect 395798 266472 395804 266484
rect 395028 266444 395804 266472
rect 395028 266432 395034 266444
rect 395798 266432 395804 266444
rect 395856 266432 395862 266484
rect 396258 266432 396264 266484
rect 396316 266472 396322 266484
rect 397270 266472 397276 266484
rect 396316 266444 397276 266472
rect 396316 266432 396322 266444
rect 397270 266432 397276 266444
rect 397328 266432 397334 266484
rect 408678 266472 408684 266484
rect 398806 266444 408684 266472
rect 398806 266404 398834 266444
rect 408678 266432 408684 266444
rect 408736 266432 408742 266484
rect 408770 266432 408776 266484
rect 408828 266472 408834 266484
rect 479518 266472 479524 266484
rect 408828 266444 479524 266472
rect 408828 266432 408834 266444
rect 479518 266432 479524 266444
rect 479576 266432 479582 266484
rect 393286 266376 398834 266404
rect 410058 266364 410064 266416
rect 410116 266404 410122 266416
rect 411070 266404 411076 266416
rect 410116 266376 411076 266404
rect 410116 266364 410122 266376
rect 411070 266364 411076 266376
rect 411128 266364 411134 266416
rect 355778 266296 355784 266348
rect 355836 266336 355842 266348
rect 499574 266336 499580 266348
rect 355836 266308 499580 266336
rect 355836 266296 355842 266308
rect 499574 266296 499580 266308
rect 499632 266296 499638 266348
rect 358446 266228 358452 266280
rect 358504 266268 358510 266280
rect 506474 266268 506480 266280
rect 358504 266240 506480 266268
rect 358504 266228 358510 266240
rect 506474 266228 506480 266240
rect 506532 266228 506538 266280
rect 361114 266160 361120 266212
rect 361172 266200 361178 266212
rect 513374 266200 513380 266212
rect 361172 266172 513380 266200
rect 361172 266160 361178 266172
rect 513374 266160 513380 266172
rect 513432 266160 513438 266212
rect 373166 266092 373172 266144
rect 373224 266132 373230 266144
rect 545114 266132 545120 266144
rect 373224 266104 545120 266132
rect 373224 266092 373230 266104
rect 545114 266092 545120 266104
rect 545172 266092 545178 266144
rect 374454 266024 374460 266076
rect 374512 266064 374518 266076
rect 549254 266064 549260 266076
rect 374512 266036 549260 266064
rect 374512 266024 374518 266036
rect 549254 266024 549260 266036
rect 549312 266024 549318 266076
rect 674650 266024 674656 266076
rect 674708 266064 674714 266076
rect 676214 266064 676220 266076
rect 674708 266036 676220 266064
rect 674708 266024 674714 266036
rect 676214 266024 676220 266036
rect 676272 266024 676278 266076
rect 375834 265956 375840 266008
rect 375892 265996 375898 266008
rect 552014 265996 552020 266008
rect 375892 265968 552020 265996
rect 375892 265956 375898 265968
rect 552014 265956 552020 265968
rect 552072 265956 552078 266008
rect 377122 265888 377128 265940
rect 377180 265928 377186 265940
rect 556154 265928 556160 265940
rect 377180 265900 556160 265928
rect 377180 265888 377186 265900
rect 556154 265888 556160 265900
rect 556212 265888 556218 265940
rect 378502 265820 378508 265872
rect 378560 265860 378566 265872
rect 558914 265860 558920 265872
rect 378560 265832 558920 265860
rect 378560 265820 378566 265832
rect 558914 265820 558920 265832
rect 558972 265820 558978 265872
rect 379790 265752 379796 265804
rect 379848 265792 379854 265804
rect 563054 265792 563060 265804
rect 379848 265764 563060 265792
rect 379848 265752 379854 265764
rect 563054 265752 563060 265764
rect 563112 265752 563118 265804
rect 382458 265684 382464 265736
rect 382516 265724 382522 265736
rect 569954 265724 569960 265736
rect 382516 265696 569960 265724
rect 382516 265684 382522 265696
rect 569954 265684 569960 265696
rect 570012 265684 570018 265736
rect 385586 265616 385592 265668
rect 385644 265656 385650 265668
rect 578234 265656 578240 265668
rect 385644 265628 578240 265656
rect 385644 265616 385650 265628
rect 578234 265616 578240 265628
rect 578292 265616 578298 265668
rect 194686 265548 194692 265600
rect 194744 265588 194750 265600
rect 195606 265588 195612 265600
rect 194744 265560 195612 265588
rect 194744 265548 194750 265560
rect 195606 265548 195612 265560
rect 195664 265548 195670 265600
rect 201586 265548 201592 265600
rect 201644 265588 201650 265600
rect 202230 265588 202236 265600
rect 201644 265560 202236 265588
rect 201644 265548 201650 265560
rect 202230 265548 202236 265560
rect 202288 265548 202294 265600
rect 223666 265548 223672 265600
rect 223724 265588 223730 265600
rect 224494 265588 224500 265600
rect 223724 265560 224500 265588
rect 223724 265548 223730 265560
rect 224494 265548 224500 265560
rect 224552 265548 224558 265600
rect 238846 265548 238852 265600
rect 238904 265588 238910 265600
rect 239674 265588 239680 265600
rect 238904 265560 239680 265588
rect 238904 265548 238910 265560
rect 239674 265548 239680 265560
rect 239732 265548 239738 265600
rect 240134 265548 240140 265600
rect 240192 265588 240198 265600
rect 240502 265588 240508 265600
rect 240192 265560 240508 265588
rect 240192 265548 240198 265560
rect 240502 265548 240508 265560
rect 240560 265548 240566 265600
rect 242986 265548 242992 265600
rect 243044 265588 243050 265600
rect 243630 265588 243636 265600
rect 243044 265560 243636 265588
rect 243044 265548 243050 265560
rect 243630 265548 243636 265560
rect 243688 265548 243694 265600
rect 244366 265548 244372 265600
rect 244424 265588 244430 265600
rect 245010 265588 245016 265600
rect 244424 265560 245016 265588
rect 244424 265548 244430 265560
rect 245010 265548 245016 265560
rect 245068 265548 245074 265600
rect 247218 265548 247224 265600
rect 247276 265588 247282 265600
rect 247678 265588 247684 265600
rect 247276 265560 247684 265588
rect 247276 265548 247282 265560
rect 247678 265548 247684 265560
rect 247736 265548 247742 265600
rect 251266 265548 251272 265600
rect 251324 265588 251330 265600
rect 251726 265588 251732 265600
rect 251324 265560 251732 265588
rect 251324 265548 251330 265560
rect 251726 265548 251732 265560
rect 251784 265548 251790 265600
rect 259638 265548 259644 265600
rect 259696 265588 259702 265600
rect 260190 265588 260196 265600
rect 259696 265560 260196 265588
rect 259696 265548 259702 265560
rect 260190 265548 260196 265560
rect 260248 265548 260254 265600
rect 262306 265548 262312 265600
rect 262364 265588 262370 265600
rect 262766 265588 262772 265600
rect 262364 265560 262772 265588
rect 262364 265548 262370 265560
rect 262766 265548 262772 265560
rect 262824 265548 262830 265600
rect 264974 265548 264980 265600
rect 265032 265588 265038 265600
rect 265894 265588 265900 265600
rect 265032 265560 265900 265588
rect 265032 265548 265038 265560
rect 265894 265548 265900 265560
rect 265952 265548 265958 265600
rect 266354 265548 266360 265600
rect 266412 265588 266418 265600
rect 267274 265588 267280 265600
rect 266412 265560 267280 265588
rect 266412 265548 266418 265560
rect 267274 265548 267280 265560
rect 267332 265548 267338 265600
rect 353110 265548 353116 265600
rect 353168 265588 353174 265600
rect 491294 265588 491300 265600
rect 353168 265560 491300 265588
rect 353168 265548 353174 265560
rect 491294 265548 491300 265560
rect 491352 265548 491358 265600
rect 336182 265480 336188 265532
rect 336240 265520 336246 265532
rect 447134 265520 447140 265532
rect 336240 265492 447140 265520
rect 336240 265480 336246 265492
rect 447134 265480 447140 265492
rect 447192 265480 447198 265532
rect 334342 265412 334348 265464
rect 334400 265452 334406 265464
rect 442994 265452 443000 265464
rect 334400 265424 443000 265452
rect 334400 265412 334406 265424
rect 442994 265412 443000 265424
rect 443052 265412 443058 265464
rect 333514 265344 333520 265396
rect 333572 265384 333578 265396
rect 440234 265384 440240 265396
rect 333572 265356 440240 265384
rect 333572 265344 333578 265356
rect 440234 265344 440240 265356
rect 440292 265344 440298 265396
rect 331674 265276 331680 265328
rect 331732 265316 331738 265328
rect 434898 265316 434904 265328
rect 331732 265288 434904 265316
rect 331732 265276 331738 265288
rect 434898 265276 434904 265288
rect 434956 265276 434962 265328
rect 327718 265208 327724 265260
rect 327776 265248 327782 265260
rect 425054 265248 425060 265260
rect 327776 265220 425060 265248
rect 327776 265208 327782 265220
rect 425054 265208 425060 265220
rect 425112 265208 425118 265260
rect 673362 265208 673368 265260
rect 673420 265248 673426 265260
rect 676214 265248 676220 265260
rect 673420 265220 676220 265248
rect 673420 265208 673426 265220
rect 676214 265208 676220 265220
rect 676272 265208 676278 265260
rect 325050 265140 325056 265192
rect 325108 265180 325114 265192
rect 418154 265180 418160 265192
rect 325108 265152 418160 265180
rect 325108 265140 325114 265152
rect 418154 265140 418160 265152
rect 418212 265140 418218 265192
rect 673270 265072 673276 265124
rect 673328 265112 673334 265124
rect 676030 265112 676036 265124
rect 673328 265084 676036 265112
rect 673328 265072 673334 265084
rect 676030 265072 676036 265084
rect 676088 265072 676094 265124
rect 673362 264936 673368 264988
rect 673420 264976 673426 264988
rect 676122 264976 676128 264988
rect 673420 264948 676128 264976
rect 673420 264936 673426 264948
rect 676122 264936 676128 264948
rect 676180 264936 676186 264988
rect 367002 264460 367008 264512
rect 367060 264500 367066 264512
rect 528554 264500 528560 264512
rect 367060 264472 528560 264500
rect 367060 264460 367066 264472
rect 528554 264460 528560 264472
rect 528612 264460 528618 264512
rect 384942 264392 384948 264444
rect 385000 264432 385006 264444
rect 575474 264432 575480 264444
rect 385000 264404 575480 264432
rect 385000 264392 385006 264404
rect 575474 264392 575480 264404
rect 575532 264392 575538 264444
rect 387610 264324 387616 264376
rect 387668 264364 387674 264376
rect 582558 264364 582564 264376
rect 387668 264336 582564 264364
rect 387668 264324 387674 264336
rect 582558 264324 582564 264336
rect 582616 264324 582622 264376
rect 393038 264256 393044 264308
rect 393096 264296 393102 264308
rect 597554 264296 597560 264308
rect 393096 264268 597560 264296
rect 393096 264256 393102 264268
rect 597554 264256 597560 264268
rect 597612 264256 597618 264308
rect 43990 264188 43996 264240
rect 44048 264228 44054 264240
rect 662414 264228 662420 264240
rect 44048 264200 662420 264228
rect 44048 264188 44054 264200
rect 662414 264188 662420 264200
rect 662472 264188 662478 264240
rect 399754 264120 399760 264172
rect 399812 264120 399818 264172
rect 401226 264120 401232 264172
rect 401284 264160 401290 264172
rect 607398 264160 607404 264172
rect 401284 264132 607404 264160
rect 401284 264120 401290 264132
rect 607398 264120 607404 264132
rect 607456 264120 607462 264172
rect 399772 264092 399800 264120
rect 615494 264092 615500 264104
rect 399772 264064 615500 264092
rect 615494 264052 615500 264064
rect 615552 264052 615558 264104
rect 673270 263576 673276 263628
rect 673328 263616 673334 263628
rect 676214 263616 676220 263628
rect 673328 263588 676220 263616
rect 673328 263576 673334 263588
rect 676214 263576 676220 263588
rect 676272 263576 676278 263628
rect 415302 262216 415308 262268
rect 415360 262256 415366 262268
rect 572714 262256 572720 262268
rect 415360 262228 572720 262256
rect 415360 262216 415366 262228
rect 572714 262216 572720 262228
rect 572772 262216 572778 262268
rect 674558 259088 674564 259140
rect 674616 259128 674622 259140
rect 676214 259128 676220 259140
rect 674616 259100 676220 259128
rect 674616 259088 674622 259100
rect 676214 259088 676220 259100
rect 676272 259088 676278 259140
rect 35802 258068 35808 258120
rect 35860 258108 35866 258120
rect 44910 258108 44916 258120
rect 35860 258080 44916 258108
rect 35860 258068 35866 258080
rect 44910 258068 44916 258080
rect 44968 258068 44974 258120
rect 179414 258068 179420 258120
rect 179472 258108 179478 258120
rect 189074 258108 189080 258120
rect 179472 258080 189080 258108
rect 179472 258068 179478 258080
rect 189074 258068 189080 258080
rect 189132 258068 189138 258120
rect 414198 258068 414204 258120
rect 414256 258108 414262 258120
rect 571518 258108 571524 258120
rect 414256 258080 571524 258108
rect 414256 258068 414262 258080
rect 571518 258068 571524 258080
rect 571576 258068 571582 258120
rect 673178 258068 673184 258120
rect 673236 258108 673242 258120
rect 676214 258108 676220 258120
rect 673236 258080 676220 258108
rect 673236 258068 673242 258080
rect 676214 258068 676220 258080
rect 676272 258068 676278 258120
rect 31662 258000 31668 258052
rect 31720 258040 31726 258052
rect 43714 258040 43720 258052
rect 31720 258012 43720 258040
rect 31720 258000 31726 258012
rect 43714 258000 43720 258012
rect 43772 258000 43778 258052
rect 31570 257864 31576 257916
rect 31628 257904 31634 257916
rect 44726 257904 44732 257916
rect 31628 257876 44732 257904
rect 31628 257864 31634 257876
rect 44726 257864 44732 257876
rect 44784 257864 44790 257916
rect 31662 257728 31668 257780
rect 31720 257768 31726 257780
rect 46198 257768 46204 257780
rect 31720 257740 46204 257768
rect 31720 257728 31726 257740
rect 46198 257728 46204 257740
rect 46256 257728 46262 257780
rect 673086 256708 673092 256760
rect 673144 256748 673150 256760
rect 683114 256748 683120 256760
rect 673144 256720 683120 256748
rect 673144 256708 673150 256720
rect 683114 256708 683120 256720
rect 683172 256708 683178 256760
rect 415302 255280 415308 255332
rect 415360 255320 415366 255332
rect 571426 255320 571432 255332
rect 415360 255292 571432 255320
rect 415360 255280 415366 255292
rect 571426 255280 571432 255292
rect 571484 255280 571490 255332
rect 414382 252560 414388 252612
rect 414440 252600 414446 252612
rect 574738 252600 574744 252612
rect 414440 252572 574744 252600
rect 414440 252560 414446 252572
rect 574738 252560 574744 252572
rect 574796 252560 574802 252612
rect 675754 252560 675760 252612
rect 675812 252600 675818 252612
rect 678238 252600 678244 252612
rect 675812 252572 678244 252600
rect 675812 252560 675818 252572
rect 678238 252560 678244 252572
rect 678296 252560 678302 252612
rect 675202 251608 675208 251660
rect 675260 251648 675266 251660
rect 676490 251648 676496 251660
rect 675260 251620 676496 251648
rect 675260 251608 675266 251620
rect 676490 251608 676496 251620
rect 676548 251608 676554 251660
rect 675018 251540 675024 251592
rect 675076 251580 675082 251592
rect 676858 251580 676864 251592
rect 675076 251552 676864 251580
rect 675076 251540 675082 251552
rect 676858 251540 676864 251552
rect 676916 251540 676922 251592
rect 676950 251540 676956 251592
rect 677008 251540 677014 251592
rect 674006 251472 674012 251524
rect 674064 251512 674070 251524
rect 676968 251512 676996 251540
rect 674064 251484 676996 251512
rect 674064 251472 674070 251484
rect 173894 251336 173900 251388
rect 173952 251376 173958 251388
rect 179414 251376 179420 251388
rect 173952 251348 179420 251376
rect 173952 251336 173958 251348
rect 179414 251336 179420 251348
rect 179472 251336 179478 251388
rect 675754 251200 675760 251252
rect 675812 251200 675818 251252
rect 675772 250980 675800 251200
rect 675754 250928 675760 250980
rect 675812 250928 675818 250980
rect 674466 249976 674472 250028
rect 674524 250016 674530 250028
rect 675202 250016 675208 250028
rect 674524 249988 675208 250016
rect 674524 249976 674530 249988
rect 675202 249976 675208 249988
rect 675260 249976 675266 250028
rect 673638 249840 673644 249892
rect 673696 249880 673702 249892
rect 674558 249880 674564 249892
rect 673696 249852 674564 249880
rect 673696 249840 673702 249852
rect 674558 249840 674564 249852
rect 674616 249840 674622 249892
rect 674558 249704 674564 249756
rect 674616 249744 674622 249756
rect 675018 249744 675024 249756
rect 674616 249716 675024 249744
rect 674616 249704 674622 249716
rect 675018 249704 675024 249716
rect 675076 249704 675082 249756
rect 171778 249296 171784 249348
rect 171836 249336 171842 249348
rect 173894 249336 173900 249348
rect 171836 249308 173900 249336
rect 171836 249296 171842 249308
rect 173894 249296 173900 249308
rect 173952 249296 173958 249348
rect 675202 248480 675208 248532
rect 675260 248480 675266 248532
rect 414198 248412 414204 248464
rect 414256 248452 414262 248464
rect 574094 248452 574100 248464
rect 414256 248424 574100 248452
rect 414256 248412 414262 248424
rect 574094 248412 574100 248424
rect 574152 248412 574158 248464
rect 675220 248328 675248 248480
rect 675202 248276 675208 248328
rect 675260 248276 675266 248328
rect 675018 247868 675024 247920
rect 675076 247908 675082 247920
rect 675478 247908 675484 247920
rect 675076 247880 675484 247908
rect 675076 247868 675082 247880
rect 675478 247868 675484 247880
rect 675536 247868 675542 247920
rect 674466 247256 674472 247308
rect 674524 247296 674530 247308
rect 675110 247296 675116 247308
rect 674524 247268 675116 247296
rect 674524 247256 674530 247268
rect 675110 247256 675116 247268
rect 675168 247256 675174 247308
rect 674558 247052 674564 247104
rect 674616 247092 674622 247104
rect 675386 247092 675392 247104
rect 674616 247064 675392 247092
rect 674616 247052 674622 247064
rect 675386 247052 675392 247064
rect 675444 247052 675450 247104
rect 674006 246508 674012 246560
rect 674064 246548 674070 246560
rect 675386 246548 675392 246560
rect 674064 246520 675392 246548
rect 674064 246508 674070 246520
rect 675386 246508 675392 246520
rect 675444 246508 675450 246560
rect 675110 246032 675116 246084
rect 675168 246072 675174 246084
rect 675386 246072 675392 246084
rect 675168 246044 675392 246072
rect 675168 246032 675174 246044
rect 675386 246032 675392 246044
rect 675444 246032 675450 246084
rect 42426 245760 42432 245812
rect 42484 245800 42490 245812
rect 42702 245800 42708 245812
rect 42484 245772 42708 245800
rect 42484 245760 42490 245772
rect 42702 245760 42708 245772
rect 42760 245760 42766 245812
rect 35802 245624 35808 245676
rect 35860 245664 35866 245676
rect 191098 245664 191104 245676
rect 35860 245636 191104 245664
rect 35860 245624 35866 245636
rect 191098 245624 191104 245636
rect 191156 245624 191162 245676
rect 415302 245624 415308 245676
rect 415360 245664 415366 245676
rect 565078 245664 565084 245676
rect 415360 245636 565084 245664
rect 415360 245624 415366 245636
rect 565078 245624 565084 245636
rect 565136 245624 565142 245676
rect 673914 243584 673920 243636
rect 673972 243624 673978 243636
rect 675294 243624 675300 243636
rect 673972 243596 675300 243624
rect 673972 243584 673978 243596
rect 675294 243584 675300 243596
rect 675352 243584 675358 243636
rect 414382 242904 414388 242956
rect 414440 242944 414446 242956
rect 623038 242944 623044 242956
rect 414440 242916 623044 242944
rect 414440 242904 414446 242916
rect 623038 242904 623044 242916
rect 623096 242904 623102 242956
rect 673638 242836 673644 242888
rect 673696 242876 673702 242888
rect 675294 242876 675300 242888
rect 673696 242848 675300 242876
rect 673696 242836 673702 242848
rect 675294 242836 675300 242848
rect 675352 242836 675358 242888
rect 171778 241544 171784 241596
rect 171836 241544 171842 241596
rect 164878 241408 164884 241460
rect 164936 241448 164942 241460
rect 171796 241448 171824 241544
rect 164936 241420 171824 241448
rect 164936 241408 164942 241420
rect 673178 241204 673184 241256
rect 673236 241244 673242 241256
rect 675294 241244 675300 241256
rect 673236 241216 675300 241244
rect 673236 241204 673242 241216
rect 675294 241204 675300 241216
rect 675352 241204 675358 241256
rect 42150 240320 42156 240372
rect 42208 240360 42214 240372
rect 42426 240360 42432 240372
rect 42208 240332 42432 240360
rect 42208 240320 42214 240332
rect 42426 240320 42432 240332
rect 42484 240320 42490 240372
rect 42702 238756 42708 238808
rect 42760 238796 42766 238808
rect 43162 238796 43168 238808
rect 42760 238768 43168 238796
rect 42760 238756 42766 238768
rect 43162 238756 43168 238768
rect 43220 238756 43226 238808
rect 185578 237396 185584 237448
rect 185636 237436 185642 237448
rect 189074 237436 189080 237448
rect 185636 237408 189080 237436
rect 185636 237396 185642 237408
rect 189074 237396 189080 237408
rect 189132 237396 189138 237448
rect 42150 235356 42156 235408
rect 42208 235396 42214 235408
rect 44542 235396 44548 235408
rect 42208 235368 44548 235396
rect 42208 235356 42214 235368
rect 44542 235356 44548 235368
rect 44600 235356 44606 235408
rect 182910 234948 182916 235000
rect 182968 234988 182974 235000
rect 185578 234988 185584 235000
rect 182968 234960 185584 234988
rect 182968 234948 182974 234960
rect 185578 234948 185584 234960
rect 185636 234948 185642 235000
rect 42150 233996 42156 234048
rect 42208 234036 42214 234048
rect 44450 234036 44456 234048
rect 42208 234008 44456 234036
rect 42208 233996 42214 234008
rect 44450 233996 44456 234008
rect 44508 233996 44514 234048
rect 178034 233452 178040 233504
rect 178092 233492 178098 233504
rect 182910 233492 182916 233504
rect 178092 233464 182916 233492
rect 178092 233452 178098 233464
rect 182910 233452 182916 233464
rect 182968 233452 182974 233504
rect 414198 232500 414204 232552
rect 414256 232540 414262 232552
rect 639138 232540 639144 232552
rect 414256 232512 639144 232540
rect 414256 232500 414262 232512
rect 639138 232500 639144 232512
rect 639196 232500 639202 232552
rect 414934 232432 414940 232484
rect 414992 232472 414998 232484
rect 638218 232472 638224 232484
rect 414992 232444 638224 232472
rect 414992 232432 414998 232444
rect 638218 232432 638224 232444
rect 638276 232432 638282 232484
rect 414290 232364 414296 232416
rect 414348 232404 414354 232416
rect 577498 232404 577504 232416
rect 414348 232376 577504 232404
rect 414348 232364 414354 232376
rect 577498 232364 577504 232376
rect 577556 232364 577562 232416
rect 190362 231684 190368 231736
rect 190420 231724 190426 231736
rect 604454 231724 604460 231736
rect 190420 231696 604460 231724
rect 190420 231684 190426 231696
rect 604454 231684 604460 231696
rect 604512 231684 604518 231736
rect 67542 231616 67548 231668
rect 67600 231656 67606 231668
rect 178034 231656 178040 231668
rect 67600 231628 178040 231656
rect 67600 231616 67606 231628
rect 178034 231616 178040 231628
rect 178092 231616 178098 231668
rect 191098 231616 191104 231668
rect 191156 231656 191162 231668
rect 663978 231656 663984 231668
rect 191156 231628 663984 231656
rect 191156 231616 191162 231628
rect 663978 231616 663984 231628
rect 664036 231616 664042 231668
rect 85022 231548 85028 231600
rect 85080 231588 85086 231600
rect 663794 231588 663800 231600
rect 85080 231560 663800 231588
rect 85080 231548 85086 231560
rect 663794 231548 663800 231560
rect 663852 231548 663858 231600
rect 84838 231480 84844 231532
rect 84896 231520 84902 231532
rect 663886 231520 663892 231532
rect 84896 231492 663892 231520
rect 84896 231480 84902 231492
rect 663886 231480 663892 231492
rect 663944 231480 663950 231532
rect 50338 231412 50344 231464
rect 50396 231452 50402 231464
rect 650638 231452 650644 231464
rect 50396 231424 650644 231452
rect 50396 231412 50402 231424
rect 650638 231412 650644 231424
rect 650696 231412 650702 231464
rect 48958 231344 48964 231396
rect 49016 231384 49022 231396
rect 649350 231384 649356 231396
rect 49016 231356 649356 231384
rect 49016 231344 49022 231356
rect 649350 231344 649356 231356
rect 649408 231344 649414 231396
rect 54478 231276 54484 231328
rect 54536 231316 54542 231328
rect 655514 231316 655520 231328
rect 54536 231288 655520 231316
rect 54536 231276 54542 231288
rect 655514 231276 655520 231288
rect 655572 231276 655578 231328
rect 51718 231208 51724 231260
rect 51776 231248 51782 231260
rect 652754 231248 652760 231260
rect 51776 231220 652760 231248
rect 51776 231208 51782 231220
rect 652754 231208 652760 231220
rect 652812 231208 652818 231260
rect 49050 231140 49056 231192
rect 49108 231180 49114 231192
rect 661034 231180 661040 231192
rect 49108 231152 661040 231180
rect 49108 231140 49114 231152
rect 661034 231140 661040 231152
rect 661092 231140 661098 231192
rect 43806 231072 43812 231124
rect 43864 231112 43870 231124
rect 662506 231112 662512 231124
rect 43864 231084 662512 231112
rect 43864 231072 43870 231084
rect 662506 231072 662512 231084
rect 662564 231072 662570 231124
rect 350166 230596 350172 230648
rect 350224 230636 350230 230648
rect 423674 230636 423680 230648
rect 350224 230608 423680 230636
rect 350224 230596 350230 230608
rect 423674 230596 423680 230608
rect 423732 230596 423738 230648
rect 385126 230528 385132 230580
rect 385184 230568 385190 230580
rect 507854 230568 507860 230580
rect 385184 230540 507860 230568
rect 385184 230528 385190 230540
rect 507854 230528 507860 230540
rect 507912 230528 507918 230580
rect 333606 230460 333612 230512
rect 333664 230500 333670 230512
rect 333664 230472 333928 230500
rect 333664 230460 333670 230472
rect 179322 230392 179328 230444
rect 179380 230432 179386 230444
rect 246114 230432 246120 230444
rect 179380 230404 246120 230432
rect 179380 230392 179386 230404
rect 246114 230392 246120 230404
rect 246172 230392 246178 230444
rect 262858 230392 262864 230444
rect 262916 230432 262922 230444
rect 269942 230432 269948 230444
rect 262916 230404 269948 230432
rect 262916 230392 262922 230404
rect 269942 230392 269948 230404
rect 270000 230392 270006 230444
rect 274634 230432 274640 230444
rect 271064 230404 274640 230432
rect 42058 230324 42064 230376
rect 42116 230364 42122 230376
rect 42978 230364 42984 230376
rect 42116 230336 42984 230364
rect 42116 230324 42122 230336
rect 42978 230324 42984 230336
rect 43036 230324 43042 230376
rect 175182 230324 175188 230376
rect 175240 230364 175246 230376
rect 244642 230364 244648 230376
rect 175240 230336 244648 230364
rect 175240 230324 175246 230336
rect 244642 230324 244648 230336
rect 244700 230324 244706 230376
rect 246942 230324 246948 230376
rect 247000 230364 247006 230376
rect 271064 230364 271092 230404
rect 274634 230392 274640 230404
rect 274692 230392 274698 230444
rect 276658 230392 276664 230444
rect 276716 230432 276722 230444
rect 277762 230432 277768 230444
rect 276716 230404 277768 230432
rect 276716 230392 276722 230404
rect 277762 230392 277768 230404
rect 277820 230392 277826 230444
rect 285306 230432 285312 230444
rect 277964 230404 285312 230432
rect 247000 230336 271092 230364
rect 247000 230324 247006 230336
rect 271138 230324 271144 230376
rect 271196 230364 271202 230376
rect 272794 230364 272800 230376
rect 271196 230336 272800 230364
rect 271196 230324 271202 230336
rect 272794 230324 272800 230336
rect 272852 230324 272858 230376
rect 169662 230256 169668 230308
rect 169720 230296 169726 230308
rect 241790 230296 241796 230308
rect 169720 230268 241796 230296
rect 169720 230256 169726 230268
rect 241790 230256 241796 230268
rect 241848 230256 241854 230308
rect 244182 230256 244188 230308
rect 244240 230296 244246 230308
rect 274266 230296 274272 230308
rect 244240 230268 274272 230296
rect 244240 230256 244246 230268
rect 274266 230256 274272 230268
rect 274324 230256 274330 230308
rect 274542 230256 274548 230308
rect 274600 230296 274606 230308
rect 277964 230296 277992 230404
rect 285306 230392 285312 230404
rect 285364 230392 285370 230444
rect 286962 230392 286968 230444
rect 287020 230432 287026 230444
rect 287020 230404 288296 230432
rect 287020 230392 287026 230404
rect 279418 230324 279424 230376
rect 279476 230364 279482 230376
rect 283190 230364 283196 230376
rect 279476 230336 283196 230364
rect 279476 230324 279482 230336
rect 283190 230324 283196 230336
rect 283248 230324 283254 230376
rect 287422 230364 287428 230376
rect 283300 230336 287428 230364
rect 274600 230268 277992 230296
rect 274600 230256 274606 230268
rect 278038 230256 278044 230308
rect 278096 230296 278102 230308
rect 283300 230296 283328 230336
rect 287422 230324 287428 230336
rect 287480 230324 287486 230376
rect 288268 230364 288296 230404
rect 288342 230392 288348 230444
rect 288400 230432 288406 230444
rect 292758 230432 292764 230444
rect 288400 230404 292764 230432
rect 288400 230392 288406 230404
rect 292758 230392 292764 230404
rect 292816 230392 292822 230444
rect 297450 230392 297456 230444
rect 297508 230432 297514 230444
rect 299934 230432 299940 230444
rect 297508 230404 299940 230432
rect 297508 230392 297514 230404
rect 299934 230392 299940 230404
rect 299992 230392 299998 230444
rect 300210 230392 300216 230444
rect 300268 230432 300274 230444
rect 303982 230432 303988 230444
rect 300268 230404 303988 230432
rect 300268 230392 300274 230404
rect 303982 230392 303988 230404
rect 304040 230392 304046 230444
rect 311710 230392 311716 230444
rect 311768 230432 311774 230444
rect 315298 230432 315304 230444
rect 311768 230404 315304 230432
rect 311768 230392 311774 230404
rect 315298 230392 315304 230404
rect 315356 230392 315362 230444
rect 323118 230392 323124 230444
rect 323176 230432 323182 230444
rect 323176 230404 325694 230432
rect 323176 230392 323182 230404
rect 291746 230364 291752 230376
rect 288268 230336 291752 230364
rect 291746 230324 291752 230336
rect 291804 230324 291810 230376
rect 292574 230324 292580 230376
rect 292632 230364 292638 230376
rect 293862 230364 293868 230376
rect 292632 230336 293868 230364
rect 292632 230324 292638 230336
rect 293862 230324 293868 230336
rect 293920 230324 293926 230376
rect 298094 230324 298100 230376
rect 298152 230364 298158 230376
rect 299290 230364 299296 230376
rect 298152 230336 299296 230364
rect 298152 230324 298158 230336
rect 299290 230324 299296 230336
rect 299348 230324 299354 230376
rect 299566 230324 299572 230376
rect 299624 230364 299630 230376
rect 300486 230364 300492 230376
rect 299624 230336 300492 230364
rect 299624 230324 299630 230336
rect 300486 230324 300492 230336
rect 300544 230324 300550 230376
rect 304166 230324 304172 230376
rect 304224 230364 304230 230376
rect 304902 230364 304908 230376
rect 304224 230336 304908 230364
rect 304224 230324 304230 230336
rect 304902 230324 304908 230336
rect 304960 230324 304966 230376
rect 305638 230324 305644 230376
rect 305696 230364 305702 230376
rect 306190 230364 306196 230376
rect 305696 230336 306196 230364
rect 305696 230324 305702 230336
rect 306190 230324 306196 230336
rect 306248 230324 306254 230376
rect 307018 230324 307024 230376
rect 307076 230364 307082 230376
rect 307570 230364 307576 230376
rect 307076 230336 307576 230364
rect 307076 230324 307082 230336
rect 307570 230324 307576 230336
rect 307628 230324 307634 230376
rect 312078 230324 312084 230376
rect 312136 230364 312142 230376
rect 313182 230364 313188 230376
rect 312136 230336 313188 230364
rect 312136 230324 312142 230336
rect 313182 230324 313188 230336
rect 313240 230324 313246 230376
rect 314930 230324 314936 230376
rect 314988 230364 314994 230376
rect 315942 230364 315948 230376
rect 314988 230336 315948 230364
rect 314988 230324 314994 230336
rect 315942 230324 315948 230336
rect 316000 230324 316006 230376
rect 316310 230324 316316 230376
rect 316368 230364 316374 230376
rect 317322 230364 317328 230376
rect 316368 230336 317328 230364
rect 316368 230324 316374 230336
rect 317322 230324 317328 230336
rect 317380 230324 317386 230376
rect 319254 230324 319260 230376
rect 319312 230364 319318 230376
rect 319898 230364 319904 230376
rect 319312 230336 319904 230364
rect 319312 230324 319318 230336
rect 319898 230324 319904 230336
rect 319956 230324 319962 230376
rect 323486 230324 323492 230376
rect 323544 230364 323550 230376
rect 324222 230364 324228 230376
rect 323544 230336 324228 230364
rect 323544 230324 323550 230336
rect 324222 230324 324228 230336
rect 324280 230324 324286 230376
rect 325666 230364 325694 230404
rect 328454 230392 328460 230444
rect 328512 230432 328518 230444
rect 329558 230432 329564 230444
rect 328512 230404 329564 230432
rect 328512 230392 328518 230404
rect 329558 230392 329564 230404
rect 329616 230392 329622 230444
rect 329834 230392 329840 230444
rect 329892 230432 329898 230444
rect 330846 230432 330852 230444
rect 329892 230404 330852 230432
rect 329892 230392 329898 230404
rect 330846 230392 330852 230404
rect 330904 230392 330910 230444
rect 331674 230392 331680 230444
rect 331732 230432 331738 230444
rect 332410 230432 332416 230444
rect 331732 230404 332416 230432
rect 331732 230392 331738 230404
rect 332410 230392 332416 230404
rect 332468 230392 332474 230444
rect 333054 230392 333060 230444
rect 333112 230432 333118 230444
rect 333790 230432 333796 230444
rect 333112 230404 333796 230432
rect 333112 230392 333118 230404
rect 333790 230392 333796 230404
rect 333848 230392 333854 230444
rect 333900 230432 333928 230472
rect 386230 230460 386236 230512
rect 386288 230500 386294 230512
rect 511258 230500 511264 230512
rect 386288 230472 511264 230500
rect 386288 230460 386294 230472
rect 511258 230460 511264 230472
rect 511316 230460 511322 230512
rect 604454 230460 604460 230512
rect 604512 230500 604518 230512
rect 605742 230500 605748 230512
rect 604512 230472 605748 230500
rect 604512 230460 604518 230472
rect 605742 230460 605748 230472
rect 605800 230500 605806 230512
rect 636838 230500 636844 230512
rect 605800 230472 636844 230500
rect 605800 230460 605806 230472
rect 636838 230460 636844 230472
rect 636896 230460 636902 230512
rect 371878 230432 371884 230444
rect 333900 230404 371884 230432
rect 371878 230392 371884 230404
rect 371936 230392 371942 230444
rect 382274 230392 382280 230444
rect 382332 230432 382338 230444
rect 383562 230432 383568 230444
rect 382332 230404 383568 230432
rect 382332 230392 382338 230404
rect 383562 230392 383568 230404
rect 383620 230392 383626 230444
rect 386874 230392 386880 230444
rect 386932 230432 386938 230444
rect 388438 230432 388444 230444
rect 386932 230404 388444 230432
rect 386932 230392 386938 230404
rect 388438 230392 388444 230404
rect 388496 230392 388502 230444
rect 393314 230392 393320 230444
rect 393372 230432 393378 230444
rect 394602 230432 394608 230444
rect 393372 230404 394608 230432
rect 393372 230392 393378 230404
rect 394602 230392 394608 230404
rect 394660 230392 394666 230444
rect 401870 230392 401876 230444
rect 401928 230432 401934 230444
rect 456150 230432 456156 230444
rect 401928 230404 456156 230432
rect 401928 230392 401934 230404
rect 456150 230392 456156 230404
rect 456208 230392 456214 230444
rect 340138 230364 340144 230376
rect 325666 230336 340144 230364
rect 340138 230324 340144 230336
rect 340196 230324 340202 230376
rect 341978 230324 341984 230376
rect 342036 230364 342042 230376
rect 380434 230364 380440 230376
rect 342036 230336 380440 230364
rect 342036 230324 342042 230336
rect 380434 230324 380440 230336
rect 380492 230324 380498 230376
rect 381170 230324 381176 230376
rect 381228 230364 381234 230376
rect 382182 230364 382188 230376
rect 381228 230336 382188 230364
rect 381228 230324 381234 230336
rect 382182 230324 382188 230336
rect 382240 230324 382246 230376
rect 382642 230324 382648 230376
rect 382700 230364 382706 230376
rect 383378 230364 383384 230376
rect 382700 230336 383384 230364
rect 382700 230324 382706 230336
rect 383378 230324 383384 230336
rect 383436 230324 383442 230376
rect 383654 230324 383660 230376
rect 383712 230364 383718 230376
rect 384942 230364 384948 230376
rect 383712 230336 384948 230364
rect 383712 230324 383718 230336
rect 384942 230324 384948 230336
rect 385000 230324 385006 230376
rect 385494 230324 385500 230376
rect 385552 230364 385558 230376
rect 386322 230364 386328 230376
rect 385552 230336 386328 230364
rect 385552 230324 385558 230336
rect 386322 230324 386328 230336
rect 386380 230324 386386 230376
rect 386506 230324 386512 230376
rect 386564 230364 386570 230376
rect 387702 230364 387708 230376
rect 386564 230336 387708 230364
rect 386564 230324 386570 230336
rect 387702 230324 387708 230336
rect 387760 230324 387766 230376
rect 387794 230324 387800 230376
rect 387852 230364 387858 230376
rect 400674 230364 400680 230376
rect 387852 230336 400680 230364
rect 387852 230324 387858 230336
rect 400674 230324 400680 230336
rect 400732 230324 400738 230376
rect 403342 230324 403348 230376
rect 403400 230364 403406 230376
rect 404170 230364 404176 230376
rect 403400 230336 404176 230364
rect 403400 230324 403406 230336
rect 404170 230324 404176 230336
rect 404228 230324 404234 230376
rect 406194 230324 406200 230376
rect 406252 230364 406258 230376
rect 407022 230364 407028 230376
rect 406252 230336 407028 230364
rect 406252 230324 406258 230336
rect 407022 230324 407028 230336
rect 407080 230324 407086 230376
rect 409046 230324 409052 230376
rect 409104 230364 409110 230376
rect 411162 230364 411168 230376
rect 409104 230336 411168 230364
rect 409104 230324 409110 230336
rect 411162 230324 411168 230336
rect 411220 230324 411226 230376
rect 411346 230324 411352 230376
rect 411404 230364 411410 230376
rect 461578 230364 461584 230376
rect 411404 230336 461584 230364
rect 411404 230324 411410 230336
rect 461578 230324 461584 230336
rect 461636 230324 461642 230376
rect 278096 230268 283328 230296
rect 278096 230256 278102 230268
rect 285582 230256 285588 230308
rect 285640 230296 285646 230308
rect 290642 230296 290648 230308
rect 285640 230268 290648 230296
rect 285640 230256 285646 230268
rect 290642 230256 290648 230268
rect 290700 230256 290706 230308
rect 310606 230256 310612 230308
rect 310664 230296 310670 230308
rect 314470 230296 314476 230308
rect 310664 230268 314476 230296
rect 310664 230256 310670 230268
rect 314470 230256 314476 230268
rect 314528 230256 314534 230308
rect 317414 230256 317420 230308
rect 317472 230296 317478 230308
rect 317472 230268 320220 230296
rect 317472 230256 317478 230268
rect 136358 230188 136364 230240
rect 136416 230228 136422 230240
rect 213270 230228 213276 230240
rect 136416 230200 213276 230228
rect 136416 230188 136422 230200
rect 213270 230188 213276 230200
rect 213328 230188 213334 230240
rect 219250 230188 219256 230240
rect 219308 230228 219314 230240
rect 263226 230228 263232 230240
rect 219308 230200 263232 230228
rect 219308 230188 219314 230200
rect 263226 230188 263232 230200
rect 263284 230188 263290 230240
rect 276750 230188 276756 230240
rect 276808 230228 276814 230240
rect 287054 230228 287060 230240
rect 276808 230200 287060 230228
rect 276808 230188 276814 230200
rect 287054 230188 287060 230200
rect 287112 230188 287118 230240
rect 298830 230188 298836 230240
rect 298888 230228 298894 230240
rect 302418 230228 302424 230240
rect 298888 230200 302424 230228
rect 298888 230188 298894 230200
rect 302418 230188 302424 230200
rect 302476 230188 302482 230240
rect 314562 230188 314568 230240
rect 314620 230228 314626 230240
rect 314620 230200 316034 230228
rect 314620 230188 314626 230200
rect 155862 230120 155868 230172
rect 155920 230160 155926 230172
rect 236086 230160 236092 230172
rect 155920 230132 236092 230160
rect 155920 230120 155926 230132
rect 236086 230120 236092 230132
rect 236144 230120 236150 230172
rect 240042 230120 240048 230172
rect 240100 230160 240106 230172
rect 271782 230160 271788 230172
rect 240100 230132 271788 230160
rect 240100 230120 240106 230132
rect 271782 230120 271788 230132
rect 271840 230120 271846 230172
rect 275370 230120 275376 230172
rect 275428 230160 275434 230172
rect 277670 230160 277676 230172
rect 275428 230132 277676 230160
rect 275428 230120 275434 230132
rect 277670 230120 277676 230132
rect 277728 230120 277734 230172
rect 277762 230120 277768 230172
rect 277820 230160 277826 230172
rect 286042 230160 286048 230172
rect 277820 230132 286048 230160
rect 277820 230120 277826 230132
rect 286042 230120 286048 230132
rect 286100 230120 286106 230172
rect 316006 230160 316034 230200
rect 317782 230188 317788 230240
rect 317840 230228 317846 230240
rect 318702 230228 318708 230240
rect 317840 230200 318708 230228
rect 317840 230188 317846 230200
rect 318702 230188 318708 230200
rect 318760 230188 318766 230240
rect 319346 230160 319352 230172
rect 316006 230132 319352 230160
rect 319346 230120 319352 230132
rect 319404 230120 319410 230172
rect 320192 230160 320220 230268
rect 320266 230256 320272 230308
rect 320324 230296 320330 230308
rect 337378 230296 337384 230308
rect 320324 230268 337384 230296
rect 320324 230256 320330 230268
rect 337378 230256 337384 230268
rect 337436 230256 337442 230308
rect 339126 230256 339132 230308
rect 339184 230296 339190 230308
rect 378962 230296 378968 230308
rect 339184 230268 378968 230296
rect 339184 230256 339190 230268
rect 378962 230256 378968 230268
rect 379020 230256 379026 230308
rect 385862 230256 385868 230308
rect 385920 230296 385926 230308
rect 391106 230296 391112 230308
rect 385920 230268 391112 230296
rect 385920 230256 385926 230268
rect 391106 230256 391112 230268
rect 391164 230256 391170 230308
rect 398650 230256 398656 230308
rect 398708 230296 398714 230308
rect 405734 230296 405740 230308
rect 398708 230268 405740 230296
rect 398708 230256 398714 230268
rect 405734 230256 405740 230268
rect 405792 230256 405798 230308
rect 405826 230256 405832 230308
rect 405884 230296 405890 230308
rect 409598 230296 409604 230308
rect 405884 230268 409604 230296
rect 405884 230256 405890 230268
rect 409598 230256 409604 230268
rect 409656 230256 409662 230308
rect 409782 230256 409788 230308
rect 409840 230296 409846 230308
rect 467098 230296 467104 230308
rect 409840 230268 467104 230296
rect 409840 230256 409846 230268
rect 467098 230256 467104 230268
rect 467156 230256 467162 230308
rect 321646 230188 321652 230240
rect 321704 230228 321710 230240
rect 338758 230228 338764 230240
rect 321704 230200 338764 230228
rect 321704 230188 321710 230200
rect 338758 230188 338764 230200
rect 338816 230188 338822 230240
rect 347682 230188 347688 230240
rect 347740 230228 347746 230240
rect 387610 230228 387616 230240
rect 347740 230200 387616 230228
rect 347740 230188 347746 230200
rect 387610 230188 387616 230200
rect 387668 230188 387674 230240
rect 389082 230188 389088 230240
rect 389140 230228 389146 230240
rect 396718 230228 396724 230240
rect 389140 230200 396724 230228
rect 389140 230188 389146 230200
rect 396718 230188 396724 230200
rect 396776 230188 396782 230240
rect 398098 230188 398104 230240
rect 398156 230228 398162 230240
rect 403066 230228 403072 230240
rect 398156 230200 403072 230228
rect 398156 230188 398162 230200
rect 403066 230188 403072 230200
rect 403124 230188 403130 230240
rect 403986 230188 403992 230240
rect 404044 230228 404050 230240
rect 406654 230228 406660 230240
rect 404044 230200 406660 230228
rect 404044 230188 404050 230200
rect 406654 230188 406660 230200
rect 406712 230188 406718 230240
rect 406838 230188 406844 230240
rect 406896 230228 406902 230240
rect 411070 230228 411076 230240
rect 406896 230200 411076 230228
rect 406896 230188 406902 230200
rect 411070 230188 411076 230200
rect 411128 230188 411134 230240
rect 411254 230188 411260 230240
rect 411312 230228 411318 230240
rect 468478 230228 468484 230240
rect 411312 230200 468484 230228
rect 411312 230188 411318 230200
rect 468478 230188 468484 230200
rect 468536 230188 468542 230240
rect 330110 230160 330116 230172
rect 320192 230132 330116 230160
rect 330110 230120 330116 230132
rect 330168 230120 330174 230172
rect 330202 230120 330208 230172
rect 330260 230160 330266 230172
rect 331030 230160 331036 230172
rect 330260 230132 331036 230160
rect 330260 230120 330266 230132
rect 331030 230120 331036 230132
rect 331088 230120 331094 230172
rect 336642 230120 336648 230172
rect 336700 230160 336706 230172
rect 376018 230160 376024 230172
rect 336700 230132 376024 230160
rect 336700 230120 336706 230132
rect 376018 230120 376024 230132
rect 376076 230120 376082 230172
rect 378318 230120 378324 230172
rect 378376 230160 378382 230172
rect 443638 230160 443644 230172
rect 378376 230132 443644 230160
rect 378376 230120 378382 230132
rect 443638 230120 443644 230132
rect 443696 230120 443702 230172
rect 146202 230052 146208 230104
rect 146260 230092 146266 230104
rect 231854 230092 231860 230104
rect 146260 230064 231860 230092
rect 146260 230052 146266 230064
rect 231854 230052 231860 230064
rect 231912 230052 231918 230104
rect 234522 230052 234528 230104
rect 234580 230092 234586 230104
rect 262858 230092 262864 230104
rect 234580 230064 262864 230092
rect 234580 230052 234586 230064
rect 262858 230052 262864 230064
rect 262916 230052 262922 230104
rect 268930 230092 268936 230104
rect 267706 230064 268936 230092
rect 139302 229984 139308 230036
rect 139360 230024 139366 230036
rect 229002 230024 229008 230036
rect 139360 229996 229008 230024
rect 139360 229984 139366 229996
rect 229002 229984 229008 229996
rect 229060 229984 229066 230036
rect 233142 229984 233148 230036
rect 233200 230024 233206 230036
rect 267706 230024 267734 230064
rect 268930 230052 268936 230064
rect 268988 230052 268994 230104
rect 271322 230052 271328 230104
rect 271380 230092 271386 230104
rect 277118 230092 277124 230104
rect 271380 230064 277124 230092
rect 271380 230052 271386 230064
rect 277118 230052 277124 230064
rect 277176 230052 277182 230104
rect 283834 230092 283840 230104
rect 277228 230064 283840 230092
rect 233200 229996 267734 230024
rect 233200 229984 233206 229996
rect 270310 229984 270316 230036
rect 270368 230024 270374 230036
rect 277228 230024 277256 230064
rect 283834 230052 283840 230064
rect 283892 230052 283898 230104
rect 315850 230052 315856 230104
rect 315908 230092 315914 230104
rect 322198 230092 322204 230104
rect 315908 230064 322204 230092
rect 315908 230052 315914 230064
rect 322198 230052 322204 230064
rect 322256 230052 322262 230104
rect 323762 230052 323768 230104
rect 323820 230092 323826 230104
rect 364518 230092 364524 230104
rect 323820 230064 364524 230092
rect 323820 230052 323826 230064
rect 364518 230052 364524 230064
rect 364576 230052 364582 230104
rect 368014 230052 368020 230104
rect 368072 230092 368078 230104
rect 387518 230092 387524 230104
rect 368072 230064 387524 230092
rect 368072 230052 368078 230064
rect 387518 230052 387524 230064
rect 387576 230052 387582 230104
rect 387978 230052 387984 230104
rect 388036 230092 388042 230104
rect 515398 230092 515404 230104
rect 388036 230064 515404 230092
rect 388036 230052 388042 230064
rect 515398 230052 515404 230064
rect 515456 230052 515462 230104
rect 270368 229996 277256 230024
rect 270368 229984 270374 229996
rect 277302 229984 277308 230036
rect 277360 230024 277366 230036
rect 282454 230024 282460 230036
rect 277360 229996 282460 230024
rect 277360 229984 277366 229996
rect 282454 229984 282460 229996
rect 282512 229984 282518 230036
rect 284202 229984 284208 230036
rect 284260 230024 284266 230036
rect 290274 230024 290280 230036
rect 284260 229996 290280 230024
rect 284260 229984 284266 229996
rect 290274 229984 290280 229996
rect 290332 229984 290338 230036
rect 312354 229984 312360 230036
rect 312412 230024 312418 230036
rect 336918 230024 336924 230036
rect 312412 229996 336924 230024
rect 312412 229984 312418 229996
rect 336918 229984 336924 229996
rect 336976 229984 336982 230036
rect 343726 229984 343732 230036
rect 343784 230024 343790 230036
rect 385678 230024 385684 230036
rect 343784 229996 385684 230024
rect 343784 229984 343790 229996
rect 385678 229984 385684 229996
rect 385736 229984 385742 230036
rect 399018 229984 399024 230036
rect 399076 230024 399082 230036
rect 400122 230024 400128 230036
rect 399076 229996 400128 230024
rect 399076 229984 399082 229996
rect 400122 229984 400128 229996
rect 400180 229984 400186 230036
rect 401134 229984 401140 230036
rect 401192 230024 401198 230036
rect 406746 230024 406752 230036
rect 401192 229996 406752 230024
rect 401192 229984 401198 229996
rect 406746 229984 406752 229996
rect 406804 229984 406810 230036
rect 407022 229984 407028 230036
rect 407080 230024 407086 230036
rect 409782 230024 409788 230036
rect 407080 229996 409788 230024
rect 407080 229984 407086 229996
rect 409782 229984 409788 229996
rect 409840 229984 409846 230036
rect 539594 230024 539600 230036
rect 409984 229996 539600 230024
rect 132402 229916 132408 229968
rect 132460 229956 132466 229968
rect 226150 229956 226156 229968
rect 132460 229928 226156 229956
rect 132460 229916 132466 229928
rect 226150 229916 226156 229928
rect 226208 229916 226214 229968
rect 226242 229916 226248 229968
rect 226300 229956 226306 229968
rect 266078 229956 266084 229968
rect 226300 229928 266084 229956
rect 226300 229916 226306 229928
rect 266078 229916 266084 229928
rect 266136 229916 266142 229968
rect 270402 229916 270408 229968
rect 270460 229956 270466 229968
rect 284570 229956 284576 229968
rect 270460 229928 284576 229956
rect 270460 229916 270466 229928
rect 284570 229916 284576 229928
rect 284628 229916 284634 229968
rect 285490 229916 285496 229968
rect 285548 229956 285554 229968
rect 291378 229956 291384 229968
rect 285548 229928 291384 229956
rect 285548 229916 285554 229928
rect 291378 229916 291384 229928
rect 291436 229916 291442 229968
rect 303522 229916 303528 229968
rect 303580 229956 303586 229968
rect 312538 229956 312544 229968
rect 303580 229928 312544 229956
rect 303580 229916 303586 229928
rect 312538 229916 312544 229928
rect 312596 229916 312602 229968
rect 313826 229916 313832 229968
rect 313884 229956 313890 229968
rect 341242 229956 341248 229968
rect 313884 229928 341248 229956
rect 313884 229916 313890 229928
rect 341242 229916 341248 229928
rect 341300 229916 341306 229968
rect 356238 229916 356244 229968
rect 356296 229956 356302 229968
rect 357066 229956 357072 229968
rect 356296 229928 357072 229956
rect 356296 229916 356302 229928
rect 357066 229916 357072 229928
rect 357124 229916 357130 229968
rect 359090 229916 359096 229968
rect 359148 229956 359154 229968
rect 360102 229956 360108 229968
rect 359148 229928 360108 229956
rect 359148 229916 359154 229928
rect 360102 229916 360108 229928
rect 360160 229916 360166 229968
rect 360562 229916 360568 229968
rect 360620 229956 360626 229968
rect 361298 229956 361304 229968
rect 360620 229928 361304 229956
rect 360620 229916 360626 229928
rect 361298 229916 361304 229928
rect 361356 229916 361362 229968
rect 361942 229916 361948 229968
rect 362000 229956 362006 229968
rect 362678 229956 362684 229968
rect 362000 229928 362684 229956
rect 362000 229916 362006 229928
rect 362678 229916 362684 229928
rect 362736 229916 362742 229968
rect 362770 229916 362776 229968
rect 362828 229956 362834 229968
rect 406470 229956 406476 229968
rect 362828 229928 406476 229956
rect 362828 229916 362834 229928
rect 406470 229916 406476 229928
rect 406528 229916 406534 229968
rect 407206 229916 407212 229968
rect 407264 229956 407270 229968
rect 407264 229928 409828 229956
rect 407264 229916 407270 229928
rect 91738 229848 91744 229900
rect 91796 229888 91802 229900
rect 203334 229888 203340 229900
rect 91796 229860 203340 229888
rect 91796 229848 91802 229860
rect 203334 229848 203340 229860
rect 203392 229848 203398 229900
rect 212442 229848 212448 229900
rect 212500 229888 212506 229900
rect 260374 229888 260380 229900
rect 212500 229860 260380 229888
rect 212500 229848 212506 229860
rect 260374 229848 260380 229860
rect 260432 229848 260438 229900
rect 263502 229848 263508 229900
rect 263560 229888 263566 229900
rect 281718 229888 281724 229900
rect 263560 229860 281724 229888
rect 263560 229848 263566 229860
rect 281718 229848 281724 229860
rect 281776 229848 281782 229900
rect 296714 229848 296720 229900
rect 296772 229888 296778 229900
rect 299566 229888 299572 229900
rect 296772 229860 299572 229888
rect 296772 229848 296778 229860
rect 299566 229848 299572 229860
rect 299624 229848 299630 229900
rect 304994 229848 305000 229900
rect 305052 229888 305058 229900
rect 311434 229888 311440 229900
rect 305052 229860 311440 229888
rect 305052 229848 305058 229860
rect 311434 229848 311440 229860
rect 311492 229848 311498 229900
rect 316678 229848 316684 229900
rect 316736 229888 316742 229900
rect 346486 229888 346492 229900
rect 316736 229860 346492 229888
rect 316736 229848 316742 229860
rect 346486 229848 346492 229860
rect 346544 229848 346550 229900
rect 352006 229848 352012 229900
rect 352064 229888 352070 229900
rect 398098 229888 398104 229900
rect 352064 229860 398104 229888
rect 352064 229848 352070 229860
rect 398098 229848 398104 229860
rect 398156 229848 398162 229900
rect 399754 229848 399760 229900
rect 399812 229888 399818 229900
rect 407758 229888 407764 229900
rect 399812 229860 407764 229888
rect 399812 229848 399818 229860
rect 407758 229848 407764 229860
rect 407816 229848 407822 229900
rect 409800 229888 409828 229928
rect 409984 229888 410012 229996
rect 539594 229984 539600 229996
rect 539652 229984 539658 230036
rect 411346 229956 411352 229968
rect 409800 229860 410012 229888
rect 410168 229928 411352 229956
rect 85390 229780 85396 229832
rect 85448 229820 85454 229832
rect 206186 229820 206192 229832
rect 85448 229792 206192 229820
rect 85448 229780 85454 229792
rect 206186 229780 206192 229792
rect 206244 229780 206250 229832
rect 206738 229780 206744 229832
rect 206796 229820 206802 229832
rect 257522 229820 257528 229832
rect 206796 229792 257528 229820
rect 206796 229780 206802 229792
rect 257522 229780 257528 229792
rect 257580 229780 257586 229832
rect 259362 229780 259368 229832
rect 259420 229820 259426 229832
rect 280338 229820 280344 229832
rect 259420 229792 280344 229820
rect 259420 229780 259426 229792
rect 280338 229780 280344 229792
rect 280396 229780 280402 229832
rect 281350 229780 281356 229832
rect 281408 229820 281414 229832
rect 289906 229820 289912 229832
rect 281408 229792 289912 229820
rect 281408 229780 281414 229792
rect 289906 229780 289912 229792
rect 289964 229780 289970 229832
rect 302050 229780 302056 229832
rect 302108 229820 302114 229832
rect 311158 229820 311164 229832
rect 302108 229792 311164 229820
rect 302108 229780 302114 229792
rect 311158 229780 311164 229792
rect 311216 229780 311222 229832
rect 318058 229780 318064 229832
rect 318116 229820 318122 229832
rect 350902 229820 350908 229832
rect 318116 229792 350908 229820
rect 318116 229780 318122 229792
rect 350902 229780 350908 229792
rect 350960 229780 350966 229832
rect 354858 229780 354864 229832
rect 354916 229820 354922 229832
rect 407114 229820 407120 229832
rect 354916 229792 407120 229820
rect 354916 229780 354922 229792
rect 407114 229780 407120 229792
rect 407172 229780 407178 229832
rect 410168 229820 410196 229928
rect 411346 229916 411352 229928
rect 411404 229916 411410 229968
rect 547138 229956 547144 229968
rect 412606 229928 547144 229956
rect 412606 229888 412634 229928
rect 547138 229916 547144 229928
rect 547196 229916 547202 229968
rect 408236 229792 410196 229820
rect 410260 229860 412634 229888
rect 71682 229712 71688 229764
rect 71740 229752 71746 229764
rect 200482 229752 200488 229764
rect 71740 229724 200488 229752
rect 71740 229712 71746 229724
rect 200482 229712 200488 229724
rect 200540 229712 200546 229764
rect 200666 229712 200672 229764
rect 200724 229752 200730 229764
rect 254670 229752 254676 229764
rect 200724 229724 254676 229752
rect 200724 229712 200730 229724
rect 254670 229712 254676 229724
rect 254728 229712 254734 229764
rect 255222 229712 255228 229764
rect 255280 229752 255286 229764
rect 278498 229752 278504 229764
rect 255280 229724 278504 229752
rect 255280 229712 255286 229724
rect 278498 229712 278504 229724
rect 278556 229712 278562 229764
rect 278682 229712 278688 229764
rect 278740 229752 278746 229764
rect 288526 229752 288532 229764
rect 278740 229724 288532 229752
rect 278740 229712 278746 229724
rect 288526 229712 288532 229724
rect 288584 229712 288590 229764
rect 315206 229712 315212 229764
rect 315264 229752 315270 229764
rect 343726 229752 343732 229764
rect 315264 229724 343732 229752
rect 315264 229712 315270 229724
rect 343726 229712 343732 229724
rect 343784 229712 343790 229764
rect 344830 229712 344836 229764
rect 344888 229752 344894 229764
rect 406378 229752 406384 229764
rect 344888 229724 406384 229752
rect 344888 229712 344894 229724
rect 406378 229712 406384 229724
rect 406436 229712 406442 229764
rect 406654 229712 406660 229764
rect 406712 229752 406718 229764
rect 408236 229752 408264 229792
rect 406712 229724 408264 229752
rect 406712 229712 406718 229724
rect 408310 229712 408316 229764
rect 408368 229752 408374 229764
rect 410260 229752 410288 229860
rect 410426 229780 410432 229832
rect 410484 229820 410490 229832
rect 563698 229820 563704 229832
rect 410484 229792 563704 229820
rect 410484 229780 410490 229792
rect 563698 229780 563704 229792
rect 563756 229780 563762 229832
rect 408368 229724 410288 229752
rect 408368 229712 408374 229724
rect 411530 229712 411536 229764
rect 411588 229752 411594 229764
rect 570598 229752 570604 229764
rect 411588 229724 570604 229752
rect 411588 229712 411594 229724
rect 570598 229712 570604 229724
rect 570656 229712 570662 229764
rect 140038 229644 140044 229696
rect 140096 229684 140102 229696
rect 205818 229684 205824 229696
rect 140096 229656 205824 229684
rect 140096 229644 140102 229656
rect 205818 229644 205824 229656
rect 205876 229644 205882 229696
rect 227530 229644 227536 229696
rect 227588 229684 227594 229696
rect 267090 229684 267096 229696
rect 227588 229656 267096 229684
rect 227588 229644 227594 229656
rect 267090 229644 267096 229656
rect 267148 229644 267154 229696
rect 268378 229644 268384 229696
rect 268436 229684 268442 229696
rect 277210 229684 277216 229696
rect 268436 229656 277216 229684
rect 268436 229644 268442 229656
rect 277210 229644 277216 229656
rect 277268 229644 277274 229696
rect 277302 229644 277308 229696
rect 277360 229684 277366 229696
rect 277486 229684 277492 229696
rect 277360 229656 277492 229684
rect 277360 229644 277366 229656
rect 277486 229644 277492 229656
rect 277544 229644 277550 229696
rect 277670 229644 277676 229696
rect 277728 229684 277734 229696
rect 285674 229684 285680 229696
rect 277728 229656 285680 229684
rect 277728 229644 277734 229656
rect 285674 229644 285680 229656
rect 285732 229644 285738 229696
rect 318794 229644 318800 229696
rect 318852 229684 318858 229696
rect 334710 229684 334716 229696
rect 318852 229656 334716 229684
rect 318852 229644 318858 229656
rect 334710 229644 334716 229656
rect 334768 229644 334774 229696
rect 340874 229644 340880 229696
rect 340932 229684 340938 229696
rect 380250 229684 380256 229696
rect 340932 229656 380256 229684
rect 340932 229644 340938 229656
rect 380250 229644 380256 229656
rect 380308 229644 380314 229696
rect 391198 229644 391204 229696
rect 391256 229684 391262 229696
rect 392578 229684 392584 229696
rect 391256 229656 392584 229684
rect 391256 229644 391262 229656
rect 392578 229644 392584 229656
rect 392636 229644 392642 229696
rect 400766 229644 400772 229696
rect 400824 229684 400830 229696
rect 453298 229684 453304 229696
rect 400824 229656 453304 229684
rect 400824 229644 400830 229656
rect 453298 229644 453304 229656
rect 453356 229644 453362 229696
rect 151814 229576 151820 229628
rect 151872 229616 151878 229628
rect 218974 229616 218980 229628
rect 151872 229588 218980 229616
rect 151872 229576 151878 229588
rect 218974 229576 218980 229588
rect 219032 229576 219038 229628
rect 248322 229576 248328 229628
rect 248380 229616 248386 229628
rect 248380 229588 258074 229616
rect 248380 229576 248386 229588
rect 149698 229508 149704 229560
rect 149756 229548 149762 229560
rect 216122 229548 216128 229560
rect 149756 229520 216128 229548
rect 149756 229508 149762 229520
rect 216122 229508 216128 229520
rect 216180 229508 216186 229560
rect 244918 229508 244924 229560
rect 244976 229548 244982 229560
rect 254302 229548 254308 229560
rect 244976 229520 254308 229548
rect 244976 229508 244982 229520
rect 254302 229508 254308 229520
rect 254360 229508 254366 229560
rect 258046 229548 258074 229588
rect 260098 229576 260104 229628
rect 260156 229616 260162 229628
rect 262582 229616 262588 229628
rect 260156 229588 262588 229616
rect 260156 229576 260162 229588
rect 262582 229576 262588 229588
rect 262640 229576 262646 229628
rect 270126 229576 270132 229628
rect 270184 229616 270190 229628
rect 271414 229616 271420 229628
rect 270184 229588 271420 229616
rect 270184 229576 270190 229588
rect 271414 229576 271420 229588
rect 271472 229576 271478 229628
rect 275646 229616 275652 229628
rect 271524 229588 275652 229616
rect 271524 229548 271552 229588
rect 275646 229576 275652 229588
rect 275704 229576 275710 229628
rect 280062 229576 280068 229628
rect 280120 229616 280126 229628
rect 288894 229616 288900 229628
rect 280120 229588 288900 229616
rect 280120 229576 280126 229588
rect 288894 229576 288900 229588
rect 288952 229576 288958 229628
rect 313458 229576 313464 229628
rect 313516 229616 313522 229628
rect 314562 229616 314568 229628
rect 313516 229588 314568 229616
rect 313516 229576 313522 229588
rect 314562 229576 314568 229588
rect 314620 229576 314626 229628
rect 328822 229576 328828 229628
rect 328880 229616 328886 229628
rect 329650 229616 329656 229628
rect 328880 229588 329656 229616
rect 328880 229576 328886 229588
rect 329650 229576 329656 229588
rect 329708 229576 329714 229628
rect 330110 229576 330116 229628
rect 330168 229616 330174 229628
rect 334618 229616 334624 229628
rect 330168 229588 334624 229616
rect 330168 229576 330174 229588
rect 334618 229576 334624 229588
rect 334676 229576 334682 229628
rect 338022 229576 338028 229628
rect 338080 229616 338086 229628
rect 338080 229588 345014 229616
rect 338080 229576 338086 229588
rect 258046 229520 271552 229548
rect 272978 229508 272984 229560
rect 273036 229548 273042 229560
rect 281074 229548 281080 229560
rect 273036 229520 281080 229548
rect 273036 229508 273042 229520
rect 281074 229508 281080 229520
rect 281132 229508 281138 229560
rect 300670 229508 300676 229560
rect 300728 229548 300734 229560
rect 305546 229548 305552 229560
rect 300728 229520 305552 229548
rect 300728 229508 300734 229520
rect 305546 229508 305552 229520
rect 305604 229508 305610 229560
rect 327350 229508 327356 229560
rect 327408 229548 327414 229560
rect 341518 229548 341524 229560
rect 327408 229520 341524 229548
rect 327408 229508 327414 229520
rect 341518 229508 341524 229520
rect 341576 229508 341582 229560
rect 344986 229548 345014 229588
rect 350534 229576 350540 229628
rect 350592 229616 350598 229628
rect 388070 229616 388076 229628
rect 350592 229588 388076 229616
rect 350592 229576 350598 229588
rect 388070 229576 388076 229588
rect 388128 229576 388134 229628
rect 397638 229576 397644 229628
rect 397696 229616 397702 229628
rect 398558 229616 398564 229628
rect 397696 229588 398564 229616
rect 397696 229576 397702 229588
rect 398558 229576 398564 229588
rect 398616 229576 398622 229628
rect 398650 229576 398656 229628
rect 398708 229616 398714 229628
rect 404354 229616 404360 229628
rect 398708 229588 404360 229616
rect 398708 229576 398714 229588
rect 404354 229576 404360 229588
rect 404412 229576 404418 229628
rect 407114 229576 407120 229628
rect 407172 229616 407178 229628
rect 407666 229616 407672 229628
rect 407172 229588 407672 229616
rect 407172 229576 407178 229588
rect 407666 229576 407672 229588
rect 407724 229576 407730 229628
rect 407758 229576 407764 229628
rect 407816 229616 407822 229628
rect 449158 229616 449164 229628
rect 407816 229588 449164 229616
rect 407816 229576 407822 229588
rect 449158 229576 449164 229588
rect 449216 229576 449222 229628
rect 352558 229548 352564 229560
rect 344986 229520 352564 229548
rect 352558 229508 352564 229520
rect 352616 229508 352622 229560
rect 366542 229508 366548 229560
rect 366600 229548 366606 229560
rect 416682 229548 416688 229560
rect 366600 229520 416688 229548
rect 366600 229508 366606 229520
rect 416682 229508 416688 229520
rect 416740 229508 416746 229560
rect 146386 229440 146392 229492
rect 146444 229480 146450 229492
rect 209038 229480 209044 229492
rect 146444 229452 209044 229480
rect 146444 229440 146450 229452
rect 209038 229440 209044 229452
rect 209096 229440 209102 229492
rect 275278 229440 275284 229492
rect 275336 229480 275342 229492
rect 283926 229480 283932 229492
rect 275336 229452 283932 229480
rect 275336 229440 275342 229452
rect 283926 229440 283932 229452
rect 283984 229440 283990 229492
rect 339494 229440 339500 229492
rect 339552 229480 339558 229492
rect 353938 229480 353944 229492
rect 339552 229452 353944 229480
rect 339552 229440 339558 229452
rect 353938 229440 353944 229452
rect 353996 229440 354002 229492
rect 355502 229440 355508 229492
rect 355560 229480 355566 229492
rect 386966 229480 386972 229492
rect 355560 229452 386972 229480
rect 355560 229440 355566 229452
rect 386966 229440 386972 229452
rect 387024 229440 387030 229492
rect 393682 229440 393688 229492
rect 393740 229480 393746 229492
rect 400950 229480 400956 229492
rect 393740 229452 400956 229480
rect 393740 229440 393746 229452
rect 400950 229440 400956 229452
rect 401008 229440 401014 229492
rect 401502 229440 401508 229492
rect 401560 229480 401566 229492
rect 404998 229480 405004 229492
rect 401560 229452 405004 229480
rect 401560 229440 401566 229452
rect 404998 229440 405004 229452
rect 405056 229440 405062 229492
rect 405734 229440 405740 229492
rect 405792 229480 405798 229492
rect 441706 229480 441712 229492
rect 405792 229452 441712 229480
rect 405792 229440 405798 229452
rect 441706 229440 441712 229452
rect 441764 229440 441770 229492
rect 186958 229372 186964 229424
rect 187016 229412 187022 229424
rect 248966 229412 248972 229424
rect 187016 229384 248972 229412
rect 187016 229372 187022 229384
rect 248966 229372 248972 229384
rect 249024 229372 249030 229424
rect 273898 229372 273904 229424
rect 273956 229412 273962 229424
rect 282822 229412 282828 229424
rect 273956 229384 282828 229412
rect 273956 229372 273962 229384
rect 282822 229372 282828 229384
rect 282880 229372 282886 229424
rect 298462 229372 298468 229424
rect 298520 229412 298526 229424
rect 301130 229412 301136 229424
rect 298520 229384 301136 229412
rect 298520 229372 298526 229384
rect 301130 229372 301136 229384
rect 301188 229372 301194 229424
rect 332686 229372 332692 229424
rect 332744 229412 332750 229424
rect 333882 229412 333888 229424
rect 332744 229384 333888 229412
rect 332744 229372 332750 229384
rect 333882 229372 333888 229384
rect 333940 229372 333946 229424
rect 334526 229372 334532 229424
rect 334584 229412 334590 229424
rect 342898 229412 342904 229424
rect 334584 229384 342904 229412
rect 334584 229372 334590 229384
rect 342898 229372 342904 229384
rect 342956 229372 342962 229424
rect 361206 229372 361212 229424
rect 361264 229412 361270 229424
rect 383102 229412 383108 229424
rect 361264 229384 383108 229412
rect 361264 229372 361270 229384
rect 383102 229372 383108 229384
rect 383160 229372 383166 229424
rect 392210 229372 392216 229424
rect 392268 229412 392274 229424
rect 430758 229412 430764 229424
rect 392268 229384 430764 229412
rect 392268 229372 392274 229384
rect 430758 229372 430764 229384
rect 430816 229372 430822 229424
rect 162854 229304 162860 229356
rect 162912 229344 162918 229356
rect 223298 229344 223304 229356
rect 162912 229316 223304 229344
rect 162912 229304 162918 229316
rect 223298 229304 223304 229316
rect 223356 229304 223362 229356
rect 277486 229304 277492 229356
rect 277544 229344 277550 229356
rect 286686 229344 286692 229356
rect 277544 229316 286692 229344
rect 277544 229304 277550 229316
rect 286686 229304 286692 229316
rect 286744 229304 286750 229356
rect 295242 229304 295248 229356
rect 295300 229344 295306 229356
rect 296898 229344 296904 229356
rect 295300 229316 296904 229344
rect 295300 229304 295306 229316
rect 296898 229304 296904 229316
rect 296956 229304 296962 229356
rect 331306 229304 331312 229356
rect 331364 229344 331370 229356
rect 332226 229344 332232 229356
rect 331364 229316 332232 229344
rect 331364 229304 331370 229316
rect 332226 229304 332232 229316
rect 332284 229304 332290 229356
rect 342346 229304 342352 229356
rect 342404 229344 342410 229356
rect 343266 229344 343272 229356
rect 342404 229316 343272 229344
rect 342404 229304 342410 229316
rect 343266 229304 343272 229316
rect 343324 229304 343330 229356
rect 371970 229304 371976 229356
rect 372028 229344 372034 229356
rect 398650 229344 398656 229356
rect 372028 229316 398656 229344
rect 372028 229304 372034 229316
rect 398650 229304 398656 229316
rect 398708 229304 398714 229356
rect 402974 229304 402980 229356
rect 403032 229344 403038 229356
rect 404262 229344 404268 229356
rect 403032 229316 404268 229344
rect 403032 229304 403038 229316
rect 404262 229304 404268 229316
rect 404320 229304 404326 229356
rect 404722 229304 404728 229356
rect 404780 229344 404786 229356
rect 409782 229344 409788 229356
rect 404780 229316 409788 229344
rect 404780 229304 404786 229316
rect 409782 229304 409788 229316
rect 409840 229304 409846 229356
rect 410058 229304 410064 229356
rect 410116 229344 410122 229356
rect 435542 229344 435548 229356
rect 410116 229316 435548 229344
rect 410116 229304 410122 229316
rect 435542 229304 435548 229316
rect 435600 229304 435606 229356
rect 180794 229236 180800 229288
rect 180852 229276 180858 229288
rect 238938 229276 238944 229288
rect 180852 229248 238944 229276
rect 180852 229236 180858 229248
rect 238938 229236 238944 229248
rect 238996 229236 239002 229288
rect 271230 229236 271236 229288
rect 271288 229276 271294 229288
rect 279970 229276 279976 229288
rect 271288 229248 279976 229276
rect 271288 229236 271294 229248
rect 279970 229236 279976 229248
rect 280028 229236 280034 229288
rect 281442 229236 281448 229288
rect 281500 229276 281506 229288
rect 288158 229276 288164 229288
rect 281500 229248 288164 229276
rect 281500 229236 281506 229248
rect 288158 229236 288164 229248
rect 288216 229236 288222 229288
rect 313090 229236 313096 229288
rect 313148 229276 313154 229288
rect 318058 229276 318064 229288
rect 313148 229248 318064 229276
rect 313148 229236 313154 229248
rect 318058 229236 318064 229248
rect 318116 229236 318122 229288
rect 357710 229236 357716 229288
rect 357768 229276 357774 229288
rect 376110 229276 376116 229288
rect 357768 229248 376116 229276
rect 357768 229236 357774 229248
rect 376110 229236 376116 229248
rect 376168 229236 376174 229288
rect 384390 229236 384396 229288
rect 384448 229276 384454 229288
rect 411346 229276 411352 229288
rect 384448 229248 411352 229276
rect 384448 229236 384454 229248
rect 411346 229236 411352 229248
rect 411404 229236 411410 229288
rect 255958 229168 255964 229220
rect 256016 229208 256022 229220
rect 260006 229208 260012 229220
rect 256016 229180 260012 229208
rect 256016 229168 256022 229180
rect 260006 229168 260012 229180
rect 260064 229168 260070 229220
rect 282822 229168 282828 229220
rect 282880 229208 282886 229220
rect 289262 229208 289268 229220
rect 282880 229180 289268 229208
rect 282880 229168 282886 229180
rect 289262 229168 289268 229180
rect 289320 229168 289326 229220
rect 296346 229168 296352 229220
rect 296404 229208 296410 229220
rect 298462 229208 298468 229220
rect 296404 229180 298468 229208
rect 296404 229168 296410 229180
rect 298462 229168 298468 229180
rect 298520 229168 298526 229220
rect 369394 229168 369400 229220
rect 369452 229208 369458 229220
rect 378594 229208 378600 229220
rect 369452 229180 378600 229208
rect 369452 229168 369458 229180
rect 378594 229168 378600 229180
rect 378652 229168 378658 229220
rect 395062 229168 395068 229220
rect 395120 229208 395126 229220
rect 408402 229208 408408 229220
rect 395120 229180 408408 229208
rect 395120 229168 395126 229180
rect 408402 229168 408408 229180
rect 408460 229168 408466 229220
rect 409322 229168 409328 229220
rect 409380 229208 409386 229220
rect 409380 229180 411392 229208
rect 409380 229168 409386 229180
rect 67542 229140 67548 229152
rect 63512 229112 67548 229140
rect 62114 229032 62120 229084
rect 62172 229072 62178 229084
rect 63512 229072 63540 229112
rect 67542 229100 67548 229112
rect 67600 229100 67606 229152
rect 257338 229100 257344 229152
rect 257396 229140 257402 229152
rect 258902 229140 258908 229152
rect 257396 229112 258908 229140
rect 257396 229100 257402 229112
rect 258902 229100 258908 229112
rect 258960 229100 258966 229152
rect 284110 229100 284116 229152
rect 284168 229140 284174 229152
rect 289538 229140 289544 229152
rect 284168 229112 289544 229140
rect 284168 229100 284174 229112
rect 289538 229100 289544 229112
rect 289596 229100 289602 229152
rect 405090 229100 405096 229152
rect 405148 229140 405154 229152
rect 411254 229140 411260 229152
rect 405148 229112 411260 229140
rect 405148 229100 405154 229112
rect 411254 229100 411260 229112
rect 411312 229100 411318 229152
rect 411364 229140 411392 229180
rect 411898 229168 411904 229220
rect 411956 229208 411962 229220
rect 420178 229208 420184 229220
rect 411956 229180 420184 229208
rect 411956 229168 411962 229180
rect 420178 229168 420184 229180
rect 420236 229168 420242 229220
rect 551278 229140 551284 229152
rect 411364 229112 551284 229140
rect 551278 229100 551284 229112
rect 551336 229100 551342 229152
rect 62172 229044 63540 229072
rect 62172 229032 62178 229044
rect 120810 229032 120816 229084
rect 120868 229072 120874 229084
rect 220814 229072 220820 229084
rect 120868 229044 220820 229072
rect 120868 229032 120874 229044
rect 220814 229032 220820 229044
rect 220872 229032 220878 229084
rect 365162 229032 365168 229084
rect 365220 229072 365226 229084
rect 460934 229072 460940 229084
rect 365220 229044 460940 229072
rect 365220 229032 365226 229044
rect 460934 229032 460940 229044
rect 460992 229032 460998 229084
rect 117222 228964 117228 229016
rect 117280 229004 117286 229016
rect 219342 229004 219348 229016
rect 117280 228976 219348 229004
rect 117280 228964 117286 228976
rect 219342 228964 219348 228976
rect 219400 228964 219406 229016
rect 332042 228964 332048 229016
rect 332100 229004 332106 229016
rect 370222 229004 370228 229016
rect 332100 228976 370228 229004
rect 332100 228964 332106 228976
rect 370222 228964 370228 228976
rect 370280 228964 370286 229016
rect 373350 228964 373356 229016
rect 373408 229004 373414 229016
rect 480254 229004 480260 229016
rect 373408 228976 480260 229004
rect 373408 228964 373414 228976
rect 480254 228964 480260 228976
rect 480312 228964 480318 229016
rect 114186 228896 114192 228948
rect 114244 228936 114250 228948
rect 217962 228936 217968 228948
rect 114244 228908 217968 228936
rect 114244 228896 114250 228908
rect 217962 228896 217968 228908
rect 218020 228896 218026 228948
rect 224034 228896 224040 228948
rect 224092 228936 224098 228948
rect 234706 228936 234712 228948
rect 224092 228908 234712 228936
rect 224092 228896 224098 228908
rect 234706 228896 234712 228908
rect 234764 228896 234770 228948
rect 329190 228896 329196 228948
rect 329248 228936 329254 228948
rect 371326 228936 371332 228948
rect 329248 228908 371332 228936
rect 329248 228896 329254 228908
rect 371326 228896 371332 228908
rect 371384 228896 371390 228948
rect 375098 228896 375104 228948
rect 375156 228936 375162 228948
rect 483474 228936 483480 228948
rect 375156 228908 483480 228936
rect 375156 228896 375162 228908
rect 483474 228896 483480 228908
rect 483532 228896 483538 228948
rect 110690 228828 110696 228880
rect 110748 228868 110754 228880
rect 216490 228868 216496 228880
rect 110748 228840 216496 228868
rect 110748 228828 110754 228840
rect 216490 228828 216496 228840
rect 216548 228828 216554 228880
rect 227714 228828 227720 228880
rect 227772 228868 227778 228880
rect 240410 228868 240416 228880
rect 227772 228840 240416 228868
rect 227772 228828 227778 228840
rect 240410 228828 240416 228840
rect 240468 228828 240474 228880
rect 327718 228828 327724 228880
rect 327776 228868 327782 228880
rect 372706 228868 372712 228880
rect 327776 228840 372712 228868
rect 327776 228828 327782 228840
rect 372706 228828 372712 228840
rect 372764 228828 372770 228880
rect 376570 228828 376576 228880
rect 376628 228868 376634 228880
rect 487706 228868 487712 228880
rect 376628 228840 487712 228868
rect 376628 228828 376634 228840
rect 487706 228828 487712 228840
rect 487764 228828 487770 228880
rect 107470 228760 107476 228812
rect 107528 228800 107534 228812
rect 215110 228800 215116 228812
rect 107528 228772 215116 228800
rect 107528 228760 107534 228772
rect 215110 228760 215116 228772
rect 215168 228760 215174 228812
rect 216674 228760 216680 228812
rect 216732 228800 216738 228812
rect 224678 228800 224684 228812
rect 216732 228772 224684 228800
rect 216732 228760 216738 228772
rect 224678 228760 224684 228772
rect 224736 228760 224742 228812
rect 230290 228760 230296 228812
rect 230348 228800 230354 228812
rect 230348 228772 230612 228800
rect 230348 228760 230354 228772
rect 103974 228692 103980 228744
rect 104032 228732 104038 228744
rect 213638 228732 213644 228744
rect 104032 228704 213644 228732
rect 104032 228692 104038 228704
rect 213638 228692 213644 228704
rect 213696 228692 213702 228744
rect 222102 228692 222108 228744
rect 222160 228732 222166 228744
rect 230382 228732 230388 228744
rect 222160 228704 230388 228732
rect 222160 228692 222166 228704
rect 230382 228692 230388 228704
rect 230440 228692 230446 228744
rect 230584 228732 230612 228772
rect 233510 228760 233516 228812
rect 233568 228800 233574 228812
rect 268194 228800 268200 228812
rect 233568 228772 268200 228800
rect 233568 228760 233574 228772
rect 268194 228760 268200 228772
rect 268252 228760 268258 228812
rect 330570 228760 330576 228812
rect 330628 228800 330634 228812
rect 375282 228800 375288 228812
rect 330628 228772 375288 228800
rect 330628 228760 330634 228772
rect 375282 228760 375288 228772
rect 375340 228760 375346 228812
rect 377950 228760 377956 228812
rect 378008 228800 378014 228812
rect 491294 228800 491300 228812
rect 378008 228772 491300 228800
rect 378008 228760 378014 228772
rect 491294 228760 491300 228772
rect 491352 228760 491358 228812
rect 266722 228732 266728 228744
rect 230584 228704 266728 228732
rect 266722 228692 266728 228704
rect 266780 228692 266786 228744
rect 328086 228692 328092 228744
rect 328144 228732 328150 228744
rect 373994 228732 374000 228744
rect 328144 228704 374000 228732
rect 328144 228692 328150 228704
rect 373994 228692 374000 228704
rect 374052 228692 374058 228744
rect 391934 228692 391940 228744
rect 391992 228732 391998 228744
rect 523034 228732 523040 228744
rect 391992 228704 523040 228732
rect 391992 228692 391998 228704
rect 523034 228692 523040 228704
rect 523092 228692 523098 228744
rect 100662 228624 100668 228676
rect 100720 228664 100726 228676
rect 212258 228664 212264 228676
rect 100720 228636 212264 228664
rect 100720 228624 100726 228636
rect 212258 228624 212264 228636
rect 212316 228624 212322 228676
rect 215110 228624 215116 228676
rect 215168 228664 215174 228676
rect 260742 228664 260748 228676
rect 215168 228636 260748 228664
rect 215168 228624 215174 228636
rect 260742 228624 260748 228636
rect 260800 228624 260806 228676
rect 334894 228624 334900 228676
rect 334952 228664 334958 228676
rect 389266 228664 389272 228676
rect 334952 228636 389272 228664
rect 334952 228624 334958 228636
rect 389266 228624 389272 228636
rect 389324 228624 389330 228676
rect 392946 228624 392952 228676
rect 393004 228664 393010 228676
rect 526346 228664 526352 228676
rect 393004 228636 526352 228664
rect 393004 228624 393010 228636
rect 526346 228624 526352 228636
rect 526404 228624 526410 228676
rect 97258 228556 97264 228608
rect 97316 228596 97322 228608
rect 210786 228596 210792 228608
rect 97316 228568 210792 228596
rect 97316 228556 97322 228568
rect 210786 228556 210792 228568
rect 210844 228556 210850 228608
rect 213822 228556 213828 228608
rect 213880 228596 213886 228608
rect 258534 228596 258540 228608
rect 213880 228568 258540 228596
rect 213880 228556 213886 228568
rect 258534 228556 258540 228568
rect 258592 228556 258598 228608
rect 336274 228556 336280 228608
rect 336332 228596 336338 228608
rect 392486 228596 392492 228608
rect 336332 228568 392492 228596
rect 336332 228556 336338 228568
rect 392486 228556 392492 228568
rect 392544 228556 392550 228608
rect 398282 228556 398288 228608
rect 398340 228596 398346 228608
rect 538214 228596 538220 228608
rect 398340 228568 538220 228596
rect 398340 228556 398346 228568
rect 538214 228556 538220 228568
rect 538272 228556 538278 228608
rect 77938 228488 77944 228540
rect 77996 228528 78002 228540
rect 91738 228528 91744 228540
rect 77996 228500 91744 228528
rect 77996 228488 78002 228500
rect 91738 228488 91744 228500
rect 91796 228488 91802 228540
rect 93762 228488 93768 228540
rect 93820 228528 93826 228540
rect 209406 228528 209412 228540
rect 93820 228500 209412 228528
rect 93820 228488 93826 228500
rect 209406 228488 209412 228500
rect 209464 228488 209470 228540
rect 209866 228488 209872 228540
rect 209924 228528 209930 228540
rect 257154 228528 257160 228540
rect 209924 228500 257160 228528
rect 209924 228488 209930 228500
rect 257154 228488 257160 228500
rect 257212 228488 257218 228540
rect 306650 228488 306656 228540
rect 306708 228528 306714 228540
rect 323670 228528 323676 228540
rect 306708 228500 323676 228528
rect 306708 228488 306714 228500
rect 323670 228488 323676 228500
rect 323728 228488 323734 228540
rect 337746 228488 337752 228540
rect 337804 228528 337810 228540
rect 396166 228528 396172 228540
rect 337804 228500 396172 228528
rect 337804 228488 337810 228500
rect 396166 228488 396172 228500
rect 396224 228488 396230 228540
rect 397270 228488 397276 228540
rect 397328 228528 397334 228540
rect 536834 228528 536840 228540
rect 397328 228500 536840 228528
rect 397328 228488 397334 228500
rect 536834 228488 536840 228500
rect 536892 228488 536898 228540
rect 54386 228420 54392 228472
rect 54444 228460 54450 228472
rect 193306 228460 193312 228472
rect 54444 228432 193312 228460
rect 54444 228420 54450 228432
rect 193306 228420 193312 228432
rect 193364 228420 193370 228472
rect 194962 228420 194968 228472
rect 195020 228460 195026 228472
rect 252186 228460 252192 228472
rect 195020 228432 252192 228460
rect 195020 228420 195026 228432
rect 252186 228420 252192 228432
rect 252244 228420 252250 228472
rect 276382 228460 276388 228472
rect 258046 228432 276388 228460
rect 53650 228352 53656 228404
rect 53708 228392 53714 228404
rect 192294 228392 192300 228404
rect 53708 228364 192300 228392
rect 53708 228352 53714 228364
rect 192294 228352 192300 228364
rect 192352 228352 192358 228404
rect 194134 228352 194140 228404
rect 194192 228392 194198 228404
rect 252830 228392 252836 228404
rect 194192 228364 252836 228392
rect 194192 228352 194198 228364
rect 252830 228352 252836 228364
rect 252888 228352 252894 228404
rect 127526 228284 127532 228336
rect 127584 228324 127590 228336
rect 223666 228324 223672 228336
rect 127584 228296 223672 228324
rect 127584 228284 127590 228296
rect 223666 228284 223672 228296
rect 223724 228284 223730 228336
rect 252002 228284 252008 228336
rect 252060 228324 252066 228336
rect 258046 228324 258074 228432
rect 276382 228420 276388 228432
rect 276440 228420 276446 228472
rect 309870 228420 309876 228472
rect 309928 228460 309934 228472
rect 327810 228460 327816 228472
rect 309928 228432 327816 228460
rect 309928 228420 309934 228432
rect 327810 228420 327816 228432
rect 327868 228420 327874 228472
rect 340598 228420 340604 228472
rect 340656 228460 340662 228472
rect 402974 228460 402980 228472
rect 340656 228432 402980 228460
rect 340656 228420 340662 228432
rect 402974 228420 402980 228432
rect 403032 228420 403038 228472
rect 409782 228420 409788 228472
rect 409840 228460 409846 228472
rect 553946 228460 553952 228472
rect 409840 228432 553952 228460
rect 409840 228420 409846 228432
rect 553946 228420 553952 228432
rect 554004 228420 554010 228472
rect 260558 228352 260564 228404
rect 260616 228392 260622 228404
rect 279602 228392 279608 228404
rect 260616 228364 279608 228392
rect 260616 228352 260622 228364
rect 279602 228352 279608 228364
rect 279660 228352 279666 228404
rect 308122 228352 308128 228404
rect 308180 228392 308186 228404
rect 327074 228392 327080 228404
rect 308180 228364 327080 228392
rect 308180 228352 308186 228364
rect 327074 228352 327080 228364
rect 327132 228352 327138 228404
rect 345198 228352 345204 228404
rect 345256 228392 345262 228404
rect 408494 228392 408500 228404
rect 345256 228364 408500 228392
rect 345256 228352 345262 228364
rect 408494 228352 408500 228364
rect 408552 228352 408558 228404
rect 410794 228352 410800 228404
rect 410852 228392 410858 228404
rect 569126 228392 569132 228404
rect 410852 228364 569132 228392
rect 410852 228352 410858 228364
rect 569126 228352 569132 228364
rect 569184 228352 569190 228404
rect 252060 228296 258074 228324
rect 252060 228284 252066 228296
rect 353386 228284 353392 228336
rect 353444 228324 353450 228336
rect 433334 228324 433340 228336
rect 353444 228296 433340 228324
rect 353444 228284 353450 228296
rect 433334 228284 433340 228296
rect 433392 228284 433398 228336
rect 131022 228216 131028 228268
rect 131080 228256 131086 228268
rect 225046 228256 225052 228268
rect 131080 228228 225052 228256
rect 131080 228216 131086 228228
rect 225046 228216 225052 228228
rect 225104 228216 225110 228268
rect 349154 228216 349160 228268
rect 349212 228256 349218 228268
rect 423030 228256 423036 228268
rect 349212 228228 423036 228256
rect 349212 228216 349218 228228
rect 423030 228216 423036 228228
rect 423088 228216 423094 228268
rect 137738 228148 137744 228200
rect 137796 228188 137802 228200
rect 227898 228188 227904 228200
rect 137796 228160 227904 228188
rect 137796 228148 137802 228160
rect 227898 228148 227904 228160
rect 227956 228148 227962 228200
rect 334158 228148 334164 228200
rect 334216 228188 334222 228200
rect 378502 228188 378508 228200
rect 334216 228160 378508 228188
rect 334216 228148 334222 228160
rect 378502 228148 378508 228160
rect 378560 228148 378566 228200
rect 378962 228148 378968 228200
rect 379020 228188 379026 228200
rect 399386 228188 399392 228200
rect 379020 228160 399392 228188
rect 379020 228148 379026 228160
rect 399386 228148 399392 228160
rect 399444 228148 399450 228200
rect 404354 228148 404360 228200
rect 404412 228188 404418 228200
rect 476114 228188 476120 228200
rect 404412 228160 476120 228188
rect 404412 228148 404418 228160
rect 476114 228148 476120 228160
rect 476172 228148 476178 228200
rect 144362 228080 144368 228132
rect 144420 228120 144426 228132
rect 230750 228120 230756 228132
rect 144420 228092 230756 228120
rect 144420 228080 144426 228092
rect 230750 228080 230756 228092
rect 230808 228080 230814 228132
rect 346302 228080 346308 228132
rect 346360 228120 346366 228132
rect 409966 228120 409972 228132
rect 346360 228092 409972 228120
rect 346360 228080 346366 228092
rect 409966 228080 409972 228092
rect 410024 228080 410030 228132
rect 420178 228080 420184 228132
rect 420236 228120 420242 228132
rect 485130 228120 485136 228132
rect 420236 228092 485136 228120
rect 420236 228080 420242 228092
rect 485130 228080 485136 228092
rect 485188 228080 485194 228132
rect 154482 228012 154488 228064
rect 154540 228052 154546 228064
rect 235074 228052 235080 228064
rect 154540 228024 235080 228052
rect 154540 228012 154546 228024
rect 235074 228012 235080 228024
rect 235132 228012 235138 228064
rect 343450 228012 343456 228064
rect 343508 228052 343514 228064
rect 387242 228052 387248 228064
rect 343508 228024 387248 228052
rect 343508 228012 343514 228024
rect 387242 228012 387248 228024
rect 387300 228012 387306 228064
rect 406470 228012 406476 228064
rect 406528 228052 406534 228064
rect 454034 228052 454040 228064
rect 406528 228024 454040 228052
rect 406528 228012 406534 228024
rect 454034 228012 454040 228024
rect 454092 228012 454098 228064
rect 161290 227944 161296 227996
rect 161348 227984 161354 227996
rect 237926 227984 237932 227996
rect 161348 227956 237932 227984
rect 161348 227944 161354 227956
rect 237926 227944 237932 227956
rect 237984 227944 237990 227996
rect 388070 227944 388076 227996
rect 388128 227984 388134 227996
rect 426434 227984 426440 227996
rect 388128 227956 426440 227984
rect 388128 227944 388134 227956
rect 426434 227944 426440 227956
rect 426492 227944 426498 227996
rect 171042 227876 171048 227928
rect 171100 227916 171106 227928
rect 242158 227916 242164 227928
rect 171100 227888 242164 227916
rect 171100 227876 171106 227888
rect 242158 227876 242164 227888
rect 242216 227876 242222 227928
rect 387610 227876 387616 227928
rect 387668 227916 387674 227928
rect 419534 227916 419540 227928
rect 387668 227888 419540 227916
rect 387668 227876 387674 227888
rect 419534 227876 419540 227888
rect 419592 227876 419598 227928
rect 403066 227808 403072 227860
rect 403124 227848 403130 227860
rect 429654 227848 429660 227860
rect 403124 227820 429660 227848
rect 403124 227808 403130 227820
rect 429654 227808 429660 227820
rect 429712 227808 429718 227860
rect 375466 227740 375472 227792
rect 375524 227780 375530 227792
rect 379698 227780 379704 227792
rect 375524 227752 379704 227780
rect 375524 227740 375530 227752
rect 379698 227740 379704 227752
rect 379756 227740 379762 227792
rect 380434 227740 380440 227792
rect 380492 227780 380498 227792
rect 406102 227780 406108 227792
rect 380492 227752 406108 227780
rect 380492 227740 380498 227752
rect 406102 227740 406108 227752
rect 406160 227740 406166 227792
rect 160370 227672 160376 227724
rect 160428 227712 160434 227724
rect 238570 227712 238576 227724
rect 160428 227684 238576 227712
rect 160428 227672 160434 227684
rect 238570 227672 238576 227684
rect 238628 227672 238634 227724
rect 364426 227672 364432 227724
rect 364484 227712 364490 227724
rect 457346 227712 457352 227724
rect 364484 227684 457352 227712
rect 364484 227672 364490 227684
rect 457346 227672 457352 227684
rect 457404 227672 457410 227724
rect 157058 227604 157064 227656
rect 157116 227644 157122 227656
rect 237190 227644 237196 227656
rect 157116 227616 237196 227644
rect 157116 227604 157122 227616
rect 237190 227604 237196 227616
rect 237248 227604 237254 227656
rect 360194 227604 360200 227656
rect 360252 227644 360258 227656
rect 447318 227644 447324 227656
rect 360252 227616 447324 227644
rect 360252 227604 360258 227616
rect 447318 227604 447324 227616
rect 447376 227604 447382 227656
rect 449158 227604 449164 227656
rect 449216 227644 449222 227656
rect 542998 227644 543004 227656
rect 449216 227616 543004 227644
rect 449216 227604 449222 227616
rect 542998 227604 543004 227616
rect 543056 227604 543062 227656
rect 153654 227536 153660 227588
rect 153712 227576 153718 227588
rect 235718 227576 235724 227588
rect 153712 227548 235724 227576
rect 153712 227536 153718 227548
rect 235718 227536 235724 227548
rect 235776 227536 235782 227588
rect 365898 227536 365904 227588
rect 365956 227576 365962 227588
rect 461210 227576 461216 227588
rect 365956 227548 461216 227576
rect 365956 227536 365962 227548
rect 461210 227536 461216 227548
rect 461268 227536 461274 227588
rect 461578 227536 461584 227588
rect 461636 227576 461642 227588
rect 552658 227576 552664 227588
rect 461636 227548 552664 227576
rect 461636 227536 461642 227548
rect 552658 227536 552664 227548
rect 552716 227536 552722 227588
rect 108206 227468 108212 227520
rect 108264 227508 108270 227520
rect 149698 227508 149704 227520
rect 108264 227480 149704 227508
rect 108264 227468 108270 227480
rect 149698 227468 149704 227480
rect 149756 227468 149762 227520
rect 150342 227468 150348 227520
rect 150400 227508 150406 227520
rect 234338 227508 234344 227520
rect 150400 227480 234344 227508
rect 150400 227468 150406 227480
rect 234338 227468 234344 227480
rect 234396 227468 234402 227520
rect 367278 227468 367284 227520
rect 367336 227508 367342 227520
rect 464154 227508 464160 227520
rect 367336 227480 464160 227508
rect 367336 227468 367342 227480
rect 464154 227468 464160 227480
rect 464212 227468 464218 227520
rect 147490 227400 147496 227452
rect 147548 227440 147554 227452
rect 232222 227440 232228 227452
rect 147548 227412 232228 227440
rect 147548 227400 147554 227412
rect 232222 227400 232228 227412
rect 232280 227400 232286 227452
rect 309502 227400 309508 227452
rect 309560 227440 309566 227452
rect 330386 227440 330392 227452
rect 309560 227412 330392 227440
rect 309560 227400 309566 227412
rect 330386 227400 330392 227412
rect 330444 227400 330450 227452
rect 368750 227400 368756 227452
rect 368808 227440 368814 227452
rect 467834 227440 467840 227452
rect 368808 227412 467840 227440
rect 368808 227400 368814 227412
rect 467834 227400 467840 227412
rect 467892 227400 467898 227452
rect 468478 227400 468484 227452
rect 468536 227440 468542 227452
rect 554958 227440 554964 227452
rect 468536 227412 554964 227440
rect 468536 227400 468542 227412
rect 554958 227400 554964 227412
rect 555016 227400 555022 227452
rect 91370 227332 91376 227384
rect 91428 227372 91434 227384
rect 146386 227372 146392 227384
rect 91428 227344 146392 227372
rect 91428 227332 91434 227344
rect 146386 227332 146392 227344
rect 146444 227332 146450 227384
rect 146938 227332 146944 227384
rect 146996 227372 147002 227384
rect 232866 227372 232872 227384
rect 146996 227344 232872 227372
rect 146996 227332 147002 227344
rect 232866 227332 232872 227344
rect 232924 227332 232930 227384
rect 315574 227332 315580 227384
rect 315632 227372 315638 227384
rect 341334 227372 341340 227384
rect 315632 227344 341340 227372
rect 315632 227332 315638 227344
rect 341334 227332 341340 227344
rect 341392 227332 341398 227384
rect 370130 227332 370136 227384
rect 370188 227372 370194 227384
rect 470870 227372 470876 227384
rect 370188 227344 470876 227372
rect 370188 227332 370194 227344
rect 470870 227332 470876 227344
rect 470928 227332 470934 227384
rect 141050 227264 141056 227316
rect 141108 227304 141114 227316
rect 229370 227304 229376 227316
rect 141108 227276 229376 227304
rect 141108 227264 141114 227276
rect 229370 227264 229376 227276
rect 229428 227264 229434 227316
rect 312722 227264 312728 227316
rect 312780 227304 312786 227316
rect 333974 227304 333980 227316
rect 312780 227276 333980 227304
rect 312780 227264 312786 227276
rect 333974 227264 333980 227276
rect 334032 227264 334038 227316
rect 335170 227264 335176 227316
rect 335228 227304 335234 227316
rect 363138 227304 363144 227316
rect 335228 227276 363144 227304
rect 335228 227264 335234 227276
rect 363138 227264 363144 227276
rect 363196 227264 363202 227316
rect 371602 227264 371608 227316
rect 371660 227304 371666 227316
rect 474182 227304 474188 227316
rect 371660 227276 474188 227304
rect 371660 227264 371666 227276
rect 474182 227264 474188 227276
rect 474240 227264 474246 227316
rect 143442 227196 143448 227248
rect 143500 227236 143506 227248
rect 231486 227236 231492 227248
rect 143500 227208 231492 227236
rect 143500 227196 143506 227208
rect 231486 227196 231492 227208
rect 231544 227196 231550 227248
rect 232774 227196 232780 227248
rect 232832 227236 232838 227248
rect 247494 227236 247500 227248
rect 232832 227208 247500 227236
rect 232832 227196 232838 227208
rect 247494 227196 247500 227208
rect 247552 227196 247558 227248
rect 318426 227196 318432 227248
rect 318484 227236 318490 227248
rect 348050 227236 348056 227248
rect 318484 227208 348056 227236
rect 318484 227196 318490 227208
rect 348050 227196 348056 227208
rect 348108 227196 348114 227248
rect 372982 227196 372988 227248
rect 373040 227236 373046 227248
rect 477586 227236 477592 227248
rect 373040 227208 477592 227236
rect 373040 227196 373046 227208
rect 477586 227196 477592 227208
rect 477644 227196 477650 227248
rect 478138 227196 478144 227248
rect 478196 227236 478202 227248
rect 489362 227236 489368 227248
rect 478196 227208 489368 227236
rect 478196 227196 478202 227208
rect 489362 227196 489368 227208
rect 489420 227196 489426 227248
rect 82722 227128 82728 227180
rect 82780 227168 82786 227180
rect 140038 227168 140044 227180
rect 82780 227140 140044 227168
rect 82780 227128 82786 227140
rect 140038 227128 140044 227140
rect 140096 227128 140102 227180
rect 140130 227128 140136 227180
rect 140188 227168 140194 227180
rect 230014 227168 230020 227180
rect 140188 227140 230020 227168
rect 140188 227128 140194 227140
rect 230014 227128 230020 227140
rect 230072 227128 230078 227180
rect 237374 227128 237380 227180
rect 237432 227168 237438 227180
rect 256050 227168 256056 227180
rect 237432 227140 256056 227168
rect 237432 227128 237438 227140
rect 256050 227128 256056 227140
rect 256108 227128 256114 227180
rect 258810 227128 258816 227180
rect 258868 227168 258874 227180
rect 279234 227168 279240 227180
rect 258868 227140 279240 227168
rect 258868 227128 258874 227140
rect 279234 227128 279240 227140
rect 279292 227128 279298 227180
rect 321278 227128 321284 227180
rect 321336 227168 321342 227180
rect 354766 227168 354772 227180
rect 321336 227140 354772 227168
rect 321336 227128 321342 227140
rect 354766 227128 354772 227140
rect 354824 227128 354830 227180
rect 374454 227128 374460 227180
rect 374512 227168 374518 227180
rect 480898 227168 480904 227180
rect 374512 227140 480904 227168
rect 374512 227128 374518 227140
rect 480898 227128 480904 227140
rect 480956 227128 480962 227180
rect 134242 227060 134248 227112
rect 134300 227100 134306 227112
rect 226518 227100 226524 227112
rect 134300 227072 226524 227100
rect 134300 227060 134306 227072
rect 226518 227060 226524 227072
rect 226576 227060 226582 227112
rect 234706 227060 234712 227112
rect 234764 227100 234770 227112
rect 253198 227100 253204 227112
rect 234764 227072 253204 227100
rect 234764 227060 234770 227072
rect 253198 227060 253204 227072
rect 253256 227060 253262 227112
rect 255130 227060 255136 227112
rect 255188 227100 255194 227112
rect 277854 227100 277860 227112
rect 255188 227072 277860 227100
rect 255188 227060 255194 227072
rect 277854 227060 277860 227072
rect 277912 227060 277918 227112
rect 325602 227060 325608 227112
rect 325660 227100 325666 227112
rect 360286 227100 360292 227112
rect 325660 227072 360292 227100
rect 325660 227060 325666 227072
rect 360286 227060 360292 227072
rect 360344 227060 360350 227112
rect 374822 227060 374828 227112
rect 374880 227100 374886 227112
rect 483106 227100 483112 227112
rect 374880 227072 483112 227100
rect 374880 227060 374886 227072
rect 483106 227060 483112 227072
rect 483164 227060 483170 227112
rect 124122 226992 124128 227044
rect 124180 227032 124186 227044
rect 222194 227032 222200 227044
rect 124180 227004 222200 227032
rect 124180 226992 124186 227004
rect 222194 226992 222200 227004
rect 222252 226992 222258 227044
rect 237006 226992 237012 227044
rect 237064 227032 237070 227044
rect 269574 227032 269580 227044
rect 237064 227004 269580 227032
rect 237064 226992 237070 227004
rect 269574 226992 269580 227004
rect 269632 226992 269638 227044
rect 305270 226992 305276 227044
rect 305328 227032 305334 227044
rect 320266 227032 320272 227044
rect 305328 227004 320272 227032
rect 305328 226992 305334 227004
rect 320266 226992 320272 227004
rect 320324 226992 320330 227044
rect 329466 226992 329472 227044
rect 329524 227032 329530 227044
rect 365346 227032 365352 227044
rect 329524 227004 365352 227032
rect 329524 226992 329530 227004
rect 365346 226992 365352 227004
rect 365404 226992 365410 227044
rect 409690 226992 409696 227044
rect 409748 227032 409754 227044
rect 565906 227032 565912 227044
rect 409748 227004 565912 227032
rect 409748 226992 409754 227004
rect 565906 226992 565912 227004
rect 565964 226992 565970 227044
rect 125042 226924 125048 226976
rect 125100 226964 125106 226976
rect 162854 226964 162860 226976
rect 125100 226936 162860 226964
rect 125100 226924 125106 226936
rect 162854 226924 162860 226936
rect 162912 226924 162918 226976
rect 163682 226924 163688 226976
rect 163740 226964 163746 226976
rect 239766 226964 239772 226976
rect 163740 226936 239772 226964
rect 163740 226924 163746 226936
rect 239766 226924 239772 226936
rect 239824 226924 239830 226976
rect 363046 226924 363052 226976
rect 363104 226964 363110 226976
rect 454126 226964 454132 226976
rect 363104 226936 454132 226964
rect 363104 226924 363110 226936
rect 454126 226924 454132 226936
rect 454184 226924 454190 226976
rect 166902 226856 166908 226908
rect 166960 226896 166966 226908
rect 241422 226896 241428 226908
rect 166960 226868 241428 226896
rect 166960 226856 166966 226868
rect 241422 226856 241428 226868
rect 241480 226856 241486 226908
rect 361574 226856 361580 226908
rect 361632 226896 361638 226908
rect 450630 226896 450636 226908
rect 361632 226868 450636 226896
rect 361632 226856 361638 226868
rect 450630 226856 450636 226868
rect 450688 226856 450694 226908
rect 164602 226788 164608 226840
rect 164660 226828 164666 226840
rect 239306 226828 239312 226840
rect 164660 226800 239312 226828
rect 164660 226788 164666 226800
rect 239306 226788 239312 226800
rect 239364 226788 239370 226840
rect 358722 226788 358728 226840
rect 358780 226828 358786 226840
rect 444374 226828 444380 226840
rect 358780 226800 444380 226828
rect 358780 226788 358786 226800
rect 444374 226788 444380 226800
rect 444432 226788 444438 226840
rect 173802 226720 173808 226772
rect 173860 226760 173866 226772
rect 244274 226760 244280 226772
rect 173860 226732 244280 226760
rect 173860 226720 173866 226732
rect 244274 226720 244280 226732
rect 244332 226720 244338 226772
rect 357342 226720 357348 226772
rect 357400 226760 357406 226772
rect 440602 226760 440608 226772
rect 357400 226732 440608 226760
rect 357400 226720 357406 226732
rect 440602 226720 440608 226732
rect 440660 226720 440666 226772
rect 42150 226652 42156 226704
rect 42208 226692 42214 226704
rect 44358 226692 44364 226704
rect 42208 226664 44364 226692
rect 42208 226652 42214 226664
rect 44358 226652 44364 226664
rect 44416 226652 44422 226704
rect 174630 226652 174636 226704
rect 174688 226692 174694 226704
rect 243630 226692 243636 226704
rect 174688 226664 243636 226692
rect 174688 226652 174694 226664
rect 243630 226652 243636 226664
rect 243688 226652 243694 226704
rect 355870 226652 355876 226704
rect 355928 226692 355934 226704
rect 437474 226692 437480 226704
rect 355928 226664 437480 226692
rect 355928 226652 355934 226664
rect 437474 226652 437480 226664
rect 437532 226652 437538 226704
rect 177206 226584 177212 226636
rect 177264 226624 177270 226636
rect 245746 226624 245752 226636
rect 177264 226596 245752 226624
rect 177264 226584 177270 226596
rect 245746 226584 245752 226596
rect 245804 226584 245810 226636
rect 354490 226584 354496 226636
rect 354548 226624 354554 226636
rect 433794 226624 433800 226636
rect 354548 226596 433800 226624
rect 354548 226584 354554 226596
rect 433794 226584 433800 226596
rect 433852 226584 433858 226636
rect 190270 226516 190276 226568
rect 190328 226556 190334 226568
rect 251450 226556 251456 226568
rect 190328 226528 251456 226556
rect 190328 226516 190334 226528
rect 251450 226516 251456 226528
rect 251508 226516 251514 226568
rect 351638 226516 351644 226568
rect 351696 226556 351702 226568
rect 427078 226556 427084 226568
rect 351696 226528 427084 226556
rect 351696 226516 351702 226528
rect 427078 226516 427084 226528
rect 427136 226516 427142 226568
rect 57606 226312 57612 226364
rect 57664 226352 57670 226364
rect 62114 226352 62120 226364
rect 57664 226324 62120 226352
rect 57664 226312 57670 226324
rect 62114 226312 62120 226324
rect 62172 226312 62178 226364
rect 116578 226244 116584 226296
rect 116636 226284 116642 226296
rect 220078 226284 220084 226296
rect 116636 226256 220084 226284
rect 116636 226244 116642 226256
rect 220078 226244 220084 226256
rect 220136 226244 220142 226296
rect 364242 226244 364248 226296
rect 364300 226284 364306 226296
rect 455690 226284 455696 226296
rect 364300 226256 455696 226284
rect 364300 226244 364306 226256
rect 455690 226244 455696 226256
rect 455748 226244 455754 226296
rect 456150 226244 456156 226296
rect 456208 226284 456214 226296
rect 548150 226284 548156 226296
rect 456208 226256 548156 226284
rect 456208 226244 456214 226256
rect 548150 226244 548156 226256
rect 548208 226244 548214 226296
rect 112990 226176 112996 226228
rect 113048 226216 113054 226228
rect 218606 226216 218612 226228
rect 113048 226188 218612 226216
rect 113048 226176 113054 226188
rect 218606 226176 218612 226188
rect 218664 226176 218670 226228
rect 223114 226176 223120 226228
rect 223172 226216 223178 226228
rect 233234 226216 233240 226228
rect 223172 226188 233240 226216
rect 223172 226176 223178 226188
rect 233234 226176 233240 226188
rect 233292 226176 233298 226228
rect 365530 226176 365536 226228
rect 365588 226216 365594 226228
rect 459554 226216 459560 226228
rect 365588 226188 459560 226216
rect 365588 226176 365594 226188
rect 459554 226176 459560 226188
rect 459612 226176 459618 226228
rect 109862 226108 109868 226160
rect 109920 226148 109926 226160
rect 217226 226148 217232 226160
rect 109920 226120 217232 226148
rect 109920 226108 109926 226120
rect 217226 226108 217232 226120
rect 217284 226108 217290 226160
rect 218054 226108 218060 226160
rect 218112 226148 218118 226160
rect 227254 226148 227260 226160
rect 218112 226120 227260 226148
rect 218112 226108 218118 226120
rect 227254 226108 227260 226120
rect 227312 226108 227318 226160
rect 227346 226108 227352 226160
rect 227404 226148 227410 226160
rect 237558 226148 237564 226160
rect 227404 226120 237564 226148
rect 227404 226108 227410 226120
rect 237558 226108 237564 226120
rect 237616 226108 237622 226160
rect 366910 226108 366916 226160
rect 366968 226148 366974 226160
rect 462406 226148 462412 226160
rect 366968 226120 462412 226148
rect 366968 226108 366974 226120
rect 462406 226108 462412 226120
rect 462464 226108 462470 226160
rect 106550 226040 106556 226092
rect 106608 226080 106614 226092
rect 215754 226080 215760 226092
rect 106608 226052 215760 226080
rect 106608 226040 106614 226052
rect 215754 226040 215760 226052
rect 215812 226040 215818 226092
rect 224954 226040 224960 226092
rect 225012 226080 225018 226092
rect 251818 226080 251824 226092
rect 225012 226052 251824 226080
rect 225012 226040 225018 226052
rect 251818 226040 251824 226052
rect 251876 226040 251882 226092
rect 253842 226040 253848 226092
rect 253900 226080 253906 226092
rect 276474 226080 276480 226092
rect 253900 226052 276480 226080
rect 253900 226040 253906 226052
rect 276474 226040 276480 226052
rect 276532 226040 276538 226092
rect 335906 226040 335912 226092
rect 335964 226080 335970 226092
rect 367738 226080 367744 226092
rect 335964 226052 367744 226080
rect 335964 226040 335970 226052
rect 367738 226040 367744 226052
rect 367796 226040 367802 226092
rect 368382 226040 368388 226092
rect 368440 226080 368446 226092
rect 465074 226080 465080 226092
rect 368440 226052 465080 226080
rect 368440 226040 368446 226052
rect 465074 226040 465080 226052
rect 465132 226040 465138 226092
rect 103238 225972 103244 226024
rect 103296 226012 103302 226024
rect 214374 226012 214380 226024
rect 103296 225984 214380 226012
rect 103296 225972 103302 225984
rect 214374 225972 214380 225984
rect 214432 225972 214438 226024
rect 220630 225972 220636 226024
rect 220688 226012 220694 226024
rect 264238 226012 264244 226024
rect 220688 225984 264244 226012
rect 220688 225972 220694 225984
rect 264238 225972 264244 225984
rect 264296 225972 264302 226024
rect 358354 225972 358360 226024
rect 358412 226012 358418 226024
rect 441614 226012 441620 226024
rect 358412 225984 441620 226012
rect 358412 225972 358418 225984
rect 441614 225972 441620 225984
rect 441672 225972 441678 226024
rect 441706 225972 441712 226024
rect 441764 226012 441770 226024
rect 540422 226012 540428 226024
rect 441764 225984 540428 226012
rect 441764 225972 441770 225984
rect 540422 225972 540428 225984
rect 540480 225972 540486 226024
rect 99834 225904 99840 225956
rect 99892 225944 99898 225956
rect 212902 225944 212908 225956
rect 99892 225916 212908 225944
rect 99892 225904 99898 225916
rect 212902 225904 212908 225916
rect 212960 225904 212966 225956
rect 215294 225904 215300 225956
rect 215352 225944 215358 225956
rect 261386 225944 261392 225956
rect 215352 225916 261392 225944
rect 215352 225904 215358 225916
rect 261386 225904 261392 225916
rect 261444 225904 261450 225956
rect 322750 225904 322756 225956
rect 322808 225944 322814 225956
rect 358170 225944 358176 225956
rect 322808 225916 358176 225944
rect 322808 225904 322814 225916
rect 358170 225904 358176 225916
rect 358228 225904 358234 225956
rect 369762 225904 369768 225956
rect 369820 225944 369826 225956
rect 469214 225944 469220 225956
rect 369820 225916 469220 225944
rect 369820 225904 369826 225916
rect 469214 225904 469220 225916
rect 469272 225904 469278 225956
rect 96522 225836 96528 225888
rect 96580 225876 96586 225888
rect 211522 225876 211528 225888
rect 96580 225848 211528 225876
rect 96580 225836 96586 225848
rect 211522 225836 211528 225848
rect 211580 225836 211586 225888
rect 211706 225836 211712 225888
rect 211764 225876 211770 225888
rect 258994 225876 259000 225888
rect 211764 225848 259000 225876
rect 211764 225836 211770 225848
rect 258994 225836 259000 225848
rect 259052 225836 259058 225888
rect 326982 225836 326988 225888
rect 327040 225876 327046 225888
rect 362954 225876 362960 225888
rect 327040 225848 362960 225876
rect 327040 225836 327046 225848
rect 362954 225836 362960 225848
rect 363012 225836 363018 225888
rect 371234 225836 371240 225888
rect 371292 225876 371298 225888
rect 471974 225876 471980 225888
rect 371292 225848 471980 225876
rect 371292 225836 371298 225848
rect 471974 225836 471980 225848
rect 472032 225836 472038 225888
rect 86310 225768 86316 225820
rect 86368 225808 86374 225820
rect 207198 225808 207204 225820
rect 86368 225780 207204 225808
rect 86368 225768 86374 225780
rect 207198 225768 207204 225780
rect 207256 225768 207262 225820
rect 208302 225768 208308 225820
rect 208360 225808 208366 225820
rect 257890 225808 257896 225820
rect 208360 225780 257896 225808
rect 208360 225768 208366 225780
rect 257890 225768 257896 225780
rect 257948 225768 257954 225820
rect 324130 225768 324136 225820
rect 324188 225808 324194 225820
rect 361574 225808 361580 225820
rect 324188 225780 361580 225808
rect 324188 225768 324194 225780
rect 361574 225768 361580 225780
rect 361632 225768 361638 225820
rect 372614 225768 372620 225820
rect 372672 225808 372678 225820
rect 476206 225808 476212 225820
rect 372672 225780 476212 225808
rect 372672 225768 372678 225780
rect 476206 225768 476212 225780
rect 476264 225768 476270 225820
rect 76282 225700 76288 225752
rect 76340 225740 76346 225752
rect 202966 225740 202972 225752
rect 76340 225712 202972 225740
rect 76340 225700 76346 225712
rect 202966 225700 202972 225712
rect 203024 225700 203030 225752
rect 206830 225700 206836 225752
rect 206888 225740 206894 225752
rect 256786 225740 256792 225752
rect 206888 225712 256792 225740
rect 206888 225700 206894 225712
rect 256786 225700 256792 225712
rect 256844 225700 256850 225752
rect 303798 225700 303804 225752
rect 303856 225740 303862 225752
rect 317414 225740 317420 225752
rect 303856 225712 317420 225740
rect 303856 225700 303862 225712
rect 317414 225700 317420 225712
rect 317472 225700 317478 225752
rect 343082 225700 343088 225752
rect 343140 225740 343146 225752
rect 407114 225740 407120 225752
rect 343140 225712 407120 225740
rect 343140 225700 343146 225712
rect 407114 225700 407120 225712
rect 407172 225700 407178 225752
rect 408402 225700 408408 225752
rect 408460 225740 408466 225752
rect 531406 225740 531412 225752
rect 408460 225712 531412 225740
rect 408460 225700 408466 225712
rect 531406 225700 531412 225712
rect 531464 225700 531470 225752
rect 539594 225700 539600 225752
rect 539652 225740 539658 225752
rect 560294 225740 560300 225752
rect 539652 225712 560300 225740
rect 539652 225700 539658 225712
rect 560294 225700 560300 225712
rect 560352 225700 560358 225752
rect 56042 225632 56048 225684
rect 56100 225672 56106 225684
rect 194410 225672 194416 225684
rect 56100 225644 194416 225672
rect 56100 225632 56106 225644
rect 194410 225632 194416 225644
rect 194468 225632 194474 225684
rect 199010 225632 199016 225684
rect 199068 225672 199074 225684
rect 200666 225672 200672 225684
rect 199068 225644 200672 225672
rect 199068 225632 199074 225644
rect 200666 225632 200672 225644
rect 200724 225632 200730 225684
rect 203242 225632 203248 225684
rect 203300 225672 203306 225684
rect 255314 225672 255320 225684
rect 203300 225644 255320 225672
rect 203300 225632 203306 225644
rect 255314 225632 255320 225644
rect 255372 225632 255378 225684
rect 263410 225632 263416 225684
rect 263468 225672 263474 225684
rect 280982 225672 280988 225684
rect 263468 225644 280988 225672
rect 263468 225632 263474 225644
rect 280982 225632 280988 225644
rect 281040 225632 281046 225684
rect 302694 225632 302700 225684
rect 302752 225672 302758 225684
rect 313550 225672 313556 225684
rect 302752 225644 313556 225672
rect 302752 225632 302758 225644
rect 313550 225632 313556 225644
rect 313608 225632 313614 225684
rect 314470 225632 314476 225684
rect 314528 225672 314534 225684
rect 331214 225672 331220 225684
rect 314528 225644 331220 225672
rect 314528 225632 314534 225644
rect 331214 225632 331220 225644
rect 331272 225632 331278 225684
rect 341610 225632 341616 225684
rect 341668 225672 341674 225684
rect 403526 225672 403532 225684
rect 341668 225644 403532 225672
rect 341668 225632 341674 225644
rect 403526 225632 403532 225644
rect 403584 225632 403590 225684
rect 403618 225632 403624 225684
rect 403676 225672 403682 225684
rect 552014 225672 552020 225684
rect 403676 225644 552020 225672
rect 403676 225632 403682 225644
rect 552014 225632 552020 225644
rect 552072 225632 552078 225684
rect 52730 225564 52736 225616
rect 52788 225604 52794 225616
rect 192662 225604 192668 225616
rect 52788 225576 192668 225604
rect 52788 225564 52794 225576
rect 192662 225564 192668 225576
rect 192720 225564 192726 225616
rect 201402 225564 201408 225616
rect 201460 225604 201466 225616
rect 255038 225604 255044 225616
rect 201460 225576 255044 225604
rect 201460 225564 201466 225576
rect 255038 225564 255044 225576
rect 255096 225564 255102 225616
rect 257062 225564 257068 225616
rect 257120 225604 257126 225616
rect 278130 225604 278136 225616
rect 257120 225576 278136 225604
rect 257120 225564 257126 225576
rect 278130 225564 278136 225576
rect 278188 225564 278194 225616
rect 310974 225564 310980 225616
rect 311032 225604 311038 225616
rect 334066 225604 334072 225616
rect 311032 225576 334072 225604
rect 311032 225564 311038 225576
rect 334066 225564 334072 225576
rect 334124 225564 334130 225616
rect 344462 225564 344468 225616
rect 344520 225604 344526 225616
rect 410242 225604 410248 225616
rect 344520 225576 410248 225604
rect 344520 225564 344526 225576
rect 410242 225564 410248 225576
rect 410300 225564 410306 225616
rect 411070 225564 411076 225616
rect 411128 225604 411134 225616
rect 559190 225604 559196 225616
rect 411128 225576 559196 225604
rect 411128 225564 411134 225576
rect 559190 225564 559196 225576
rect 559248 225564 559254 225616
rect 119890 225496 119896 225548
rect 119948 225536 119954 225548
rect 221182 225536 221188 225548
rect 119948 225508 221188 225536
rect 119948 225496 119954 225508
rect 221182 225496 221188 225508
rect 221240 225496 221246 225548
rect 362862 225496 362868 225548
rect 362920 225536 362926 225548
rect 452654 225536 452660 225548
rect 362920 225508 452660 225536
rect 362920 225496 362926 225508
rect 452654 225496 452660 225508
rect 452712 225496 452718 225548
rect 123386 225428 123392 225480
rect 123444 225468 123450 225480
rect 222930 225468 222936 225480
rect 123444 225440 222936 225468
rect 123444 225428 123450 225440
rect 222930 225428 222936 225440
rect 222988 225428 222994 225480
rect 359826 225428 359832 225480
rect 359884 225468 359890 225480
rect 445754 225468 445760 225480
rect 359884 225440 445760 225468
rect 359884 225428 359890 225440
rect 445754 225428 445760 225440
rect 445812 225428 445818 225480
rect 126790 225360 126796 225412
rect 126848 225400 126854 225412
rect 224310 225400 224316 225412
rect 126848 225372 224316 225400
rect 126848 225360 126854 225372
rect 224310 225360 224316 225372
rect 224368 225360 224374 225412
rect 356974 225360 356980 225412
rect 357032 225400 357038 225412
rect 438854 225400 438860 225412
rect 357032 225372 438860 225400
rect 357032 225360 357038 225372
rect 438854 225360 438860 225372
rect 438912 225360 438918 225412
rect 130102 225292 130108 225344
rect 130160 225332 130166 225344
rect 225782 225332 225788 225344
rect 130160 225304 225788 225332
rect 130160 225292 130166 225304
rect 225782 225292 225788 225304
rect 225840 225292 225846 225344
rect 348786 225292 348792 225344
rect 348844 225332 348850 225344
rect 420362 225332 420368 225344
rect 348844 225304 420368 225332
rect 348844 225292 348850 225304
rect 420362 225292 420368 225304
rect 420420 225292 420426 225344
rect 133506 225224 133512 225276
rect 133564 225264 133570 225276
rect 227162 225264 227168 225276
rect 133564 225236 227168 225264
rect 133564 225224 133570 225236
rect 227162 225224 227168 225236
rect 227220 225224 227226 225276
rect 345934 225224 345940 225276
rect 345992 225264 345998 225276
rect 414014 225264 414020 225276
rect 345992 225236 414020 225264
rect 345992 225224 345998 225236
rect 414014 225224 414020 225236
rect 414072 225224 414078 225276
rect 170490 225156 170496 225208
rect 170548 225196 170554 225208
rect 242894 225196 242900 225208
rect 170548 225168 242900 225196
rect 170548 225156 170554 225168
rect 242894 225156 242900 225168
rect 242952 225156 242958 225208
rect 339034 225156 339040 225208
rect 339092 225196 339098 225208
rect 382274 225196 382280 225208
rect 339092 225168 382280 225196
rect 339092 225156 339098 225168
rect 382274 225156 382280 225168
rect 382332 225156 382338 225208
rect 383102 225156 383108 225208
rect 383160 225196 383166 225208
rect 448974 225196 448980 225208
rect 383160 225168 448980 225196
rect 383160 225156 383166 225168
rect 448974 225156 448980 225168
rect 449032 225156 449038 225208
rect 180610 225088 180616 225140
rect 180668 225128 180674 225140
rect 247126 225128 247132 225140
rect 180668 225100 247132 225128
rect 180668 225088 180674 225100
rect 247126 225088 247132 225100
rect 247184 225088 247190 225140
rect 340230 225088 340236 225140
rect 340288 225128 340294 225140
rect 385678 225128 385684 225140
rect 340288 225100 385684 225128
rect 340288 225088 340294 225100
rect 385678 225088 385684 225100
rect 385736 225088 385742 225140
rect 386966 225088 386972 225140
rect 387024 225128 387030 225140
rect 434714 225128 434720 225140
rect 387024 225100 434720 225128
rect 387024 225088 387030 225100
rect 434714 225088 434720 225100
rect 434772 225088 434778 225140
rect 192846 224952 192852 225004
rect 192904 224992 192910 225004
rect 197630 224992 197636 225004
rect 192904 224964 197636 224992
rect 192904 224952 192910 224964
rect 197630 224952 197636 224964
rect 197688 224952 197694 225004
rect 162762 224884 162768 224936
rect 162820 224924 162826 224936
rect 238202 224924 238208 224936
rect 162820 224896 238208 224924
rect 162820 224884 162826 224896
rect 238202 224884 238208 224896
rect 238260 224884 238266 224936
rect 374086 224884 374092 224936
rect 374144 224924 374150 224936
rect 479242 224924 479248 224936
rect 374144 224896 479248 224924
rect 374144 224884 374150 224896
rect 479242 224884 479248 224896
rect 479300 224884 479306 224936
rect 159542 224816 159548 224868
rect 159600 224856 159606 224868
rect 236822 224856 236828 224868
rect 159600 224828 236828 224856
rect 159600 224816 159606 224828
rect 236822 224816 236828 224828
rect 236880 224816 236886 224868
rect 370866 224816 370872 224868
rect 370924 224856 370930 224868
rect 475010 224856 475016 224868
rect 370924 224828 475016 224856
rect 370924 224816 370930 224828
rect 475010 224816 475016 224828
rect 475068 224816 475074 224868
rect 155770 224748 155776 224800
rect 155828 224788 155834 224800
rect 235350 224788 235356 224800
rect 155828 224760 235356 224788
rect 155828 224748 155834 224760
rect 235350 224748 235356 224760
rect 235408 224748 235414 224800
rect 372246 224748 372252 224800
rect 372304 224788 372310 224800
rect 478966 224788 478972 224800
rect 372304 224760 478972 224788
rect 372304 224748 372310 224760
rect 478966 224748 478972 224760
rect 479024 224748 479030 224800
rect 114922 224680 114928 224732
rect 114980 224720 114986 224732
rect 151814 224720 151820 224732
rect 114980 224692 151820 224720
rect 114980 224680 114986 224692
rect 151814 224680 151820 224692
rect 151872 224680 151878 224732
rect 152918 224680 152924 224732
rect 152976 224720 152982 224732
rect 233970 224720 233976 224732
rect 152976 224692 233976 224720
rect 152976 224680 152982 224692
rect 233970 224680 233976 224692
rect 234028 224680 234034 224732
rect 332318 224680 332324 224732
rect 332376 224720 332382 224732
rect 372614 224720 372620 224732
rect 332376 224692 372620 224720
rect 332376 224680 332382 224692
rect 372614 224680 372620 224692
rect 372672 224680 372678 224732
rect 373718 224680 373724 224732
rect 373776 224720 373782 224732
rect 481818 224720 481824 224732
rect 373776 224692 481824 224720
rect 373776 224680 373782 224692
rect 481818 224680 481824 224692
rect 481876 224680 481882 224732
rect 149422 224612 149428 224664
rect 149480 224652 149486 224664
rect 232314 224652 232320 224664
rect 149480 224624 232320 224652
rect 149480 224612 149486 224624
rect 232314 224612 232320 224624
rect 232372 224612 232378 224664
rect 338390 224612 338396 224664
rect 338448 224652 338454 224664
rect 380158 224652 380164 224664
rect 338448 224624 380164 224652
rect 338448 224612 338454 224624
rect 380158 224612 380164 224624
rect 380216 224612 380222 224664
rect 388714 224612 388720 224664
rect 388772 224652 388778 224664
rect 516226 224652 516232 224664
rect 388772 224624 516232 224652
rect 388772 224612 388778 224624
rect 516226 224612 516232 224624
rect 516284 224612 516290 224664
rect 146110 224544 146116 224596
rect 146168 224584 146174 224596
rect 231118 224584 231124 224596
rect 146168 224556 231124 224584
rect 146168 224544 146174 224556
rect 231118 224544 231124 224556
rect 231176 224544 231182 224596
rect 337010 224544 337016 224596
rect 337068 224584 337074 224596
rect 378686 224584 378692 224596
rect 337068 224556 378692 224584
rect 337068 224544 337074 224556
rect 378686 224544 378692 224556
rect 378744 224544 378750 224596
rect 389726 224544 389732 224596
rect 389784 224584 389790 224596
rect 518894 224584 518900 224596
rect 389784 224556 518900 224584
rect 389784 224544 389790 224556
rect 518894 224544 518900 224556
rect 518952 224544 518958 224596
rect 142706 224476 142712 224528
rect 142764 224516 142770 224528
rect 229646 224516 229652 224528
rect 142764 224488 229652 224516
rect 142764 224476 142770 224488
rect 229646 224476 229652 224488
rect 229704 224476 229710 224528
rect 342714 224476 342720 224528
rect 342772 224516 342778 224528
rect 405918 224516 405924 224528
rect 342772 224488 405924 224516
rect 342772 224476 342778 224488
rect 405918 224476 405924 224488
rect 405976 224476 405982 224528
rect 406746 224476 406752 224528
rect 406804 224516 406810 224528
rect 545758 224516 545764 224528
rect 406804 224488 545764 224516
rect 406804 224476 406810 224488
rect 545758 224476 545764 224488
rect 545816 224476 545822 224528
rect 139210 224408 139216 224460
rect 139268 224448 139274 224460
rect 228266 224448 228272 224460
rect 139268 224420 228272 224448
rect 139268 224408 139274 224420
rect 228266 224408 228272 224420
rect 228324 224408 228330 224460
rect 234614 224408 234620 224460
rect 234672 224448 234678 224460
rect 250346 224448 250352 224460
rect 234672 224420 250352 224448
rect 234672 224408 234678 224420
rect 250346 224408 250352 224420
rect 250404 224408 250410 224460
rect 268930 224408 268936 224460
rect 268988 224448 268994 224460
rect 283558 224448 283564 224460
rect 268988 224420 283564 224448
rect 268988 224408 268994 224420
rect 283558 224408 283564 224420
rect 283616 224408 283622 224460
rect 333698 224408 333704 224460
rect 333756 224448 333762 224460
rect 378042 224448 378048 224460
rect 333756 224420 378048 224448
rect 333756 224408 333762 224420
rect 378042 224408 378048 224420
rect 378100 224408 378106 224460
rect 400030 224408 400036 224460
rect 400088 224448 400094 224460
rect 543182 224448 543188 224460
rect 400088 224420 543188 224448
rect 400088 224408 400094 224420
rect 543182 224408 543188 224420
rect 543240 224408 543246 224460
rect 135990 224340 135996 224392
rect 136048 224380 136054 224392
rect 226794 224380 226800 224392
rect 136048 224352 226800 224380
rect 136048 224340 136054 224352
rect 226794 224340 226800 224352
rect 226852 224340 226858 224392
rect 246850 224340 246856 224392
rect 246908 224380 246914 224392
rect 273622 224380 273628 224392
rect 246908 224352 273628 224380
rect 246908 224340 246914 224352
rect 273622 224340 273628 224352
rect 273680 224340 273686 224392
rect 307754 224340 307760 224392
rect 307812 224380 307818 224392
rect 325694 224380 325700 224392
rect 307812 224352 325700 224380
rect 307812 224340 307818 224352
rect 325694 224340 325700 224352
rect 325752 224340 325758 224392
rect 339862 224340 339868 224392
rect 339920 224380 339926 224392
rect 386966 224380 386972 224392
rect 339920 224352 386972 224380
rect 339920 224340 339926 224352
rect 386966 224340 386972 224352
rect 387024 224340 387030 224392
rect 402238 224340 402244 224392
rect 402296 224380 402302 224392
rect 548242 224380 548248 224392
rect 402296 224352 548248 224380
rect 402296 224340 402302 224352
rect 548242 224340 548248 224352
rect 548300 224340 548306 224392
rect 101490 224272 101496 224324
rect 101548 224312 101554 224324
rect 136358 224312 136364 224324
rect 101548 224284 136364 224312
rect 101548 224272 101554 224284
rect 136358 224272 136364 224284
rect 136416 224272 136422 224324
rect 136450 224272 136456 224324
rect 136508 224312 136514 224324
rect 228634 224312 228640 224324
rect 136508 224284 228640 224312
rect 136508 224272 136514 224284
rect 228634 224272 228640 224284
rect 228692 224272 228698 224324
rect 232406 224272 232412 224324
rect 232464 224312 232470 224324
rect 243262 224312 243268 224324
rect 232464 224284 243268 224312
rect 232464 224272 232470 224284
rect 243262 224272 243268 224284
rect 243320 224272 243326 224324
rect 243630 224272 243636 224324
rect 243688 224312 243694 224324
rect 272242 224312 272248 224324
rect 243688 224284 272248 224312
rect 243688 224272 243694 224284
rect 272242 224272 272248 224284
rect 272300 224272 272306 224324
rect 309226 224272 309232 224324
rect 309284 224312 309290 224324
rect 328730 224312 328736 224324
rect 309284 224284 328736 224312
rect 309284 224272 309290 224284
rect 328730 224272 328736 224284
rect 328788 224272 328794 224324
rect 341426 224272 341432 224324
rect 341484 224312 341490 224324
rect 401870 224312 401876 224324
rect 341484 224284 401876 224312
rect 341484 224272 341490 224284
rect 401870 224272 401876 224284
rect 401928 224272 401934 224324
rect 408678 224272 408684 224324
rect 408736 224312 408742 224324
rect 408736 224284 412220 224312
rect 408736 224272 408742 224284
rect 88150 224204 88156 224256
rect 88208 224244 88214 224256
rect 207566 224244 207572 224256
rect 88208 224216 207572 224244
rect 88208 224204 88214 224216
rect 207566 224204 207572 224216
rect 207624 224204 207630 224256
rect 239950 224204 239956 224256
rect 240008 224244 240014 224256
rect 271046 224244 271052 224256
rect 240008 224216 271052 224244
rect 240008 224204 240014 224216
rect 271046 224204 271052 224216
rect 271104 224204 271110 224256
rect 292574 224204 292580 224256
rect 292632 224244 292638 224256
rect 293494 224244 293500 224256
rect 292632 224216 293500 224244
rect 292632 224204 292638 224216
rect 293494 224204 293500 224216
rect 293552 224204 293558 224256
rect 311342 224204 311348 224256
rect 311400 224244 311406 224256
rect 331306 224244 331312 224256
rect 311400 224216 331312 224244
rect 311400 224204 311406 224216
rect 331306 224204 331312 224216
rect 331364 224204 331370 224256
rect 344094 224204 344100 224256
rect 344152 224244 344158 224256
rect 408586 224244 408592 224256
rect 344152 224216 408592 224244
rect 344152 224204 344158 224216
rect 408586 224204 408592 224216
rect 408644 224204 408650 224256
rect 411346 224204 411352 224256
rect 411404 224244 411410 224256
rect 412192 224244 412220 224284
rect 412266 224272 412272 224324
rect 412324 224312 412330 224324
rect 556154 224312 556160 224324
rect 412324 224284 556160 224312
rect 412324 224272 412330 224284
rect 556154 224272 556160 224284
rect 556212 224272 556218 224324
rect 563606 224244 563612 224256
rect 411404 224216 412128 224244
rect 412192 224216 563612 224244
rect 411404 224204 411410 224216
rect 166258 224136 166264 224188
rect 166316 224176 166322 224188
rect 239674 224176 239680 224188
rect 166316 224148 239680 224176
rect 166316 224136 166322 224148
rect 239674 224136 239680 224148
rect 239732 224136 239738 224188
rect 345566 224136 345572 224188
rect 345624 224176 345630 224188
rect 411990 224176 411996 224188
rect 345624 224148 411996 224176
rect 345624 224136 345630 224148
rect 411990 224136 411996 224148
rect 412048 224136 412054 224188
rect 412100 224176 412128 224216
rect 563606 224204 563612 224216
rect 563664 224204 563670 224256
rect 506474 224176 506480 224188
rect 412100 224148 506480 224176
rect 506474 224136 506480 224148
rect 506532 224136 506538 224188
rect 169570 224068 169576 224120
rect 169628 224108 169634 224120
rect 241054 224108 241060 224120
rect 169628 224080 241060 224108
rect 169628 224068 169634 224080
rect 241054 224068 241060 224080
rect 241112 224068 241118 224120
rect 335538 224068 335544 224120
rect 335596 224108 335602 224120
rect 377306 224108 377312 224120
rect 335596 224080 377312 224108
rect 335596 224068 335602 224080
rect 377306 224068 377312 224080
rect 377364 224068 377370 224120
rect 378594 224068 378600 224120
rect 378652 224108 378658 224120
rect 472066 224108 472072 224120
rect 378652 224080 472072 224108
rect 378652 224068 378658 224080
rect 472066 224068 472072 224080
rect 472124 224068 472130 224120
rect 172974 224000 172980 224052
rect 173032 224040 173038 224052
rect 242526 224040 242532 224052
rect 173032 224012 242532 224040
rect 173032 224000 173038 224012
rect 242526 224000 242532 224012
rect 242584 224000 242590 224052
rect 387518 224000 387524 224052
rect 387576 224040 387582 224052
rect 468294 224040 468300 224052
rect 387576 224012 468300 224040
rect 387576 224000 387582 224012
rect 468294 224000 468300 224012
rect 468352 224000 468358 224052
rect 176470 223932 176476 223984
rect 176528 223972 176534 223984
rect 243906 223972 243912 223984
rect 176528 223944 243912 223972
rect 176528 223932 176534 223944
rect 243906 223932 243912 223944
rect 243964 223932 243970 223984
rect 349798 223932 349804 223984
rect 349856 223972 349862 223984
rect 422386 223972 422392 223984
rect 349856 223944 422392 223972
rect 349856 223932 349862 223944
rect 422386 223932 422392 223944
rect 422444 223932 422450 223984
rect 179690 223864 179696 223916
rect 179748 223904 179754 223916
rect 245378 223904 245384 223916
rect 179748 223876 245384 223904
rect 179748 223864 179754 223876
rect 245378 223864 245384 223876
rect 245436 223864 245442 223916
rect 347314 223864 347320 223916
rect 347372 223904 347378 223916
rect 417050 223904 417056 223916
rect 347372 223876 417056 223904
rect 347372 223864 347378 223876
rect 417050 223864 417056 223876
rect 417108 223864 417114 223916
rect 183186 223796 183192 223848
rect 183244 223836 183250 223848
rect 246758 223836 246764 223848
rect 183244 223808 246764 223836
rect 183244 223796 183250 223808
rect 246758 223796 246764 223808
rect 246816 223796 246822 223848
rect 348418 223796 348424 223848
rect 348476 223836 348482 223848
rect 418706 223836 418712 223848
rect 348476 223808 418712 223836
rect 348476 223796 348482 223808
rect 418706 223796 418712 223808
rect 418764 223796 418770 223848
rect 186222 223728 186228 223780
rect 186280 223768 186286 223780
rect 248230 223768 248236 223780
rect 186280 223740 248236 223768
rect 186280 223728 186286 223740
rect 248230 223728 248236 223740
rect 248288 223728 248294 223780
rect 346946 223728 346952 223780
rect 347004 223768 347010 223780
rect 415486 223768 415492 223780
rect 347004 223740 415492 223768
rect 347004 223728 347010 223740
rect 415486 223728 415492 223740
rect 415544 223728 415550 223780
rect 416682 223728 416688 223780
rect 416740 223768 416746 223780
rect 465166 223768 465172 223780
rect 416740 223740 465172 223768
rect 416740 223728 416746 223740
rect 465166 223728 465172 223740
rect 465224 223728 465230 223780
rect 405458 223660 405464 223712
rect 405516 223700 405522 223712
rect 412266 223700 412272 223712
rect 405516 223672 412272 223700
rect 405516 223660 405522 223672
rect 412266 223660 412272 223672
rect 412324 223660 412330 223712
rect 125870 223524 125876 223576
rect 125928 223564 125934 223576
rect 222562 223564 222568 223576
rect 125928 223536 222568 223564
rect 125928 223524 125934 223536
rect 222562 223524 222568 223536
rect 222620 223524 222626 223576
rect 357986 223524 357992 223576
rect 358044 223564 358050 223576
rect 444742 223564 444748 223576
rect 358044 223536 444748 223564
rect 358044 223524 358050 223536
rect 444742 223524 444748 223536
rect 444800 223524 444806 223576
rect 115750 223456 115756 223508
rect 115808 223496 115814 223508
rect 210418 223496 210424 223508
rect 115808 223468 210424 223496
rect 115808 223456 115814 223468
rect 210418 223456 210424 223468
rect 210476 223456 210482 223508
rect 213914 223456 213920 223508
rect 213972 223496 213978 223508
rect 221826 223496 221832 223508
rect 213972 223468 221832 223496
rect 213972 223456 213978 223468
rect 221826 223456 221832 223468
rect 221884 223456 221890 223508
rect 359458 223456 359464 223508
rect 359516 223496 359522 223508
rect 448606 223496 448612 223508
rect 359516 223468 448612 223496
rect 359516 223456 359522 223468
rect 448606 223456 448612 223468
rect 448664 223456 448670 223508
rect 108850 223388 108856 223440
rect 108908 223428 108914 223440
rect 215386 223428 215392 223440
rect 108908 223400 215392 223428
rect 108908 223388 108914 223400
rect 215386 223388 215392 223400
rect 215444 223388 215450 223440
rect 361114 223388 361120 223440
rect 361172 223428 361178 223440
rect 451458 223428 451464 223440
rect 361172 223400 451464 223428
rect 361172 223388 361178 223400
rect 451458 223388 451464 223400
rect 451516 223388 451522 223440
rect 105722 223320 105728 223372
rect 105780 223360 105786 223372
rect 214006 223360 214012 223372
rect 105780 223332 214012 223360
rect 105780 223320 105786 223332
rect 214006 223320 214012 223332
rect 214064 223320 214070 223372
rect 352282 223320 352288 223372
rect 352340 223360 352346 223372
rect 431310 223360 431316 223372
rect 352340 223332 431316 223360
rect 352340 223320 352346 223332
rect 431310 223320 431316 223332
rect 431368 223320 431374 223372
rect 431402 223320 431408 223372
rect 431460 223360 431466 223372
rect 525058 223360 525064 223372
rect 431460 223332 525064 223360
rect 431460 223320 431466 223332
rect 525058 223320 525064 223332
rect 525116 223320 525122 223372
rect 101950 223252 101956 223304
rect 102008 223292 102014 223304
rect 102008 223264 209820 223292
rect 102008 223252 102014 223264
rect 95602 223184 95608 223236
rect 95660 223224 95666 223236
rect 209792 223224 209820 223264
rect 210418 223252 210424 223304
rect 210476 223292 210482 223304
rect 218238 223292 218244 223304
rect 210476 223264 218244 223292
rect 210476 223252 210482 223264
rect 218238 223252 218244 223264
rect 218296 223252 218302 223304
rect 390094 223252 390100 223304
rect 390152 223292 390158 223304
rect 395706 223292 395712 223304
rect 390152 223264 395712 223292
rect 390152 223252 390158 223264
rect 395706 223252 395712 223264
rect 395764 223252 395770 223304
rect 396350 223252 396356 223304
rect 396408 223292 396414 223304
rect 523126 223292 523132 223304
rect 396408 223264 523132 223292
rect 396408 223252 396414 223264
rect 523126 223252 523132 223264
rect 523184 223252 523190 223304
rect 212534 223224 212540 223236
rect 95660 223196 205634 223224
rect 209792 223196 212540 223224
rect 95660 223184 95666 223196
rect 82170 223116 82176 223168
rect 82228 223156 82234 223168
rect 203978 223156 203984 223168
rect 82228 223128 203984 223156
rect 82228 223116 82234 223128
rect 203978 223116 203984 223128
rect 204036 223116 204042 223168
rect 205606 223156 205634 223196
rect 212534 223184 212540 223196
rect 212592 223184 212598 223236
rect 314194 223184 314200 223236
rect 314252 223224 314258 223236
rect 338114 223224 338120 223236
rect 314252 223196 338120 223224
rect 314252 223184 314258 223196
rect 338114 223184 338120 223196
rect 338172 223184 338178 223236
rect 353754 223184 353760 223236
rect 353812 223224 353818 223236
rect 434806 223224 434812 223236
rect 353812 223196 434812 223224
rect 353812 223184 353818 223196
rect 434806 223184 434812 223196
rect 434864 223184 434870 223236
rect 435542 223184 435548 223236
rect 435600 223224 435606 223236
rect 567194 223224 567200 223236
rect 435600 223196 567200 223224
rect 435600 223184 435606 223196
rect 567194 223184 567200 223196
rect 567252 223184 567258 223236
rect 209682 223156 209688 223168
rect 205606 223128 209688 223156
rect 209682 223116 209688 223128
rect 209740 223116 209746 223168
rect 250346 223116 250352 223168
rect 250404 223156 250410 223168
rect 275094 223156 275100 223168
rect 250404 223128 275100 223156
rect 250404 223116 250410 223128
rect 275094 223116 275100 223128
rect 275152 223116 275158 223168
rect 317046 223116 317052 223168
rect 317104 223156 317110 223168
rect 345014 223156 345020 223168
rect 317104 223128 345020 223156
rect 317104 223116 317110 223128
rect 345014 223116 345020 223128
rect 345072 223116 345078 223168
rect 395798 223116 395804 223168
rect 395856 223156 395862 223168
rect 395856 223128 396488 223156
rect 395856 223116 395862 223128
rect 75362 223048 75368 223100
rect 75420 223088 75426 223100
rect 201126 223088 201132 223100
rect 75420 223060 201132 223088
rect 75420 223048 75426 223060
rect 201126 223048 201132 223060
rect 201184 223048 201190 223100
rect 204898 223048 204904 223100
rect 204956 223088 204962 223100
rect 256418 223088 256424 223100
rect 204956 223060 256424 223088
rect 204956 223048 204962 223060
rect 256418 223048 256424 223060
rect 256476 223048 256482 223100
rect 319254 223048 319260 223100
rect 319312 223088 319318 223100
rect 350626 223088 350632 223100
rect 319312 223060 350632 223088
rect 319312 223048 319318 223060
rect 350626 223048 350632 223060
rect 350684 223048 350690 223100
rect 391566 223048 391572 223100
rect 391624 223088 391630 223100
rect 396350 223088 396356 223100
rect 391624 223060 396356 223088
rect 391624 223048 391630 223060
rect 396350 223048 396356 223060
rect 396408 223048 396414 223100
rect 396460 223088 396488 223128
rect 398834 223116 398840 223168
rect 398892 223156 398898 223168
rect 530578 223156 530584 223168
rect 398892 223128 530584 223156
rect 398892 223116 398898 223128
rect 530578 223116 530584 223128
rect 530636 223116 530642 223168
rect 671430 223116 671436 223168
rect 671488 223156 671494 223168
rect 675938 223156 675944 223168
rect 671488 223128 675944 223156
rect 671488 223116 671494 223128
rect 675938 223116 675944 223128
rect 675996 223116 676002 223168
rect 533062 223088 533068 223100
rect 396460 223060 533068 223088
rect 533062 223048 533068 223060
rect 533120 223048 533126 223100
rect 68738 222980 68744 223032
rect 68796 223020 68802 223032
rect 68796 222992 197032 223020
rect 68796 222980 68802 222992
rect 65334 222912 65340 222964
rect 65392 222952 65398 222964
rect 196894 222952 196900 222964
rect 65392 222924 196900 222952
rect 65392 222912 65398 222924
rect 196894 222912 196900 222924
rect 196952 222912 196958 222964
rect 197004 222952 197032 222992
rect 198182 222980 198188 223032
rect 198240 223020 198246 223032
rect 253566 223020 253572 223032
rect 198240 222992 253572 223020
rect 198240 222980 198246 222992
rect 253566 222980 253572 222992
rect 253624 222980 253630 223032
rect 311434 222980 311440 223032
rect 311492 223020 311498 223032
rect 318886 223020 318892 223032
rect 311492 222992 318892 223020
rect 311492 222980 311498 222992
rect 318886 222980 318892 222992
rect 318944 222980 318950 223032
rect 330938 222980 330944 223032
rect 330996 223020 331002 223032
rect 365990 223020 365996 223032
rect 330996 222992 365996 223020
rect 330996 222980 331002 222992
rect 365990 222980 365996 222992
rect 366048 222980 366054 223032
rect 397914 222980 397920 223032
rect 397972 223020 397978 223032
rect 538306 223020 538312 223032
rect 397972 222992 538312 223020
rect 397972 222980 397978 222992
rect 538306 222980 538312 222992
rect 538364 222980 538370 223032
rect 198274 222952 198280 222964
rect 197004 222924 198280 222952
rect 198274 222912 198280 222924
rect 198332 222912 198338 222964
rect 199930 222912 199936 222964
rect 199988 222952 199994 222964
rect 253934 222952 253940 222964
rect 199988 222924 253940 222952
rect 199988 222912 199994 222924
rect 253934 222912 253940 222924
rect 253992 222912 253998 222964
rect 265526 222912 265532 222964
rect 265584 222952 265590 222964
rect 282086 222952 282092 222964
rect 265584 222924 282092 222952
rect 265584 222912 265590 222924
rect 282086 222912 282092 222924
rect 282144 222912 282150 222964
rect 306374 222912 306380 222964
rect 306432 222952 306438 222964
rect 321922 222952 321928 222964
rect 306432 222924 321928 222952
rect 306432 222912 306438 222924
rect 321922 222912 321928 222924
rect 321980 222912 321986 222964
rect 326614 222912 326620 222964
rect 326672 222952 326678 222964
rect 371234 222952 371240 222964
rect 326672 222924 371240 222952
rect 326672 222912 326678 222924
rect 371234 222912 371240 222924
rect 371292 222912 371298 222964
rect 379790 222912 379796 222964
rect 379848 222952 379854 222964
rect 389174 222952 389180 222964
rect 379848 222924 389180 222952
rect 379848 222912 379854 222924
rect 389174 222912 389180 222924
rect 389232 222912 389238 222964
rect 394786 222912 394792 222964
rect 394844 222952 394850 222964
rect 398834 222952 398840 222964
rect 394844 222924 398840 222952
rect 394844 222912 394850 222924
rect 398834 222912 398840 222924
rect 398892 222912 398898 222964
rect 404630 222912 404636 222964
rect 404688 222952 404694 222964
rect 553670 222952 553676 222964
rect 404688 222924 553676 222952
rect 404688 222912 404694 222924
rect 553670 222912 553676 222924
rect 553728 222912 553734 222964
rect 66070 222844 66076 222896
rect 66128 222884 66134 222896
rect 198366 222884 198372 222896
rect 66128 222856 198372 222884
rect 66128 222844 66134 222856
rect 198366 222844 198372 222856
rect 198424 222844 198430 222896
rect 200758 222844 200764 222896
rect 200816 222884 200822 222896
rect 255682 222884 255688 222896
rect 200816 222856 255688 222884
rect 200816 222844 200822 222856
rect 255682 222844 255688 222856
rect 255740 222844 255746 222896
rect 262122 222844 262128 222896
rect 262180 222884 262186 222896
rect 280706 222884 280712 222896
rect 262180 222856 280712 222884
rect 262180 222844 262186 222856
rect 280706 222844 280712 222856
rect 280764 222844 280770 222896
rect 308490 222844 308496 222896
rect 308548 222884 308554 222896
rect 324498 222884 324504 222896
rect 308548 222856 324504 222884
rect 308548 222844 308554 222856
rect 324498 222844 324504 222856
rect 324556 222844 324562 222896
rect 337654 222844 337660 222896
rect 337712 222884 337718 222896
rect 390646 222884 390652 222896
rect 337712 222856 390652 222884
rect 337712 222844 337718 222856
rect 390646 222844 390652 222856
rect 390704 222844 390710 222896
rect 407574 222844 407580 222896
rect 407632 222884 407638 222896
rect 560938 222884 560944 222896
rect 407632 222856 560944 222884
rect 407632 222844 407638 222856
rect 560938 222844 560944 222856
rect 560996 222844 561002 222896
rect 132310 222776 132316 222828
rect 132368 222816 132374 222828
rect 225414 222816 225420 222828
rect 132368 222788 225420 222816
rect 132368 222776 132374 222788
rect 225414 222776 225420 222788
rect 225472 222776 225478 222828
rect 356606 222776 356612 222828
rect 356664 222816 356670 222828
rect 441706 222816 441712 222828
rect 356664 222788 441712 222816
rect 356664 222776 356670 222788
rect 441706 222776 441712 222788
rect 441764 222776 441770 222828
rect 177850 222708 177856 222760
rect 177908 222748 177914 222760
rect 245010 222748 245016 222760
rect 177908 222720 245016 222748
rect 177908 222708 177914 222720
rect 245010 222708 245016 222720
rect 245068 222708 245074 222760
rect 355134 222708 355140 222760
rect 355192 222748 355198 222760
rect 438026 222748 438032 222760
rect 355192 222720 438032 222748
rect 355192 222708 355198 222720
rect 438026 222708 438032 222720
rect 438084 222708 438090 222760
rect 674374 222708 674380 222760
rect 674432 222748 674438 222760
rect 675938 222748 675944 222760
rect 674432 222720 675944 222748
rect 674432 222708 674438 222720
rect 675938 222708 675944 222720
rect 675996 222708 676002 222760
rect 162026 222640 162032 222692
rect 162084 222680 162090 222692
rect 180794 222680 180800 222692
rect 162084 222652 180800 222680
rect 162084 222640 162090 222652
rect 180794 222640 180800 222652
rect 180852 222640 180858 222692
rect 181346 222640 181352 222692
rect 181404 222680 181410 222692
rect 246482 222680 246488 222692
rect 181404 222652 246488 222680
rect 181404 222640 181410 222652
rect 246482 222640 246488 222652
rect 246540 222640 246546 222692
rect 352650 222640 352656 222692
rect 352708 222680 352714 222692
rect 429286 222680 429292 222692
rect 352708 222652 429292 222680
rect 352708 222640 352714 222652
rect 429286 222640 429292 222652
rect 429344 222640 429350 222692
rect 187326 222572 187332 222624
rect 187384 222612 187390 222624
rect 249978 222612 249984 222624
rect 187384 222584 249984 222612
rect 187384 222572 187390 222584
rect 249978 222572 249984 222584
rect 250036 222572 250042 222624
rect 351178 222572 351184 222624
rect 351236 222612 351242 222624
rect 427906 222612 427912 222624
rect 351236 222584 427912 222612
rect 351236 222572 351242 222584
rect 427906 222572 427912 222584
rect 427964 222572 427970 222624
rect 428642 222572 428648 222624
rect 428700 222612 428706 222624
rect 488534 222612 488540 222624
rect 428700 222584 488540 222612
rect 428700 222572 428706 222584
rect 488534 222572 488540 222584
rect 488592 222572 488598 222624
rect 184750 222504 184756 222556
rect 184808 222544 184814 222556
rect 247862 222544 247868 222556
rect 184808 222516 247868 222544
rect 184808 222504 184814 222516
rect 247862 222504 247868 222516
rect 247920 222504 247926 222556
rect 349430 222504 349436 222556
rect 349488 222544 349494 222556
rect 425054 222544 425060 222556
rect 349488 222516 425060 222544
rect 349488 222504 349494 222516
rect 425054 222504 425060 222516
rect 425112 222504 425118 222556
rect 188154 222436 188160 222488
rect 188212 222476 188218 222488
rect 249334 222476 249340 222488
rect 188212 222448 249340 222476
rect 188212 222436 188218 222448
rect 249334 222436 249340 222448
rect 249392 222436 249398 222488
rect 348142 222436 348148 222488
rect 348200 222476 348206 222488
rect 421190 222476 421196 222488
rect 348200 222448 421196 222476
rect 348200 222436 348206 222448
rect 421190 222436 421196 222448
rect 421248 222436 421254 222488
rect 191558 222368 191564 222420
rect 191616 222408 191622 222420
rect 250714 222408 250720 222420
rect 191616 222380 250720 222408
rect 191616 222368 191622 222380
rect 250714 222368 250720 222380
rect 250772 222368 250778 222420
rect 346670 222368 346676 222420
rect 346728 222408 346734 222420
rect 415302 222408 415308 222420
rect 346728 222380 415308 222408
rect 346728 222368 346734 222380
rect 415302 222368 415308 222380
rect 415360 222368 415366 222420
rect 196526 222300 196532 222352
rect 196584 222340 196590 222352
rect 252278 222340 252284 222352
rect 196584 222312 252284 222340
rect 196584 222300 196590 222312
rect 252278 222300 252284 222312
rect 252336 222300 252342 222352
rect 664530 222164 664536 222216
rect 664588 222204 664594 222216
rect 676030 222204 676036 222216
rect 664588 222176 676036 222204
rect 664588 222164 664594 222176
rect 676030 222164 676036 222176
rect 676088 222164 676094 222216
rect 122466 222096 122472 222148
rect 122524 222136 122530 222148
rect 220998 222136 221004 222148
rect 122524 222108 221004 222136
rect 122524 222096 122530 222108
rect 220998 222096 221004 222108
rect 221056 222096 221062 222148
rect 228450 222096 228456 222148
rect 228508 222136 228514 222148
rect 266446 222136 266452 222148
rect 228508 222108 266452 222136
rect 228508 222096 228514 222108
rect 266446 222096 266452 222108
rect 266504 222096 266510 222148
rect 311158 222096 311164 222148
rect 311216 222136 311222 222148
rect 311986 222136 311992 222148
rect 311216 222108 311992 222136
rect 311216 222096 311222 222108
rect 311986 222096 311992 222108
rect 312044 222096 312050 222148
rect 312538 222096 312544 222148
rect 312596 222136 312602 222148
rect 315298 222136 315304 222148
rect 312596 222108 315304 222136
rect 312596 222096 312602 222108
rect 315298 222096 315304 222108
rect 315356 222096 315362 222148
rect 318702 222096 318708 222148
rect 318760 222136 318766 222148
rect 349154 222136 349160 222148
rect 318760 222108 349160 222136
rect 318760 222096 318766 222108
rect 349154 222096 349160 222108
rect 349212 222096 349218 222148
rect 362678 222096 362684 222148
rect 362736 222136 362742 222148
rect 453206 222136 453212 222148
rect 362736 222108 453212 222136
rect 362736 222096 362742 222108
rect 453206 222096 453212 222108
rect 453264 222096 453270 222148
rect 453298 222096 453304 222148
rect 453356 222136 453362 222148
rect 545206 222136 545212 222148
rect 453356 222108 545212 222136
rect 453356 222096 453362 222108
rect 545206 222096 545212 222108
rect 545264 222096 545270 222148
rect 119154 222028 119160 222080
rect 119212 222068 119218 222080
rect 219526 222068 219532 222080
rect 119212 222040 219532 222068
rect 119212 222028 119218 222040
rect 219526 222028 219532 222040
rect 219584 222028 219590 222080
rect 226794 222028 226800 222080
rect 226852 222068 226858 222080
rect 265158 222068 265164 222080
rect 226852 222040 265164 222068
rect 226852 222028 226858 222040
rect 265158 222028 265164 222040
rect 265216 222028 265222 222080
rect 320818 222028 320824 222080
rect 320876 222068 320882 222080
rect 356054 222068 356060 222080
rect 320876 222040 356060 222068
rect 320876 222028 320882 222040
rect 356054 222028 356060 222040
rect 356112 222028 356118 222080
rect 363598 222028 363604 222080
rect 363656 222068 363662 222080
rect 456794 222068 456800 222080
rect 363656 222040 456800 222068
rect 363656 222028 363662 222040
rect 456794 222028 456800 222040
rect 456852 222028 456858 222080
rect 100754 221960 100760 222012
rect 100812 222000 100818 222012
rect 204438 222000 204444 222012
rect 100812 221972 204444 222000
rect 100812 221960 100818 221972
rect 204438 221960 204444 221972
rect 204496 221960 204502 222012
rect 224862 221960 224868 222012
rect 224920 222000 224926 222012
rect 265066 222000 265072 222012
rect 224920 221972 265072 222000
rect 224920 221960 224926 221972
rect 265066 221960 265072 221972
rect 265124 221960 265130 222012
rect 322290 221960 322296 222012
rect 322348 222000 322354 222012
rect 359090 222000 359096 222012
rect 322348 221972 359096 222000
rect 322348 221960 322354 221972
rect 359090 221960 359096 221972
rect 359148 221960 359154 222012
rect 365070 221960 365076 222012
rect 365128 222000 365134 222012
rect 460014 222000 460020 222012
rect 365128 221972 460020 222000
rect 365128 221960 365134 221972
rect 460014 221960 460020 221972
rect 460072 221960 460078 222012
rect 112438 221892 112444 221944
rect 112496 221932 112502 221944
rect 216766 221932 216772 221944
rect 112496 221904 216772 221932
rect 112496 221892 112502 221904
rect 216766 221892 216772 221904
rect 216824 221892 216830 221944
rect 223482 221892 223488 221944
rect 223540 221932 223546 221944
rect 263778 221932 263784 221944
rect 223540 221904 263784 221932
rect 223540 221892 223546 221904
rect 263778 221892 263784 221904
rect 263836 221892 263842 221944
rect 321186 221892 321192 221944
rect 321244 221932 321250 221944
rect 357526 221932 357532 221944
rect 321244 221904 357532 221932
rect 321244 221892 321250 221904
rect 357526 221892 357532 221904
rect 357584 221892 357590 221944
rect 363966 221892 363972 221944
rect 364024 221932 364030 221944
rect 458358 221932 458364 221944
rect 364024 221904 458364 221932
rect 364024 221892 364030 221904
rect 458358 221892 458364 221904
rect 458416 221892 458422 221944
rect 88886 221824 88892 221876
rect 88944 221864 88950 221876
rect 88944 221836 205312 221864
rect 88944 221824 88950 221836
rect 85482 221756 85488 221808
rect 85540 221796 85546 221808
rect 205174 221796 205180 221808
rect 85540 221768 205180 221796
rect 85540 221756 85546 221768
rect 205174 221756 205180 221768
rect 205232 221756 205238 221808
rect 205284 221796 205312 221836
rect 205542 221824 205548 221876
rect 205600 221864 205606 221876
rect 206738 221864 206744 221876
rect 205600 221836 206744 221864
rect 205600 221824 205606 221836
rect 206738 221824 206744 221836
rect 206796 221824 206802 221876
rect 220078 221824 220084 221876
rect 220136 221864 220142 221876
rect 262306 221864 262312 221876
rect 220136 221836 262312 221864
rect 220136 221824 220142 221836
rect 262306 221824 262312 221836
rect 262364 221824 262370 221876
rect 322658 221824 322664 221876
rect 322716 221864 322722 221876
rect 360746 221864 360752 221876
rect 322716 221836 360752 221864
rect 322716 221824 322722 221836
rect 360746 221824 360752 221836
rect 360804 221824 360810 221876
rect 366450 221824 366456 221876
rect 366508 221864 366514 221876
rect 463694 221864 463700 221876
rect 366508 221836 463700 221864
rect 366508 221824 366514 221836
rect 463694 221824 463700 221836
rect 463752 221824 463758 221876
rect 672626 221824 672632 221876
rect 672684 221864 672690 221876
rect 676030 221864 676036 221876
rect 672684 221836 676036 221864
rect 672684 221824 672690 221836
rect 676030 221824 676036 221836
rect 676088 221824 676094 221876
rect 206646 221796 206652 221808
rect 205284 221768 206652 221796
rect 206646 221756 206652 221768
rect 206704 221756 206710 221808
rect 208210 221756 208216 221808
rect 208268 221796 208274 221808
rect 220170 221796 220176 221808
rect 208268 221768 220176 221796
rect 208268 221756 208274 221768
rect 220170 221756 220176 221768
rect 220228 221756 220234 221808
rect 221734 221756 221740 221808
rect 221792 221796 221798 221808
rect 263686 221796 263692 221808
rect 221792 221768 263692 221796
rect 221792 221756 221798 221768
rect 263686 221756 263692 221768
rect 263744 221756 263750 221808
rect 324222 221756 324228 221808
rect 324280 221796 324286 221808
rect 362402 221796 362408 221808
rect 324280 221768 362408 221796
rect 324280 221756 324286 221768
rect 362402 221756 362408 221768
rect 362460 221756 362466 221808
rect 367922 221756 367928 221808
rect 367980 221796 367986 221808
rect 466730 221796 466736 221808
rect 367980 221768 466736 221796
rect 367980 221756 367986 221768
rect 466730 221756 466736 221768
rect 466788 221756 466794 221808
rect 467098 221756 467104 221808
rect 467156 221796 467162 221808
rect 557810 221796 557816 221808
rect 467156 221768 557816 221796
rect 467156 221756 467162 221768
rect 557810 221756 557816 221768
rect 557868 221756 557874 221808
rect 83826 221688 83832 221740
rect 83884 221728 83890 221740
rect 204806 221728 204812 221740
rect 83884 221700 204812 221728
rect 83884 221688 83890 221700
rect 204806 221688 204812 221700
rect 204864 221688 204870 221740
rect 206922 221688 206928 221740
rect 206980 221728 206986 221740
rect 217318 221728 217324 221740
rect 206980 221700 217324 221728
rect 206980 221688 206986 221700
rect 217318 221688 217324 221700
rect 217376 221688 217382 221740
rect 218422 221688 218428 221740
rect 218480 221728 218486 221740
rect 261846 221728 261852 221740
rect 218480 221700 261852 221728
rect 218480 221688 218486 221700
rect 261846 221688 261852 221700
rect 261904 221688 261910 221740
rect 325142 221688 325148 221740
rect 325200 221728 325206 221740
rect 365806 221728 365812 221740
rect 325200 221700 365812 221728
rect 325200 221688 325206 221700
rect 365806 221688 365812 221700
rect 365864 221688 365870 221740
rect 369302 221688 369308 221740
rect 369360 221728 369366 221740
rect 470134 221728 470140 221740
rect 369360 221700 470140 221728
rect 369360 221688 369366 221700
rect 470134 221688 470140 221700
rect 470192 221688 470198 221740
rect 80422 221620 80428 221672
rect 80480 221660 80486 221672
rect 203426 221660 203432 221672
rect 80480 221632 203432 221660
rect 80480 221620 80486 221632
rect 203426 221620 203432 221632
rect 203484 221620 203490 221672
rect 203702 221620 203708 221672
rect 203760 221660 203766 221672
rect 214466 221660 214472 221672
rect 203760 221632 214472 221660
rect 203760 221620 203766 221632
rect 214466 221620 214472 221632
rect 214524 221620 214530 221672
rect 216582 221620 216588 221672
rect 216640 221660 216646 221672
rect 261018 221660 261024 221672
rect 216640 221632 261024 221660
rect 216640 221620 216646 221632
rect 261018 221620 261024 221632
rect 261076 221620 261082 221672
rect 326522 221620 326528 221672
rect 326580 221660 326586 221672
rect 369118 221660 369124 221672
rect 326580 221632 369124 221660
rect 326580 221620 326586 221632
rect 369118 221620 369124 221632
rect 369176 221620 369182 221672
rect 370774 221620 370780 221672
rect 370832 221660 370838 221672
rect 473538 221660 473544 221672
rect 370832 221632 473544 221660
rect 370832 221620 370838 221632
rect 473538 221620 473544 221632
rect 473596 221620 473602 221672
rect 551278 221620 551284 221672
rect 551336 221660 551342 221672
rect 565446 221660 565452 221672
rect 551336 221632 565452 221660
rect 551336 221620 551342 221632
rect 565446 221620 565452 221632
rect 565504 221620 565510 221672
rect 77018 221552 77024 221604
rect 77076 221592 77082 221604
rect 201954 221592 201960 221604
rect 77076 221564 201960 221592
rect 77076 221552 77082 221564
rect 201954 221552 201960 221564
rect 202012 221552 202018 221604
rect 202414 221552 202420 221604
rect 202472 221592 202478 221604
rect 210142 221592 210148 221604
rect 202472 221564 210148 221592
rect 202472 221552 202478 221564
rect 210142 221552 210148 221564
rect 210200 221552 210206 221604
rect 213362 221552 213368 221604
rect 213420 221592 213426 221604
rect 259638 221592 259644 221604
rect 213420 221564 259644 221592
rect 213420 221552 213426 221564
rect 259638 221552 259644 221564
rect 259696 221552 259702 221604
rect 325510 221552 325516 221604
rect 325568 221592 325574 221604
rect 367462 221592 367468 221604
rect 325568 221564 367468 221592
rect 325568 221552 325574 221564
rect 367462 221552 367468 221564
rect 367520 221552 367526 221604
rect 400122 221552 400128 221604
rect 400180 221592 400186 221604
rect 541434 221592 541440 221604
rect 400180 221564 541440 221592
rect 400180 221552 400186 221564
rect 541434 221552 541440 221564
rect 541492 221552 541498 221604
rect 547138 221552 547144 221604
rect 547196 221592 547202 221604
rect 561766 221592 561772 221604
rect 547196 221564 561772 221592
rect 547196 221552 547202 221564
rect 561766 221552 561772 221564
rect 561824 221552 561830 221604
rect 63402 221484 63408 221536
rect 63460 221524 63466 221536
rect 196250 221524 196256 221536
rect 63460 221496 196256 221524
rect 63460 221484 63466 221496
rect 196250 221484 196256 221496
rect 196308 221484 196314 221536
rect 197262 221484 197268 221536
rect 197320 221524 197326 221536
rect 244918 221524 244924 221536
rect 197320 221496 244924 221524
rect 197320 221484 197326 221496
rect 244918 221484 244924 221496
rect 244976 221484 244982 221536
rect 245286 221484 245292 221536
rect 245344 221524 245350 221536
rect 273438 221524 273444 221536
rect 245344 221496 273444 221524
rect 245344 221484 245350 221496
rect 273438 221484 273444 221496
rect 273496 221484 273502 221536
rect 275554 221484 275560 221536
rect 275612 221524 275618 221536
rect 286134 221524 286140 221536
rect 275612 221496 286140 221524
rect 275612 221484 275618 221496
rect 286134 221484 286140 221496
rect 286192 221484 286198 221536
rect 319438 221484 319444 221536
rect 319496 221524 319502 221536
rect 352374 221524 352380 221536
rect 319496 221496 352380 221524
rect 319496 221484 319502 221496
rect 352374 221484 352380 221496
rect 352432 221484 352438 221536
rect 352558 221484 352564 221536
rect 352616 221524 352622 221536
rect 397730 221524 397736 221536
rect 352616 221496 397736 221524
rect 352616 221484 352622 221496
rect 397730 221484 397736 221496
rect 397788 221484 397794 221536
rect 404170 221484 404176 221536
rect 404228 221524 404234 221536
rect 551278 221524 551284 221536
rect 404228 221496 551284 221524
rect 404228 221484 404234 221496
rect 551278 221484 551284 221496
rect 551336 221484 551342 221536
rect 674650 221484 674656 221536
rect 674708 221524 674714 221536
rect 676030 221524 676036 221536
rect 674708 221496 676036 221524
rect 674708 221484 674714 221496
rect 676030 221484 676036 221496
rect 676088 221484 676094 221536
rect 60274 221416 60280 221468
rect 60332 221456 60338 221468
rect 194870 221456 194876 221468
rect 60332 221428 194876 221456
rect 60332 221416 60338 221428
rect 194870 221416 194876 221428
rect 194928 221416 194934 221468
rect 209682 221416 209688 221468
rect 209740 221456 209746 221468
rect 258258 221456 258264 221468
rect 209740 221428 258264 221456
rect 209740 221416 209746 221428
rect 258258 221416 258264 221428
rect 258316 221416 258322 221468
rect 272242 221416 272248 221468
rect 272300 221456 272306 221468
rect 284662 221456 284668 221468
rect 272300 221428 284668 221456
rect 272300 221416 272306 221428
rect 284662 221416 284668 221428
rect 284720 221416 284726 221468
rect 301222 221416 301228 221468
rect 301280 221456 301286 221468
rect 310514 221456 310520 221468
rect 301280 221428 310520 221456
rect 301280 221416 301286 221428
rect 310514 221416 310520 221428
rect 310572 221416 310578 221468
rect 319806 221416 319812 221468
rect 319864 221456 319870 221468
rect 354030 221456 354036 221468
rect 319864 221428 354036 221456
rect 319864 221416 319870 221428
rect 354030 221416 354036 221428
rect 354088 221416 354094 221468
rect 401134 221456 401140 221468
rect 354646 221428 401140 221456
rect 129274 221348 129280 221400
rect 129332 221388 129338 221400
rect 223758 221388 223764 221400
rect 129332 221360 223764 221388
rect 129332 221348 129338 221360
rect 223758 221348 223764 221360
rect 223816 221348 223822 221400
rect 231670 221348 231676 221400
rect 231728 221388 231734 221400
rect 267826 221388 267832 221400
rect 231728 221360 267832 221388
rect 231728 221348 231734 221360
rect 267826 221348 267832 221360
rect 267884 221348 267890 221400
rect 317322 221348 317328 221400
rect 317380 221388 317386 221400
rect 345566 221388 345572 221400
rect 317380 221360 345572 221388
rect 317380 221348 317386 221360
rect 345566 221348 345572 221360
rect 345624 221348 345630 221400
rect 151078 221280 151084 221332
rect 151136 221320 151142 221332
rect 233418 221320 233424 221332
rect 151136 221292 233424 221320
rect 151136 221280 151142 221292
rect 233418 221280 233424 221292
rect 233476 221280 233482 221332
rect 235258 221280 235264 221332
rect 235316 221320 235322 221332
rect 269206 221320 269212 221332
rect 235316 221292 269212 221320
rect 235316 221280 235322 221292
rect 269206 221280 269212 221292
rect 269264 221280 269270 221332
rect 315942 221280 315948 221332
rect 316000 221320 316006 221332
rect 342254 221320 342260 221332
rect 316000 221292 342260 221320
rect 316000 221280 316006 221292
rect 342254 221280 342260 221292
rect 342312 221280 342318 221332
rect 353938 221280 353944 221332
rect 353996 221320 354002 221332
rect 354646 221320 354674 221428
rect 401134 221416 401140 221428
rect 401192 221416 401198 221468
rect 406286 221416 406292 221468
rect 406344 221456 406350 221468
rect 558454 221456 558460 221468
rect 406344 221428 558460 221456
rect 406344 221416 406350 221428
rect 558454 221416 558460 221428
rect 558512 221416 558518 221468
rect 565078 221416 565084 221468
rect 565136 221456 565142 221468
rect 573542 221456 573548 221468
rect 565136 221428 573548 221456
rect 565136 221416 565142 221428
rect 573542 221416 573548 221428
rect 573600 221416 573606 221468
rect 361298 221348 361304 221400
rect 361356 221388 361362 221400
rect 449894 221388 449900 221400
rect 361356 221360 449900 221388
rect 361356 221348 361362 221360
rect 449894 221348 449900 221360
rect 449952 221348 449958 221400
rect 353996 221292 354674 221320
rect 353996 221280 354002 221292
rect 360102 221280 360108 221332
rect 360160 221320 360166 221332
rect 446582 221320 446588 221332
rect 360160 221292 446588 221320
rect 360160 221280 360166 221292
rect 446582 221280 446588 221292
rect 446640 221280 446646 221332
rect 157794 221212 157800 221264
rect 157852 221252 157858 221264
rect 236178 221252 236184 221264
rect 157852 221224 236184 221252
rect 157852 221212 157858 221224
rect 236178 221212 236184 221224
rect 236236 221212 236242 221264
rect 238570 221212 238576 221264
rect 238628 221252 238634 221264
rect 270678 221252 270684 221264
rect 238628 221224 270684 221252
rect 238628 221212 238634 221224
rect 270678 221212 270684 221224
rect 270736 221212 270742 221264
rect 314562 221212 314568 221264
rect 314620 221252 314626 221264
rect 338850 221252 338856 221264
rect 314620 221224 338856 221252
rect 314620 221212 314626 221224
rect 338850 221212 338856 221224
rect 338908 221212 338914 221264
rect 357066 221212 357072 221264
rect 357124 221252 357130 221264
rect 439774 221252 439780 221264
rect 357124 221224 439780 221252
rect 357124 221212 357130 221224
rect 439774 221212 439780 221224
rect 439832 221212 439838 221264
rect 443638 221212 443644 221264
rect 443696 221252 443702 221264
rect 491386 221252 491392 221264
rect 443696 221224 491392 221252
rect 443696 221212 443702 221224
rect 491386 221212 491392 221224
rect 491444 221212 491450 221264
rect 167914 221144 167920 221196
rect 167972 221184 167978 221196
rect 240502 221184 240508 221196
rect 167972 221156 240508 221184
rect 167972 221144 167978 221156
rect 240502 221144 240508 221156
rect 240560 221144 240566 221196
rect 241974 221144 241980 221196
rect 242032 221184 242038 221196
rect 271966 221184 271972 221196
rect 242032 221156 271972 221184
rect 242032 221144 242038 221156
rect 271966 221144 271972 221156
rect 272024 221144 272030 221196
rect 313182 221144 313188 221196
rect 313240 221184 313246 221196
rect 335538 221184 335544 221196
rect 313240 221156 335544 221184
rect 313240 221144 313246 221156
rect 335538 221144 335544 221156
rect 335596 221144 335602 221196
rect 351546 221144 351552 221196
rect 351604 221184 351610 221196
rect 425514 221184 425520 221196
rect 351604 221156 425520 221184
rect 351604 221144 351610 221156
rect 425514 221144 425520 221156
rect 425572 221144 425578 221196
rect 183922 221076 183928 221128
rect 183980 221116 183986 221128
rect 248506 221116 248512 221128
rect 183980 221088 248512 221116
rect 183980 221076 183986 221088
rect 248506 221076 248512 221088
rect 248564 221076 248570 221128
rect 248690 221076 248696 221128
rect 248748 221116 248754 221128
rect 274818 221116 274824 221128
rect 248748 221088 274824 221116
rect 248748 221076 248754 221088
rect 274818 221076 274824 221088
rect 274876 221076 274882 221128
rect 376110 221076 376116 221128
rect 376168 221116 376174 221128
rect 443178 221116 443184 221128
rect 376168 221088 443184 221116
rect 376168 221076 376174 221088
rect 443178 221076 443184 221088
rect 443236 221076 443242 221128
rect 189810 221008 189816 221060
rect 189868 221048 189874 221060
rect 249426 221048 249432 221060
rect 189868 221020 249432 221048
rect 189868 221008 189874 221020
rect 249426 221008 249432 221020
rect 249484 221008 249490 221060
rect 343266 221008 343272 221060
rect 343324 221048 343330 221060
rect 407850 221048 407856 221060
rect 343324 221020 407856 221048
rect 343324 221008 343330 221020
rect 407850 221008 407856 221020
rect 407908 221008 407914 221060
rect 436462 221048 436468 221060
rect 412606 221020 436468 221048
rect 192938 220940 192944 220992
rect 192996 220980 193002 220992
rect 250806 220980 250812 220992
rect 192996 220952 250812 220980
rect 192996 220940 193002 220952
rect 250806 220940 250812 220952
rect 250864 220940 250870 220992
rect 385770 220940 385776 220992
rect 385828 220980 385834 220992
rect 411254 220980 411260 220992
rect 385828 220952 411260 220980
rect 385828 220940 385834 220952
rect 411254 220940 411260 220952
rect 411312 220940 411318 220992
rect 195146 220872 195152 220924
rect 195204 220912 195210 220924
rect 211614 220912 211620 220924
rect 195204 220884 211620 220912
rect 195204 220872 195210 220884
rect 211614 220872 211620 220884
rect 211672 220872 211678 220924
rect 380250 220872 380256 220924
rect 380308 220912 380314 220924
rect 404446 220912 404452 220924
rect 380308 220884 404452 220912
rect 380308 220872 380314 220884
rect 404446 220872 404452 220884
rect 404504 220872 404510 220924
rect 407666 220872 407672 220924
rect 407724 220912 407730 220924
rect 412606 220912 412634 221020
rect 436462 221008 436468 221020
rect 436520 221008 436526 221060
rect 672534 221008 672540 221060
rect 672592 221048 672598 221060
rect 676030 221048 676036 221060
rect 672592 221020 676036 221048
rect 672592 221008 672598 221020
rect 676030 221008 676036 221020
rect 676088 221008 676094 221060
rect 563606 220940 563612 220992
rect 563664 220980 563670 220992
rect 563664 220952 568068 220980
rect 563664 220940 563670 220952
rect 407724 220884 412634 220912
rect 407724 220872 407730 220884
rect 563698 220872 563704 220924
rect 563756 220912 563762 220924
rect 567930 220912 567936 220924
rect 563756 220884 567936 220912
rect 563756 220872 563762 220884
rect 567930 220872 567936 220884
rect 567988 220872 567994 220924
rect 568040 220912 568068 220952
rect 569126 220940 569132 220992
rect 569184 220980 569190 220992
rect 621198 220980 621204 220992
rect 569184 220952 621204 220980
rect 569184 220940 569190 220952
rect 621198 220940 621204 220952
rect 621256 220940 621262 220992
rect 619818 220912 619824 220924
rect 568040 220884 619824 220912
rect 619818 220872 619824 220884
rect 619876 220872 619882 220924
rect 57606 220844 57612 220856
rect 55186 220816 57612 220844
rect 52454 220736 52460 220788
rect 52512 220776 52518 220788
rect 55186 220776 55214 220816
rect 57606 220804 57612 220816
rect 57664 220804 57670 220856
rect 269592 220816 270540 220844
rect 52512 220748 55214 220776
rect 52512 220736 52518 220748
rect 71222 220736 71228 220788
rect 71280 220776 71286 220788
rect 71682 220776 71688 220788
rect 71280 220748 71688 220776
rect 71280 220736 71286 220748
rect 71682 220736 71688 220748
rect 71740 220736 71746 220788
rect 84654 220736 84660 220788
rect 84712 220776 84718 220788
rect 85390 220776 85396 220788
rect 84712 220748 85396 220776
rect 84712 220736 84718 220748
rect 85390 220736 85396 220748
rect 85448 220736 85454 220788
rect 131758 220736 131764 220788
rect 131816 220776 131822 220788
rect 132402 220776 132408 220788
rect 131816 220748 132408 220776
rect 131816 220736 131822 220748
rect 132402 220736 132408 220748
rect 132460 220736 132466 220788
rect 138474 220736 138480 220788
rect 138532 220776 138538 220788
rect 139302 220776 139308 220788
rect 138532 220748 139308 220776
rect 138532 220736 138538 220748
rect 139302 220736 139308 220748
rect 139360 220736 139366 220788
rect 141878 220736 141884 220788
rect 141936 220776 141942 220788
rect 222102 220776 222108 220788
rect 141936 220748 222108 220776
rect 141936 220736 141942 220748
rect 222102 220736 222108 220748
rect 222160 220736 222166 220788
rect 232682 220736 232688 220788
rect 232740 220776 232746 220788
rect 233142 220776 233148 220788
rect 232740 220748 233148 220776
rect 232740 220736 232746 220748
rect 233142 220736 233148 220748
rect 233200 220736 233206 220788
rect 239398 220736 239404 220788
rect 239456 220776 239462 220788
rect 240042 220776 240048 220788
rect 239456 220748 240048 220776
rect 239456 220736 239462 220748
rect 240042 220736 240048 220748
rect 240100 220736 240106 220788
rect 241146 220736 241152 220788
rect 241204 220776 241210 220788
rect 269592 220776 269620 220816
rect 241204 220748 269620 220776
rect 241204 220736 241210 220748
rect 269666 220736 269672 220788
rect 269724 220776 269730 220788
rect 270402 220776 270408 220788
rect 269724 220748 270408 220776
rect 269724 220736 269730 220748
rect 270402 220736 270408 220748
rect 270460 220736 270466 220788
rect 270512 220776 270540 220816
rect 305546 220804 305552 220856
rect 305604 220844 305610 220856
rect 308582 220844 308588 220856
rect 305604 220816 308588 220844
rect 305604 220804 305610 220816
rect 308582 220804 308588 220816
rect 308640 220804 308646 220856
rect 558454 220804 558460 220856
rect 558512 220844 558518 220856
rect 618806 220844 618812 220856
rect 558512 220816 618812 220844
rect 558512 220804 558518 220816
rect 618806 220804 618812 220816
rect 618864 220804 618870 220856
rect 271138 220776 271144 220788
rect 270512 220748 271144 220776
rect 271138 220736 271144 220748
rect 271196 220736 271202 220788
rect 273898 220736 273904 220788
rect 273956 220776 273962 220788
rect 274542 220776 274548 220788
rect 273956 220748 274548 220776
rect 273956 220736 273962 220748
rect 274542 220736 274548 220748
rect 274600 220736 274606 220788
rect 278130 220736 278136 220788
rect 278188 220776 278194 220788
rect 278682 220776 278688 220788
rect 278188 220748 278688 220776
rect 278188 220736 278194 220748
rect 278682 220736 278688 220748
rect 278740 220736 278746 220788
rect 282362 220736 282368 220788
rect 282420 220776 282426 220788
rect 282822 220776 282828 220788
rect 282420 220748 282828 220776
rect 282420 220736 282426 220748
rect 282822 220736 282828 220748
rect 282880 220736 282886 220788
rect 286502 220736 286508 220788
rect 286560 220776 286566 220788
rect 286962 220776 286968 220788
rect 286560 220748 286968 220776
rect 286560 220736 286566 220748
rect 286962 220736 286968 220748
rect 287020 220736 287026 220788
rect 287330 220736 287336 220788
rect 287388 220776 287394 220788
rect 290642 220776 290648 220788
rect 287388 220748 290648 220776
rect 287388 220736 287394 220748
rect 290642 220736 290648 220748
rect 290700 220736 290706 220788
rect 290734 220736 290740 220788
rect 290792 220776 290798 220788
rect 292206 220776 292212 220788
rect 290792 220748 292212 220776
rect 290792 220736 290798 220748
rect 292206 220736 292212 220748
rect 292264 220736 292270 220788
rect 292482 220736 292488 220788
rect 292540 220776 292546 220788
rect 293218 220776 293224 220788
rect 292540 220748 293224 220776
rect 292540 220736 292546 220748
rect 293218 220736 293224 220748
rect 293276 220736 293282 220788
rect 294966 220736 294972 220788
rect 295024 220776 295030 220788
rect 295518 220776 295524 220788
rect 295024 220748 295524 220776
rect 295024 220736 295030 220748
rect 295518 220736 295524 220748
rect 295576 220736 295582 220788
rect 298002 220736 298008 220788
rect 298060 220776 298066 220788
rect 302234 220776 302240 220788
rect 298060 220748 302240 220776
rect 298060 220736 298066 220748
rect 302234 220736 302240 220748
rect 302292 220736 302298 220788
rect 324774 220736 324780 220788
rect 324832 220776 324838 220788
rect 363230 220776 363236 220788
rect 324832 220748 363236 220776
rect 324832 220736 324838 220748
rect 363230 220736 363236 220748
rect 363288 220736 363294 220788
rect 365990 220736 365996 220788
rect 366048 220776 366054 220788
rect 380894 220776 380900 220788
rect 366048 220748 380900 220776
rect 366048 220736 366054 220748
rect 380894 220736 380900 220748
rect 380952 220736 380958 220788
rect 383378 220736 383384 220788
rect 383436 220776 383442 220788
rect 502426 220776 502432 220788
rect 383436 220748 502432 220776
rect 383436 220736 383442 220748
rect 502426 220736 502432 220748
rect 502484 220736 502490 220788
rect 505002 220736 505008 220788
rect 505060 220776 505066 220788
rect 623866 220776 623872 220788
rect 505060 220748 623872 220776
rect 505060 220736 505066 220748
rect 623866 220736 623872 220748
rect 623924 220736 623930 220788
rect 134978 220668 134984 220720
rect 135036 220708 135042 220720
rect 135036 220680 210464 220708
rect 135036 220668 135042 220680
rect 57606 220600 57612 220652
rect 57664 220640 57670 220652
rect 58618 220640 58624 220652
rect 57664 220612 58624 220640
rect 57664 220600 57670 220612
rect 58618 220600 58624 220612
rect 58676 220600 58682 220652
rect 128170 220600 128176 220652
rect 128228 220640 128234 220652
rect 210436 220640 210464 220680
rect 214190 220668 214196 220720
rect 214248 220708 214254 220720
rect 215294 220708 215300 220720
rect 214248 220680 215300 220708
rect 214248 220668 214254 220680
rect 215294 220668 215300 220680
rect 215352 220668 215358 220720
rect 237742 220668 237748 220720
rect 237800 220708 237806 220720
rect 270126 220708 270132 220720
rect 237800 220680 270132 220708
rect 237800 220668 237806 220680
rect 270126 220668 270132 220680
rect 270184 220668 270190 220720
rect 274450 220668 274456 220720
rect 274508 220708 274514 220720
rect 276750 220708 276756 220720
rect 274508 220680 276756 220708
rect 274508 220668 274514 220680
rect 276750 220668 276756 220680
rect 276808 220668 276814 220720
rect 289078 220668 289084 220720
rect 289136 220708 289142 220720
rect 291838 220708 291844 220720
rect 289136 220680 291844 220708
rect 289136 220668 289142 220680
rect 291838 220668 291844 220680
rect 291896 220668 291902 220720
rect 303062 220668 303068 220720
rect 303120 220708 303126 220720
rect 311158 220708 311164 220720
rect 303120 220680 311164 220708
rect 303120 220668 303126 220680
rect 311158 220668 311164 220680
rect 311216 220668 311222 220720
rect 326246 220668 326252 220720
rect 326304 220708 326310 220720
rect 366634 220708 366640 220720
rect 326304 220680 366640 220708
rect 326304 220668 326310 220680
rect 366634 220668 366640 220680
rect 366692 220668 366698 220720
rect 367738 220668 367744 220720
rect 367796 220708 367802 220720
rect 390554 220708 390560 220720
rect 367796 220680 390560 220708
rect 367796 220668 367802 220680
rect 390554 220668 390560 220680
rect 390612 220668 390618 220720
rect 396718 220668 396724 220720
rect 396776 220708 396782 220720
rect 517514 220708 517520 220720
rect 396776 220680 517520 220708
rect 396776 220668 396782 220680
rect 517514 220668 517520 220680
rect 517572 220668 517578 220720
rect 525058 220668 525064 220720
rect 525116 220708 525122 220720
rect 577222 220708 577228 220720
rect 525116 220680 577228 220708
rect 525116 220668 525122 220680
rect 577222 220668 577228 220680
rect 577280 220668 577286 220720
rect 673362 220668 673368 220720
rect 673420 220708 673426 220720
rect 676030 220708 676036 220720
rect 673420 220680 676036 220708
rect 673420 220668 673426 220680
rect 676030 220668 676036 220680
rect 676088 220668 676094 220720
rect 218054 220640 218060 220652
rect 128228 220612 206416 220640
rect 210436 220612 218060 220640
rect 128228 220600 128234 220612
rect 118326 220532 118332 220584
rect 118384 220572 118390 220584
rect 206388 220572 206416 220612
rect 218054 220600 218060 220612
rect 218112 220600 218118 220652
rect 235902 220600 235908 220652
rect 235960 220640 235966 220652
rect 270034 220640 270040 220652
rect 235960 220612 270040 220640
rect 235960 220600 235966 220612
rect 270034 220600 270040 220612
rect 270092 220600 270098 220652
rect 271414 220600 271420 220652
rect 271472 220640 271478 220652
rect 275370 220640 275376 220652
rect 271472 220612 275376 220640
rect 271472 220600 271478 220612
rect 275370 220600 275376 220612
rect 275428 220600 275434 220652
rect 303430 220600 303436 220652
rect 303488 220640 303494 220652
rect 312814 220640 312820 220652
rect 303488 220612 312820 220640
rect 303488 220600 303494 220612
rect 312814 220600 312820 220612
rect 312872 220600 312878 220652
rect 329558 220600 329564 220652
rect 329616 220640 329622 220652
rect 371694 220640 371700 220652
rect 329616 220612 371700 220640
rect 329616 220600 329622 220612
rect 371694 220600 371700 220612
rect 371752 220600 371758 220652
rect 371878 220600 371884 220652
rect 371936 220640 371942 220652
rect 385954 220640 385960 220652
rect 371936 220612 385960 220640
rect 371936 220600 371942 220612
rect 385954 220600 385960 220612
rect 386012 220600 386018 220652
rect 388438 220600 388444 220652
rect 388496 220640 388502 220652
rect 512822 220640 512828 220652
rect 388496 220612 512828 220640
rect 388496 220600 388502 220612
rect 512822 220600 512828 220612
rect 512880 220600 512886 220652
rect 552658 220600 552664 220652
rect 552716 220640 552722 220652
rect 632330 220640 632336 220652
rect 552716 220612 632336 220640
rect 552716 220600 552722 220612
rect 632330 220600 632336 220612
rect 632388 220600 632394 220652
rect 216674 220572 216680 220584
rect 118384 220544 206324 220572
rect 206388 220544 216680 220572
rect 118384 220532 118390 220544
rect 121270 220464 121276 220516
rect 121328 220504 121334 220516
rect 206186 220504 206192 220516
rect 121328 220476 206192 220504
rect 121328 220464 121334 220476
rect 206186 220464 206192 220476
rect 206244 220464 206250 220516
rect 206296 220504 206324 220544
rect 216674 220532 216680 220544
rect 216732 220532 216738 220584
rect 231026 220532 231032 220584
rect 231084 220572 231090 220584
rect 268286 220572 268292 220584
rect 231084 220544 268292 220572
rect 231084 220532 231090 220544
rect 268286 220532 268292 220544
rect 268344 220532 268350 220584
rect 273070 220532 273076 220584
rect 273128 220572 273134 220584
rect 276658 220572 276664 220584
rect 273128 220544 276664 220572
rect 273128 220532 273134 220544
rect 276658 220532 276664 220544
rect 276716 220532 276722 220584
rect 293218 220532 293224 220584
rect 293276 220572 293282 220584
rect 294322 220572 294328 220584
rect 293276 220544 294328 220572
rect 293276 220532 293282 220544
rect 294322 220532 294328 220544
rect 294380 220532 294386 220584
rect 299290 220532 299296 220584
rect 299348 220572 299354 220584
rect 303614 220572 303620 220584
rect 299348 220544 303620 220572
rect 299348 220532 299354 220544
rect 303614 220532 303620 220544
rect 303672 220532 303678 220584
rect 306190 220532 306196 220584
rect 306248 220572 306254 220584
rect 317874 220572 317880 220584
rect 306248 220544 317880 220572
rect 306248 220532 306254 220544
rect 317874 220532 317880 220544
rect 317932 220532 317938 220584
rect 329650 220532 329656 220584
rect 329708 220572 329714 220584
rect 373350 220572 373356 220584
rect 329708 220544 373356 220572
rect 329708 220532 329714 220544
rect 373350 220532 373356 220544
rect 373408 220532 373414 220584
rect 375282 220532 375288 220584
rect 375340 220572 375346 220584
rect 379514 220572 379520 220584
rect 375340 220544 379520 220572
rect 375340 220532 375346 220544
rect 379514 220532 379520 220544
rect 379572 220532 379578 220584
rect 379606 220532 379612 220584
rect 379664 220572 379670 220584
rect 394694 220572 394700 220584
rect 379664 220544 394700 220572
rect 379664 220532 379670 220544
rect 394694 220532 394700 220544
rect 394752 220532 394758 220584
rect 395706 220532 395712 220584
rect 395764 220572 395770 220584
rect 519998 220572 520004 220584
rect 395764 220544 520004 220572
rect 395764 220532 395770 220544
rect 519998 220532 520004 220544
rect 520056 220572 520062 220584
rect 520056 220544 572714 220572
rect 520056 220532 520062 220544
rect 208210 220504 208216 220516
rect 206296 220476 208216 220504
rect 208210 220464 208216 220476
rect 208268 220464 208274 220516
rect 224954 220504 224960 220516
rect 219406 220476 224960 220504
rect 111610 220396 111616 220448
rect 111668 220436 111674 220448
rect 206922 220436 206928 220448
rect 111668 220408 206928 220436
rect 111668 220396 111674 220408
rect 206922 220396 206928 220408
rect 206980 220396 206986 220448
rect 145190 220328 145196 220380
rect 145248 220368 145254 220380
rect 146202 220368 146208 220380
rect 145248 220340 146208 220368
rect 145248 220328 145254 220340
rect 146202 220328 146208 220340
rect 146260 220328 146266 220380
rect 155310 220328 155316 220380
rect 155368 220368 155374 220380
rect 155862 220368 155868 220380
rect 155368 220340 155868 220368
rect 155368 220328 155374 220340
rect 155862 220328 155868 220340
rect 155920 220328 155926 220380
rect 168742 220328 168748 220380
rect 168800 220368 168806 220380
rect 169662 220368 169668 220380
rect 168800 220340 169668 220368
rect 168800 220328 168806 220340
rect 169662 220328 169668 220340
rect 169720 220328 169726 220380
rect 178862 220328 178868 220380
rect 178920 220368 178926 220380
rect 179322 220368 179328 220380
rect 178920 220340 179328 220368
rect 178920 220328 178926 220340
rect 179322 220328 179328 220340
rect 179380 220328 179386 220380
rect 192294 220328 192300 220380
rect 192352 220368 192358 220380
rect 219406 220368 219434 220476
rect 224954 220464 224960 220476
rect 225012 220464 225018 220516
rect 229370 220464 229376 220516
rect 229428 220504 229434 220516
rect 262582 220504 262588 220516
rect 229428 220476 262588 220504
rect 229428 220464 229434 220476
rect 262582 220464 262588 220476
rect 262640 220464 262646 220516
rect 262950 220464 262956 220516
rect 263008 220504 263014 220516
rect 263502 220504 263508 220516
rect 263008 220476 263508 220504
rect 263008 220464 263014 220476
rect 263502 220464 263508 220476
rect 263560 220464 263566 220516
rect 304810 220464 304816 220516
rect 304868 220504 304874 220516
rect 316126 220504 316132 220516
rect 304868 220476 316132 220504
rect 304868 220464 304874 220476
rect 316126 220464 316132 220476
rect 316184 220464 316190 220516
rect 322198 220464 322204 220516
rect 322256 220504 322262 220516
rect 342990 220504 342996 220516
rect 322256 220476 342996 220504
rect 322256 220464 322262 220476
rect 342990 220464 342996 220476
rect 343048 220464 343054 220516
rect 343082 220464 343088 220516
rect 343140 220504 343146 220516
rect 386782 220504 386788 220516
rect 343140 220476 386788 220504
rect 343140 220464 343146 220476
rect 386782 220464 386788 220476
rect 386840 220464 386846 220516
rect 392578 220464 392584 220516
rect 392636 220504 392642 220516
rect 522574 220504 522580 220516
rect 392636 220476 522580 220504
rect 392636 220464 392642 220476
rect 522574 220464 522580 220476
rect 522632 220504 522638 220516
rect 560570 220504 560576 220516
rect 522632 220476 560576 220504
rect 522632 220464 522638 220476
rect 560570 220464 560576 220476
rect 560628 220464 560634 220516
rect 572686 220504 572714 220544
rect 574738 220532 574744 220584
rect 574796 220572 574802 220584
rect 575474 220572 575480 220584
rect 574796 220544 575480 220572
rect 574796 220532 574802 220544
rect 575474 220532 575480 220544
rect 575532 220532 575538 220584
rect 576394 220504 576400 220516
rect 572686 220476 576400 220504
rect 576394 220464 576400 220476
rect 576452 220464 576458 220516
rect 577130 220504 577136 220516
rect 576826 220476 577136 220504
rect 222562 220396 222568 220448
rect 222620 220436 222626 220448
rect 264330 220436 264336 220448
rect 222620 220408 264336 220436
rect 222620 220396 222626 220408
rect 264330 220396 264336 220408
rect 264388 220396 264394 220448
rect 299382 220396 299388 220448
rect 299440 220436 299446 220448
rect 305270 220436 305276 220448
rect 299440 220408 305276 220436
rect 299440 220396 299446 220408
rect 305270 220396 305276 220408
rect 305328 220396 305334 220448
rect 306098 220396 306104 220448
rect 306156 220436 306162 220448
rect 319530 220436 319536 220448
rect 306156 220408 319536 220436
rect 306156 220396 306162 220408
rect 319530 220396 319536 220408
rect 319588 220396 319594 220448
rect 330846 220396 330852 220448
rect 330904 220436 330910 220448
rect 375374 220436 375380 220448
rect 330904 220408 375380 220436
rect 330904 220396 330910 220408
rect 375374 220396 375380 220408
rect 375432 220396 375438 220448
rect 376018 220396 376024 220448
rect 376076 220436 376082 220448
rect 376076 220408 377260 220436
rect 376076 220396 376082 220408
rect 192352 220340 219434 220368
rect 192352 220328 192358 220340
rect 224310 220328 224316 220380
rect 224368 220368 224374 220380
rect 265434 220368 265440 220380
rect 224368 220340 265440 220368
rect 224368 220328 224374 220340
rect 265434 220328 265440 220340
rect 265492 220328 265498 220380
rect 307570 220328 307576 220380
rect 307628 220368 307634 220380
rect 321554 220368 321560 220380
rect 307628 220340 321560 220368
rect 307628 220328 307634 220340
rect 321554 220328 321560 220340
rect 321612 220328 321618 220380
rect 332226 220328 332232 220380
rect 332284 220368 332290 220380
rect 376202 220368 376208 220380
rect 332284 220340 376208 220368
rect 332284 220328 332290 220340
rect 376202 220328 376208 220340
rect 376260 220328 376266 220380
rect 377232 220368 377260 220408
rect 377306 220396 377312 220448
rect 377364 220436 377370 220448
rect 388530 220436 388536 220448
rect 377364 220408 388536 220436
rect 377364 220396 377370 220408
rect 388530 220396 388536 220408
rect 388588 220396 388594 220448
rect 394602 220396 394608 220448
rect 394660 220436 394666 220448
rect 527266 220436 527272 220448
rect 394660 220408 527272 220436
rect 394660 220396 394666 220408
rect 527266 220396 527272 220408
rect 527324 220436 527330 220448
rect 527324 220408 528554 220436
rect 527324 220396 527330 220408
rect 379606 220368 379612 220380
rect 377232 220340 379612 220368
rect 379606 220328 379612 220340
rect 379664 220328 379670 220380
rect 395614 220328 395620 220380
rect 395672 220368 395678 220380
rect 395672 220340 402974 220368
rect 395672 220328 395678 220340
rect 79594 220260 79600 220312
rect 79652 220300 79658 220312
rect 100754 220300 100760 220312
rect 79652 220272 100760 220300
rect 79652 220260 79658 220272
rect 100754 220260 100760 220272
rect 100812 220260 100818 220312
rect 104710 220260 104716 220312
rect 104768 220300 104774 220312
rect 203702 220300 203708 220312
rect 104768 220272 203708 220300
rect 104768 220260 104774 220272
rect 203702 220260 203708 220272
rect 203760 220260 203766 220312
rect 206186 220260 206192 220312
rect 206244 220300 206250 220312
rect 213914 220300 213920 220312
rect 206244 220272 213920 220300
rect 206244 220260 206250 220272
rect 213914 220260 213920 220272
rect 213972 220260 213978 220312
rect 217594 220260 217600 220312
rect 217652 220300 217658 220312
rect 260098 220300 260104 220312
rect 217652 220272 260104 220300
rect 217652 220260 217658 220272
rect 260098 220260 260104 220272
rect 260156 220260 260162 220312
rect 264698 220260 264704 220312
rect 264756 220300 264762 220312
rect 273806 220300 273812 220312
rect 264756 220272 273812 220300
rect 264756 220260 264762 220272
rect 273806 220260 273812 220272
rect 273864 220260 273870 220312
rect 283190 220260 283196 220312
rect 283248 220300 283254 220312
rect 284202 220300 284208 220312
rect 283248 220272 284208 220300
rect 283248 220260 283254 220272
rect 284202 220260 284208 220272
rect 284260 220260 284266 220312
rect 291562 220260 291568 220312
rect 291620 220300 291626 220312
rect 293954 220300 293960 220312
rect 291620 220272 293960 220300
rect 291620 220260 291626 220272
rect 293954 220260 293960 220272
rect 294012 220260 294018 220312
rect 307386 220260 307392 220312
rect 307444 220300 307450 220312
rect 322934 220300 322940 220312
rect 307444 220272 322940 220300
rect 307444 220260 307450 220272
rect 322934 220260 322940 220272
rect 322992 220260 322998 220312
rect 331030 220260 331036 220312
rect 331088 220300 331094 220312
rect 376938 220300 376944 220312
rect 331088 220272 376944 220300
rect 331088 220260 331094 220272
rect 376938 220260 376944 220272
rect 376996 220260 377002 220312
rect 378686 220260 378692 220312
rect 378744 220300 378750 220312
rect 391934 220300 391940 220312
rect 378744 220272 391940 220300
rect 378744 220260 378750 220272
rect 391934 220260 391940 220272
rect 391992 220260 391998 220312
rect 396810 220260 396816 220312
rect 396868 220300 396874 220312
rect 402946 220300 402974 220340
rect 415302 220328 415308 220380
rect 415360 220368 415366 220380
rect 418154 220368 418160 220380
rect 415360 220340 418160 220368
rect 415360 220328 415366 220340
rect 418154 220328 418160 220340
rect 418212 220328 418218 220380
rect 528526 220368 528554 220408
rect 560266 220408 569954 220436
rect 560266 220368 560294 220408
rect 528526 220340 560294 220368
rect 569926 220368 569954 220408
rect 574186 220368 574192 220380
rect 569926 220340 574192 220368
rect 574186 220328 574192 220340
rect 574244 220328 574250 220380
rect 532694 220300 532700 220312
rect 396868 220272 397040 220300
rect 402946 220272 532700 220300
rect 396868 220260 396874 220272
rect 94774 220192 94780 220244
rect 94832 220232 94838 220244
rect 202414 220232 202420 220244
rect 94832 220204 202420 220232
rect 94832 220192 94838 220204
rect 202414 220192 202420 220204
rect 202472 220192 202478 220244
rect 204530 220232 204536 220244
rect 202524 220204 204536 220232
rect 81250 220124 81256 220176
rect 81308 220164 81314 220176
rect 202524 220164 202552 220204
rect 204530 220192 204536 220204
rect 204588 220192 204594 220244
rect 207474 220192 207480 220244
rect 207532 220232 207538 220244
rect 213822 220232 213828 220244
rect 207532 220204 213828 220232
rect 207532 220192 207538 220204
rect 213822 220192 213828 220204
rect 213880 220192 213886 220244
rect 215846 220192 215852 220244
rect 215904 220232 215910 220244
rect 261478 220232 261484 220244
rect 215904 220204 261484 220232
rect 215904 220192 215910 220204
rect 261478 220192 261484 220204
rect 261536 220192 261542 220244
rect 262582 220192 262588 220244
rect 262640 220232 262646 220244
rect 267182 220232 267188 220244
rect 262640 220204 267188 220232
rect 262640 220192 262646 220204
rect 267182 220192 267188 220204
rect 267240 220192 267246 220244
rect 304902 220192 304908 220244
rect 304960 220232 304966 220244
rect 314654 220232 314660 220244
rect 304960 220204 314660 220232
rect 304960 220192 304966 220204
rect 314654 220192 314660 220204
rect 314712 220192 314718 220244
rect 315390 220192 315396 220244
rect 315448 220232 315454 220244
rect 332962 220232 332968 220244
rect 315448 220204 332968 220232
rect 315448 220192 315454 220204
rect 332962 220192 332968 220204
rect 333020 220192 333026 220244
rect 333882 220192 333888 220244
rect 333940 220232 333946 220244
rect 381814 220232 381820 220244
rect 333940 220204 381820 220232
rect 333940 220192 333946 220204
rect 381814 220192 381820 220204
rect 381872 220192 381878 220244
rect 382274 220192 382280 220244
rect 382332 220232 382338 220244
rect 396902 220232 396908 220244
rect 382332 220204 396908 220232
rect 382332 220192 382338 220204
rect 396902 220192 396908 220204
rect 396960 220192 396966 220244
rect 397012 220232 397040 220272
rect 532694 220260 532700 220272
rect 532752 220260 532758 220312
rect 560570 220260 560576 220312
rect 560628 220300 560634 220312
rect 576826 220300 576854 220476
rect 577130 220464 577136 220476
rect 577188 220464 577194 220516
rect 560628 220272 576854 220300
rect 560628 220260 560634 220272
rect 535362 220232 535368 220244
rect 397012 220204 535368 220232
rect 535362 220192 535368 220204
rect 535420 220232 535426 220244
rect 605926 220232 605932 220244
rect 535420 220204 605932 220232
rect 535420 220192 535426 220204
rect 605926 220192 605932 220204
rect 605984 220192 605990 220244
rect 674650 220192 674656 220244
rect 674708 220232 674714 220244
rect 676030 220232 676036 220244
rect 674708 220204 676036 220232
rect 674708 220192 674714 220204
rect 676030 220192 676036 220204
rect 676088 220192 676094 220244
rect 81308 220136 202552 220164
rect 81308 220124 81314 220136
rect 204070 220124 204076 220176
rect 204128 220164 204134 220176
rect 209866 220164 209872 220176
rect 204128 220136 209872 220164
rect 204128 220124 204134 220136
rect 209866 220124 209872 220136
rect 209924 220124 209930 220176
rect 210786 220124 210792 220176
rect 210844 220164 210850 220176
rect 210844 220136 252232 220164
rect 210844 220124 210850 220136
rect 64506 220056 64512 220108
rect 64564 220096 64570 220108
rect 192846 220096 192852 220108
rect 64564 220068 192852 220096
rect 64564 220056 64570 220068
rect 192846 220056 192852 220068
rect 192904 220056 192910 220108
rect 209130 220056 209136 220108
rect 209188 220096 209194 220108
rect 252094 220096 252100 220108
rect 209188 220068 252100 220096
rect 209188 220056 209194 220068
rect 252094 220056 252100 220068
rect 252152 220056 252158 220108
rect 252204 220096 252232 220136
rect 254578 220124 254584 220176
rect 254636 220164 254642 220176
rect 255222 220164 255228 220176
rect 254636 220136 255228 220164
rect 254636 220124 254642 220136
rect 255222 220124 255228 220136
rect 255280 220124 255286 220176
rect 257890 220124 257896 220176
rect 257948 220164 257954 220176
rect 271230 220164 271236 220176
rect 257948 220136 271236 220164
rect 257948 220124 257954 220136
rect 271230 220124 271236 220136
rect 271288 220124 271294 220176
rect 279418 220164 279424 220176
rect 277366 220136 279424 220164
rect 255958 220096 255964 220108
rect 252204 220068 255964 220096
rect 255958 220056 255964 220068
rect 256016 220056 256022 220108
rect 266170 220056 266176 220108
rect 266228 220096 266234 220108
rect 277366 220096 277394 220136
rect 279418 220124 279424 220136
rect 279476 220124 279482 220176
rect 280614 220124 280620 220176
rect 280672 220164 280678 220176
rect 281442 220164 281448 220176
rect 280672 220136 281448 220164
rect 280672 220124 280678 220136
rect 281442 220124 281448 220136
rect 281500 220124 281506 220176
rect 287514 220164 287520 220176
rect 281552 220136 287520 220164
rect 266228 220068 277394 220096
rect 266228 220056 266234 220068
rect 278590 220056 278596 220108
rect 278648 220096 278654 220108
rect 281552 220096 281580 220136
rect 287514 220124 287520 220136
rect 287572 220124 287578 220176
rect 308766 220124 308772 220176
rect 308824 220164 308830 220176
rect 326246 220164 326252 220176
rect 308824 220136 326252 220164
rect 308824 220124 308830 220136
rect 326246 220124 326252 220136
rect 326304 220124 326310 220176
rect 332410 220124 332416 220176
rect 332468 220164 332474 220176
rect 380066 220164 380072 220176
rect 332468 220136 380072 220164
rect 332468 220124 332474 220136
rect 380066 220124 380072 220136
rect 380124 220124 380130 220176
rect 380158 220124 380164 220176
rect 380216 220164 380222 220176
rect 395246 220164 395252 220176
rect 380216 220136 395252 220164
rect 380216 220124 380222 220136
rect 395246 220124 395252 220136
rect 395304 220124 395310 220176
rect 398558 220124 398564 220176
rect 398616 220164 398622 220176
rect 537386 220164 537392 220176
rect 398616 220136 537392 220164
rect 398616 220124 398622 220136
rect 537386 220124 537392 220136
rect 537444 220124 537450 220176
rect 548150 220124 548156 220176
rect 548208 220164 548214 220176
rect 615494 220164 615500 220176
rect 548208 220136 615500 220164
rect 548208 220124 548214 220136
rect 615494 220124 615500 220136
rect 615552 220124 615558 220176
rect 278648 220068 281580 220096
rect 278648 220056 278654 220068
rect 284846 220056 284852 220108
rect 284904 220096 284910 220108
rect 285490 220096 285496 220108
rect 284904 220068 285496 220096
rect 284904 220056 284910 220068
rect 285490 220056 285496 220068
rect 285548 220056 285554 220108
rect 301958 220056 301964 220108
rect 302016 220096 302022 220108
rect 309410 220096 309416 220108
rect 302016 220068 309416 220096
rect 302016 220056 302022 220068
rect 309410 220056 309416 220068
rect 309468 220056 309474 220108
rect 310238 220056 310244 220108
rect 310296 220096 310302 220108
rect 329834 220096 329840 220108
rect 310296 220068 329840 220096
rect 310296 220056 310302 220068
rect 329834 220056 329840 220068
rect 329892 220056 329898 220108
rect 333790 220056 333796 220108
rect 333848 220096 333854 220108
rect 383654 220096 383660 220108
rect 333848 220068 383660 220096
rect 333848 220056 333854 220068
rect 383654 220056 383660 220068
rect 383712 220056 383718 220108
rect 385678 220056 385684 220108
rect 385736 220096 385742 220108
rect 400306 220096 400312 220108
rect 385736 220068 400312 220096
rect 385736 220056 385742 220068
rect 400306 220056 400312 220068
rect 400364 220056 400370 220108
rect 404262 220056 404268 220108
rect 404320 220096 404326 220108
rect 549990 220096 549996 220108
rect 404320 220068 549996 220096
rect 404320 220056 404326 220068
rect 549990 220056 549996 220068
rect 550048 220056 550054 220108
rect 551278 220056 551284 220108
rect 551336 220096 551342 220108
rect 609606 220096 609612 220108
rect 551336 220068 609612 220096
rect 551336 220056 551342 220068
rect 609606 220056 609612 220068
rect 609664 220056 609670 220108
rect 148594 219988 148600 220040
rect 148652 220028 148658 220040
rect 223114 220028 223120 220040
rect 148652 220000 223120 220028
rect 148652 219988 148658 220000
rect 223114 219988 223120 220000
rect 223172 219988 223178 220040
rect 247862 219988 247868 220040
rect 247920 220028 247926 220040
rect 248322 220028 248328 220040
rect 247920 220000 248328 220028
rect 247920 219988 247926 220000
rect 248322 219988 248328 220000
rect 248380 219988 248386 220040
rect 272886 220028 272892 220040
rect 249536 220000 272892 220028
rect 151722 219920 151728 219972
rect 151780 219960 151786 219972
rect 224034 219960 224040 219972
rect 151780 219932 224040 219960
rect 151780 219920 151786 219932
rect 224034 219920 224040 219932
rect 224092 219920 224098 219972
rect 246114 219920 246120 219972
rect 246172 219960 246178 219972
rect 246942 219960 246948 219972
rect 246172 219932 246948 219960
rect 246172 219920 246178 219932
rect 246942 219920 246948 219932
rect 247000 219920 247006 219972
rect 249536 219960 249564 220000
rect 272886 219988 272892 220000
rect 272944 219988 272950 220040
rect 289630 219988 289636 220040
rect 289688 220028 289694 220040
rect 292850 220028 292856 220040
rect 289688 220000 292856 220028
rect 289688 219988 289694 220000
rect 292850 219988 292856 220000
rect 292908 219988 292914 220040
rect 319346 219988 319352 220040
rect 319404 220028 319410 220040
rect 339678 220028 339684 220040
rect 319404 220000 339684 220028
rect 319404 219988 319410 220000
rect 339678 219988 339684 220000
rect 339736 219988 339742 220040
rect 341518 219988 341524 220040
rect 341576 220028 341582 220040
rect 370038 220028 370044 220040
rect 341576 220000 370044 220028
rect 341576 219988 341582 220000
rect 370038 219988 370044 220000
rect 370096 219988 370102 220040
rect 370222 219988 370228 220040
rect 370280 220028 370286 220040
rect 382642 220028 382648 220040
rect 370280 220000 382648 220028
rect 370280 219988 370286 220000
rect 382642 219988 382648 220000
rect 382700 219988 382706 220040
rect 384942 219988 384948 220040
rect 385000 220028 385006 220040
rect 505002 220028 505008 220040
rect 385000 220000 505008 220028
rect 385000 219988 385006 220000
rect 505002 219988 505008 220000
rect 505060 219988 505066 220040
rect 542998 219988 543004 220040
rect 543056 220028 543062 220040
rect 614114 220028 614120 220040
rect 543056 220000 614120 220028
rect 543056 219988 543062 220000
rect 614114 219988 614120 220000
rect 614172 219988 614178 220040
rect 276198 219960 276204 219972
rect 248386 219932 249564 219960
rect 249628 219932 276204 219960
rect 158622 219852 158628 219904
rect 158680 219892 158686 219904
rect 227346 219892 227352 219904
rect 158680 219864 227352 219892
rect 158680 219852 158686 219864
rect 227346 219852 227352 219864
rect 227404 219852 227410 219904
rect 242802 219852 242808 219904
rect 242860 219892 242866 219904
rect 248386 219892 248414 219932
rect 242860 219864 248414 219892
rect 242860 219852 242866 219864
rect 249518 219852 249524 219904
rect 249576 219892 249582 219904
rect 249628 219892 249656 219932
rect 276198 219920 276204 219932
rect 276256 219920 276262 219972
rect 318058 219920 318064 219972
rect 318116 219960 318122 219972
rect 336734 219960 336740 219972
rect 318116 219932 336740 219960
rect 318116 219920 318122 219932
rect 336734 219920 336740 219932
rect 336792 219920 336798 219972
rect 340138 219920 340144 219972
rect 340196 219960 340202 219972
rect 360194 219960 360200 219972
rect 340196 219932 360200 219960
rect 340196 219920 340202 219932
rect 360194 219920 360200 219932
rect 360252 219920 360258 219972
rect 363138 219920 363144 219972
rect 363196 219960 363202 219972
rect 391014 219960 391020 219972
rect 363196 219932 391020 219960
rect 363196 219920 363202 219932
rect 391014 219920 391020 219932
rect 391072 219920 391078 219972
rect 391106 219920 391112 219972
rect 391164 219960 391170 219972
rect 509878 219960 509884 219972
rect 391164 219932 509884 219960
rect 391164 219920 391170 219932
rect 509878 219920 509884 219932
rect 509936 219920 509942 219972
rect 540422 219920 540428 219972
rect 540480 219960 540486 219972
rect 613378 219960 613384 219972
rect 540480 219932 613384 219960
rect 540480 219920 540486 219932
rect 613378 219920 613384 219932
rect 613436 219920 613442 219972
rect 249576 219864 249656 219892
rect 249576 219852 249582 219864
rect 252922 219852 252928 219904
rect 252980 219892 252986 219904
rect 277578 219892 277584 219904
rect 252980 219864 277584 219892
rect 252980 219852 252986 219864
rect 277578 219852 277584 219864
rect 277636 219852 277642 219904
rect 338758 219852 338764 219904
rect 338816 219892 338822 219904
rect 356514 219892 356520 219904
rect 338816 219864 356520 219892
rect 338816 219852 338822 219864
rect 356514 219852 356520 219864
rect 356572 219852 356578 219904
rect 365346 219852 365352 219904
rect 365404 219892 365410 219904
rect 377582 219892 377588 219904
rect 365404 219864 377588 219892
rect 365404 219852 365410 219864
rect 377582 219852 377588 219864
rect 377640 219852 377646 219904
rect 386966 219852 386972 219904
rect 387024 219892 387030 219904
rect 398834 219892 398840 219904
rect 387024 219864 398840 219892
rect 387024 219852 387030 219864
rect 398834 219852 398840 219864
rect 398892 219852 398898 219904
rect 400674 219852 400680 219904
rect 400732 219892 400738 219904
rect 513834 219892 513840 219904
rect 400732 219864 513840 219892
rect 400732 219852 400738 219864
rect 513834 219852 513840 219864
rect 513892 219852 513898 219904
rect 517514 219852 517520 219904
rect 517572 219892 517578 219904
rect 574830 219892 574836 219904
rect 517572 219864 574836 219892
rect 517572 219852 517578 219864
rect 574830 219852 574836 219864
rect 574888 219852 574894 219904
rect 673270 219852 673276 219904
rect 673328 219892 673334 219904
rect 676030 219892 676036 219904
rect 673328 219864 676036 219892
rect 673328 219852 673334 219864
rect 676030 219852 676036 219864
rect 676088 219852 676094 219904
rect 165430 219784 165436 219836
rect 165488 219824 165494 219836
rect 227714 219824 227720 219836
rect 165488 219796 227720 219824
rect 165488 219784 165494 219796
rect 227714 219784 227720 219796
rect 227772 219784 227778 219836
rect 256234 219784 256240 219836
rect 256292 219824 256298 219836
rect 278958 219824 278964 219836
rect 256292 219796 278964 219824
rect 256292 219784 256298 219796
rect 278958 219784 278964 219796
rect 279016 219784 279022 219836
rect 337378 219784 337384 219836
rect 337436 219824 337442 219836
rect 353294 219824 353300 219836
rect 337436 219796 353300 219824
rect 337436 219784 337442 219796
rect 353294 219784 353300 219796
rect 353352 219784 353358 219836
rect 362954 219784 362960 219836
rect 363012 219824 363018 219836
rect 368474 219824 368480 219836
rect 363012 219796 368480 219824
rect 363012 219784 363018 219796
rect 368474 219784 368480 219796
rect 368532 219784 368538 219836
rect 376202 219784 376208 219836
rect 376260 219824 376266 219836
rect 378410 219824 378416 219836
rect 376260 219796 378416 219824
rect 376260 219784 376266 219796
rect 378410 219784 378416 219796
rect 378468 219784 378474 219836
rect 379698 219784 379704 219836
rect 379756 219824 379762 219836
rect 484394 219824 484400 219836
rect 379756 219796 484400 219824
rect 379756 219784 379762 219796
rect 484394 219784 484400 219796
rect 484452 219784 484458 219836
rect 529934 219784 529940 219836
rect 529992 219824 529998 219836
rect 611998 219824 612004 219836
rect 529992 219796 612004 219824
rect 529992 219784 529998 219796
rect 611998 219784 612004 219796
rect 612056 219784 612062 219836
rect 172146 219716 172152 219768
rect 172204 219756 172210 219768
rect 232406 219756 232412 219768
rect 172204 219728 232412 219756
rect 172204 219716 172210 219728
rect 232406 219716 232412 219728
rect 232464 219716 232470 219768
rect 250990 219716 250996 219768
rect 251048 219756 251054 219768
rect 271322 219756 271328 219768
rect 251048 219728 271328 219756
rect 251048 219716 251054 219728
rect 271322 219716 271328 219728
rect 271380 219716 271386 219768
rect 334710 219716 334716 219768
rect 334768 219756 334774 219768
rect 349798 219756 349804 219768
rect 334768 219728 349804 219756
rect 334768 219716 334774 219728
rect 349798 219716 349804 219728
rect 349856 219716 349862 219768
rect 372614 219716 372620 219768
rect 372672 219756 372678 219768
rect 384298 219756 384304 219768
rect 372672 219728 384304 219756
rect 372672 219716 372678 219728
rect 384298 219716 384304 219728
rect 384356 219716 384362 219768
rect 387242 219716 387248 219768
rect 387300 219756 387306 219768
rect 409874 219756 409880 219768
rect 387300 219728 409880 219756
rect 387300 219716 387306 219728
rect 409874 219716 409880 219728
rect 409932 219716 409938 219768
rect 409966 219716 409972 219768
rect 410024 219756 410030 219768
rect 416222 219756 416228 219768
rect 410024 219728 416228 219756
rect 410024 219716 410030 219728
rect 416222 219716 416228 219728
rect 416280 219716 416286 219768
rect 515398 219716 515404 219768
rect 515456 219756 515462 219768
rect 625246 219756 625252 219768
rect 515456 219728 625252 219756
rect 515456 219716 515462 219728
rect 625246 219716 625252 219728
rect 625304 219716 625310 219768
rect 185578 219648 185584 219700
rect 185636 219688 185642 219700
rect 186958 219688 186964 219700
rect 185636 219660 186964 219688
rect 185636 219648 185642 219660
rect 186958 219648 186964 219660
rect 187016 219648 187022 219700
rect 232774 219688 232780 219700
rect 187068 219660 232780 219688
rect 181990 219580 181996 219632
rect 182048 219620 182054 219632
rect 187068 219620 187096 219660
rect 232774 219648 232780 219660
rect 232832 219648 232838 219700
rect 252094 219648 252100 219700
rect 252152 219688 252158 219700
rect 257338 219688 257344 219700
rect 252152 219660 257344 219688
rect 252152 219648 252158 219660
rect 257338 219648 257344 219660
rect 257396 219648 257402 219700
rect 268010 219648 268016 219700
rect 268068 219688 268074 219700
rect 275278 219688 275284 219700
rect 268068 219660 275284 219688
rect 268068 219648 268074 219660
rect 275278 219648 275284 219660
rect 275336 219648 275342 219700
rect 334618 219648 334624 219700
rect 334676 219688 334682 219700
rect 346486 219688 346492 219700
rect 334676 219660 346492 219688
rect 334676 219648 334682 219660
rect 346486 219648 346492 219660
rect 346544 219648 346550 219700
rect 378042 219648 378048 219700
rect 378100 219688 378106 219700
rect 387794 219688 387800 219700
rect 378100 219660 387800 219688
rect 378100 219648 378106 219660
rect 387794 219648 387800 219660
rect 387852 219648 387858 219700
rect 512822 219648 512828 219700
rect 512880 219688 512886 219700
rect 625522 219688 625528 219700
rect 512880 219660 625528 219688
rect 512880 219648 512886 219660
rect 625522 219648 625528 219660
rect 625580 219648 625586 219700
rect 182048 219592 187096 219620
rect 182048 219580 182054 219592
rect 188890 219580 188896 219632
rect 188948 219620 188954 219632
rect 234614 219620 234620 219632
rect 188948 219592 234620 219620
rect 188948 219580 188954 219592
rect 234614 219580 234620 219592
rect 234672 219580 234678 219632
rect 261294 219580 261300 219632
rect 261352 219620 261358 219632
rect 272978 219620 272984 219632
rect 261352 219592 272984 219620
rect 261352 219580 261358 219592
rect 272978 219580 272984 219592
rect 273036 219580 273042 219632
rect 300486 219580 300492 219632
rect 300544 219620 300550 219632
rect 306926 219620 306932 219632
rect 300544 219592 306932 219620
rect 300544 219580 300550 219592
rect 306926 219580 306932 219592
rect 306984 219580 306990 219632
rect 406378 219580 406384 219632
rect 406436 219620 406442 219632
rect 412910 219620 412916 219632
rect 406436 219592 412916 219620
rect 406436 219580 406442 219592
rect 412910 219580 412916 219592
rect 412968 219580 412974 219632
rect 509878 219580 509884 219632
rect 509936 219620 509942 219632
rect 623774 219620 623780 219632
rect 509936 219592 623780 219620
rect 509936 219580 509942 219592
rect 623774 219580 623780 219592
rect 623832 219580 623838 219632
rect 61102 219512 61108 219564
rect 61160 219552 61166 219564
rect 66898 219552 66904 219564
rect 61160 219524 66904 219552
rect 61160 219512 61166 219524
rect 66898 219512 66904 219524
rect 66956 219512 66962 219564
rect 97810 219512 97816 219564
rect 97868 219552 97874 219564
rect 97868 219524 103514 219552
rect 97868 219512 97874 219524
rect 103486 219484 103514 219524
rect 195698 219512 195704 219564
rect 195756 219552 195762 219564
rect 234706 219552 234712 219564
rect 195756 219524 234712 219552
rect 195756 219512 195762 219524
rect 234706 219512 234712 219524
rect 234764 219512 234770 219564
rect 301590 219512 301596 219564
rect 301648 219552 301654 219564
rect 307754 219552 307760 219564
rect 301648 219524 307760 219552
rect 301648 219512 301654 219524
rect 307754 219512 307760 219524
rect 307812 219512 307818 219564
rect 408494 219512 408500 219564
rect 408552 219552 408558 219564
rect 414566 219552 414572 219564
rect 408552 219524 414572 219552
rect 408552 219512 408558 219524
rect 414566 219512 414572 219524
rect 414624 219512 414630 219564
rect 502426 219512 502432 219564
rect 502484 219552 502490 219564
rect 622946 219552 622952 219564
rect 502484 219524 622952 219552
rect 502484 219512 502490 219524
rect 622946 219512 622952 219524
rect 623004 219512 623010 219564
rect 195146 219484 195152 219496
rect 103486 219456 195152 219484
rect 195146 219444 195152 219456
rect 195204 219444 195210 219496
rect 202414 219444 202420 219496
rect 202472 219484 202478 219496
rect 237374 219484 237380 219496
rect 202472 219456 237380 219484
rect 202472 219444 202478 219456
rect 237374 219444 237380 219456
rect 237432 219444 237438 219496
rect 267182 219444 267188 219496
rect 267240 219484 267246 219496
rect 268378 219484 268384 219496
rect 267240 219456 268384 219484
rect 267240 219444 267246 219456
rect 268378 219444 268384 219456
rect 268436 219444 268442 219496
rect 276474 219444 276480 219496
rect 276532 219484 276538 219496
rect 278038 219484 278044 219496
rect 276532 219456 278044 219484
rect 276532 219444 276538 219456
rect 278038 219444 278044 219456
rect 278096 219444 278102 219496
rect 300578 219444 300584 219496
rect 300636 219484 300642 219496
rect 306374 219484 306380 219496
rect 300636 219456 306380 219484
rect 300636 219444 300642 219456
rect 306374 219444 306380 219456
rect 306432 219444 306438 219496
rect 360286 219444 360292 219496
rect 360344 219484 360350 219496
rect 364978 219484 364984 219496
rect 360344 219456 364984 219484
rect 360344 219444 360350 219456
rect 364978 219444 364984 219456
rect 365036 219444 365042 219496
rect 371326 219444 371332 219496
rect 371384 219484 371390 219496
rect 375926 219484 375932 219496
rect 371384 219456 375932 219484
rect 371384 219444 371390 219456
rect 375926 219444 375932 219456
rect 375984 219444 375990 219496
rect 378502 219444 378508 219496
rect 378560 219484 378566 219496
rect 385126 219484 385132 219496
rect 378560 219456 385132 219484
rect 378560 219444 378566 219456
rect 385126 219444 385132 219456
rect 385184 219444 385190 219496
rect 390646 219444 390652 219496
rect 390704 219484 390710 219496
rect 393590 219484 393596 219496
rect 390704 219456 393596 219484
rect 390704 219444 390710 219456
rect 393590 219444 393596 219456
rect 393648 219444 393654 219496
rect 394510 219444 394516 219496
rect 394568 219484 394574 219496
rect 529934 219484 529940 219496
rect 394568 219456 529940 219484
rect 394568 219444 394574 219456
rect 529934 219444 529940 219456
rect 529992 219444 529998 219496
rect 565446 219444 565452 219496
rect 565504 219484 565510 219496
rect 577038 219484 577044 219496
rect 565504 219456 574692 219484
rect 565504 219444 565510 219456
rect 354398 219376 354404 219428
rect 354456 219416 354462 219428
rect 432230 219416 432236 219428
rect 354456 219388 432236 219416
rect 354456 219376 354462 219388
rect 432230 219376 432236 219388
rect 432288 219376 432294 219428
rect 574664 219416 574692 219456
rect 575584 219456 577044 219484
rect 575584 219416 575612 219456
rect 577038 219444 577044 219456
rect 577096 219444 577102 219496
rect 574664 219388 575612 219416
rect 353202 219308 353208 219360
rect 353260 219348 353266 219360
rect 430574 219348 430580 219360
rect 353260 219320 430580 219348
rect 353260 219308 353266 219320
rect 430574 219308 430580 219320
rect 430632 219308 430638 219360
rect 379422 219240 379428 219292
rect 379480 219280 379486 219292
rect 494514 219280 494520 219292
rect 379480 219252 494520 219280
rect 379480 219240 379486 219252
rect 494514 219240 494520 219252
rect 494572 219240 494578 219292
rect 380802 219172 380808 219224
rect 380860 219212 380866 219224
rect 498194 219212 498200 219224
rect 380860 219184 498200 219212
rect 380860 219172 380866 219184
rect 498194 219172 498200 219184
rect 498252 219172 498258 219224
rect 567930 219172 567936 219224
rect 567988 219212 567994 219224
rect 616782 219212 616788 219224
rect 567988 219184 616788 219212
rect 567988 219172 567994 219184
rect 616782 219172 616788 219184
rect 616840 219172 616846 219224
rect 383562 219104 383568 219156
rect 383620 219144 383626 219156
rect 501230 219144 501236 219156
rect 383620 219116 501236 219144
rect 383620 219104 383626 219116
rect 501230 219104 501236 219116
rect 501288 219104 501294 219156
rect 545758 219104 545764 219156
rect 545816 219144 545822 219156
rect 576302 219144 576308 219156
rect 545816 219116 576308 219144
rect 545816 219104 545822 219116
rect 576302 219104 576308 219116
rect 576360 219104 576366 219156
rect 383470 219036 383476 219088
rect 383528 219076 383534 219088
rect 503714 219076 503720 219088
rect 383528 219048 503720 219076
rect 383528 219036 383534 219048
rect 503714 219036 503720 219048
rect 503772 219036 503778 219088
rect 543182 219036 543188 219088
rect 543240 219076 543246 219088
rect 543642 219076 543648 219088
rect 543240 219048 543648 219076
rect 543240 219036 543246 219048
rect 543642 219036 543648 219048
rect 543700 219076 543706 219088
rect 576210 219076 576216 219088
rect 543700 219048 576216 219076
rect 543700 219036 543706 219048
rect 576210 219036 576216 219048
rect 576268 219036 576274 219088
rect 386322 218968 386328 219020
rect 386380 219008 386386 219020
rect 508774 219008 508780 219020
rect 386380 218980 508780 219008
rect 386380 218968 386386 218980
rect 508774 218968 508780 218980
rect 508832 218968 508838 219020
rect 541434 218968 541440 219020
rect 541492 219008 541498 219020
rect 576118 219008 576124 219020
rect 541492 218980 576124 219008
rect 541492 218968 541498 218980
rect 576118 218968 576124 218980
rect 576176 218968 576182 219020
rect 35710 218900 35716 218952
rect 35768 218940 35774 218952
rect 55950 218940 55956 218952
rect 35768 218912 55956 218940
rect 35768 218900 35774 218912
rect 55950 218900 55956 218912
rect 56008 218900 56014 218952
rect 387702 218900 387708 218952
rect 387760 218940 387766 218952
rect 511350 218940 511356 218952
rect 387760 218912 511356 218940
rect 387760 218900 387766 218912
rect 511350 218900 511356 218912
rect 511408 218900 511414 218952
rect 570598 218900 570604 218952
rect 570656 218940 570662 218952
rect 617518 218940 617524 218952
rect 570656 218912 617524 218940
rect 570656 218900 570662 218912
rect 617518 218900 617524 218912
rect 617576 218900 617582 218952
rect 47578 218832 47584 218884
rect 47636 218872 47642 218884
rect 647142 218872 647148 218884
rect 47636 218844 647148 218872
rect 47636 218832 47642 218844
rect 647142 218832 647148 218844
rect 647200 218832 647206 218884
rect 55858 218764 55864 218816
rect 55916 218804 55922 218816
rect 656894 218804 656900 218816
rect 55916 218776 656900 218804
rect 55916 218764 55922 218776
rect 656894 218764 656900 218776
rect 656952 218764 656958 218816
rect 45002 218696 45008 218748
rect 45060 218736 45066 218748
rect 662506 218736 662512 218748
rect 45060 218708 662512 218736
rect 45060 218696 45066 218708
rect 662506 218696 662512 218708
rect 662564 218696 662570 218748
rect 553670 218628 553676 218680
rect 553728 218668 553734 218680
rect 576026 218668 576032 218680
rect 553728 218640 576032 218668
rect 553728 218628 553734 218640
rect 576026 218628 576032 218640
rect 576084 218628 576090 218680
rect 518158 218560 518164 218612
rect 518216 218600 518222 218612
rect 518434 218600 518440 218612
rect 518216 218572 518440 218600
rect 518216 218560 518222 218572
rect 518434 218560 518440 218572
rect 518492 218600 518498 218612
rect 575934 218600 575940 218612
rect 518492 218572 575940 218600
rect 518492 218560 518498 218572
rect 575934 218560 575940 218572
rect 575992 218560 575998 218612
rect 515490 218492 515496 218544
rect 515548 218532 515554 218544
rect 516042 218532 516048 218544
rect 515548 218504 516048 218532
rect 515548 218492 515554 218504
rect 516042 218492 516048 218504
rect 516100 218532 516106 218544
rect 608410 218532 608416 218544
rect 516100 218504 608416 218532
rect 516100 218492 516106 218504
rect 608410 218492 608416 218504
rect 608468 218492 608474 218544
rect 511258 218424 511264 218476
rect 511316 218464 511322 218476
rect 609882 218464 609888 218476
rect 511316 218436 609888 218464
rect 511316 218424 511322 218436
rect 609882 218424 609888 218436
rect 609940 218424 609946 218476
rect 487798 218356 487804 218408
rect 487856 218396 487862 218408
rect 606662 218396 606668 218408
rect 487856 218368 606668 218396
rect 487856 218356 487862 218368
rect 606662 218356 606668 218368
rect 606720 218356 606726 218408
rect 489362 218288 489368 218340
rect 489420 218328 489426 218340
rect 489822 218328 489828 218340
rect 489420 218300 489828 218328
rect 489420 218288 489426 218300
rect 489822 218288 489828 218300
rect 489880 218328 489886 218340
rect 620278 218328 620284 218340
rect 489880 218300 620284 218328
rect 489880 218288 489886 218300
rect 620278 218288 620284 218300
rect 620336 218288 620342 218340
rect 499666 218220 499672 218272
rect 499724 218260 499730 218272
rect 500218 218260 500224 218272
rect 499724 218232 500224 218260
rect 499724 218220 499730 218232
rect 500218 218220 500224 218232
rect 500276 218260 500282 218272
rect 636010 218260 636016 218272
rect 500276 218232 636016 218260
rect 500276 218220 500282 218232
rect 636010 218220 636016 218232
rect 636068 218220 636074 218272
rect 493410 218152 493416 218204
rect 493468 218192 493474 218204
rect 629938 218192 629944 218204
rect 493468 218164 629944 218192
rect 493468 218152 493474 218164
rect 629938 218152 629944 218164
rect 629996 218152 630002 218204
rect 486418 218084 486424 218136
rect 486476 218124 486482 218136
rect 486476 218096 489914 218124
rect 486476 218084 486482 218096
rect 487522 218016 487528 218068
rect 487580 218056 487586 218068
rect 487798 218056 487804 218068
rect 487580 218028 487804 218056
rect 487580 218016 487586 218028
rect 487798 218016 487804 218028
rect 487856 218016 487862 218068
rect 489886 218056 489914 218096
rect 496078 218084 496084 218136
rect 496136 218124 496142 218136
rect 636102 218124 636108 218136
rect 496136 218096 636108 218124
rect 496136 218084 496142 218096
rect 636102 218084 636108 218096
rect 636160 218084 636166 218136
rect 638310 218056 638316 218068
rect 489886 218028 638316 218056
rect 638310 218016 638316 218028
rect 638368 218016 638374 218068
rect 523034 217880 523040 217932
rect 523092 217920 523098 217932
rect 523954 217920 523960 217932
rect 523092 217892 523960 217920
rect 523092 217880 523098 217892
rect 523954 217880 523960 217892
rect 524012 217880 524018 217932
rect 538214 217880 538220 217932
rect 538272 217920 538278 217932
rect 539042 217920 539048 217932
rect 538272 217892 539048 217920
rect 538272 217880 538278 217892
rect 539042 217880 539048 217892
rect 539100 217880 539106 217932
rect 296714 217812 296720 217864
rect 296772 217852 296778 217864
rect 297634 217852 297640 217864
rect 296772 217824 297640 217852
rect 296772 217812 296778 217824
rect 297634 217812 297640 217824
rect 297692 217812 297698 217864
rect 299566 217812 299572 217864
rect 299624 217852 299630 217864
rect 300210 217852 300216 217864
rect 299624 217824 300216 217852
rect 299624 217812 299630 217824
rect 300210 217812 300216 217824
rect 300268 217812 300274 217864
rect 331214 217812 331220 217864
rect 331272 217852 331278 217864
rect 332134 217852 332140 217864
rect 331272 217824 332140 217852
rect 331272 217812 331278 217824
rect 332134 217812 332140 217824
rect 332192 217812 332198 217864
rect 333974 217812 333980 217864
rect 334032 217852 334038 217864
rect 334710 217852 334716 217864
rect 334032 217824 334716 217852
rect 334032 217812 334038 217824
rect 334710 217812 334716 217824
rect 334768 217812 334774 217864
rect 350626 217812 350632 217864
rect 350684 217852 350690 217864
rect 351454 217852 351460 217864
rect 350684 217824 351460 217852
rect 350684 217812 350690 217824
rect 351454 217812 351460 217824
rect 351512 217812 351518 217864
rect 434714 217812 434720 217864
rect 434772 217852 434778 217864
rect 435634 217852 435640 217864
rect 434772 217824 435640 217852
rect 434772 217812 434778 217824
rect 435634 217812 435640 217824
rect 435692 217812 435698 217864
rect 441614 217812 441620 217864
rect 441672 217852 441678 217864
rect 442350 217852 442356 217864
rect 441672 217824 442356 217852
rect 441672 217812 441678 217824
rect 442350 217812 442356 217824
rect 442408 217812 442414 217864
rect 454034 217812 454040 217864
rect 454092 217852 454098 217864
rect 454954 217852 454960 217864
rect 454092 217824 454960 217852
rect 454092 217812 454098 217824
rect 454954 217812 454960 217824
rect 455012 217812 455018 217864
rect 460934 217812 460940 217864
rect 460992 217852 460998 217864
rect 461670 217852 461676 217864
rect 460992 217824 461676 217852
rect 460992 217812 460998 217824
rect 461670 217812 461676 217824
rect 461728 217812 461734 217864
rect 465074 217812 465080 217864
rect 465132 217852 465138 217864
rect 465902 217852 465908 217864
rect 465132 217824 465908 217852
rect 465132 217812 465138 217824
rect 465902 217812 465908 217824
rect 465960 217812 465966 217864
rect 471974 217812 471980 217864
rect 472032 217852 472038 217864
rect 472618 217852 472624 217864
rect 472032 217824 472624 217852
rect 472032 217812 472038 217824
rect 472618 217812 472624 217824
rect 472676 217812 472682 217864
rect 476114 217812 476120 217864
rect 476172 217852 476178 217864
rect 476850 217852 476856 217864
rect 476172 217824 476856 217852
rect 476172 217812 476178 217824
rect 476850 217812 476856 217824
rect 476908 217812 476914 217864
rect 491386 217812 491392 217864
rect 491444 217852 491450 217864
rect 492582 217852 492588 217864
rect 491444 217824 492588 217852
rect 491444 217812 491450 217824
rect 492582 217812 492588 217824
rect 492640 217852 492646 217864
rect 619910 217852 619916 217864
rect 492640 217824 619916 217852
rect 492640 217812 492646 217824
rect 619910 217812 619916 217824
rect 619968 217812 619974 217864
rect 508406 217744 508412 217796
rect 508464 217784 508470 217796
rect 575842 217784 575848 217796
rect 508464 217756 575848 217784
rect 508464 217744 508470 217756
rect 575842 217744 575848 217756
rect 575900 217744 575906 217796
rect 561766 217676 561772 217728
rect 561824 217716 561830 217728
rect 562870 217716 562876 217728
rect 561824 217688 562876 217716
rect 561824 217676 561830 217688
rect 562870 217676 562876 217688
rect 562928 217716 562934 217728
rect 634538 217716 634544 217728
rect 562928 217688 634544 217716
rect 562928 217676 562934 217688
rect 634538 217676 634544 217688
rect 634596 217676 634602 217728
rect 560294 217608 560300 217660
rect 560352 217648 560358 217660
rect 634078 217648 634084 217660
rect 560352 217620 634084 217648
rect 560352 217608 560358 217620
rect 634078 217608 634084 217620
rect 634136 217608 634142 217660
rect 557810 217540 557816 217592
rect 557868 217580 557874 217592
rect 633618 217580 633624 217592
rect 557868 217552 633624 217580
rect 557868 217540 557874 217552
rect 633618 217540 633624 217552
rect 633676 217540 633682 217592
rect 545206 217472 545212 217524
rect 545264 217512 545270 217524
rect 621014 217512 621020 217524
rect 545264 217484 621020 217512
rect 545264 217472 545270 217484
rect 621014 217472 621020 217484
rect 621072 217472 621078 217524
rect 555694 217404 555700 217456
rect 555752 217444 555758 217456
rect 633158 217444 633164 217456
rect 555752 217416 633164 217444
rect 555752 217404 555758 217416
rect 633158 217404 633164 217416
rect 633216 217404 633222 217456
rect 499574 217336 499580 217388
rect 499632 217376 499638 217388
rect 500862 217376 500868 217388
rect 499632 217348 500868 217376
rect 499632 217336 499638 217348
rect 500862 217336 500868 217348
rect 500920 217376 500926 217388
rect 576946 217376 576952 217388
rect 500920 217348 576952 217376
rect 500920 217336 500926 217348
rect 576946 217336 576952 217348
rect 577004 217336 577010 217388
rect 35618 217268 35624 217320
rect 35676 217308 35682 217320
rect 46290 217308 46296 217320
rect 35676 217280 46296 217308
rect 35676 217268 35682 217280
rect 46290 217268 46296 217280
rect 46348 217268 46354 217320
rect 52178 217268 52184 217320
rect 52236 217308 52242 217320
rect 164878 217308 164884 217320
rect 52236 217280 164884 217308
rect 52236 217268 52242 217280
rect 164878 217268 164884 217280
rect 164936 217268 164942 217320
rect 550542 217268 550548 217320
rect 550600 217308 550606 217320
rect 629202 217308 629208 217320
rect 550600 217280 629208 217308
rect 550600 217268 550606 217280
rect 629202 217268 629208 217280
rect 629260 217268 629266 217320
rect 497642 217200 497648 217252
rect 497700 217240 497706 217252
rect 575750 217240 575756 217252
rect 497700 217212 575756 217240
rect 497700 217200 497706 217212
rect 575750 217200 575756 217212
rect 575808 217200 575814 217252
rect 537846 217132 537852 217184
rect 537904 217172 537910 217184
rect 618990 217172 618996 217184
rect 537904 217144 618996 217172
rect 537904 217132 537910 217144
rect 618990 217132 618996 217144
rect 619048 217132 619054 217184
rect 532970 217064 532976 217116
rect 533028 217104 533034 217116
rect 618162 217104 618168 217116
rect 533028 217076 618168 217104
rect 533028 217064 533034 217076
rect 618162 217064 618168 217076
rect 618220 217064 618226 217116
rect 513650 216996 513656 217048
rect 513708 217036 513714 217048
rect 610802 217036 610808 217048
rect 513708 217008 610808 217036
rect 513708 216996 513714 217008
rect 610802 216996 610808 217008
rect 610860 216996 610866 217048
rect 506106 216928 506112 216980
rect 506164 216968 506170 216980
rect 607490 216968 607496 216980
rect 506164 216940 607496 216968
rect 506164 216928 506170 216940
rect 607490 216928 607496 216940
rect 607548 216928 607554 216980
rect 502518 216860 502524 216912
rect 502576 216900 502582 216912
rect 503530 216900 503536 216912
rect 502576 216872 503536 216900
rect 502576 216860 502582 216872
rect 503530 216860 503536 216872
rect 503588 216900 503594 216912
rect 608502 216900 608508 216912
rect 503588 216872 608508 216900
rect 503588 216860 503594 216872
rect 608502 216860 608508 216872
rect 608560 216860 608566 216912
rect 494330 216792 494336 216844
rect 494388 216832 494394 216844
rect 607582 216832 607588 216844
rect 494388 216804 607588 216832
rect 494388 216792 494394 216804
rect 607582 216792 607588 216804
rect 607640 216792 607646 216844
rect 499114 216724 499120 216776
rect 499172 216764 499178 216776
rect 622578 216764 622584 216776
rect 499172 216736 622584 216764
rect 499172 216724 499178 216736
rect 622578 216724 622584 216736
rect 622636 216724 622642 216776
rect 566642 216656 566648 216708
rect 566700 216696 566706 216708
rect 575658 216696 575664 216708
rect 566700 216668 575664 216696
rect 566700 216656 566706 216668
rect 575658 216656 575664 216668
rect 575716 216656 575722 216708
rect 553366 216464 556660 216492
rect 490926 216384 490932 216436
rect 490984 216424 490990 216436
rect 490984 216396 499574 216424
rect 490984 216384 490990 216396
rect 499546 215336 499574 216396
rect 521194 216384 521200 216436
rect 521252 216424 521258 216436
rect 521252 216396 523356 216424
rect 521252 216384 521258 216396
rect 523328 215404 523356 216396
rect 523770 216384 523776 216436
rect 523828 216424 523834 216436
rect 523828 216396 525104 216424
rect 523828 216384 523834 216396
rect 525076 215472 525104 216396
rect 526254 216384 526260 216436
rect 526312 216424 526318 216436
rect 526312 216396 526806 216424
rect 526312 216384 526318 216396
rect 526778 215540 526806 216396
rect 528554 216384 528560 216436
rect 528612 216424 528618 216436
rect 528612 216396 528692 216424
rect 528612 216384 528618 216396
rect 528664 215608 528692 216396
rect 531222 216384 531228 216436
rect 531280 216424 531286 216436
rect 531280 216396 533292 216424
rect 531280 216384 531286 216396
rect 533264 215676 533292 216396
rect 533798 216384 533804 216436
rect 533856 216424 533862 216436
rect 533856 216396 534856 216424
rect 533856 216384 533862 216396
rect 534828 215744 534856 216396
rect 536374 216384 536380 216436
rect 536432 216424 536438 216436
rect 536432 216396 538214 216424
rect 536432 216384 536438 216396
rect 538186 215812 538214 216396
rect 538858 216384 538864 216436
rect 538916 216424 538922 216436
rect 538916 216396 547874 216424
rect 538916 216384 538922 216396
rect 547846 215880 547874 216396
rect 548978 216384 548984 216436
rect 549036 216384 549042 216436
rect 548996 216356 549024 216384
rect 553366 216356 553394 216464
rect 556522 216384 556528 216436
rect 556580 216384 556586 216436
rect 548996 216328 553394 216356
rect 556540 216016 556568 216384
rect 556632 216084 556660 216464
rect 560266 216464 569954 216492
rect 560266 216084 560294 216464
rect 561582 216384 561588 216436
rect 561640 216424 561646 216436
rect 561640 216396 564204 216424
rect 561640 216384 561646 216396
rect 556632 216056 560294 216084
rect 564176 216016 564204 216396
rect 569926 216152 569954 216464
rect 615494 216452 615500 216504
rect 615552 216492 615558 216504
rect 631778 216492 631784 216504
rect 615552 216464 631784 216492
rect 615552 216452 615558 216464
rect 631778 216452 631784 216464
rect 631836 216452 631842 216504
rect 574186 216384 574192 216436
rect 574244 216424 574250 216436
rect 574244 216396 574324 216424
rect 574244 216384 574250 216396
rect 574296 216152 574324 216396
rect 574830 216384 574836 216436
rect 574888 216384 574894 216436
rect 613378 216384 613384 216436
rect 613436 216424 613442 216436
rect 630398 216424 630404 216436
rect 613436 216396 630404 216424
rect 613436 216384 613442 216396
rect 630398 216384 630404 216396
rect 630456 216384 630462 216436
rect 574848 216220 574876 216384
rect 611998 216316 612004 216368
rect 612056 216356 612062 216368
rect 628466 216356 628472 216368
rect 612056 216328 628472 216356
rect 612056 216316 612062 216328
rect 628466 216316 628472 216328
rect 628524 216316 628530 216368
rect 614114 216248 614120 216300
rect 614172 216288 614178 216300
rect 630858 216288 630864 216300
rect 614172 216260 630864 216288
rect 614172 216248 614178 216260
rect 630858 216248 630864 216260
rect 630916 216248 630922 216300
rect 626166 216220 626172 216232
rect 574848 216192 626172 216220
rect 626166 216180 626172 216192
rect 626224 216180 626230 216232
rect 628006 216152 628012 216164
rect 569926 216124 572714 216152
rect 574296 216124 628012 216152
rect 572686 216084 572714 216124
rect 628006 216112 628012 216124
rect 628064 216112 628070 216164
rect 674374 216112 674380 216164
rect 674432 216152 674438 216164
rect 676030 216152 676036 216164
rect 674432 216124 676036 216152
rect 674432 216112 674438 216124
rect 676030 216112 676036 216124
rect 676088 216112 676094 216164
rect 577866 216084 577872 216096
rect 572686 216056 577872 216084
rect 577866 216044 577872 216056
rect 577924 216044 577930 216096
rect 605926 216044 605932 216096
rect 605984 216084 605990 216096
rect 629478 216084 629484 216096
rect 605984 216056 629484 216084
rect 605984 216044 605990 216056
rect 629478 216044 629484 216056
rect 629536 216044 629542 216096
rect 619634 216016 619640 216028
rect 556540 215988 563054 216016
rect 564176 215988 619640 216016
rect 563026 215948 563054 215988
rect 619634 215976 619640 215988
rect 619692 215976 619698 216028
rect 618714 215948 618720 215960
rect 563026 215920 618720 215948
rect 618714 215908 618720 215920
rect 618772 215908 618778 215960
rect 676214 215908 676220 215960
rect 676272 215948 676278 215960
rect 676858 215948 676864 215960
rect 676272 215920 676864 215948
rect 676272 215908 676278 215920
rect 676858 215908 676864 215920
rect 676916 215908 676922 215960
rect 615494 215880 615500 215892
rect 547846 215852 615500 215880
rect 615494 215840 615500 215852
rect 615552 215840 615558 215892
rect 615034 215812 615040 215824
rect 538186 215784 615040 215812
rect 615034 215772 615040 215784
rect 615092 215772 615098 215824
rect 614574 215744 614580 215756
rect 534828 215716 614580 215744
rect 614574 215704 614580 215716
rect 614632 215704 614638 215756
rect 674466 215704 674472 215756
rect 674524 215744 674530 215756
rect 676030 215744 676036 215756
rect 674524 215716 676036 215744
rect 674524 215704 674530 215716
rect 676030 215704 676036 215716
rect 676088 215704 676094 215756
rect 614022 215676 614028 215688
rect 533264 215648 614028 215676
rect 614022 215636 614028 215648
rect 614080 215636 614086 215688
rect 613562 215608 613568 215620
rect 528664 215580 613568 215608
rect 613562 215568 613568 215580
rect 613620 215568 613626 215620
rect 613102 215540 613108 215552
rect 526778 215512 613108 215540
rect 613102 215500 613108 215512
rect 613160 215500 613166 215552
rect 612642 215472 612648 215484
rect 525076 215444 612648 215472
rect 612642 215432 612648 215444
rect 612700 215432 612706 215484
rect 612182 215404 612188 215416
rect 523328 215376 612188 215404
rect 612182 215364 612188 215376
rect 612240 215364 612246 215416
rect 607122 215336 607128 215348
rect 499546 215308 607128 215336
rect 607122 215296 607128 215308
rect 607180 215296 607186 215348
rect 577130 214820 577136 214872
rect 577188 214860 577194 214872
rect 627086 214860 627092 214872
rect 577188 214832 627092 214860
rect 577188 214820 577194 214832
rect 627086 214820 627092 214832
rect 627144 214820 627150 214872
rect 577222 214684 577228 214736
rect 577280 214724 577286 214736
rect 627546 214724 627552 214736
rect 577280 214696 627552 214724
rect 577280 214684 577286 214696
rect 627546 214684 627552 214696
rect 627604 214684 627610 214736
rect 576394 214616 576400 214668
rect 576452 214656 576458 214668
rect 626626 214656 626632 214668
rect 576452 214628 626632 214656
rect 576452 214616 576458 214628
rect 626626 214616 626632 214628
rect 626684 214616 626690 214668
rect 35802 214548 35808 214600
rect 35860 214588 35866 214600
rect 43622 214588 43628 214600
rect 35860 214560 43628 214588
rect 35860 214548 35866 214560
rect 43622 214548 43628 214560
rect 43680 214548 43686 214600
rect 577038 214548 577044 214600
rect 577096 214588 577102 214600
rect 634998 214588 635004 214600
rect 577096 214560 635004 214588
rect 577096 214548 577102 214560
rect 634998 214548 635004 214560
rect 635056 214548 635062 214600
rect 48958 214344 48964 214396
rect 49016 214384 49022 214396
rect 665266 214384 665272 214396
rect 49016 214356 665272 214384
rect 49016 214344 49022 214356
rect 665266 214344 665272 214356
rect 665324 214344 665330 214396
rect 46566 214276 46572 214328
rect 46624 214316 46630 214328
rect 668946 214316 668952 214328
rect 46624 214288 668952 214316
rect 46624 214276 46630 214288
rect 668946 214276 668952 214288
rect 669004 214276 669010 214328
rect 40862 214208 40868 214260
rect 40920 214248 40926 214260
rect 666186 214248 666192 214260
rect 40920 214220 666192 214248
rect 40920 214208 40926 214220
rect 666186 214208 666192 214220
rect 666244 214208 666250 214260
rect 42794 214140 42800 214192
rect 42852 214180 42858 214192
rect 668118 214180 668124 214192
rect 42852 214152 668124 214180
rect 42852 214140 42858 214152
rect 668118 214140 668124 214152
rect 668176 214140 668182 214192
rect 40678 214072 40684 214124
rect 40736 214112 40742 214124
rect 665726 214112 665732 214124
rect 40736 214084 665732 214112
rect 40736 214072 40742 214084
rect 665726 214072 665732 214084
rect 665784 214072 665790 214124
rect 673178 214072 673184 214124
rect 673236 214112 673242 214124
rect 676030 214112 676036 214124
rect 673236 214084 676036 214112
rect 673236 214072 673242 214084
rect 676030 214072 676036 214084
rect 676088 214072 676094 214124
rect 41782 214004 41788 214056
rect 41840 214044 41846 214056
rect 668854 214044 668860 214056
rect 41840 214016 668860 214044
rect 41840 214004 41846 214016
rect 668854 214004 668860 214016
rect 668912 214004 668918 214056
rect 41322 213936 41328 213988
rect 41380 213976 41386 213988
rect 668762 213976 668768 213988
rect 41380 213948 668768 213976
rect 41380 213936 41386 213948
rect 668762 213936 668768 213948
rect 668820 213936 668826 213988
rect 576946 213868 576952 213920
rect 577004 213908 577010 213920
rect 608502 213908 608508 213920
rect 577004 213880 608508 213908
rect 577004 213868 577010 213880
rect 608502 213868 608508 213880
rect 608560 213868 608566 213920
rect 636102 213868 636108 213920
rect 636160 213908 636166 213920
rect 637390 213908 637396 213920
rect 636160 213880 637396 213908
rect 636160 213868 636166 213880
rect 637390 213868 637396 213880
rect 637448 213868 637454 213920
rect 638218 213868 638224 213920
rect 638276 213908 638282 213920
rect 640610 213908 640616 213920
rect 638276 213880 640616 213908
rect 638276 213868 638282 213880
rect 640610 213868 640616 213880
rect 640668 213868 640674 213920
rect 575750 213800 575756 213852
rect 575808 213840 575814 213852
rect 608042 213840 608048 213852
rect 575808 213812 608048 213840
rect 575808 213800 575814 213812
rect 608042 213800 608048 213812
rect 608100 213800 608106 213852
rect 609606 213800 609612 213852
rect 609664 213840 609670 213852
rect 617794 213840 617800 213852
rect 609664 213812 617800 213840
rect 609664 213800 609670 213812
rect 617794 213800 617800 213812
rect 617852 213800 617858 213852
rect 619910 213800 619916 213852
rect 619968 213840 619974 213852
rect 622026 213840 622032 213852
rect 619968 213812 622032 213840
rect 619968 213800 619974 213812
rect 622026 213800 622032 213812
rect 622084 213800 622090 213852
rect 629938 213800 629944 213852
rect 629996 213840 630002 213852
rect 636562 213840 636568 213852
rect 629996 213812 636568 213840
rect 629996 213800 630002 213812
rect 636562 213800 636568 213812
rect 636620 213800 636626 213852
rect 636838 213800 636844 213852
rect 636896 213840 636902 213852
rect 639230 213840 639236 213852
rect 636896 213812 639236 213840
rect 636896 213800 636902 213812
rect 639230 213800 639236 213812
rect 639288 213800 639294 213852
rect 575842 213732 575848 213784
rect 575900 213772 575906 213784
rect 609882 213772 609888 213784
rect 575900 213744 609888 213772
rect 575900 213732 575906 213744
rect 609882 213732 609888 213744
rect 609940 213732 609946 213784
rect 610342 213732 610348 213784
rect 610400 213772 610406 213784
rect 621474 213772 621480 213784
rect 610400 213744 621480 213772
rect 610400 213732 610406 213744
rect 621474 213732 621480 213744
rect 621532 213732 621538 213784
rect 636010 213732 636016 213784
rect 636068 213772 636074 213784
rect 637850 213772 637856 213784
rect 636068 213744 637856 213772
rect 636068 213732 636074 213744
rect 637850 213732 637856 213744
rect 637908 213732 637914 213784
rect 575934 213664 575940 213716
rect 575992 213704 575998 213716
rect 611722 213704 611728 213716
rect 575992 213676 611728 213704
rect 575992 213664 575998 213676
rect 611722 213664 611728 213676
rect 611780 213664 611786 213716
rect 621014 213664 621020 213716
rect 621072 213704 621078 213716
rect 631318 213704 631324 213716
rect 621072 213676 631324 213704
rect 621072 213664 621078 213676
rect 631318 213664 631324 213676
rect 631376 213664 631382 213716
rect 674558 213664 674564 213716
rect 674616 213704 674622 213716
rect 676030 213704 676036 213716
rect 674616 213676 676036 213704
rect 674616 213664 674622 213676
rect 676030 213664 676036 213676
rect 676088 213664 676094 213716
rect 577866 213596 577872 213648
rect 577924 213636 577930 213648
rect 617334 213636 617340 213648
rect 577924 213608 617340 213636
rect 577924 213596 577930 213608
rect 617334 213596 617340 213608
rect 617392 213596 617398 213648
rect 618162 213596 618168 213648
rect 618220 213636 618226 213648
rect 628926 213636 628932 213648
rect 618220 213608 628932 213636
rect 618220 213596 618226 213608
rect 628926 213596 628932 213608
rect 628984 213596 628990 213648
rect 629202 213596 629208 213648
rect 629260 213636 629266 213648
rect 632238 213636 632244 213648
rect 629260 213608 632244 213636
rect 629260 213596 629266 213608
rect 632238 213596 632244 213608
rect 632296 213596 632302 213648
rect 576118 213528 576124 213580
rect 576176 213568 576182 213580
rect 615954 213568 615960 213580
rect 576176 213540 615960 213568
rect 576176 213528 576182 213540
rect 615954 213528 615960 213540
rect 616012 213528 616018 213580
rect 618990 213528 618996 213580
rect 619048 213568 619054 213580
rect 629938 213568 629944 213580
rect 619048 213540 629944 213568
rect 619048 213528 619054 213540
rect 629938 213528 629944 213540
rect 629996 213528 630002 213580
rect 576210 213460 576216 213512
rect 576268 213500 576274 213512
rect 616414 213500 616420 213512
rect 576268 213472 616420 213500
rect 576268 213460 576274 213472
rect 616414 213460 616420 213472
rect 616472 213460 616478 213512
rect 616782 213460 616788 213512
rect 616840 213500 616846 213512
rect 635458 213500 635464 213512
rect 616840 213472 635464 213500
rect 616840 213460 616846 213472
rect 635458 213460 635464 213472
rect 635516 213460 635522 213512
rect 576302 213392 576308 213444
rect 576360 213432 576366 213444
rect 616874 213432 616880 213444
rect 576360 213404 616880 213432
rect 576360 213392 576366 213404
rect 616874 213392 616880 213404
rect 616932 213392 616938 213444
rect 617518 213392 617524 213444
rect 617576 213432 617582 213444
rect 635918 213432 635924 213444
rect 617576 213404 635924 213432
rect 617576 213392 617582 213404
rect 635918 213392 635924 213404
rect 635976 213392 635982 213444
rect 576026 213324 576032 213376
rect 576084 213364 576090 213376
rect 618254 213364 618260 213376
rect 576084 213336 618260 213364
rect 576084 213324 576090 213336
rect 618254 213324 618260 213336
rect 618312 213324 618318 213376
rect 620278 213324 620284 213376
rect 620336 213364 620342 213376
rect 636378 213364 636384 213376
rect 620336 213336 636384 213364
rect 620336 213324 620342 213336
rect 636378 213324 636384 213336
rect 636436 213324 636442 213376
rect 575658 213256 575664 213308
rect 575716 213296 575722 213308
rect 620554 213296 620560 213308
rect 575716 213268 620560 213296
rect 575716 213256 575722 213268
rect 620554 213256 620560 213268
rect 620612 213256 620618 213308
rect 623038 213256 623044 213308
rect 623096 213296 623102 213308
rect 641070 213296 641076 213308
rect 623096 213268 641076 213296
rect 623096 213256 623102 213268
rect 641070 213256 641076 213268
rect 641128 213256 641134 213308
rect 642726 213256 642732 213308
rect 642784 213296 642790 213308
rect 649994 213296 650000 213308
rect 642784 213268 650000 213296
rect 642784 213256 642790 213268
rect 649994 213256 650000 213268
rect 650052 213256 650058 213308
rect 577498 213188 577504 213240
rect 577556 213228 577562 213240
rect 640150 213228 640156 213240
rect 577556 213200 640156 213228
rect 577556 213188 577562 213200
rect 640150 213188 640156 213200
rect 640208 213188 640214 213240
rect 643830 213188 643836 213240
rect 643888 213228 643894 213240
rect 651374 213228 651380 213240
rect 643888 213200 651380 213228
rect 643888 213188 643894 213200
rect 651374 213188 651380 213200
rect 651432 213188 651438 213240
rect 607490 213120 607496 213172
rect 607548 213160 607554 213172
rect 609422 213160 609428 213172
rect 607548 213132 609428 213160
rect 607548 213120 607554 213132
rect 609422 213120 609428 213132
rect 609480 213120 609486 213172
rect 608410 213052 608416 213104
rect 608468 213092 608474 213104
rect 611262 213092 611268 213104
rect 608468 213064 611268 213092
rect 608468 213052 608474 213064
rect 611262 213052 611268 213064
rect 611320 213052 611326 213104
rect 646958 212984 646964 213036
rect 647016 213024 647022 213036
rect 651466 213024 651472 213036
rect 647016 212996 651472 213024
rect 647016 212984 647022 212996
rect 651466 212984 651472 212996
rect 651524 212984 651530 213036
rect 645578 212576 645584 212628
rect 645636 212616 645642 212628
rect 650086 212616 650092 212628
rect 645636 212588 650092 212616
rect 645636 212576 645642 212588
rect 650086 212576 650092 212588
rect 650144 212576 650150 212628
rect 623774 212372 623780 212424
rect 623832 212412 623838 212424
rect 624418 212412 624424 212424
rect 623832 212384 624424 212412
rect 623832 212372 623838 212384
rect 624418 212372 624424 212384
rect 624476 212372 624482 212424
rect 625246 212372 625252 212424
rect 625304 212412 625310 212424
rect 625706 212412 625712 212424
rect 625304 212384 625712 212412
rect 625304 212372 625310 212384
rect 625706 212372 625712 212384
rect 625764 212372 625770 212424
rect 663794 212372 663800 212424
rect 663852 212412 663858 212424
rect 664438 212412 664444 212424
rect 663852 212384 664444 212412
rect 663852 212372 663858 212384
rect 664438 212372 664444 212384
rect 664496 212372 664502 212424
rect 663886 212304 663892 212356
rect 663944 212344 663950 212356
rect 664346 212344 664352 212356
rect 663944 212316 664352 212344
rect 663944 212304 663950 212316
rect 664346 212304 664352 212316
rect 664404 212304 664410 212356
rect 671430 211148 671436 211200
rect 671488 211188 671494 211200
rect 676030 211188 676036 211200
rect 671488 211160 676036 211188
rect 671488 211148 671494 211160
rect 676030 211148 676036 211160
rect 676088 211148 676094 211200
rect 662414 210536 662420 210588
rect 662472 210576 662478 210588
rect 663058 210576 663064 210588
rect 662472 210548 663064 210576
rect 662472 210536 662478 210548
rect 663058 210536 663064 210548
rect 663116 210536 663122 210588
rect 652018 210400 652024 210452
rect 652076 210440 652082 210452
rect 667198 210440 667204 210452
rect 652076 210412 667204 210440
rect 652076 210400 652082 210412
rect 667198 210400 667204 210412
rect 667256 210400 667262 210452
rect 580258 209788 580264 209840
rect 580316 209828 580322 209840
rect 638402 209828 638408 209840
rect 580316 209800 638408 209828
rect 580316 209788 580322 209800
rect 638402 209788 638408 209800
rect 638460 209788 638466 209840
rect 579062 209720 579068 209772
rect 579120 209760 579126 209772
rect 603166 209760 603172 209772
rect 579120 209732 603172 209760
rect 579120 209720 579126 209732
rect 603166 209720 603172 209732
rect 603224 209720 603230 209772
rect 578878 209652 578884 209704
rect 578936 209692 578942 209704
rect 603074 209692 603080 209704
rect 578936 209664 603080 209692
rect 578936 209652 578942 209664
rect 603074 209652 603080 209664
rect 603132 209652 603138 209704
rect 665450 209652 665456 209704
rect 665508 209692 665514 209704
rect 666922 209692 666928 209704
rect 665508 209664 666928 209692
rect 665508 209652 665514 209664
rect 666922 209652 666928 209664
rect 666980 209652 666986 209704
rect 578970 208292 578976 208344
rect 579028 208332 579034 208344
rect 603074 208332 603080 208344
rect 579028 208304 603080 208332
rect 579028 208292 579034 208304
rect 603074 208292 603080 208304
rect 603132 208292 603138 208344
rect 578418 206932 578424 206984
rect 578476 206972 578482 206984
rect 603074 206972 603080 206984
rect 578476 206944 603080 206972
rect 578476 206932 578482 206944
rect 603074 206932 603080 206944
rect 603132 206932 603138 206984
rect 578510 205572 578516 205624
rect 578568 205612 578574 205624
rect 603074 205612 603080 205624
rect 578568 205584 603080 205612
rect 578568 205572 578574 205584
rect 603074 205572 603080 205584
rect 603132 205572 603138 205624
rect 579522 205504 579528 205556
rect 579580 205544 579586 205556
rect 603166 205544 603172 205556
rect 579580 205516 603172 205544
rect 579580 205504 579586 205516
rect 603166 205504 603172 205516
rect 603224 205504 603230 205556
rect 578786 204212 578792 204264
rect 578844 204252 578850 204264
rect 603074 204252 603080 204264
rect 578844 204224 603080 204252
rect 578844 204212 578850 204224
rect 603074 204212 603080 204224
rect 603132 204212 603138 204264
rect 35802 202852 35808 202904
rect 35860 202892 35866 202904
rect 48958 202892 48964 202904
rect 35860 202864 48964 202892
rect 35860 202852 35866 202864
rect 48958 202852 48964 202864
rect 49016 202852 49022 202904
rect 579430 202784 579436 202836
rect 579488 202824 579494 202836
rect 603074 202824 603080 202836
rect 579488 202796 603080 202824
rect 579488 202784 579494 202796
rect 603074 202784 603080 202796
rect 603132 202784 603138 202836
rect 674374 201832 674380 201884
rect 674432 201872 674438 201884
rect 675386 201872 675392 201884
rect 674432 201844 675392 201872
rect 674432 201832 674438 201844
rect 675386 201832 675392 201844
rect 675444 201832 675450 201884
rect 579246 201424 579252 201476
rect 579304 201464 579310 201476
rect 603166 201464 603172 201476
rect 579304 201436 603172 201464
rect 579304 201424 579310 201436
rect 603166 201424 603172 201436
rect 603224 201424 603230 201476
rect 674466 201424 674472 201476
rect 674524 201464 674530 201476
rect 675386 201464 675392 201476
rect 674524 201436 675392 201464
rect 674524 201424 674530 201436
rect 675386 201424 675392 201436
rect 675444 201424 675450 201476
rect 578878 201356 578884 201408
rect 578936 201396 578942 201408
rect 603074 201396 603080 201408
rect 578936 201368 603080 201396
rect 578936 201356 578942 201368
rect 603074 201356 603080 201368
rect 603132 201356 603138 201408
rect 675110 200676 675116 200728
rect 675168 200716 675174 200728
rect 675386 200716 675392 200728
rect 675168 200688 675392 200716
rect 675168 200676 675174 200688
rect 675386 200676 675392 200688
rect 675444 200676 675450 200728
rect 578234 200064 578240 200116
rect 578292 200104 578298 200116
rect 603074 200104 603080 200116
rect 578292 200076 603080 200104
rect 578292 200064 578298 200076
rect 603074 200064 603080 200076
rect 603132 200064 603138 200116
rect 578418 198636 578424 198688
rect 578476 198676 578482 198688
rect 603074 198676 603080 198688
rect 578476 198648 603080 198676
rect 578476 198636 578482 198648
rect 603074 198636 603080 198648
rect 603132 198636 603138 198688
rect 673178 197412 673184 197464
rect 673236 197452 673242 197464
rect 675478 197452 675484 197464
rect 673236 197424 675484 197452
rect 673236 197412 673242 197424
rect 675478 197412 675484 197424
rect 675536 197412 675542 197464
rect 579062 197276 579068 197328
rect 579120 197316 579126 197328
rect 603166 197316 603172 197328
rect 579120 197288 603172 197316
rect 579120 197276 579126 197288
rect 603166 197276 603172 197288
rect 603224 197276 603230 197328
rect 674834 197004 674840 197056
rect 674892 197044 674898 197056
rect 675386 197044 675392 197056
rect 674892 197016 675392 197044
rect 674892 197004 674898 197016
rect 675386 197004 675392 197016
rect 675444 197004 675450 197056
rect 579522 196596 579528 196648
rect 579580 196636 579586 196648
rect 603074 196636 603080 196648
rect 579580 196608 603080 196636
rect 579580 196596 579586 196608
rect 603074 196596 603080 196608
rect 603132 196596 603138 196648
rect 674558 196528 674564 196580
rect 674616 196568 674622 196580
rect 675386 196568 675392 196580
rect 674616 196540 675392 196568
rect 674616 196528 674622 196540
rect 675386 196528 675392 196540
rect 675444 196528 675450 196580
rect 579522 195236 579528 195288
rect 579580 195276 579586 195288
rect 603074 195276 603080 195288
rect 579580 195248 603080 195276
rect 579580 195236 579586 195248
rect 603074 195236 603080 195248
rect 603132 195236 603138 195288
rect 579522 193808 579528 193860
rect 579580 193848 579586 193860
rect 603074 193848 603080 193860
rect 579580 193820 603080 193848
rect 579580 193808 579586 193820
rect 603074 193808 603080 193820
rect 603132 193808 603138 193860
rect 42058 193128 42064 193180
rect 42116 193168 42122 193180
rect 44450 193168 44456 193180
rect 42116 193140 44456 193168
rect 42116 193128 42122 193140
rect 44450 193128 44456 193140
rect 44508 193128 44514 193180
rect 579522 192448 579528 192500
rect 579580 192488 579586 192500
rect 603074 192488 603080 192500
rect 579580 192460 603080 192488
rect 579580 192448 579586 192460
rect 603074 192448 603080 192460
rect 603132 192448 603138 192500
rect 674834 192448 674840 192500
rect 674892 192488 674898 192500
rect 675386 192488 675392 192500
rect 674892 192460 675392 192488
rect 674892 192448 674898 192460
rect 675386 192448 675392 192460
rect 675444 192448 675450 192500
rect 579246 191836 579252 191888
rect 579304 191876 579310 191888
rect 603074 191876 603080 191888
rect 579304 191848 603080 191876
rect 579304 191836 579310 191848
rect 603074 191836 603080 191848
rect 603132 191836 603138 191888
rect 42058 191632 42064 191684
rect 42116 191672 42122 191684
rect 42978 191672 42984 191684
rect 42116 191644 42984 191672
rect 42116 191632 42122 191644
rect 42978 191632 42984 191644
rect 43036 191632 43042 191684
rect 42150 191564 42156 191616
rect 42208 191604 42214 191616
rect 44358 191604 44364 191616
rect 42208 191576 44364 191604
rect 42208 191564 42214 191576
rect 44358 191564 44364 191576
rect 44416 191564 44422 191616
rect 42150 190816 42156 190868
rect 42208 190856 42214 190868
rect 43070 190856 43076 190868
rect 42208 190828 43076 190856
rect 42208 190816 42214 190828
rect 43070 190816 43076 190828
rect 43128 190816 43134 190868
rect 675754 190612 675760 190664
rect 675812 190612 675818 190664
rect 578234 190476 578240 190528
rect 578292 190516 578298 190528
rect 603074 190516 603080 190528
rect 578292 190488 603080 190516
rect 578292 190476 578298 190488
rect 603074 190476 603080 190488
rect 603132 190476 603138 190528
rect 675772 190392 675800 190612
rect 675754 190340 675760 190392
rect 675812 190340 675818 190392
rect 579522 189116 579528 189168
rect 579580 189156 579586 189168
rect 603074 189156 603080 189168
rect 579580 189128 603080 189156
rect 579580 189116 579586 189128
rect 603074 189116 603080 189128
rect 603132 189116 603138 189168
rect 579246 189048 579252 189100
rect 579304 189088 579310 189100
rect 603166 189088 603172 189100
rect 579304 189060 603172 189088
rect 579304 189048 579310 189060
rect 603166 189048 603172 189060
rect 603224 189048 603230 189100
rect 578786 187688 578792 187740
rect 578844 187728 578850 187740
rect 603074 187728 603080 187740
rect 578844 187700 603080 187728
rect 578844 187688 578850 187700
rect 603074 187688 603080 187700
rect 603132 187688 603138 187740
rect 42150 187620 42156 187672
rect 42208 187660 42214 187672
rect 44266 187660 44272 187672
rect 42208 187632 44272 187660
rect 42208 187620 42214 187632
rect 44266 187620 44272 187632
rect 44324 187620 44330 187672
rect 579338 186328 579344 186380
rect 579396 186368 579402 186380
rect 603074 186368 603080 186380
rect 579396 186340 603080 186368
rect 579396 186328 579402 186340
rect 603074 186328 603080 186340
rect 603132 186328 603138 186380
rect 42058 186260 42064 186312
rect 42116 186300 42122 186312
rect 42886 186300 42892 186312
rect 42116 186272 42892 186300
rect 42116 186260 42122 186272
rect 42886 186260 42892 186272
rect 42944 186260 42950 186312
rect 42150 185852 42156 185904
rect 42208 185892 42214 185904
rect 42794 185892 42800 185904
rect 42208 185864 42800 185892
rect 42208 185852 42214 185864
rect 42794 185852 42800 185864
rect 42852 185852 42858 185904
rect 578970 184968 578976 185020
rect 579028 185008 579034 185020
rect 603074 185008 603080 185020
rect 579028 184980 603080 185008
rect 579028 184968 579034 184980
rect 603074 184968 603080 184980
rect 603132 184968 603138 185020
rect 579062 184900 579068 184952
rect 579120 184940 579126 184952
rect 603166 184940 603172 184952
rect 579120 184912 603172 184940
rect 579120 184900 579126 184912
rect 603166 184900 603172 184912
rect 603224 184900 603230 184952
rect 668302 184152 668308 184204
rect 668360 184192 668366 184204
rect 671338 184192 671344 184204
rect 668360 184164 671344 184192
rect 668360 184152 668366 184164
rect 671338 184152 671344 184164
rect 671396 184152 671402 184204
rect 579246 183540 579252 183592
rect 579304 183580 579310 183592
rect 603074 183580 603080 183592
rect 579304 183552 603080 183580
rect 579304 183540 579310 183552
rect 603074 183540 603080 183552
rect 603132 183540 603138 183592
rect 42150 183404 42156 183456
rect 42208 183444 42214 183456
rect 44174 183444 44180 183456
rect 42208 183416 44180 183444
rect 42208 183404 42214 183416
rect 44174 183404 44180 183416
rect 44232 183404 44238 183456
rect 578234 182180 578240 182232
rect 578292 182220 578298 182232
rect 603074 182220 603080 182232
rect 578292 182192 603080 182220
rect 578292 182180 578298 182192
rect 603074 182180 603080 182192
rect 603132 182180 603138 182232
rect 578326 180888 578332 180940
rect 578384 180928 578390 180940
rect 603166 180928 603172 180940
rect 578384 180900 603172 180928
rect 578384 180888 578390 180900
rect 603166 180888 603172 180900
rect 603224 180888 603230 180940
rect 578418 180820 578424 180872
rect 578476 180860 578482 180872
rect 603074 180860 603080 180872
rect 578476 180832 603080 180860
rect 578476 180820 578482 180832
rect 603074 180820 603080 180832
rect 603132 180820 603138 180872
rect 578786 179392 578792 179444
rect 578844 179432 578850 179444
rect 603074 179432 603080 179444
rect 578844 179404 603080 179432
rect 578844 179392 578850 179404
rect 603074 179392 603080 179404
rect 603132 179392 603138 179444
rect 667934 178780 667940 178832
rect 667992 178820 667998 178832
rect 670050 178820 670056 178832
rect 667992 178792 670056 178820
rect 667992 178780 667998 178792
rect 670050 178780 670056 178792
rect 670108 178780 670114 178832
rect 672994 178168 673000 178220
rect 673052 178208 673058 178220
rect 676030 178208 676036 178220
rect 673052 178180 676036 178208
rect 673052 178168 673058 178180
rect 676030 178168 676036 178180
rect 676088 178168 676094 178220
rect 578694 178032 578700 178084
rect 578752 178072 578758 178084
rect 603074 178072 603080 178084
rect 578752 178044 603080 178072
rect 578752 178032 578758 178044
rect 603074 178032 603080 178044
rect 603132 178032 603138 178084
rect 674098 178032 674104 178084
rect 674156 178072 674162 178084
rect 676030 178072 676036 178084
rect 674156 178044 676036 178072
rect 674156 178032 674162 178044
rect 676030 178032 676036 178044
rect 676088 178032 676094 178084
rect 672626 176944 672632 176996
rect 672684 176984 672690 176996
rect 676030 176984 676036 176996
rect 672684 176956 676036 176984
rect 672684 176944 672690 176956
rect 676030 176944 676036 176956
rect 676088 176944 676094 176996
rect 671614 176808 671620 176860
rect 671672 176848 671678 176860
rect 675938 176848 675944 176860
rect 671672 176820 675944 176848
rect 671672 176808 671678 176820
rect 675938 176808 675944 176820
rect 675996 176808 676002 176860
rect 579430 176740 579436 176792
rect 579488 176780 579494 176792
rect 603166 176780 603172 176792
rect 579488 176752 603172 176780
rect 579488 176740 579494 176752
rect 603166 176740 603172 176752
rect 603224 176740 603230 176792
rect 674006 176740 674012 176792
rect 674064 176780 674070 176792
rect 676030 176780 676036 176792
rect 674064 176752 676036 176780
rect 674064 176740 674070 176752
rect 676030 176740 676036 176752
rect 676088 176740 676094 176792
rect 579246 176672 579252 176724
rect 579304 176712 579310 176724
rect 603074 176712 603080 176724
rect 579304 176684 603080 176712
rect 579304 176672 579310 176684
rect 603074 176672 603080 176684
rect 603132 176672 603138 176724
rect 672534 176468 672540 176520
rect 672592 176508 672598 176520
rect 676030 176508 676036 176520
rect 672592 176480 676036 176508
rect 672592 176468 672598 176480
rect 676030 176468 676036 176480
rect 676088 176468 676094 176520
rect 674558 175992 674564 176044
rect 674616 176032 674622 176044
rect 676030 176032 676036 176044
rect 674616 176004 676036 176032
rect 674616 175992 674622 176004
rect 676030 175992 676036 176004
rect 676088 175992 676094 176044
rect 674650 175652 674656 175704
rect 674708 175692 674714 175704
rect 676030 175692 676036 175704
rect 674708 175664 676036 175692
rect 674708 175652 674714 175664
rect 676030 175652 676036 175664
rect 676088 175652 676094 175704
rect 581638 175244 581644 175296
rect 581696 175284 581702 175296
rect 603074 175284 603080 175296
rect 581696 175256 603080 175284
rect 581696 175244 581702 175256
rect 603074 175244 603080 175256
rect 603132 175244 603138 175296
rect 674558 175176 674564 175228
rect 674616 175216 674622 175228
rect 676030 175216 676036 175228
rect 674616 175188 676036 175216
rect 674616 175176 674622 175188
rect 676030 175176 676036 175188
rect 676088 175176 676094 175228
rect 673362 174360 673368 174412
rect 673420 174400 673426 174412
rect 676030 174400 676036 174412
rect 673420 174372 676036 174400
rect 673420 174360 673426 174372
rect 676030 174360 676036 174372
rect 676088 174360 676094 174412
rect 580350 173884 580356 173936
rect 580408 173924 580414 173936
rect 603074 173924 603080 173936
rect 580408 173896 603080 173924
rect 580408 173884 580414 173896
rect 603074 173884 603080 173896
rect 603132 173884 603138 173936
rect 667934 173612 667940 173664
rect 667992 173652 667998 173664
rect 670142 173652 670148 173664
rect 667992 173624 670148 173652
rect 667992 173612 667998 173624
rect 670142 173612 670148 173624
rect 670200 173612 670206 173664
rect 579154 172524 579160 172576
rect 579212 172564 579218 172576
rect 603074 172564 603080 172576
rect 579212 172536 603080 172564
rect 579212 172524 579218 172536
rect 603074 172524 603080 172536
rect 603132 172524 603138 172576
rect 674834 172524 674840 172576
rect 674892 172564 674898 172576
rect 676030 172564 676036 172576
rect 674892 172536 676036 172564
rect 674892 172524 674898 172536
rect 676030 172524 676036 172536
rect 676088 172524 676094 172576
rect 579338 171096 579344 171148
rect 579396 171136 579402 171148
rect 603074 171136 603080 171148
rect 579396 171108 603080 171136
rect 579396 171096 579402 171108
rect 603074 171096 603080 171108
rect 603132 171096 603138 171148
rect 674466 170280 674472 170332
rect 674524 170320 674530 170332
rect 676030 170320 676036 170332
rect 674524 170292 676036 170320
rect 674524 170280 674530 170292
rect 676030 170280 676036 170292
rect 676088 170280 676094 170332
rect 578970 169804 578976 169856
rect 579028 169844 579034 169856
rect 603074 169844 603080 169856
rect 579028 169816 603080 169844
rect 579028 169804 579034 169816
rect 603074 169804 603080 169816
rect 603132 169804 603138 169856
rect 579062 169736 579068 169788
rect 579120 169776 579126 169788
rect 603166 169776 603172 169788
rect 579120 169748 603172 169776
rect 579120 169736 579126 169748
rect 603166 169736 603172 169748
rect 603224 169736 603230 169788
rect 673178 169464 673184 169516
rect 673236 169504 673242 169516
rect 676030 169504 676036 169516
rect 673236 169476 676036 169504
rect 673236 169464 673242 169476
rect 676030 169464 676036 169476
rect 676088 169464 676094 169516
rect 674374 169056 674380 169108
rect 674432 169096 674438 169108
rect 676030 169096 676036 169108
rect 674432 169068 676036 169096
rect 674432 169056 674438 169068
rect 676030 169056 676036 169068
rect 676088 169056 676094 169108
rect 673270 168648 673276 168700
rect 673328 168688 673334 168700
rect 676030 168688 676036 168700
rect 673328 168660 676036 168688
rect 673328 168648 673334 168660
rect 676030 168648 676036 168660
rect 676088 168648 676094 168700
rect 578878 168376 578884 168428
rect 578936 168416 578942 168428
rect 603074 168416 603080 168428
rect 578936 168388 603080 168416
rect 578936 168376 578942 168388
rect 603074 168376 603080 168388
rect 603132 168376 603138 168428
rect 674098 168240 674104 168292
rect 674156 168280 674162 168292
rect 676030 168280 676036 168292
rect 674156 168252 676036 168280
rect 674156 168240 674162 168252
rect 676030 168240 676036 168252
rect 676088 168240 676094 168292
rect 672994 167832 673000 167884
rect 673052 167872 673058 167884
rect 676030 167872 676036 167884
rect 673052 167844 676036 167872
rect 673052 167832 673058 167844
rect 676030 167832 676036 167844
rect 676088 167832 676094 167884
rect 583110 167016 583116 167068
rect 583168 167056 583174 167068
rect 603074 167056 603080 167068
rect 583168 167028 603080 167056
rect 583168 167016 583174 167028
rect 603074 167016 603080 167028
rect 603132 167016 603138 167068
rect 671338 167016 671344 167068
rect 671396 167056 671402 167068
rect 676030 167056 676036 167068
rect 671396 167028 676036 167056
rect 671396 167016 671402 167028
rect 676030 167016 676036 167028
rect 676088 167016 676094 167068
rect 578694 166676 578700 166728
rect 578752 166716 578758 166728
rect 581638 166716 581644 166728
rect 578752 166688 581644 166716
rect 578752 166676 578758 166688
rect 581638 166676 581644 166688
rect 581696 166676 581702 166728
rect 581730 165588 581736 165640
rect 581788 165628 581794 165640
rect 603074 165628 603080 165640
rect 581788 165600 603080 165628
rect 581788 165588 581794 165600
rect 603074 165588 603080 165600
rect 603132 165588 603138 165640
rect 578234 164568 578240 164620
rect 578292 164608 578298 164620
rect 580350 164608 580356 164620
rect 578292 164580 580356 164608
rect 578292 164568 578298 164580
rect 580350 164568 580356 164580
rect 580408 164568 580414 164620
rect 581638 164228 581644 164280
rect 581696 164268 581702 164280
rect 603074 164268 603080 164280
rect 581696 164240 603080 164268
rect 581696 164228 581702 164240
rect 603074 164228 603080 164240
rect 603132 164228 603138 164280
rect 579522 164160 579528 164212
rect 579580 164200 579586 164212
rect 603718 164200 603724 164212
rect 579580 164172 603724 164200
rect 579580 164160 579586 164172
rect 603718 164160 603724 164172
rect 603776 164160 603782 164212
rect 668394 163956 668400 164008
rect 668452 163996 668458 164008
rect 672718 163996 672724 164008
rect 668452 163968 672724 163996
rect 668452 163956 668458 163968
rect 672718 163956 672724 163968
rect 672776 163956 672782 164008
rect 580350 162868 580356 162920
rect 580408 162908 580414 162920
rect 603074 162908 603080 162920
rect 580408 162880 603080 162908
rect 580408 162868 580414 162880
rect 603074 162868 603080 162880
rect 603132 162868 603138 162920
rect 583018 161440 583024 161492
rect 583076 161480 583082 161492
rect 603074 161480 603080 161492
rect 583076 161452 603080 161480
rect 583076 161440 583082 161452
rect 603074 161440 603080 161452
rect 603132 161440 603138 161492
rect 674834 160760 674840 160812
rect 674892 160800 674898 160812
rect 675478 160800 675484 160812
rect 674892 160772 675484 160800
rect 674892 160760 674898 160772
rect 675478 160760 675484 160772
rect 675536 160760 675542 160812
rect 579430 160080 579436 160132
rect 579488 160120 579494 160132
rect 603074 160120 603080 160132
rect 579488 160092 603080 160120
rect 579488 160080 579494 160092
rect 603074 160080 603080 160092
rect 603132 160080 603138 160132
rect 579338 158720 579344 158772
rect 579396 158760 579402 158772
rect 603074 158760 603080 158772
rect 579396 158732 603080 158760
rect 579396 158720 579402 158732
rect 603074 158720 603080 158732
rect 603132 158720 603138 158772
rect 585870 157428 585876 157480
rect 585928 157468 585934 157480
rect 603074 157468 603080 157480
rect 585928 157440 603080 157468
rect 585928 157428 585934 157440
rect 603074 157428 603080 157440
rect 603132 157428 603138 157480
rect 584398 157360 584404 157412
rect 584456 157400 584462 157412
rect 603166 157400 603172 157412
rect 584456 157372 603172 157400
rect 584456 157360 584462 157372
rect 603166 157360 603172 157372
rect 603224 157360 603230 157412
rect 587250 155932 587256 155984
rect 587308 155972 587314 155984
rect 603074 155972 603080 155984
rect 587308 155944 603080 155972
rect 587308 155932 587314 155944
rect 603074 155932 603080 155944
rect 603132 155932 603138 155984
rect 673178 155456 673184 155508
rect 673236 155496 673242 155508
rect 675478 155496 675484 155508
rect 673236 155468 675484 155496
rect 673236 155456 673242 155468
rect 675478 155456 675484 155468
rect 675536 155456 675542 155508
rect 578510 154640 578516 154692
rect 578568 154680 578574 154692
rect 583110 154680 583116 154692
rect 578568 154652 583116 154680
rect 578568 154640 578574 154652
rect 583110 154640 583116 154652
rect 583168 154640 583174 154692
rect 579154 154572 579160 154624
rect 579212 154612 579218 154624
rect 603074 154612 603080 154624
rect 579212 154584 603080 154612
rect 579212 154572 579218 154584
rect 603074 154572 603080 154584
rect 603132 154572 603138 154624
rect 579062 153280 579068 153332
rect 579120 153320 579126 153332
rect 603166 153320 603172 153332
rect 579120 153292 603172 153320
rect 579120 153280 579126 153292
rect 603166 153280 603172 153292
rect 603224 153280 603230 153332
rect 578970 153212 578976 153264
rect 579028 153252 579034 153264
rect 603074 153252 603080 153264
rect 579028 153224 603080 153252
rect 579028 153212 579034 153224
rect 603074 153212 603080 153224
rect 603132 153212 603138 153264
rect 579246 153076 579252 153128
rect 579304 153116 579310 153128
rect 581730 153116 581736 153128
rect 579304 153088 581736 153116
rect 579304 153076 579310 153088
rect 581730 153076 581736 153088
rect 581788 153076 581794 153128
rect 579246 152940 579252 152992
rect 579304 152980 579310 152992
rect 579430 152980 579436 152992
rect 579304 152952 579436 152980
rect 579304 152940 579310 152952
rect 579430 152940 579436 152952
rect 579488 152940 579494 152992
rect 674374 152532 674380 152584
rect 674432 152572 674438 152584
rect 675386 152572 675392 152584
rect 674432 152544 675392 152572
rect 674432 152532 674438 152544
rect 675386 152532 675392 152544
rect 675444 152532 675450 152584
rect 587158 151784 587164 151836
rect 587216 151824 587222 151836
rect 603074 151824 603080 151836
rect 587216 151796 603080 151824
rect 587216 151784 587222 151796
rect 603074 151784 603080 151796
rect 603132 151784 603138 151836
rect 579522 151716 579528 151768
rect 579580 151756 579586 151768
rect 603810 151756 603816 151768
rect 579580 151728 603816 151756
rect 579580 151716 579586 151728
rect 603810 151716 603816 151728
rect 603868 151716 603874 151768
rect 673270 151376 673276 151428
rect 673328 151416 673334 151428
rect 675386 151416 675392 151428
rect 673328 151388 675392 151416
rect 673328 151376 673334 151388
rect 675386 151376 675392 151388
rect 675444 151376 675450 151428
rect 578878 150424 578884 150476
rect 578936 150464 578942 150476
rect 603074 150464 603080 150476
rect 578936 150436 603080 150464
rect 578936 150424 578942 150436
rect 603074 150424 603080 150436
rect 603132 150424 603138 150476
rect 674466 150356 674472 150408
rect 674524 150396 674530 150408
rect 675386 150396 675392 150408
rect 674524 150368 675392 150396
rect 674524 150356 674530 150368
rect 675386 150356 675392 150368
rect 675444 150356 675450 150408
rect 579430 150220 579436 150272
rect 579488 150260 579494 150272
rect 581638 150260 581644 150272
rect 579488 150232 581644 150260
rect 579488 150220 579494 150232
rect 581638 150220 581644 150232
rect 581696 150220 581702 150272
rect 592770 149132 592776 149184
rect 592828 149172 592834 149184
rect 603074 149172 603080 149184
rect 592828 149144 603080 149172
rect 592828 149132 592834 149144
rect 603074 149132 603080 149144
rect 603132 149132 603138 149184
rect 589918 149064 589924 149116
rect 589976 149104 589982 149116
rect 603166 149104 603172 149116
rect 589976 149076 603172 149104
rect 589976 149064 589982 149076
rect 603166 149064 603172 149076
rect 603224 149064 603230 149116
rect 578510 148656 578516 148708
rect 578568 148696 578574 148708
rect 580350 148696 580356 148708
rect 578568 148668 580356 148696
rect 578568 148656 578574 148668
rect 580350 148656 580356 148668
rect 580408 148656 580414 148708
rect 668302 148520 668308 148572
rect 668360 148560 668366 148572
rect 674190 148560 674196 148572
rect 668360 148532 674196 148560
rect 668360 148520 668366 148532
rect 674190 148520 674196 148532
rect 674248 148520 674254 148572
rect 584582 147636 584588 147688
rect 584640 147676 584646 147688
rect 603074 147676 603080 147688
rect 584640 147648 603080 147676
rect 584640 147636 584646 147648
rect 603074 147636 603080 147648
rect 603132 147636 603138 147688
rect 578510 147296 578516 147348
rect 578568 147336 578574 147348
rect 580258 147336 580264 147348
rect 578568 147308 580264 147336
rect 578568 147296 578574 147308
rect 580258 147296 580264 147308
rect 580316 147296 580322 147348
rect 588538 146276 588544 146328
rect 588596 146316 588602 146328
rect 603074 146316 603080 146328
rect 588596 146288 603080 146316
rect 588596 146276 588602 146288
rect 603074 146276 603080 146288
rect 603132 146276 603138 146328
rect 579522 146072 579528 146124
rect 579580 146112 579586 146124
rect 583018 146112 583024 146124
rect 579580 146084 583024 146112
rect 579580 146072 579586 146084
rect 583018 146072 583024 146084
rect 583076 146072 583082 146124
rect 583110 144916 583116 144968
rect 583168 144956 583174 144968
rect 603166 144956 603172 144968
rect 583168 144928 603172 144956
rect 583168 144916 583174 144928
rect 603166 144916 603172 144928
rect 603224 144916 603230 144968
rect 578602 144848 578608 144900
rect 578660 144888 578666 144900
rect 603718 144888 603724 144900
rect 578660 144860 603724 144888
rect 578660 144848 578666 144860
rect 603718 144848 603724 144860
rect 603776 144848 603782 144900
rect 580350 143556 580356 143608
rect 580408 143596 580414 143608
rect 603074 143596 603080 143608
rect 580408 143568 603080 143596
rect 580408 143556 580414 143568
rect 603074 143556 603080 143568
rect 603132 143556 603138 143608
rect 667934 143284 667940 143336
rect 667992 143324 667998 143336
rect 670234 143324 670240 143336
rect 667992 143296 670240 143324
rect 667992 143284 667998 143296
rect 670234 143284 670240 143296
rect 670292 143284 670298 143336
rect 579522 142604 579528 142656
rect 579580 142644 579586 142656
rect 584398 142644 584404 142656
rect 579580 142616 584404 142644
rect 579580 142604 579586 142616
rect 584398 142604 584404 142616
rect 584456 142604 584462 142656
rect 585778 142128 585784 142180
rect 585836 142168 585842 142180
rect 603074 142168 603080 142180
rect 585836 142140 603080 142168
rect 585836 142128 585842 142140
rect 603074 142128 603080 142140
rect 603132 142128 603138 142180
rect 591298 140768 591304 140820
rect 591356 140808 591362 140820
rect 603074 140808 603080 140820
rect 591356 140780 603080 140808
rect 591356 140768 591362 140780
rect 603074 140768 603080 140780
rect 603132 140768 603138 140820
rect 584398 139408 584404 139460
rect 584456 139448 584462 139460
rect 603074 139448 603080 139460
rect 584456 139420 603080 139448
rect 584456 139408 584462 139420
rect 603074 139408 603080 139420
rect 603132 139408 603138 139460
rect 668026 138184 668032 138236
rect 668084 138224 668090 138236
rect 672810 138224 672816 138236
rect 668084 138196 672816 138224
rect 668084 138184 668090 138196
rect 672810 138184 672816 138196
rect 672868 138184 672874 138236
rect 598290 138048 598296 138100
rect 598348 138088 598354 138100
rect 603166 138088 603172 138100
rect 598348 138060 603172 138088
rect 598348 138048 598354 138060
rect 603166 138048 603172 138060
rect 603224 138048 603230 138100
rect 583018 137980 583024 138032
rect 583076 138020 583082 138032
rect 603074 138020 603080 138032
rect 583076 137992 603080 138020
rect 583076 137980 583082 137992
rect 603074 137980 603080 137992
rect 603132 137980 603138 138032
rect 579522 137912 579528 137964
rect 579580 137952 579586 137964
rect 587250 137952 587256 137964
rect 579580 137924 587256 137952
rect 579580 137912 579586 137924
rect 587250 137912 587256 137924
rect 587308 137912 587314 137964
rect 581638 136620 581644 136672
rect 581696 136660 581702 136672
rect 603074 136660 603080 136672
rect 581696 136632 603080 136660
rect 581696 136620 581702 136632
rect 603074 136620 603080 136632
rect 603132 136620 603138 136672
rect 579522 136484 579528 136536
rect 579580 136524 579586 136536
rect 585870 136524 585876 136536
rect 579580 136496 585876 136524
rect 579580 136484 579586 136496
rect 585870 136484 585876 136496
rect 585928 136484 585934 136536
rect 587342 135260 587348 135312
rect 587400 135300 587406 135312
rect 603074 135300 603080 135312
rect 587400 135272 603080 135300
rect 587400 135260 587406 135272
rect 603074 135260 603080 135272
rect 603132 135260 603138 135312
rect 580258 133900 580264 133952
rect 580316 133940 580322 133952
rect 603074 133940 603080 133952
rect 580316 133912 603080 133940
rect 580316 133900 580322 133912
rect 603074 133900 603080 133912
rect 603132 133900 603138 133952
rect 668578 132948 668584 133000
rect 668636 132988 668642 133000
rect 674282 132988 674288 133000
rect 668636 132960 674288 132988
rect 668636 132948 668642 132960
rect 674282 132948 674288 132960
rect 674340 132948 674346 133000
rect 672902 132880 672908 132932
rect 672960 132920 672966 132932
rect 676030 132920 676036 132932
rect 672960 132892 676036 132920
rect 672960 132880 672966 132892
rect 676030 132880 676036 132892
rect 676088 132880 676094 132932
rect 671522 132744 671528 132796
rect 671580 132784 671586 132796
rect 676214 132784 676220 132796
rect 671580 132756 676220 132784
rect 671580 132744 671586 132756
rect 676214 132744 676220 132756
rect 676272 132744 676278 132796
rect 667198 132608 667204 132660
rect 667256 132648 667262 132660
rect 676122 132648 676128 132660
rect 667256 132620 676128 132648
rect 667256 132608 667262 132620
rect 676122 132608 676128 132620
rect 676180 132608 676186 132660
rect 590010 132472 590016 132524
rect 590068 132512 590074 132524
rect 603074 132512 603080 132524
rect 590068 132484 603080 132512
rect 590068 132472 590074 132484
rect 603074 132472 603080 132484
rect 603132 132472 603138 132524
rect 674006 132268 674012 132320
rect 674064 132308 674070 132320
rect 676214 132308 676220 132320
rect 674064 132280 676220 132308
rect 674064 132268 674070 132280
rect 676214 132268 676220 132280
rect 676272 132268 676278 132320
rect 588630 131724 588636 131776
rect 588688 131764 588694 131776
rect 603166 131764 603172 131776
rect 588688 131736 603172 131764
rect 588688 131724 588694 131736
rect 603166 131724 603172 131736
rect 603224 131724 603230 131776
rect 674650 131316 674656 131368
rect 674708 131356 674714 131368
rect 676030 131356 676036 131368
rect 674708 131328 676036 131356
rect 674708 131316 674714 131328
rect 676030 131316 676036 131328
rect 676088 131316 676094 131368
rect 596910 131112 596916 131164
rect 596968 131152 596974 131164
rect 603074 131152 603080 131164
rect 596968 131124 603080 131152
rect 596968 131112 596974 131124
rect 603074 131112 603080 131124
rect 603132 131112 603138 131164
rect 668670 131112 668676 131164
rect 668728 131152 668734 131164
rect 668946 131152 668952 131164
rect 668728 131124 668952 131152
rect 668728 131112 668734 131124
rect 668946 131112 668952 131124
rect 669004 131152 669010 131164
rect 676214 131152 676220 131164
rect 669004 131124 676220 131152
rect 669004 131112 669010 131124
rect 676214 131112 676220 131124
rect 676272 131112 676278 131164
rect 579246 131044 579252 131096
rect 579304 131084 579310 131096
rect 587158 131084 587164 131096
rect 579304 131056 587164 131084
rect 579304 131044 579310 131056
rect 587158 131044 587164 131056
rect 587216 131044 587222 131096
rect 674558 130500 674564 130552
rect 674616 130540 674622 130552
rect 676030 130540 676036 130552
rect 674616 130512 676036 130540
rect 674616 130500 674622 130512
rect 676030 130500 676036 130512
rect 676088 130500 676094 130552
rect 672718 129888 672724 129940
rect 672776 129928 672782 129940
rect 676214 129928 676220 129940
rect 672776 129900 676220 129928
rect 672776 129888 672782 129900
rect 676214 129888 676220 129900
rect 676272 129888 676278 129940
rect 585870 129752 585876 129804
rect 585928 129792 585934 129804
rect 603074 129792 603080 129804
rect 585928 129764 603080 129792
rect 585928 129752 585934 129764
rect 603074 129752 603080 129764
rect 603132 129752 603138 129804
rect 668578 129752 668584 129804
rect 668636 129792 668642 129804
rect 668854 129792 668860 129804
rect 668636 129764 668860 129792
rect 668636 129752 668642 129764
rect 668854 129752 668860 129764
rect 668912 129792 668918 129804
rect 676214 129792 676220 129804
rect 668912 129764 676220 129792
rect 668912 129752 668918 129764
rect 676214 129752 676220 129764
rect 676272 129752 676278 129804
rect 581730 129004 581736 129056
rect 581788 129044 581794 129056
rect 603902 129044 603908 129056
rect 581788 129016 603908 129044
rect 581788 129004 581794 129016
rect 603902 129004 603908 129016
rect 603960 129004 603966 129056
rect 673362 128528 673368 128580
rect 673420 128568 673426 128580
rect 676122 128568 676128 128580
rect 673420 128540 676128 128568
rect 673420 128528 673426 128540
rect 676122 128528 676128 128540
rect 676180 128528 676186 128580
rect 594058 128324 594064 128376
rect 594116 128364 594122 128376
rect 603074 128364 603080 128376
rect 594116 128336 603080 128364
rect 594116 128324 594122 128336
rect 603074 128324 603080 128336
rect 603132 128324 603138 128376
rect 668762 128324 668768 128376
rect 668820 128364 668826 128376
rect 676214 128364 676220 128376
rect 668820 128336 676220 128364
rect 668820 128324 668826 128336
rect 676214 128324 676220 128336
rect 676272 128324 676278 128376
rect 578878 128256 578884 128308
rect 578936 128296 578942 128308
rect 584582 128296 584588 128308
rect 578936 128268 584588 128296
rect 578936 128256 578942 128268
rect 584582 128256 584588 128268
rect 584640 128256 584646 128308
rect 668026 128120 668032 128172
rect 668084 128160 668090 128172
rect 673086 128160 673092 128172
rect 668084 128132 673092 128160
rect 668084 128120 668090 128132
rect 673086 128120 673092 128132
rect 673144 128120 673150 128172
rect 584490 126964 584496 127016
rect 584548 127004 584554 127016
rect 603074 127004 603080 127016
rect 584548 126976 603080 127004
rect 584548 126964 584554 126976
rect 603074 126964 603080 126976
rect 603132 126964 603138 127016
rect 675110 126964 675116 127016
rect 675168 127004 675174 127016
rect 676030 127004 676036 127016
rect 675168 126976 676036 127004
rect 675168 126964 675174 126976
rect 676030 126964 676036 126976
rect 676088 126964 676094 127016
rect 579062 126896 579068 126948
rect 579120 126936 579126 126948
rect 592770 126936 592776 126948
rect 579120 126908 592776 126936
rect 579120 126896 579126 126908
rect 592770 126896 592776 126908
rect 592828 126896 592834 126948
rect 601050 125672 601056 125724
rect 601108 125712 601114 125724
rect 603074 125712 603080 125724
rect 601108 125684 603080 125712
rect 601108 125672 601114 125684
rect 603074 125672 603080 125684
rect 603132 125672 603138 125724
rect 592678 125604 592684 125656
rect 592736 125644 592742 125656
rect 603166 125644 603172 125656
rect 592736 125616 603172 125644
rect 592736 125604 592742 125616
rect 603166 125604 603172 125616
rect 603224 125604 603230 125656
rect 578418 125536 578424 125588
rect 578476 125576 578482 125588
rect 589918 125576 589924 125588
rect 578476 125548 589924 125576
rect 578476 125536 578482 125548
rect 589918 125536 589924 125548
rect 589976 125536 589982 125588
rect 591390 124176 591396 124228
rect 591448 124216 591454 124228
rect 603074 124216 603080 124228
rect 591448 124188 603080 124216
rect 591448 124176 591454 124188
rect 603074 124176 603080 124188
rect 603132 124176 603138 124228
rect 579246 124108 579252 124160
rect 579304 124148 579310 124160
rect 588538 124148 588544 124160
rect 579304 124120 588544 124148
rect 579304 124108 579310 124120
rect 588538 124108 588544 124120
rect 588596 124108 588602 124160
rect 667934 123836 667940 123888
rect 667992 123876 667998 123888
rect 671430 123876 671436 123888
rect 667992 123848 671436 123876
rect 667992 123836 667998 123848
rect 671430 123836 671436 123848
rect 671488 123836 671494 123888
rect 673362 122952 673368 123004
rect 673420 122992 673426 123004
rect 676214 122992 676220 123004
rect 673420 122964 676220 122992
rect 673420 122952 673426 122964
rect 676214 122952 676220 122964
rect 676272 122952 676278 123004
rect 589918 122816 589924 122868
rect 589976 122856 589982 122868
rect 603074 122856 603080 122868
rect 589976 122828 603080 122856
rect 589976 122816 589982 122828
rect 603074 122816 603080 122828
rect 603132 122816 603138 122868
rect 668854 122816 668860 122868
rect 668912 122856 668918 122868
rect 676214 122856 676220 122868
rect 668912 122828 676220 122856
rect 668912 122816 668918 122828
rect 676214 122816 676220 122828
rect 676272 122816 676278 122868
rect 587250 121456 587256 121508
rect 587308 121496 587314 121508
rect 603074 121496 603080 121508
rect 587308 121468 603080 121496
rect 587308 121456 587314 121468
rect 603074 121456 603080 121468
rect 603132 121456 603138 121508
rect 670142 121456 670148 121508
rect 670200 121496 670206 121508
rect 676122 121496 676128 121508
rect 670200 121468 676128 121496
rect 670200 121456 670206 121468
rect 676122 121456 676128 121468
rect 676180 121456 676186 121508
rect 579522 121388 579528 121440
rect 579580 121428 579586 121440
rect 583110 121428 583116 121440
rect 579580 121400 583116 121428
rect 579580 121388 579586 121400
rect 583110 121388 583116 121400
rect 583168 121388 583174 121440
rect 670050 120708 670056 120760
rect 670108 120748 670114 120760
rect 676214 120748 676220 120760
rect 670108 120720 676220 120748
rect 670108 120708 670114 120720
rect 676214 120708 676220 120720
rect 676272 120708 676278 120760
rect 588538 120096 588544 120148
rect 588596 120136 588602 120148
rect 603074 120136 603080 120148
rect 588596 120108 603080 120136
rect 588596 120096 588602 120108
rect 603074 120096 603080 120108
rect 603132 120096 603138 120148
rect 579246 120028 579252 120080
rect 579304 120068 579310 120080
rect 581730 120068 581736 120080
rect 579304 120040 581736 120068
rect 579304 120028 579310 120040
rect 581730 120028 581736 120040
rect 581788 120028 581794 120080
rect 579154 118668 579160 118720
rect 579212 118708 579218 118720
rect 603074 118708 603080 118720
rect 579212 118680 603080 118708
rect 579212 118668 579218 118680
rect 603074 118668 603080 118680
rect 603132 118668 603138 118720
rect 578602 118396 578608 118448
rect 578660 118436 578666 118448
rect 580350 118436 580356 118448
rect 578660 118408 580356 118436
rect 578660 118396 578666 118408
rect 580350 118396 580356 118408
rect 580408 118396 580414 118448
rect 669222 117784 669228 117836
rect 669280 117824 669286 117836
rect 674098 117824 674104 117836
rect 669280 117796 674104 117824
rect 669280 117784 669286 117796
rect 674098 117784 674104 117796
rect 674156 117784 674162 117836
rect 579062 117308 579068 117360
rect 579120 117348 579126 117360
rect 603074 117348 603080 117360
rect 579120 117320 603080 117348
rect 579120 117308 579126 117320
rect 603074 117308 603080 117320
rect 603132 117308 603138 117360
rect 579522 117240 579528 117292
rect 579580 117280 579586 117292
rect 603718 117280 603724 117292
rect 579580 117252 603724 117280
rect 579580 117240 579586 117252
rect 603718 117240 603724 117252
rect 603776 117240 603782 117292
rect 668486 117240 668492 117292
rect 668544 117280 668550 117292
rect 672994 117280 673000 117292
rect 668544 117252 673000 117280
rect 668544 117240 668550 117252
rect 672994 117240 673000 117252
rect 673052 117240 673058 117292
rect 675202 116560 675208 116612
rect 675260 116600 675266 116612
rect 683298 116600 683304 116612
rect 675260 116572 683304 116600
rect 675260 116560 675266 116572
rect 683298 116560 683304 116572
rect 683356 116560 683362 116612
rect 674650 116220 674656 116272
rect 674708 116260 674714 116272
rect 677594 116260 677600 116272
rect 674708 116232 677600 116260
rect 674708 116220 674714 116232
rect 677594 116220 677600 116232
rect 677652 116220 677658 116272
rect 678238 116192 678244 116204
rect 675036 116164 678244 116192
rect 600958 115948 600964 116000
rect 601016 115988 601022 116000
rect 603442 115988 603448 116000
rect 601016 115960 603448 115988
rect 601016 115948 601022 115960
rect 603442 115948 603448 115960
rect 603500 115948 603506 116000
rect 579522 115540 579528 115592
rect 579580 115580 579586 115592
rect 585778 115580 585784 115592
rect 579580 115552 585784 115580
rect 579580 115540 579586 115552
rect 585778 115540 585784 115552
rect 585836 115540 585842 115592
rect 675036 115444 675064 116164
rect 678238 116152 678244 116164
rect 678296 116152 678302 116204
rect 675110 115540 675116 115592
rect 675168 115580 675174 115592
rect 675386 115580 675392 115592
rect 675168 115552 675392 115580
rect 675168 115540 675174 115552
rect 675386 115540 675392 115552
rect 675444 115540 675450 115592
rect 675110 115444 675116 115456
rect 675036 115416 675116 115444
rect 675110 115404 675116 115416
rect 675168 115404 675174 115456
rect 675202 114792 675208 114844
rect 675260 114832 675266 114844
rect 675386 114832 675392 114844
rect 675260 114804 675392 114832
rect 675260 114792 675266 114804
rect 675386 114792 675392 114804
rect 675444 114792 675450 114844
rect 599578 114588 599584 114640
rect 599636 114628 599642 114640
rect 603166 114628 603172 114640
rect 599636 114600 603172 114628
rect 599636 114588 599642 114600
rect 603166 114588 603172 114600
rect 603224 114588 603230 114640
rect 674650 114588 674656 114640
rect 674708 114628 674714 114640
rect 675110 114628 675116 114640
rect 674708 114600 675116 114628
rect 674708 114588 674714 114600
rect 675110 114588 675116 114600
rect 675168 114588 675174 114640
rect 578970 114520 578976 114572
rect 579028 114560 579034 114572
rect 603074 114560 603080 114572
rect 579028 114532 603080 114560
rect 579028 114520 579034 114532
rect 603074 114520 603080 114532
rect 603132 114520 603138 114572
rect 579246 114452 579252 114504
rect 579304 114492 579310 114504
rect 591298 114492 591304 114504
rect 579304 114464 591304 114492
rect 579304 114452 579310 114464
rect 591298 114452 591304 114464
rect 591356 114452 591362 114504
rect 668486 114316 668492 114368
rect 668544 114356 668550 114368
rect 671338 114356 671344 114368
rect 668544 114328 671344 114356
rect 668544 114316 668550 114328
rect 671338 114316 671344 114328
rect 671396 114316 671402 114368
rect 578878 113160 578884 113212
rect 578936 113200 578942 113212
rect 603074 113200 603080 113212
rect 578936 113172 603080 113200
rect 578936 113160 578942 113172
rect 603074 113160 603080 113172
rect 603132 113160 603138 113212
rect 578418 112616 578424 112668
rect 578476 112656 578482 112668
rect 584398 112656 584404 112668
rect 578476 112628 584404 112656
rect 578476 112616 578482 112628
rect 584398 112616 584404 112628
rect 584456 112616 584462 112668
rect 583110 112412 583116 112464
rect 583168 112452 583174 112464
rect 603810 112452 603816 112464
rect 583168 112424 603816 112452
rect 583168 112412 583174 112424
rect 603810 112412 603816 112424
rect 603868 112412 603874 112464
rect 598198 111800 598204 111852
rect 598256 111840 598262 111852
rect 603074 111840 603080 111852
rect 598256 111812 603080 111840
rect 598256 111800 598262 111812
rect 603074 111800 603080 111812
rect 603132 111800 603138 111852
rect 578694 111732 578700 111784
rect 578752 111772 578758 111784
rect 598290 111772 598296 111784
rect 578752 111744 598296 111772
rect 578752 111732 578758 111744
rect 598290 111732 598296 111744
rect 598348 111732 598354 111784
rect 667934 111256 667940 111308
rect 667992 111296 667998 111308
rect 670142 111296 670148 111308
rect 667992 111268 670148 111296
rect 667992 111256 667998 111268
rect 670142 111256 670148 111268
rect 670200 111256 670206 111308
rect 675202 111120 675208 111172
rect 675260 111160 675266 111172
rect 675386 111160 675392 111172
rect 675260 111132 675392 111160
rect 675260 111120 675266 111132
rect 675386 111120 675392 111132
rect 675444 111120 675450 111172
rect 675110 110644 675116 110696
rect 675168 110684 675174 110696
rect 675386 110684 675392 110696
rect 675168 110656 675392 110684
rect 675168 110644 675174 110656
rect 675386 110644 675392 110656
rect 675444 110644 675450 110696
rect 595438 110440 595444 110492
rect 595496 110480 595502 110492
rect 603074 110480 603080 110492
rect 595496 110452 603080 110480
rect 595496 110440 595502 110452
rect 603074 110440 603080 110452
rect 603132 110440 603138 110492
rect 667934 110304 667940 110356
rect 667992 110344 667998 110356
rect 670050 110344 670056 110356
rect 667992 110316 670056 110344
rect 667992 110304 667998 110316
rect 670050 110304 670056 110316
rect 670108 110304 670114 110356
rect 579430 109556 579436 109608
rect 579488 109596 579494 109608
rect 583018 109596 583024 109608
rect 579488 109568 583024 109596
rect 579488 109556 579494 109568
rect 583018 109556 583024 109568
rect 583076 109556 583082 109608
rect 587158 109012 587164 109064
rect 587216 109052 587222 109064
rect 603074 109052 603080 109064
rect 587216 109024 603080 109052
rect 587216 109012 587222 109024
rect 603074 109012 603080 109024
rect 603132 109012 603138 109064
rect 579246 108740 579252 108792
rect 579304 108780 579310 108792
rect 581638 108780 581644 108792
rect 579304 108752 581644 108780
rect 579304 108740 579310 108752
rect 581638 108740 581644 108752
rect 581696 108740 581702 108792
rect 581730 107652 581736 107704
rect 581788 107692 581794 107704
rect 603074 107692 603080 107704
rect 581788 107664 603080 107692
rect 581788 107652 581794 107664
rect 603074 107652 603080 107664
rect 603132 107652 603138 107704
rect 579522 107584 579528 107636
rect 579580 107624 579586 107636
rect 587342 107624 587348 107636
rect 579580 107596 587348 107624
rect 579580 107584 579586 107596
rect 587342 107584 587348 107596
rect 587400 107584 587406 107636
rect 675110 106972 675116 107024
rect 675168 107012 675174 107024
rect 675386 107012 675392 107024
rect 675168 106984 675392 107012
rect 675168 106972 675174 106984
rect 675386 106972 675392 106984
rect 675444 106972 675450 107024
rect 675478 106564 675484 106616
rect 675536 106564 675542 106616
rect 585778 106292 585784 106344
rect 585836 106332 585842 106344
rect 603074 106332 603080 106344
rect 585836 106304 603080 106332
rect 585836 106292 585842 106304
rect 603074 106292 603080 106304
rect 603132 106292 603138 106344
rect 673362 106292 673368 106344
rect 673420 106332 673426 106344
rect 675496 106332 675524 106564
rect 673420 106304 675524 106332
rect 673420 106292 673426 106304
rect 579522 106224 579528 106276
rect 579580 106264 579586 106276
rect 588630 106264 588636 106276
rect 579580 106236 588636 106264
rect 579580 106224 579586 106236
rect 588630 106224 588636 106236
rect 588688 106224 588694 106276
rect 674742 106224 674748 106276
rect 674800 106264 674806 106276
rect 675386 106264 675392 106276
rect 674800 106236 675392 106264
rect 674800 106224 674806 106236
rect 675386 106224 675392 106236
rect 675444 106224 675450 106276
rect 669222 106088 669228 106140
rect 669280 106128 669286 106140
rect 672718 106128 672724 106140
rect 669280 106100 672724 106128
rect 669280 106088 669286 106100
rect 672718 106088 672724 106100
rect 672776 106088 672782 106140
rect 584398 104864 584404 104916
rect 584456 104904 584462 104916
rect 603074 104904 603080 104916
rect 584456 104876 603080 104904
rect 584456 104864 584462 104876
rect 603074 104864 603080 104876
rect 603132 104864 603138 104916
rect 596818 103912 596824 103964
rect 596876 103952 596882 103964
rect 603166 103952 603172 103964
rect 596876 103924 603172 103952
rect 596876 103912 596882 103924
rect 603166 103912 603172 103924
rect 603224 103912 603230 103964
rect 578510 103436 578516 103488
rect 578568 103476 578574 103488
rect 580258 103476 580264 103488
rect 578568 103448 580264 103476
rect 578568 103436 578574 103448
rect 580258 103436 580264 103448
rect 580316 103436 580322 103488
rect 583018 102212 583024 102264
rect 583076 102252 583082 102264
rect 603166 102252 603172 102264
rect 583076 102224 603172 102252
rect 583076 102212 583082 102224
rect 603166 102212 603172 102224
rect 603224 102212 603230 102264
rect 581638 102144 581644 102196
rect 581696 102184 581702 102196
rect 603074 102184 603080 102196
rect 581696 102156 603080 102184
rect 581696 102144 581702 102156
rect 603074 102144 603080 102156
rect 603132 102144 603138 102196
rect 578326 102076 578332 102128
rect 578384 102116 578390 102128
rect 590010 102116 590016 102128
rect 578384 102088 590016 102116
rect 578384 102076 578390 102088
rect 590010 102076 590016 102088
rect 590068 102076 590074 102128
rect 580258 100716 580264 100768
rect 580316 100756 580322 100768
rect 603074 100756 603080 100768
rect 580316 100728 603080 100756
rect 580316 100716 580322 100728
rect 603074 100716 603080 100728
rect 603132 100716 603138 100768
rect 578694 100648 578700 100700
rect 578752 100688 578758 100700
rect 596910 100688 596916 100700
rect 578752 100660 596916 100688
rect 578752 100648 578758 100660
rect 596910 100648 596916 100660
rect 596968 100648 596974 100700
rect 591298 99356 591304 99408
rect 591356 99396 591362 99408
rect 603074 99396 603080 99408
rect 591356 99368 603080 99396
rect 591356 99356 591362 99368
rect 603074 99356 603080 99368
rect 603132 99356 603138 99408
rect 579522 98880 579528 98932
rect 579580 98920 579586 98932
rect 585870 98920 585876 98932
rect 579580 98892 585876 98920
rect 579580 98880 579586 98892
rect 585870 98880 585876 98892
rect 585928 98880 585934 98932
rect 580350 98608 580356 98660
rect 580408 98648 580414 98660
rect 603810 98648 603816 98660
rect 580408 98620 603816 98648
rect 580408 98608 580414 98620
rect 603810 98608 603816 98620
rect 603868 98608 603874 98660
rect 625062 97928 625068 97980
rect 625120 97968 625126 97980
rect 625982 97968 625988 97980
rect 625120 97940 625988 97968
rect 625120 97928 625126 97940
rect 625982 97928 625988 97940
rect 626040 97928 626046 97980
rect 634446 97928 634452 97980
rect 634504 97968 634510 97980
rect 637574 97968 637580 97980
rect 634504 97940 637580 97968
rect 634504 97928 634510 97940
rect 637574 97928 637580 97940
rect 637632 97928 637638 97980
rect 638310 97928 638316 97980
rect 638368 97968 638374 97980
rect 644658 97968 644664 97980
rect 638368 97940 644664 97968
rect 638368 97928 638374 97940
rect 644658 97928 644664 97940
rect 644716 97928 644722 97980
rect 663058 97928 663064 97980
rect 663116 97968 663122 97980
rect 665358 97968 665364 97980
rect 663116 97940 665364 97968
rect 663116 97928 663122 97940
rect 665358 97928 665364 97940
rect 665416 97928 665422 97980
rect 624602 97860 624608 97912
rect 624660 97900 624666 97912
rect 625798 97900 625804 97912
rect 624660 97872 625804 97900
rect 624660 97860 624666 97872
rect 625798 97860 625804 97872
rect 625856 97860 625862 97912
rect 633066 97860 633072 97912
rect 633124 97900 633130 97912
rect 635274 97900 635280 97912
rect 633124 97872 635280 97900
rect 633124 97860 633130 97872
rect 635274 97860 635280 97872
rect 635332 97860 635338 97912
rect 633802 97792 633808 97844
rect 633860 97832 633866 97844
rect 636378 97832 636384 97844
rect 633860 97804 636384 97832
rect 633860 97792 633866 97804
rect 636378 97792 636384 97804
rect 636436 97792 636442 97844
rect 647510 97792 647516 97844
rect 647568 97832 647574 97844
rect 654778 97832 654784 97844
rect 647568 97804 654784 97832
rect 647568 97792 647574 97804
rect 654778 97792 654784 97804
rect 654836 97792 654842 97844
rect 637022 97724 637028 97776
rect 637080 97764 637086 97776
rect 642174 97764 642180 97776
rect 637080 97736 642180 97764
rect 637080 97724 637086 97736
rect 642174 97724 642180 97736
rect 642232 97724 642238 97776
rect 632422 97656 632428 97708
rect 632480 97696 632486 97708
rect 634078 97696 634084 97708
rect 632480 97668 634084 97696
rect 632480 97656 632486 97668
rect 634078 97656 634084 97668
rect 634136 97656 634142 97708
rect 635734 97656 635740 97708
rect 635792 97696 635798 97708
rect 639874 97696 639880 97708
rect 635792 97668 639880 97696
rect 635792 97656 635798 97668
rect 639874 97656 639880 97668
rect 639932 97656 639938 97708
rect 579522 97588 579528 97640
rect 579580 97628 579586 97640
rect 583110 97628 583116 97640
rect 579580 97600 583116 97628
rect 579580 97588 579586 97600
rect 583110 97588 583116 97600
rect 583168 97588 583174 97640
rect 631134 97588 631140 97640
rect 631192 97628 631198 97640
rect 632146 97628 632152 97640
rect 631192 97600 632152 97628
rect 631192 97588 631198 97600
rect 632146 97588 632152 97600
rect 632204 97588 632210 97640
rect 637482 97588 637488 97640
rect 637540 97628 637546 97640
rect 644566 97628 644572 97640
rect 637540 97600 644572 97628
rect 637540 97588 637546 97600
rect 644566 97588 644572 97600
rect 644624 97588 644630 97640
rect 635090 97520 635096 97572
rect 635148 97560 635154 97572
rect 639046 97560 639052 97572
rect 635148 97532 639052 97560
rect 635148 97520 635154 97532
rect 639046 97520 639052 97532
rect 639104 97520 639110 97572
rect 614850 97452 614856 97504
rect 614908 97492 614914 97504
rect 621658 97492 621664 97504
rect 614908 97464 621664 97492
rect 614908 97452 614914 97464
rect 621658 97452 621664 97464
rect 621716 97452 621722 97504
rect 643554 97452 643560 97504
rect 643612 97492 643618 97504
rect 660390 97492 660396 97504
rect 643612 97464 660396 97492
rect 643612 97452 643618 97464
rect 660390 97452 660396 97464
rect 660448 97452 660454 97504
rect 620738 97384 620744 97436
rect 620796 97424 620802 97436
rect 646038 97424 646044 97436
rect 620796 97396 646044 97424
rect 620796 97384 620802 97396
rect 646038 97384 646044 97396
rect 646096 97384 646102 97436
rect 649442 97384 649448 97436
rect 649500 97424 649506 97436
rect 658826 97424 658832 97436
rect 649500 97396 658832 97424
rect 649500 97384 649506 97396
rect 658826 97384 658832 97396
rect 658884 97384 658890 97436
rect 648154 97316 648160 97368
rect 648212 97356 648218 97368
rect 660114 97356 660120 97368
rect 648212 97328 660120 97356
rect 648212 97316 648218 97328
rect 660114 97316 660120 97328
rect 660172 97316 660178 97368
rect 622026 97248 622032 97300
rect 622084 97288 622090 97300
rect 648798 97288 648804 97300
rect 622084 97260 648804 97288
rect 622084 97248 622090 97260
rect 648798 97248 648804 97260
rect 648856 97248 648862 97300
rect 652018 97248 652024 97300
rect 652076 97288 652082 97300
rect 661954 97288 661960 97300
rect 652076 97260 661960 97288
rect 652076 97248 652082 97260
rect 661954 97248 661960 97260
rect 662012 97248 662018 97300
rect 621382 97180 621388 97232
rect 621440 97220 621446 97232
rect 647418 97220 647424 97232
rect 621440 97192 647424 97220
rect 621440 97180 621446 97192
rect 647418 97180 647424 97192
rect 647476 97180 647482 97232
rect 654686 97180 654692 97232
rect 654744 97220 654750 97232
rect 658366 97220 658372 97232
rect 654744 97192 658372 97220
rect 654744 97180 654750 97192
rect 658366 97180 658372 97192
rect 658424 97180 658430 97232
rect 659194 97180 659200 97232
rect 659252 97220 659258 97232
rect 662506 97220 662512 97232
rect 659252 97192 662512 97220
rect 659252 97180 659258 97192
rect 662506 97180 662512 97192
rect 662564 97180 662570 97232
rect 623682 97112 623688 97164
rect 623740 97152 623746 97164
rect 624418 97152 624424 97164
rect 623740 97124 624424 97152
rect 623740 97112 623746 97124
rect 624418 97112 624424 97124
rect 624476 97112 624482 97164
rect 657722 97112 657728 97164
rect 657780 97152 657786 97164
rect 660666 97152 660672 97164
rect 657780 97124 660672 97152
rect 657780 97112 657786 97124
rect 660666 97112 660672 97124
rect 660724 97112 660730 97164
rect 662322 97112 662328 97164
rect 662380 97152 662386 97164
rect 663978 97152 663984 97164
rect 662380 97124 663984 97152
rect 662380 97112 662386 97124
rect 663978 97112 663984 97124
rect 664036 97112 664042 97164
rect 610066 96908 610072 96960
rect 610124 96948 610130 96960
rect 610894 96948 610900 96960
rect 610124 96920 610900 96948
rect 610124 96908 610130 96920
rect 610894 96908 610900 96920
rect 610952 96908 610958 96960
rect 616138 96908 616144 96960
rect 616196 96948 616202 96960
rect 616782 96948 616788 96960
rect 616196 96920 616788 96948
rect 616196 96908 616202 96920
rect 616782 96908 616788 96920
rect 616840 96908 616846 96960
rect 617426 96908 617432 96960
rect 617484 96948 617490 96960
rect 618162 96948 618168 96960
rect 617484 96920 618168 96948
rect 617484 96908 617490 96920
rect 618162 96908 618168 96920
rect 618220 96908 618226 96960
rect 622670 96908 622676 96960
rect 622728 96948 622734 96960
rect 623590 96948 623596 96960
rect 622728 96920 623596 96948
rect 622728 96908 622734 96920
rect 623590 96908 623596 96920
rect 623648 96908 623654 96960
rect 625890 96908 625896 96960
rect 625948 96948 625954 96960
rect 626442 96948 626448 96960
rect 625948 96920 626448 96948
rect 625948 96908 625954 96920
rect 626442 96908 626448 96920
rect 626500 96908 626506 96960
rect 644842 96908 644848 96960
rect 644900 96948 644906 96960
rect 646498 96948 646504 96960
rect 644900 96920 646504 96948
rect 644900 96908 644906 96920
rect 646498 96908 646504 96920
rect 646556 96908 646562 96960
rect 650730 96908 650736 96960
rect 650788 96948 650794 96960
rect 651190 96948 651196 96960
rect 650788 96920 651196 96948
rect 650788 96908 650794 96920
rect 651190 96908 651196 96920
rect 651248 96908 651254 96960
rect 655422 96908 655428 96960
rect 655480 96948 655486 96960
rect 659286 96948 659292 96960
rect 655480 96920 659292 96948
rect 655480 96908 655486 96920
rect 659286 96908 659292 96920
rect 659344 96908 659350 96960
rect 618714 96840 618720 96892
rect 618772 96880 618778 96892
rect 619542 96880 619548 96892
rect 618772 96852 619548 96880
rect 618772 96840 618778 96852
rect 619542 96840 619548 96852
rect 619600 96840 619606 96892
rect 620002 96840 620008 96892
rect 620060 96880 620066 96892
rect 620922 96880 620928 96892
rect 620060 96852 620928 96880
rect 620060 96840 620066 96852
rect 620922 96840 620928 96852
rect 620980 96840 620986 96892
rect 640978 96840 640984 96892
rect 641036 96880 641042 96892
rect 643278 96880 643284 96892
rect 641036 96852 643284 96880
rect 641036 96840 641042 96852
rect 643278 96840 643284 96852
rect 643336 96840 643342 96892
rect 660574 96840 660580 96892
rect 660632 96880 660638 96892
rect 661402 96880 661408 96892
rect 660632 96852 661408 96880
rect 660632 96840 660638 96852
rect 661402 96840 661408 96852
rect 661460 96840 661466 96892
rect 655974 96772 655980 96824
rect 656032 96812 656038 96824
rect 659562 96812 659568 96824
rect 656032 96784 659568 96812
rect 656032 96772 656038 96784
rect 659562 96772 659568 96784
rect 659620 96772 659626 96824
rect 631778 96704 631784 96756
rect 631836 96744 631842 96756
rect 632974 96744 632980 96756
rect 631836 96716 632980 96744
rect 631836 96704 631842 96716
rect 632974 96704 632980 96716
rect 633032 96704 633038 96756
rect 636102 96704 636108 96756
rect 636160 96744 636166 96756
rect 640978 96744 640984 96756
rect 636160 96716 640984 96744
rect 636160 96704 636166 96716
rect 640978 96704 640984 96716
rect 641036 96704 641042 96756
rect 661862 96704 661868 96756
rect 661920 96744 661926 96756
rect 663058 96744 663064 96756
rect 661920 96716 663064 96744
rect 661920 96704 661926 96716
rect 663058 96704 663064 96716
rect 663116 96704 663122 96756
rect 578602 96568 578608 96620
rect 578660 96608 578666 96620
rect 594058 96608 594064 96620
rect 578660 96580 594064 96608
rect 578660 96568 578666 96580
rect 594058 96568 594064 96580
rect 594116 96568 594122 96620
rect 640242 96568 640248 96620
rect 640300 96608 640306 96620
rect 643186 96608 643192 96620
rect 640300 96580 643192 96608
rect 640300 96568 640306 96580
rect 643186 96568 643192 96580
rect 643244 96568 643250 96620
rect 656802 96568 656808 96620
rect 656860 96608 656866 96620
rect 658274 96608 658280 96620
rect 656860 96580 658280 96608
rect 656860 96568 656866 96580
rect 658274 96568 658280 96580
rect 658332 96568 658338 96620
rect 638862 96500 638868 96552
rect 638920 96540 638926 96552
rect 643094 96540 643100 96552
rect 638920 96512 643100 96540
rect 638920 96500 638926 96512
rect 643094 96500 643100 96512
rect 643152 96500 643158 96552
rect 656618 96160 656624 96212
rect 656676 96200 656682 96212
rect 663886 96200 663892 96212
rect 656676 96172 663892 96200
rect 656676 96160 656682 96172
rect 663886 96160 663892 96172
rect 663944 96160 663950 96212
rect 646774 96024 646780 96076
rect 646832 96064 646838 96076
rect 663794 96064 663800 96076
rect 646832 96036 663800 96064
rect 646832 96024 646838 96036
rect 663794 96024 663800 96036
rect 663852 96024 663858 96076
rect 653306 95956 653312 96008
rect 653364 95996 653370 96008
rect 665266 95996 665272 96008
rect 653364 95968 665272 95996
rect 653364 95956 653370 95968
rect 665266 95956 665272 95968
rect 665324 95956 665330 96008
rect 639598 95888 639604 95940
rect 639656 95928 639662 95940
rect 644474 95928 644480 95940
rect 639656 95900 644480 95928
rect 639656 95888 639662 95900
rect 644474 95888 644480 95900
rect 644532 95888 644538 95940
rect 646130 95888 646136 95940
rect 646188 95928 646194 95940
rect 665174 95928 665180 95940
rect 646188 95900 665180 95928
rect 646188 95888 646194 95900
rect 665174 95888 665180 95900
rect 665232 95888 665238 95940
rect 641622 95820 641628 95872
rect 641680 95860 641686 95872
rect 645854 95860 645860 95872
rect 641680 95832 645860 95860
rect 641680 95820 641686 95832
rect 645854 95820 645860 95832
rect 645912 95820 645918 95872
rect 607214 95480 607220 95532
rect 607272 95520 607278 95532
rect 607674 95520 607680 95532
rect 607272 95492 607680 95520
rect 607272 95480 607278 95492
rect 607674 95480 607680 95492
rect 607732 95480 607738 95532
rect 657262 95208 657268 95260
rect 657320 95248 657326 95260
rect 664070 95248 664076 95260
rect 657320 95220 664076 95248
rect 657320 95208 657326 95220
rect 664070 95208 664076 95220
rect 664128 95208 664134 95260
rect 578694 95140 578700 95192
rect 578752 95180 578758 95192
rect 584490 95180 584496 95192
rect 578752 95152 584496 95180
rect 578752 95140 578758 95152
rect 584490 95140 584496 95152
rect 584548 95140 584554 95192
rect 579522 93780 579528 93832
rect 579580 93820 579586 93832
rect 592678 93820 592684 93832
rect 579580 93792 592684 93820
rect 579580 93780 579586 93792
rect 592678 93780 592684 93792
rect 592736 93780 592742 93832
rect 646498 93100 646504 93152
rect 646556 93140 646562 93152
rect 654870 93140 654876 93152
rect 646556 93112 654876 93140
rect 646556 93100 646562 93112
rect 654870 93100 654876 93112
rect 654928 93100 654934 93152
rect 579522 92420 579528 92472
rect 579580 92460 579586 92472
rect 601050 92460 601056 92472
rect 579580 92432 601056 92460
rect 579580 92420 579586 92432
rect 601050 92420 601056 92432
rect 601108 92420 601114 92472
rect 644382 92420 644388 92472
rect 644440 92460 644446 92472
rect 654318 92460 654324 92472
rect 644440 92432 654324 92460
rect 644440 92420 644446 92432
rect 654318 92420 654324 92432
rect 654376 92420 654382 92472
rect 579522 90992 579528 91044
rect 579580 91032 579586 91044
rect 591390 91032 591396 91044
rect 579580 91004 591396 91032
rect 579580 90992 579586 91004
rect 591390 90992 591396 91004
rect 591448 90992 591454 91044
rect 579522 89632 579528 89684
rect 579580 89672 579586 89684
rect 602430 89672 602436 89684
rect 579580 89644 602436 89672
rect 579580 89632 579586 89644
rect 602430 89632 602436 89644
rect 602488 89632 602494 89684
rect 616690 89632 616696 89684
rect 616748 89672 616754 89684
rect 626442 89672 626448 89684
rect 616748 89644 626448 89672
rect 616748 89632 616754 89644
rect 626442 89632 626448 89644
rect 626500 89632 626506 89684
rect 656802 88816 656808 88868
rect 656860 88856 656866 88868
rect 658090 88856 658096 88868
rect 656860 88828 658096 88856
rect 656860 88816 656866 88828
rect 658090 88816 658096 88828
rect 658148 88816 658154 88868
rect 662322 88816 662328 88868
rect 662380 88856 662386 88868
rect 663978 88856 663984 88868
rect 662380 88828 663984 88856
rect 662380 88816 662386 88828
rect 663978 88816 663984 88828
rect 664036 88816 664042 88868
rect 616782 88272 616788 88324
rect 616840 88312 616846 88324
rect 626442 88312 626448 88324
rect 616840 88284 626448 88312
rect 616840 88272 616846 88284
rect 626442 88272 626448 88284
rect 626500 88272 626506 88324
rect 659470 88272 659476 88324
rect 659528 88312 659534 88324
rect 663150 88312 663156 88324
rect 659528 88284 663156 88312
rect 659528 88272 659534 88284
rect 663150 88272 663156 88284
rect 663208 88272 663214 88324
rect 620922 88204 620928 88256
rect 620980 88244 620986 88256
rect 626350 88244 626356 88256
rect 620980 88216 626356 88244
rect 620980 88204 620986 88216
rect 626350 88204 626356 88216
rect 626408 88204 626414 88256
rect 579522 86912 579528 86964
rect 579580 86952 579586 86964
rect 589918 86952 589924 86964
rect 579580 86924 589924 86952
rect 579580 86912 579586 86924
rect 589918 86912 589924 86924
rect 589976 86912 589982 86964
rect 651282 86844 651288 86896
rect 651340 86884 651346 86896
rect 657170 86884 657176 86896
rect 651340 86856 657176 86884
rect 651340 86844 651346 86856
rect 657170 86844 657176 86856
rect 657228 86844 657234 86896
rect 649902 86776 649908 86828
rect 649960 86816 649966 86828
rect 660666 86816 660672 86828
rect 649960 86788 660672 86816
rect 649960 86776 649966 86788
rect 660666 86776 660672 86788
rect 660724 86776 660730 86828
rect 651190 86708 651196 86760
rect 651248 86748 651254 86760
rect 657722 86748 657728 86760
rect 651248 86720 657728 86748
rect 651248 86708 651254 86720
rect 657722 86708 657728 86720
rect 657780 86708 657786 86760
rect 652662 86640 652668 86692
rect 652720 86680 652726 86692
rect 662506 86680 662512 86692
rect 652720 86652 662512 86680
rect 652720 86640 652726 86652
rect 662506 86640 662512 86652
rect 662564 86640 662570 86692
rect 645670 86572 645676 86624
rect 645728 86612 645734 86624
rect 660114 86612 660120 86624
rect 645728 86584 660120 86612
rect 645728 86572 645734 86584
rect 660114 86572 660120 86584
rect 660172 86572 660178 86624
rect 648522 86504 648528 86556
rect 648580 86544 648586 86556
rect 661402 86544 661408 86556
rect 648580 86516 661408 86544
rect 648580 86504 648586 86516
rect 661402 86504 661408 86516
rect 661460 86504 661466 86556
rect 653950 86436 653956 86488
rect 654008 86476 654014 86488
rect 658826 86476 658832 86488
rect 654008 86448 658832 86476
rect 654008 86436 654014 86448
rect 658826 86436 658832 86448
rect 658884 86436 658890 86488
rect 619450 86232 619456 86284
rect 619508 86272 619514 86284
rect 626442 86272 626448 86284
rect 619508 86244 626448 86272
rect 619508 86232 619514 86244
rect 626442 86232 626448 86244
rect 626500 86232 626506 86284
rect 579522 85484 579528 85536
rect 579580 85524 579586 85536
rect 587250 85524 587256 85536
rect 579580 85496 587256 85524
rect 579580 85484 579586 85496
rect 587250 85484 587256 85496
rect 587308 85484 587314 85536
rect 619542 85484 619548 85536
rect 619600 85524 619606 85536
rect 626442 85524 626448 85536
rect 619600 85496 626448 85524
rect 619600 85484 619606 85496
rect 626442 85484 626448 85496
rect 626500 85484 626506 85536
rect 579522 84124 579528 84176
rect 579580 84164 579586 84176
rect 588538 84164 588544 84176
rect 579580 84136 588544 84164
rect 579580 84124 579586 84136
rect 588538 84124 588544 84136
rect 588596 84124 588602 84176
rect 618070 84124 618076 84176
rect 618128 84164 618134 84176
rect 625614 84164 625620 84176
rect 618128 84136 625620 84164
rect 618128 84124 618134 84136
rect 625614 84124 625620 84136
rect 625672 84124 625678 84176
rect 618162 84056 618168 84108
rect 618220 84096 618226 84108
rect 626442 84096 626448 84108
rect 618220 84068 626448 84096
rect 618220 84056 618226 84068
rect 626442 84056 626448 84068
rect 626500 84056 626506 84108
rect 578510 81336 578516 81388
rect 578568 81376 578574 81388
rect 602338 81376 602344 81388
rect 578568 81348 602344 81376
rect 578568 81336 578574 81348
rect 602338 81336 602344 81348
rect 602396 81336 602402 81388
rect 579522 78616 579528 78668
rect 579580 78656 579586 78668
rect 600958 78656 600964 78668
rect 579580 78628 600964 78656
rect 579580 78616 579586 78628
rect 600958 78616 600964 78628
rect 601016 78616 601022 78668
rect 626442 78140 626448 78192
rect 626500 78180 626506 78192
rect 642450 78180 642456 78192
rect 626500 78152 642456 78180
rect 626500 78140 626506 78152
rect 642450 78140 642456 78152
rect 642508 78140 642514 78192
rect 631042 78072 631048 78124
rect 631100 78112 631106 78124
rect 638954 78112 638960 78124
rect 631100 78084 638960 78112
rect 631100 78072 631106 78084
rect 638954 78072 638960 78084
rect 639012 78072 639018 78124
rect 629202 78004 629208 78056
rect 629260 78044 629266 78056
rect 645302 78044 645308 78056
rect 629260 78016 645308 78044
rect 629260 78004 629266 78016
rect 645302 78004 645308 78016
rect 645360 78004 645366 78056
rect 605742 77936 605748 77988
rect 605800 77976 605806 77988
rect 636746 77976 636752 77988
rect 605800 77948 636752 77976
rect 605800 77936 605806 77948
rect 636746 77936 636752 77948
rect 636804 77936 636810 77988
rect 628374 77596 628380 77648
rect 628432 77636 628438 77648
rect 631502 77636 631508 77648
rect 628432 77608 631508 77636
rect 628432 77596 628438 77608
rect 631502 77596 631508 77608
rect 631560 77596 631566 77648
rect 579062 77324 579068 77376
rect 579120 77364 579126 77376
rect 628374 77364 628380 77376
rect 579120 77336 628380 77364
rect 579120 77324 579126 77336
rect 628374 77324 628380 77336
rect 628432 77324 628438 77376
rect 576118 77256 576124 77308
rect 576176 77296 576182 77308
rect 631042 77296 631048 77308
rect 576176 77268 631048 77296
rect 576176 77256 576182 77268
rect 631042 77256 631048 77268
rect 631100 77256 631106 77308
rect 623590 76576 623596 76628
rect 623648 76616 623654 76628
rect 646314 76616 646320 76628
rect 623648 76588 646320 76616
rect 623648 76576 623654 76588
rect 646314 76576 646320 76588
rect 646372 76576 646378 76628
rect 624418 76508 624424 76560
rect 624476 76548 624482 76560
rect 646958 76548 646964 76560
rect 624476 76520 646964 76548
rect 624476 76508 624482 76520
rect 646958 76508 646964 76520
rect 647016 76508 647022 76560
rect 579522 75828 579528 75880
rect 579580 75868 579586 75880
rect 599578 75868 599584 75880
rect 579580 75840 599584 75868
rect 579580 75828 579586 75840
rect 599578 75828 599584 75840
rect 599636 75828 599642 75880
rect 623682 75216 623688 75268
rect 623740 75256 623746 75268
rect 646130 75256 646136 75268
rect 623740 75228 646136 75256
rect 623740 75216 623746 75228
rect 646130 75216 646136 75228
rect 646188 75216 646194 75268
rect 615402 75148 615408 75200
rect 615460 75188 615466 75200
rect 646866 75188 646872 75200
rect 615460 75160 646872 75188
rect 615460 75148 615466 75160
rect 646866 75148 646872 75160
rect 646924 75148 646930 75200
rect 646314 74468 646320 74520
rect 646372 74508 646378 74520
rect 647234 74508 647240 74520
rect 646372 74480 647240 74508
rect 646372 74468 646378 74480
rect 647234 74468 647240 74480
rect 647292 74468 647298 74520
rect 579522 71680 579528 71732
rect 579580 71720 579586 71732
rect 598198 71720 598204 71732
rect 579580 71692 598204 71720
rect 579580 71680 579586 71692
rect 598198 71680 598204 71692
rect 598256 71680 598262 71732
rect 623038 70388 623044 70440
rect 623096 70428 623102 70440
rect 623774 70428 623780 70440
rect 623096 70400 623780 70428
rect 623096 70388 623102 70400
rect 623774 70388 623780 70400
rect 623832 70388 623838 70440
rect 579522 70320 579528 70372
rect 579580 70360 579586 70372
rect 595438 70360 595444 70372
rect 579580 70332 595444 70360
rect 579580 70320 579586 70332
rect 595438 70320 595444 70332
rect 595496 70320 595502 70372
rect 578326 68892 578332 68944
rect 578384 68932 578390 68944
rect 580350 68932 580356 68944
rect 578384 68904 580356 68932
rect 578384 68892 578390 68904
rect 580350 68892 580356 68904
rect 580408 68892 580414 68944
rect 579522 67532 579528 67584
rect 579580 67572 579586 67584
rect 587158 67572 587164 67584
rect 579580 67544 587164 67572
rect 579580 67532 579586 67544
rect 587158 67532 587164 67544
rect 587216 67532 587222 67584
rect 579246 65764 579252 65816
rect 579304 65804 579310 65816
rect 581730 65804 581736 65816
rect 579304 65776 581736 65804
rect 579304 65764 579310 65776
rect 581730 65764 581736 65776
rect 581788 65764 581794 65816
rect 579522 64268 579528 64320
rect 579580 64308 579586 64320
rect 585778 64308 585784 64320
rect 579580 64280 585784 64308
rect 579580 64268 579586 64280
rect 585778 64268 585784 64280
rect 585836 64268 585842 64320
rect 579522 63452 579528 63504
rect 579580 63492 579586 63504
rect 596818 63492 596824 63504
rect 579580 63464 596824 63492
rect 579580 63452 579586 63464
rect 596818 63452 596824 63464
rect 596876 63452 596882 63504
rect 578694 61344 578700 61396
rect 578752 61384 578758 61396
rect 584398 61384 584404 61396
rect 578752 61356 584404 61384
rect 578752 61344 578758 61356
rect 584398 61344 584404 61356
rect 584456 61344 584462 61396
rect 578970 60664 578976 60716
rect 579028 60704 579034 60716
rect 603718 60704 603724 60716
rect 579028 60676 603724 60704
rect 579028 60664 579034 60676
rect 603718 60664 603724 60676
rect 603776 60664 603782 60716
rect 618898 59848 618904 59900
rect 618956 59888 618962 59900
rect 623038 59888 623044 59900
rect 618956 59860 623044 59888
rect 618956 59848 618962 59860
rect 623038 59848 623044 59860
rect 623096 59848 623102 59900
rect 578878 58760 578884 58812
rect 578936 58800 578942 58812
rect 583018 58800 583024 58812
rect 578936 58772 583024 58800
rect 578936 58760 578942 58772
rect 583018 58760 583024 58772
rect 583076 58760 583082 58812
rect 621658 58624 621664 58676
rect 621716 58664 621722 58676
rect 662414 58664 662420 58676
rect 621716 58636 662420 58664
rect 621716 58624 621722 58636
rect 662414 58624 662420 58636
rect 662472 58624 662478 58676
rect 578878 57876 578884 57928
rect 578936 57916 578942 57928
rect 581638 57916 581644 57928
rect 578936 57888 581644 57916
rect 578936 57876 578942 57888
rect 581638 57876 581644 57888
rect 581696 57876 581702 57928
rect 578326 57196 578332 57248
rect 578384 57236 578390 57248
rect 591298 57236 591304 57248
rect 578384 57208 591304 57236
rect 578384 57196 578390 57208
rect 591298 57196 591304 57208
rect 591356 57196 591362 57248
rect 578234 55632 578240 55684
rect 578292 55672 578298 55684
rect 580258 55672 580264 55684
rect 578292 55644 580264 55672
rect 578292 55632 578298 55644
rect 580258 55632 580264 55644
rect 580316 55632 580322 55684
rect 616322 53796 616328 53848
rect 616380 53836 616386 53848
rect 618898 53836 618904 53848
rect 616380 53808 618904 53836
rect 616380 53796 616386 53808
rect 618898 53796 618904 53808
rect 618956 53796 618962 53848
rect 52270 53116 52276 53168
rect 52328 53156 52334 53168
rect 346302 53156 346308 53168
rect 52328 53128 346308 53156
rect 52328 53116 52334 53128
rect 346302 53116 346308 53128
rect 346360 53116 346366 53168
rect 145374 53048 145380 53100
rect 145432 53088 145438 53100
rect 579062 53088 579068 53100
rect 145432 53060 579068 53088
rect 145432 53048 145438 53060
rect 579062 53048 579068 53060
rect 579120 53048 579126 53100
rect 347130 52368 347136 52420
rect 347188 52408 347194 52420
rect 616322 52408 616328 52420
rect 347188 52380 616328 52408
rect 347188 52368 347194 52380
rect 616322 52368 616328 52380
rect 616380 52368 616386 52420
rect 52178 51688 52184 51740
rect 52236 51728 52242 51740
rect 60734 51728 60740 51740
rect 52236 51700 60740 51728
rect 52236 51688 52242 51700
rect 60734 51688 60740 51700
rect 60792 51688 60798 51740
rect 60734 51008 60740 51060
rect 60792 51048 60798 51060
rect 150342 51048 150348 51060
rect 60792 51020 150348 51048
rect 60792 51008 60798 51020
rect 150342 51008 150348 51020
rect 150400 51048 150406 51060
rect 189074 51048 189080 51060
rect 150400 51020 189080 51048
rect 150400 51008 150406 51020
rect 189074 51008 189080 51020
rect 189132 51008 189138 51060
rect 478138 49716 478144 49768
rect 478196 49756 478202 49768
rect 478782 49756 478788 49768
rect 478196 49728 478788 49756
rect 478196 49716 478202 49728
rect 478782 49716 478788 49728
rect 478840 49716 478846 49768
rect 664438 49036 664444 49088
rect 664496 49076 664502 49088
rect 669958 49076 669964 49088
rect 664496 49048 669964 49076
rect 664496 49036 664502 49048
rect 669958 49036 669964 49048
rect 670016 49036 670022 49088
rect 648104 47126 649670 47188
rect 648104 46658 648157 47126
rect 649617 46738 649670 47126
rect 649617 46658 650160 46738
rect 648104 46598 650160 46658
rect 648104 46590 649670 46598
rect 241514 44956 241520 45008
rect 241572 44996 241578 45008
rect 246114 44996 246120 45008
rect 241572 44968 246120 44996
rect 241572 44956 241578 44968
rect 246114 44956 246120 44968
rect 246172 44956 246178 45008
rect 251082 44888 251088 44940
rect 251140 44928 251146 44940
rect 255866 44928 255872 44940
rect 251140 44900 255872 44928
rect 251140 44888 251146 44900
rect 255866 44888 255872 44900
rect 255924 44888 255930 44940
rect 241514 44820 241520 44872
rect 241572 44860 241578 44872
rect 246114 44860 246120 44872
rect 241572 44832 246120 44860
rect 241572 44820 241578 44832
rect 246114 44820 246120 44832
rect 246172 44820 246178 44872
rect 405550 44820 405556 44872
rect 405608 44860 405614 44872
rect 608778 44860 608784 44872
rect 405608 44832 608784 44860
rect 405608 44820 405614 44832
rect 608778 44820 608784 44832
rect 608836 44820 608842 44872
rect 251082 44752 251088 44804
rect 251140 44792 251146 44804
rect 255866 44792 255872 44804
rect 251140 44764 255872 44792
rect 251140 44752 251146 44764
rect 255866 44752 255872 44764
rect 255924 44752 255930 44804
rect 473170 42476 473176 42528
rect 473228 42476 473234 42528
<< via1 >>
rect 146944 1007088 146996 1007140
rect 154580 1007088 154632 1007140
rect 195428 1006952 195480 1007004
rect 203892 1006952 203944 1007004
rect 300308 1006952 300360 1007004
rect 308956 1006952 309008 1007004
rect 426348 1006884 426400 1006936
rect 429568 1006884 429620 1006936
rect 261024 1006816 261076 1006868
rect 268384 1006816 268436 1006868
rect 427176 1006816 427228 1006868
rect 440884 1006816 440936 1006868
rect 425152 1006748 425204 1006800
rect 469864 1006748 469916 1006800
rect 427544 1006680 427596 1006732
rect 443644 1006680 443696 1006732
rect 428004 1006612 428056 1006664
rect 448612 1006612 448664 1006664
rect 198004 1006544 198056 1006596
rect 203524 1006544 203576 1006596
rect 429568 1006544 429620 1006596
rect 441620 1006544 441672 1006596
rect 95884 1006476 95936 1006528
rect 103612 1006476 103664 1006528
rect 145748 1006476 145800 1006528
rect 94504 1006408 94556 1006460
rect 103152 1006408 103204 1006460
rect 144184 1006408 144236 1006460
rect 151636 1006408 151688 1006460
rect 423496 1006476 423548 1006528
rect 446404 1006476 446456 1006528
rect 154120 1006408 154172 1006460
rect 428464 1006408 428516 1006460
rect 457444 1006408 457496 1006460
rect 508688 1006408 508740 1006460
rect 515404 1006408 515456 1006460
rect 100116 1006340 100168 1006392
rect 104348 1006340 104400 1006392
rect 150440 1006340 150492 1006392
rect 177304 1006340 177356 1006392
rect 93308 1006272 93360 1006324
rect 100668 1006272 100720 1006324
rect 93124 1006204 93176 1006256
rect 101956 1006204 102008 1006256
rect 102784 1006204 102836 1006256
rect 108856 1006272 108908 1006324
rect 195152 1006272 195204 1006324
rect 204720 1006272 204772 1006324
rect 108488 1006204 108540 1006256
rect 113824 1006204 113876 1006256
rect 97264 1006136 97316 1006188
rect 104808 1006136 104860 1006188
rect 145564 1006136 145616 1006188
rect 156144 1006136 156196 1006188
rect 196624 1006136 196676 1006188
rect 205548 1006136 205600 1006188
rect 98276 1006068 98328 1006120
rect 99104 1006068 99156 1006120
rect 149704 1006068 149756 1006120
rect 150440 1006068 150492 1006120
rect 126244 1006000 126296 1006052
rect 145656 1006000 145708 1006052
rect 157432 1006068 157484 1006120
rect 159088 1006068 159140 1006120
rect 166264 1006068 166316 1006120
rect 195244 1006068 195296 1006120
rect 204352 1006068 204404 1006120
rect 228364 1006272 228416 1006324
rect 254676 1006272 254728 1006324
rect 258172 1006272 258224 1006324
rect 301504 1006340 301556 1006392
rect 310152 1006340 310204 1006392
rect 425980 1006340 426032 1006392
rect 451924 1006340 451976 1006392
rect 551928 1006340 551980 1006392
rect 574744 1006340 574796 1006392
rect 280804 1006272 280856 1006324
rect 300216 1006272 300268 1006324
rect 308128 1006272 308180 1006324
rect 423864 1006272 423916 1006324
rect 454684 1006272 454736 1006324
rect 501328 1006272 501380 1006324
rect 517520 1006272 517572 1006324
rect 553952 1006272 554004 1006324
rect 563796 1006272 563848 1006324
rect 252468 1006204 252520 1006256
rect 253296 1006204 253348 1006256
rect 300124 1006204 300176 1006256
rect 250444 1006136 250496 1006188
rect 256516 1006136 256568 1006188
rect 298744 1006136 298796 1006188
rect 306104 1006136 306156 1006188
rect 154488 1006000 154540 1006052
rect 160652 1006000 160704 1006052
rect 201040 1006000 201092 1006052
rect 201868 1006000 201920 1006052
rect 209596 1006068 209648 1006120
rect 216036 1006068 216088 1006120
rect 247684 1006068 247736 1006120
rect 258540 1006068 258592 1006120
rect 263048 1006068 263100 1006120
rect 269764 1006068 269816 1006120
rect 298928 1006068 298980 1006120
rect 305644 1006068 305696 1006120
rect 204904 1006000 204956 1006052
rect 208768 1006000 208820 1006052
rect 249064 1006000 249116 1006052
rect 255320 1006000 255372 1006052
rect 257344 1006000 257396 1006052
rect 259000 1006000 259052 1006052
rect 262680 1006000 262732 1006052
rect 268476 1006000 268528 1006052
rect 303528 1006000 303580 1006052
rect 304080 1006000 304132 1006052
rect 304908 1006000 304960 1006052
rect 357348 1006204 357400 1006256
rect 374644 1006204 374696 1006256
rect 430028 1006204 430080 1006256
rect 468484 1006204 468536 1006256
rect 505836 1006204 505888 1006256
rect 514760 1006204 514812 1006256
rect 555976 1006204 556028 1006256
rect 570604 1006204 570656 1006256
rect 361396 1006136 361448 1006188
rect 369216 1006136 369268 1006188
rect 424692 1006136 424744 1006188
rect 460204 1006136 460256 1006188
rect 358544 1006068 358596 1006120
rect 371884 1006068 371936 1006120
rect 425520 1006068 425572 1006120
rect 464988 1006068 465040 1006120
rect 498108 1006068 498160 1006120
rect 499672 1006068 499724 1006120
rect 504548 1006068 504600 1006120
rect 520832 1006136 520884 1006188
rect 557172 1006136 557224 1006188
rect 306472 1006000 306524 1006052
rect 307024 1006000 307076 1006052
rect 310612 1006000 310664 1006052
rect 314660 1006000 314712 1006052
rect 330484 1006000 330536 1006052
rect 353116 1006000 353168 1006052
rect 354496 1006000 354548 1006052
rect 356060 1006000 356112 1006052
rect 360844 1006000 360896 1006052
rect 420736 1006000 420788 1006052
rect 422668 1006000 422720 1006052
rect 505376 1006000 505428 1006052
rect 522304 1006068 522356 1006120
rect 549168 1006068 549220 1006120
rect 550272 1006068 550324 1006120
rect 551100 1006068 551152 1006120
rect 556804 1006068 556856 1006120
rect 553124 1006000 553176 1006052
rect 556712 1006000 556764 1006052
rect 573364 1006068 573416 1006120
rect 563704 1006000 563756 1006052
rect 143724 1005388 143776 1005440
rect 152556 1005388 152608 1005440
rect 428832 1005388 428884 1005440
rect 448520 1005388 448572 1005440
rect 360568 1005320 360620 1005372
rect 380164 1005320 380216 1005372
rect 432880 1005320 432932 1005372
rect 462320 1005320 462372 1005372
rect 509884 1005320 509936 1005372
rect 520924 1005320 520976 1005372
rect 215208 1005252 215260 1005304
rect 219440 1005252 219492 1005304
rect 356520 1005252 356572 1005304
rect 377404 1005252 377456 1005304
rect 432512 1005252 432564 1005304
rect 467104 1005252 467156 1005304
rect 502892 1005252 502944 1005304
rect 517612 1005252 517664 1005304
rect 564348 1005252 564400 1005304
rect 571984 1005252 572036 1005304
rect 149704 1004912 149756 1004964
rect 152924 1004912 152976 1004964
rect 160652 1004912 160704 1004964
rect 162860 1004912 162912 1004964
rect 208400 1004844 208452 1004896
rect 209780 1004844 209832 1004896
rect 304448 1004844 304500 1004896
rect 307300 1004844 307352 1004896
rect 363420 1004844 363472 1004896
rect 366364 1004844 366416 1004896
rect 151084 1004776 151136 1004828
rect 153752 1004776 153804 1004828
rect 159456 1004776 159508 1004828
rect 161480 1004776 161532 1004828
rect 304264 1004776 304316 1004828
rect 306932 1004776 306984 1004828
rect 361764 1004776 361816 1004828
rect 364984 1004776 365036 1004828
rect 499212 1004776 499264 1004828
rect 501696 1004776 501748 1004828
rect 150348 1004708 150400 1004760
rect 152096 1004708 152148 1004760
rect 160284 1004708 160336 1004760
rect 163504 1004708 163556 1004760
rect 208768 1004708 208820 1004760
rect 211804 1004708 211856 1004760
rect 305828 1004708 305880 1004760
rect 308588 1004708 308640 1004760
rect 364248 1004708 364300 1004760
rect 366548 1004708 366600 1004760
rect 499488 1004708 499540 1004760
rect 94596 1004640 94648 1004692
rect 103152 1004640 103204 1004692
rect 151268 1004640 151320 1004692
rect 153292 1004640 153344 1004692
rect 159824 1004640 159876 1004692
rect 162124 1004640 162176 1004692
rect 199384 1004640 199436 1004692
rect 202328 1004640 202380 1004692
rect 305644 1004640 305696 1004692
rect 307760 1004640 307812 1004692
rect 354588 1004640 354640 1004692
rect 362592 1004640 362644 1004692
rect 365168 1004640 365220 1004692
rect 356520 1004572 356572 1004624
rect 500500 1004708 500552 1004760
rect 504364 1004708 504416 1004760
rect 556344 1004708 556396 1004760
rect 559748 1004708 559800 1004760
rect 557632 1004640 557684 1004692
rect 559564 1004640 559616 1004692
rect 500500 1004572 500552 1004624
rect 499396 1004504 499448 1004556
rect 501328 1004504 501380 1004556
rect 514760 1004096 514812 1004148
rect 517980 1004096 518032 1004148
rect 358084 1003892 358136 1003944
rect 378324 1003892 378376 1003944
rect 448612 1003892 448664 1003944
rect 464804 1003892 464856 1003944
rect 499488 1003484 499540 1003536
rect 500960 1003484 501012 1003536
rect 106832 1002328 106884 1002380
rect 109868 1002328 109920 1002380
rect 106188 1002260 106240 1002312
rect 108488 1002260 108540 1002312
rect 97356 1002192 97408 1002244
rect 100300 1002192 100352 1002244
rect 106004 1002192 106056 1002244
rect 108304 1002192 108356 1002244
rect 95976 1002124 96028 1002176
rect 99472 1002124 99524 1002176
rect 107660 1002124 107712 1002176
rect 109684 1002124 109736 1002176
rect 158260 1002124 158312 1002176
rect 161112 1002124 161164 1002176
rect 98828 1002056 98880 1002108
rect 101496 1002056 101548 1002108
rect 105636 1002056 105688 1002108
rect 107752 1002056 107804 1002108
rect 144092 1002056 144144 1002108
rect 150348 1002056 150400 1002108
rect 155776 1002056 155828 1002108
rect 157340 1002056 157392 1002108
rect 157432 1002056 157484 1002108
rect 159364 1002056 159416 1002108
rect 98644 1001988 98696 1002040
rect 101128 1001988 101180 1002040
rect 104348 1001988 104400 1002040
rect 106648 1001988 106700 1002040
rect 107200 1001988 107252 1002040
rect 109040 1001988 109092 1002040
rect 148324 1001988 148376 1002040
rect 151728 1001988 151780 1002040
rect 158628 1001988 158680 1002040
rect 160192 1001988 160244 1002040
rect 97540 1001920 97592 1001972
rect 99932 1001920 99984 1001972
rect 100024 1001920 100076 1001972
rect 102324 1001920 102376 1001972
rect 106464 1001920 106516 1001972
rect 107936 1001920 107988 1001972
rect 108028 1001920 108080 1001972
rect 110512 1001920 110564 1001972
rect 148508 1001920 148560 1001972
rect 150900 1001920 150952 1001972
rect 156972 1001920 157024 1001972
rect 158720 1001920 158772 1001972
rect 207204 1002532 207256 1002584
rect 210424 1002192 210476 1002244
rect 213184 1002192 213236 1002244
rect 210056 1002124 210108 1002176
rect 212540 1002124 212592 1002176
rect 202144 1002056 202196 1002108
rect 205180 1002056 205232 1002108
rect 206744 1002056 206796 1002108
rect 208400 1002056 208452 1002108
rect 211252 1002056 211304 1002108
rect 213368 1002056 213420 1002108
rect 200764 1001988 200816 1002040
rect 202696 1001988 202748 1002040
rect 211712 1001988 211764 1002040
rect 215944 1001988 215996 1002040
rect 200948 1001920 201000 1001972
rect 203064 1001920 203116 1001972
rect 203524 1001920 203576 1001972
rect 205916 1001920 205968 1001972
rect 212080 1001920 212132 1001972
rect 213920 1001920 213972 1001972
rect 253664 1002600 253716 1002652
rect 552756 1002600 552808 1002652
rect 565912 1002600 565964 1002652
rect 246672 1002532 246724 1002584
rect 254952 1002532 255004 1002584
rect 552296 1002532 552348 1002584
rect 568672 1002532 568724 1002584
rect 559196 1002260 559248 1002312
rect 562324 1002260 562376 1002312
rect 260196 1002192 260248 1002244
rect 262864 1002192 262916 1002244
rect 559656 1002192 559708 1002244
rect 561772 1002192 561824 1002244
rect 253204 1002124 253256 1002176
rect 256148 1002124 256200 1002176
rect 261852 1002124 261904 1002176
rect 264244 1002124 264296 1002176
rect 558460 1002124 558512 1002176
rect 560944 1002124 560996 1002176
rect 561312 1002124 561364 1002176
rect 566464 1002124 566516 1002176
rect 253388 1002056 253440 1002108
rect 255688 1002056 255740 1002108
rect 261484 1002056 261536 1002108
rect 263600 1002056 263652 1002108
rect 502524 1002056 502576 1002108
rect 505100 1002056 505152 1002108
rect 553216 1002056 553268 1002108
rect 554780 1002056 554832 1002108
rect 560024 1002056 560076 1002108
rect 562508 1002056 562560 1002108
rect 251916 1001988 251968 1002040
rect 254492 1001988 254544 1002040
rect 254584 1001988 254636 1002040
rect 256976 1001988 257028 1002040
rect 260656 1001988 260708 1002040
rect 262220 1001988 262272 1002040
rect 311440 1001988 311492 1002040
rect 313372 1001988 313424 1002040
rect 357072 1001988 357124 1002040
rect 358912 1001988 358964 1002040
rect 361028 1001988 361080 1002040
rect 363604 1001988 363656 1002040
rect 365076 1001988 365128 1002040
rect 370504 1001988 370556 1002040
rect 500868 1001988 500920 1002040
rect 503352 1001988 503404 1002040
rect 551744 1001988 551796 1002040
rect 553952 1001988 554004 1002040
rect 558000 1001988 558052 1002040
rect 560392 1001988 560444 1002040
rect 560852 1001988 560904 1002040
rect 565084 1001988 565136 1002040
rect 249156 1001920 249208 1001972
rect 254124 1001920 254176 1001972
rect 254768 1001920 254820 1001972
rect 257804 1001920 257856 1001972
rect 259828 1001920 259880 1001972
rect 260932 1001920 260984 1001972
rect 263508 1001920 263560 1001972
rect 265624 1001920 265676 1001972
rect 302884 1001920 302936 1001972
rect 305276 1001920 305328 1001972
rect 310152 1001920 310204 1001972
rect 311900 1001920 311952 1001972
rect 355784 1001920 355836 1001972
rect 358544 1001920 358596 1001972
rect 358728 1001920 358780 1001972
rect 359372 1001920 359424 1001972
rect 360200 1001920 360252 1001972
rect 362224 1001920 362276 1001972
rect 365444 1001920 365496 1001972
rect 367744 1001920 367796 1001972
rect 420736 1001920 420788 1001972
rect 421472 1001920 421524 1001972
rect 424324 1001920 424376 1001972
rect 425704 1001920 425756 1001972
rect 464988 1001920 465040 1001972
rect 472532 1001920 472584 1001972
rect 502156 1001920 502208 1001972
rect 502892 1001920 502944 1001972
rect 505008 1001920 505060 1001972
rect 506664 1001920 506716 1001972
rect 550548 1001920 550600 1001972
rect 553124 1001920 553176 1001972
rect 558828 1001920 558880 1001972
rect 560300 1001920 560352 1001972
rect 560484 1001920 560536 1001972
rect 563060 1001920 563112 1001972
rect 195152 1001852 195204 1001904
rect 195336 1001852 195388 1001904
rect 206928 1001852 206980 1001904
rect 207572 1001852 207624 1001904
rect 246580 1001852 246632 1001904
rect 195152 1001580 195204 1001632
rect 247040 1001240 247092 1001292
rect 251916 1001240 251968 1001292
rect 92296 1001172 92348 1001224
rect 95976 1001172 96028 1001224
rect 247132 1001172 247184 1001224
rect 253388 1001172 253440 1001224
rect 425704 1001172 425756 1001224
rect 438768 1001172 438820 1001224
rect 251548 1000560 251600 1000612
rect 254676 1000560 254728 1000612
rect 250444 1000492 250496 1000544
rect 253204 1000492 253256 1000544
rect 612740 1000492 612792 1000544
rect 625528 1000492 625580 1000544
rect 197360 1000356 197412 1000408
rect 200948 1000356 201000 1000408
rect 563796 1000084 563848 1000136
rect 565820 1000084 565872 1000136
rect 565912 1000016 565964 1000068
rect 568764 1000016 568816 1000068
rect 426348 999744 426400 999796
rect 446312 999744 446364 999796
rect 499396 999744 499448 999796
rect 504272 999744 504324 999796
rect 505100 999744 505152 999796
rect 515956 999744 516008 999796
rect 551744 999744 551796 999796
rect 562232 999744 562284 999796
rect 563704 999744 563756 999796
rect 572720 999744 572772 999796
rect 95976 999676 96028 999728
rect 98828 999676 98880 999728
rect 94780 999336 94832 999388
rect 97540 999336 97592 999388
rect 251364 999132 251416 999184
rect 254768 999132 254820 999184
rect 298192 999132 298244 999184
rect 327540 999132 327592 999184
rect 618168 999132 618220 999184
rect 625436 999132 625488 999184
rect 92296 999064 92348 999116
rect 94596 999064 94648 999116
rect 446404 999064 446456 999116
rect 448612 999064 448664 999116
rect 357348 998724 357400 998776
rect 360200 998724 360252 998776
rect 464804 998724 464856 998776
rect 472440 998724 472492 998776
rect 360844 998588 360896 998640
rect 367376 998588 367428 998640
rect 380164 998588 380216 998640
rect 383568 998588 383620 998640
rect 550548 998588 550600 998640
rect 556160 998588 556212 998640
rect 358728 998520 358780 998572
rect 372436 998520 372488 998572
rect 355784 998452 355836 998504
rect 383384 998452 383436 998504
rect 448520 998452 448572 998504
rect 472348 998520 472400 998572
rect 500868 998452 500920 998504
rect 513288 998452 513340 998504
rect 517612 998452 517664 998504
rect 523868 998452 523920 998504
rect 92388 998384 92440 998436
rect 100116 998384 100168 998436
rect 195980 998384 196032 998436
rect 206284 998384 206336 998436
rect 246764 998384 246816 998436
rect 254584 998384 254636 998436
rect 354588 998384 354640 998436
rect 383568 998384 383620 998436
rect 441620 998384 441672 998436
rect 369216 998316 369268 998368
rect 372344 998316 372396 998368
rect 502156 998384 502208 998436
rect 516048 998384 516100 998436
rect 517520 998384 517572 998436
rect 523776 998384 523828 998436
rect 472624 998316 472676 998368
rect 202420 998248 202472 998300
rect 206928 998248 206980 998300
rect 506664 998248 506716 998300
rect 516692 998248 516744 998300
rect 430856 998112 430908 998164
rect 436744 998112 436796 998164
rect 429660 998044 429712 998096
rect 431960 998044 432012 998096
rect 507032 998044 507084 998096
rect 510068 998044 510120 998096
rect 195428 997976 195480 998028
rect 199384 997976 199436 998028
rect 428464 997976 428516 998028
rect 430856 997976 430908 998028
rect 431684 997976 431736 998028
rect 433984 997976 434036 998028
rect 508228 997976 508280 998028
rect 510896 997976 510948 998028
rect 614120 997976 614172 998028
rect 625620 997976 625672 998028
rect 312176 997908 312228 997960
rect 314936 997908 314988 997960
rect 430396 997908 430448 997960
rect 432144 997908 432196 997960
rect 507860 997908 507912 997960
rect 509884 997908 509936 997960
rect 313832 997840 313884 997892
rect 316040 997840 316092 997892
rect 429200 997840 429252 997892
rect 431224 997840 431276 997892
rect 432052 997840 432104 997892
rect 433432 997840 433484 997892
rect 506204 997840 506256 997892
rect 508504 997840 508556 997892
rect 509056 997840 509108 997892
rect 510712 997840 510764 997892
rect 143724 997772 143776 997824
rect 145748 997772 145800 997824
rect 195336 997772 195388 997824
rect 196624 997772 196676 997824
rect 246856 997772 246908 997824
rect 279332 997772 279384 997824
rect 303252 997772 303304 997824
rect 305828 997772 305880 997824
rect 313004 997772 313056 997824
rect 314752 997772 314804 997824
rect 315120 997772 315172 997824
rect 319444 997772 319496 997824
rect 400128 997772 400180 997824
rect 143816 997704 143868 997756
rect 161480 997704 161532 997756
rect 195244 997704 195296 997756
rect 211252 997704 211304 997756
rect 246580 997704 246632 997756
rect 261852 997704 261904 997756
rect 298376 997704 298428 997756
rect 316040 997704 316092 997756
rect 399944 997704 399996 997756
rect 433432 997704 433484 997756
rect 507400 997772 507452 997824
rect 509240 997772 509292 997824
rect 509516 997772 509568 997824
rect 514024 997772 514076 997824
rect 540336 997772 540388 997824
rect 575572 997772 575624 997824
rect 607128 997772 607180 997824
rect 625712 997908 625764 997960
rect 440240 997704 440292 997756
rect 488908 997704 488960 997756
rect 510712 997704 510764 997756
rect 559748 997704 559800 997756
rect 625804 997772 625856 997824
rect 143908 997636 143960 997688
rect 155776 997636 155828 997688
rect 400036 997636 400088 997688
rect 432052 997636 432104 997688
rect 540888 997636 540940 997688
rect 563060 997636 563112 997688
rect 565820 997636 565872 997688
rect 623688 997636 623740 997688
rect 554320 997568 554372 997620
rect 607128 997568 607180 997620
rect 92664 997500 92716 997552
rect 95976 997500 96028 997552
rect 554688 997500 554740 997552
rect 561496 997500 561548 997552
rect 562232 997500 562284 997552
rect 614120 997500 614172 997552
rect 553216 997432 553268 997484
rect 561588 997432 561640 997484
rect 568764 997432 568816 997484
rect 618168 997432 618220 997484
rect 154580 997364 154632 997416
rect 157340 997364 157392 997416
rect 573364 997364 573416 997416
rect 612740 997364 612792 997416
rect 215760 997296 215812 997348
rect 218888 997296 218940 997348
rect 369216 997296 369268 997348
rect 372344 997296 372396 997348
rect 113824 997228 113876 997280
rect 116124 997228 116176 997280
rect 164424 997228 164476 997280
rect 167552 997228 167604 997280
rect 268476 997228 268528 997280
rect 270316 997228 270368 997280
rect 436560 997228 436612 997280
rect 439688 997228 439740 997280
rect 515404 997228 515456 997280
rect 516692 997228 516744 997280
rect 564992 997228 565044 997280
rect 568120 997228 568172 997280
rect 572720 997228 572772 997280
rect 575204 997160 575256 997212
rect 580908 997160 580960 997212
rect 585140 997228 585192 997280
rect 590936 997228 590988 997280
rect 620284 997160 620336 997212
rect 92480 997092 92532 997144
rect 97356 997092 97408 997144
rect 112996 997092 113048 997144
rect 116124 997092 116176 997144
rect 164424 997092 164476 997144
rect 167552 997092 167604 997144
rect 195244 997092 195296 997144
rect 198004 997092 198056 997144
rect 200212 997092 200264 997144
rect 204904 997092 204956 997144
rect 319444 997092 319496 997144
rect 332600 997092 332652 997144
rect 556712 997092 556764 997144
rect 605932 997092 605984 997144
rect 92572 997024 92624 997076
rect 100024 997024 100076 997076
rect 327540 997024 327592 997076
rect 367836 997024 367888 997076
rect 570604 997024 570656 997076
rect 622400 997024 622452 997076
rect 365168 996956 365220 997008
rect 372344 996956 372396 997008
rect 564992 996888 565044 996940
rect 568120 996888 568172 996940
rect 575480 996820 575532 996872
rect 580724 996820 580776 996872
rect 585508 996820 585560 996872
rect 590568 996820 590620 996872
rect 298284 996616 298336 996668
rect 300216 996616 300268 996668
rect 144828 996344 144880 996396
rect 149704 996344 149756 996396
rect 299020 996344 299072 996396
rect 301504 996344 301556 996396
rect 159364 996140 159416 996192
rect 209780 996140 209832 996192
rect 213184 996140 213236 996192
rect 263600 996140 263652 996192
rect 264244 996140 264296 996192
rect 314752 996140 314804 996192
rect 431224 996140 431276 996192
rect 506572 996140 506624 996192
rect 508504 996140 508556 996192
rect 560392 996140 560444 996192
rect 108304 996072 108356 996124
rect 158720 996072 158772 996124
rect 211804 996072 211856 996124
rect 260932 996072 260984 996124
rect 262864 996072 262916 996124
rect 313372 996072 313424 996124
rect 366364 996072 366416 996124
rect 428464 996072 428516 996124
rect 509884 996072 509936 996124
rect 561772 996072 561824 996124
rect 109684 996004 109736 996056
rect 160192 996004 160244 996056
rect 166264 996004 166316 996056
rect 212540 996004 212592 996056
rect 216036 996004 216088 996056
rect 262220 996004 262272 996056
rect 268384 996004 268436 996056
rect 314936 996004 314988 996056
rect 367376 996004 367428 996056
rect 381544 996004 381596 996056
rect 468484 996004 468536 996056
rect 509240 996004 509292 996056
rect 510068 996004 510120 996056
rect 560300 996004 560352 996056
rect 89628 995800 89680 995852
rect 92388 995800 92440 995852
rect 137376 995800 137428 995852
rect 144092 995936 144144 995988
rect 144000 995868 144052 995920
rect 195428 995868 195480 995920
rect 137928 995800 137980 995852
rect 139216 995800 139268 995852
rect 91560 995732 91612 995784
rect 92296 995732 92348 995784
rect 141056 995732 141108 995784
rect 142896 995800 142948 995852
rect 143724 995800 143776 995852
rect 189448 995800 189500 995852
rect 194324 995800 194376 995852
rect 195336 995800 195388 995852
rect 240876 995800 240928 995852
rect 246488 995800 246540 995852
rect 284392 995800 284444 995852
rect 307024 995936 307076 995988
rect 364984 995936 365036 995988
rect 382096 995936 382148 995988
rect 382280 995936 382332 995988
rect 431960 995936 432012 995988
rect 436744 995936 436796 995988
rect 510896 995936 510948 995988
rect 625436 995936 625488 995988
rect 381544 995868 381596 995920
rect 294880 995800 294932 995852
rect 298192 995800 298244 995852
rect 383384 995800 383436 995852
rect 385040 995800 385092 995852
rect 523868 995868 523920 995920
rect 625896 995868 625948 995920
rect 393596 995800 393648 995852
rect 396632 995800 396684 995852
rect 400128 995800 400180 995852
rect 472532 995800 472584 995852
rect 477684 995800 477736 995852
rect 520832 995800 520884 995852
rect 527916 995800 527968 995852
rect 528560 995800 528612 995852
rect 536840 995800 536892 995852
rect 540336 995800 540388 995852
rect 625804 995800 625856 995852
rect 626540 995800 626592 995852
rect 630864 995800 630916 995852
rect 631508 995800 631560 995852
rect 86592 995664 86644 995716
rect 92204 995664 92256 995716
rect 143632 995732 143684 995784
rect 192484 995732 192536 995784
rect 195152 995732 195204 995784
rect 240048 995732 240100 995784
rect 246672 995732 246724 995784
rect 297272 995732 297324 995784
rect 298008 995732 298060 995784
rect 383660 995732 383712 995784
rect 384396 995732 384448 995784
rect 472624 995732 472676 995784
rect 474004 995732 474056 995784
rect 516048 995732 516100 995784
rect 516692 995732 516744 995784
rect 524052 995732 524104 995784
rect 524788 995732 524840 995784
rect 625712 995732 625764 995784
rect 627184 995732 627236 995784
rect 143908 995664 143960 995716
rect 190644 995664 190696 995716
rect 195704 995664 195756 995716
rect 245568 995664 245620 995716
rect 246764 995664 246816 995716
rect 383476 995664 383528 995716
rect 385684 995664 385736 995716
rect 472440 995664 472492 995716
rect 473360 995664 473412 995716
rect 523776 995664 523828 995716
rect 529756 995664 529808 995716
rect 625620 995664 625672 995716
rect 630220 995664 630272 995716
rect 55864 995596 55916 995648
rect 107752 995596 107804 995648
rect 243268 995596 243320 995648
rect 246856 995596 246908 995648
rect 279332 995596 279384 995648
rect 316408 995596 316460 995648
rect 472716 995596 472768 995648
rect 476396 995596 476448 995648
rect 515956 995596 516008 995648
rect 516692 995596 516744 995648
rect 559564 995596 559616 995648
rect 661684 995596 661736 995648
rect 472348 995528 472400 995580
rect 474740 995528 474792 995580
rect 625528 995528 625580 995580
rect 627920 995528 627972 995580
rect 369216 995460 369268 995512
rect 372344 995460 372396 995512
rect 513288 995460 513340 995512
rect 516692 995460 516744 995512
rect 370780 995324 370832 995376
rect 372344 995324 372396 995376
rect 438768 995324 438820 995376
rect 439688 995324 439740 995376
rect 515220 995324 515272 995376
rect 516692 995324 516744 995376
rect 522304 995256 522356 995308
rect 537392 995256 537444 995308
rect 81348 995188 81400 995240
rect 92664 995188 92716 995240
rect 183514 995188 183566 995240
rect 195520 995188 195572 995240
rect 239266 995188 239318 995240
rect 249156 995188 249208 995240
rect 370780 995188 370832 995240
rect 372344 995188 372396 995240
rect 77668 995120 77720 995172
rect 92572 995120 92624 995172
rect 133420 995120 133472 995172
rect 144184 995120 144236 995172
rect 180156 995120 180208 995172
rect 195980 995120 196032 995172
rect 235908 995120 235960 995172
rect 247132 995120 247184 995172
rect 287152 995120 287204 995172
rect 304448 995120 304500 995172
rect 504272 995120 504324 995172
rect 515220 995120 515272 995172
rect 516692 995120 516744 995172
rect 574744 995188 574796 995240
rect 636154 995188 636206 995240
rect 533712 995120 533764 995172
rect 620284 995120 620336 995172
rect 638960 995120 639012 995172
rect 78312 995052 78364 995104
rect 97264 995052 97316 995104
rect 128452 995052 128504 995104
rect 154580 995052 154632 995104
rect 180616 995052 180668 995104
rect 202144 995052 202196 995104
rect 217416 995052 217468 995104
rect 218888 995052 218940 995104
rect 231584 995052 231636 995104
rect 251548 995052 251600 995104
rect 286508 995052 286560 995104
rect 305644 995052 305696 995104
rect 460204 995052 460256 995104
rect 482284 995052 482336 995104
rect 504364 995052 504416 995104
rect 534356 995052 534408 995104
rect 568672 995052 568724 995104
rect 634820 995052 634872 995104
rect 77024 994984 77076 995036
rect 106648 994984 106700 995036
rect 165988 994984 166040 995036
rect 167552 994984 167604 995036
rect 183284 994984 183336 995036
rect 208400 994984 208452 995036
rect 232872 994984 232924 995036
rect 257344 994984 257396 995036
rect 282828 994984 282880 995036
rect 311900 994984 311952 995036
rect 357072 994984 357124 995036
rect 398840 994984 398892 995036
rect 457444 994984 457496 995036
rect 485964 994984 486016 995036
rect 499212 994984 499264 995036
rect 535552 994984 535604 995036
rect 556160 994984 556212 995036
rect 637028 994984 637080 995036
rect 440240 994236 440292 994288
rect 446128 994236 446180 994288
rect 562508 993012 562560 993064
rect 660304 993012 660356 993064
rect 88340 992944 88392 992996
rect 111800 992944 111852 992996
rect 498016 992944 498068 992996
rect 666652 992944 666704 992996
rect 46204 992876 46256 992928
rect 110512 992876 110564 992928
rect 245660 992876 245712 992928
rect 251456 992876 251508 992928
rect 353116 992876 353168 992928
rect 666836 992876 666888 992928
rect 560944 991652 560996 991704
rect 658924 991652 658976 991704
rect 549168 991584 549220 991636
rect 666560 991584 666612 991636
rect 367836 991516 367888 991568
rect 381636 991516 381688 991568
rect 420736 991516 420788 991568
rect 666744 991516 666796 991568
rect 44824 991448 44876 991500
rect 107936 991448 107988 991500
rect 203156 991448 203208 991500
rect 213920 991448 213972 991500
rect 215944 991448 215996 991500
rect 235632 991448 235684 991500
rect 303528 991448 303580 991500
rect 665456 991448 665508 991500
rect 47584 990088 47636 990140
rect 109040 990088 109092 990140
rect 138296 990088 138348 990140
rect 162860 990088 162912 990140
rect 269764 990088 269816 990140
rect 300492 990088 300544 990140
rect 370504 990088 370556 990140
rect 430304 990088 430356 990140
rect 435364 990088 435416 990140
rect 478972 990088 479024 990140
rect 514024 990088 514076 990140
rect 560116 990088 560168 990140
rect 562324 990088 562376 990140
rect 663064 990088 663116 990140
rect 566464 988728 566516 988780
rect 592500 988728 592552 988780
rect 330484 987368 330536 987420
rect 365444 987368 365496 987420
rect 512644 987368 512696 987420
rect 543832 987368 543884 987420
rect 565084 987368 565136 987420
rect 624976 987368 625028 987420
rect 88340 986620 88392 986672
rect 89628 986620 89680 986672
rect 265624 986620 265676 986672
rect 268108 986620 268160 986672
rect 367744 986008 367796 986060
rect 397828 986008 397880 986060
rect 73436 985940 73488 985992
rect 102784 985940 102836 985992
rect 267004 985940 267056 985992
rect 284300 985940 284352 985992
rect 318064 985940 318116 985992
rect 349160 985940 349212 985992
rect 369124 985940 369176 985992
rect 414112 985940 414164 985992
rect 467104 985940 467156 985992
rect 495164 985940 495216 985992
rect 571984 985940 572036 985992
rect 608784 985940 608836 985992
rect 163504 985872 163556 985924
rect 170772 985872 170824 985924
rect 520924 985736 520976 985788
rect 527640 985736 527692 985788
rect 280804 984784 280856 984836
rect 650000 984784 650052 984836
rect 228364 984716 228416 984768
rect 651380 984716 651432 984768
rect 177304 984648 177356 984700
rect 650092 984648 650144 984700
rect 126244 984580 126296 984632
rect 651472 984580 651524 984632
rect 42708 975672 42760 975724
rect 62120 975672 62172 975724
rect 651656 975672 651708 975724
rect 672724 975672 672776 975724
rect 42156 967240 42208 967292
rect 42708 967240 42760 967292
rect 42156 963976 42208 964028
rect 42800 963976 42852 964028
rect 42156 962820 42208 962872
rect 42892 962820 42944 962872
rect 44916 961868 44968 961920
rect 62120 961868 62172 961920
rect 669964 961868 670016 961920
rect 674840 961868 674892 961920
rect 675024 961324 675076 961376
rect 675392 961324 675444 961376
rect 42064 959692 42116 959744
rect 44180 959692 44232 959744
rect 42156 959080 42208 959132
rect 42984 959080 43036 959132
rect 674748 958196 674800 958248
rect 675392 958196 675444 958248
rect 659016 957788 659068 957840
rect 675024 957788 675076 957840
rect 673368 956972 673420 957024
rect 675392 956972 675444 957024
rect 673184 956088 673236 956140
rect 675484 956088 675536 956140
rect 675024 955476 675076 955528
rect 675484 955476 675536 955528
rect 42156 955340 42208 955392
rect 42340 955340 42392 955392
rect 41788 954592 41840 954644
rect 41788 954388 41840 954440
rect 32404 952824 32456 952876
rect 41788 952824 41840 952876
rect 37924 952212 37976 952264
rect 42340 952212 42392 952264
rect 675760 952008 675812 952060
rect 675760 951736 675812 951788
rect 675760 949424 675812 949476
rect 678244 949424 678296 949476
rect 651564 948064 651616 948116
rect 674196 948064 674248 948116
rect 27620 947316 27672 947368
rect 62120 947316 62172 947368
rect 35808 943236 35860 943288
rect 45744 943236 45796 943288
rect 35716 943168 35768 943220
rect 44916 943168 44968 943220
rect 652024 939768 652076 939820
rect 676036 939768 676088 939820
rect 674196 939156 674248 939208
rect 676036 939156 676088 939208
rect 672724 938680 672776 938732
rect 676220 938680 676272 938732
rect 660304 938544 660356 938596
rect 676036 938544 676088 938596
rect 674656 938272 674708 938324
rect 676036 938272 676088 938324
rect 673828 937456 673880 937508
rect 676036 937456 676088 937508
rect 663064 937320 663116 937372
rect 676220 937320 676272 937372
rect 658924 937184 658976 937236
rect 676220 937184 676272 937236
rect 45744 936980 45796 937032
rect 62120 936980 62172 937032
rect 651564 936980 651616 937032
rect 659016 936980 659068 937032
rect 672356 935756 672408 935808
rect 676036 935756 676088 935808
rect 672816 935688 672868 935740
rect 676128 935688 676180 935740
rect 661684 935620 661736 935672
rect 676220 935620 676272 935672
rect 39948 932356 40000 932408
rect 41696 932356 41748 932408
rect 41696 932152 41748 932204
rect 47584 932152 47636 932204
rect 673184 931608 673236 931660
rect 676036 931608 676088 931660
rect 674748 930724 674800 930776
rect 676220 930724 676272 930776
rect 673368 930248 673420 930300
rect 676220 930248 676272 930300
rect 671344 927392 671396 927444
rect 683120 927392 683172 927444
rect 47676 923244 47728 923296
rect 62120 923244 62172 923296
rect 651564 921816 651616 921868
rect 670056 921816 670108 921868
rect 54484 909440 54536 909492
rect 62120 909440 62172 909492
rect 651564 909440 651616 909492
rect 661684 909440 661736 909492
rect 51724 896996 51776 897048
rect 62120 896996 62172 897048
rect 651564 895636 651616 895688
rect 660304 895636 660356 895688
rect 48964 884620 49016 884672
rect 62120 884620 62172 884672
rect 674472 873536 674524 873588
rect 675392 873536 675444 873588
rect 673184 872652 673236 872704
rect 675392 872652 675444 872704
rect 674564 872176 674616 872228
rect 675392 872176 675444 872228
rect 44824 870816 44876 870868
rect 62120 870816 62172 870868
rect 674288 869796 674340 869848
rect 675392 869796 675444 869848
rect 673000 869660 673052 869712
rect 675392 869660 675444 869712
rect 673092 869592 673144 869644
rect 674932 869592 674984 869644
rect 651564 869388 651616 869440
rect 671436 869388 671488 869440
rect 674932 868708 674984 868760
rect 675392 868708 675444 868760
rect 652024 868640 652076 868692
rect 674932 868572 674984 868624
rect 674380 868504 674432 868556
rect 675484 868504 675536 868556
rect 674932 866192 674984 866244
rect 675392 866192 675444 866244
rect 672908 862792 672960 862844
rect 675484 862792 675536 862844
rect 43628 858372 43680 858424
rect 62120 858372 62172 858424
rect 651564 855584 651616 855636
rect 664444 855584 664496 855636
rect 53104 844568 53156 844620
rect 62120 844568 62172 844620
rect 651564 841780 651616 841832
rect 663064 841780 663116 841832
rect 50344 832124 50396 832176
rect 62120 832124 62172 832176
rect 651564 829404 651616 829456
rect 658924 829404 658976 829456
rect 43536 818320 43588 818372
rect 62120 818320 62172 818372
rect 41328 817504 41380 817556
rect 48964 817504 49016 817556
rect 41236 817368 41288 817420
rect 51724 817368 51776 817420
rect 651564 815600 651616 815652
rect 665824 815600 665876 815652
rect 40776 811520 40828 811572
rect 41788 811520 41840 811572
rect 39856 807236 39908 807288
rect 41788 807236 41840 807288
rect 49056 805944 49108 805996
rect 62120 805944 62172 805996
rect 42156 803836 42208 803888
rect 42616 803836 42668 803888
rect 42064 803768 42116 803820
rect 42708 803768 42760 803820
rect 651564 803156 651616 803208
rect 672724 803156 672776 803208
rect 35164 801116 35216 801168
rect 43076 801116 43128 801168
rect 32404 801048 32456 801100
rect 42892 801048 42944 801100
rect 40776 800504 40828 800556
rect 42984 800504 43036 800556
rect 42156 799960 42208 800012
rect 42340 799960 42392 800012
rect 43168 799008 43220 799060
rect 47676 799008 47728 799060
rect 42156 798124 42208 798176
rect 42616 798124 42668 798176
rect 42156 797240 42208 797292
rect 43168 797240 43220 797292
rect 42156 796288 42208 796340
rect 42708 796288 42760 796340
rect 42708 796152 42760 796204
rect 42892 796152 42944 796204
rect 42156 794996 42208 795048
rect 42432 794996 42484 795048
rect 42892 794928 42944 794980
rect 44364 794928 44416 794980
rect 42432 794860 42484 794912
rect 42984 794860 43036 794912
rect 42156 794248 42208 794300
rect 42708 794248 42760 794300
rect 42708 794112 42760 794164
rect 43076 794112 43128 794164
rect 42156 793772 42208 793824
rect 42892 793772 42944 793824
rect 54484 793500 54536 793552
rect 62120 793500 62172 793552
rect 42156 793160 42208 793212
rect 42432 793160 42484 793212
rect 42432 793024 42484 793076
rect 42800 793024 42852 793076
rect 42156 790644 42208 790696
rect 42800 790644 42852 790696
rect 42156 790100 42208 790152
rect 42432 790100 42484 790152
rect 42156 789420 42208 789472
rect 42340 789420 42392 789472
rect 651656 789352 651708 789404
rect 661776 789352 661828 789404
rect 42156 788808 42208 788860
rect 42708 788808 42760 788860
rect 670608 787992 670660 788044
rect 675392 787992 675444 788044
rect 674196 787312 674248 787364
rect 675392 787312 675444 787364
rect 42156 786972 42208 787024
rect 42432 786972 42484 787024
rect 672632 786700 672684 786752
rect 675392 786700 675444 786752
rect 42156 785612 42208 785664
rect 42708 785612 42760 785664
rect 674012 784252 674064 784304
rect 675392 784252 675444 784304
rect 673276 782892 673328 782944
rect 675484 782892 675536 782944
rect 672540 780716 672592 780768
rect 675484 780716 675536 780768
rect 673644 779968 673696 780020
rect 675484 779968 675536 780020
rect 51724 779696 51776 779748
rect 62120 779696 62172 779748
rect 658924 778948 658976 779000
rect 674748 778948 674800 779000
rect 673920 778608 673972 778660
rect 675484 778608 675536 778660
rect 672448 777316 672500 777368
rect 675392 777316 675444 777368
rect 674748 777044 674800 777096
rect 675392 777044 675444 777096
rect 651564 775548 651616 775600
rect 658924 775548 658976 775600
rect 35808 774188 35860 774240
rect 53104 774188 53156 774240
rect 672172 773576 672224 773628
rect 675484 773576 675536 773628
rect 46204 767320 46256 767372
rect 62120 767320 62172 767372
rect 651564 763172 651616 763224
rect 664536 763172 664588 763224
rect 41512 761744 41564 761796
rect 48964 761744 49016 761796
rect 670056 760792 670108 760844
rect 676220 760792 676272 760844
rect 661684 760656 661736 760708
rect 676128 760656 676180 760708
rect 660304 760520 660356 760572
rect 676036 760520 676088 760572
rect 674656 760316 674708 760368
rect 676036 760316 676088 760368
rect 31024 759636 31076 759688
rect 41880 759636 41932 759688
rect 673828 759500 673880 759552
rect 676036 759500 676088 759552
rect 673368 759092 673420 759144
rect 676220 759092 676272 759144
rect 672264 759024 672316 759076
rect 676036 759024 676088 759076
rect 33784 758480 33836 758532
rect 42432 758480 42484 758532
rect 32496 758344 32548 758396
rect 42708 758344 42760 758396
rect 32404 758276 32456 758328
rect 43168 758276 43220 758328
rect 674656 758208 674708 758260
rect 676036 758208 676088 758260
rect 41880 756984 41932 757036
rect 41880 756712 41932 756764
rect 43260 756236 43312 756288
rect 44824 756236 44876 756288
rect 674288 755556 674340 755608
rect 676220 755556 676272 755608
rect 42432 755488 42484 755540
rect 42156 755420 42208 755472
rect 42616 755216 42668 755268
rect 43168 755216 43220 755268
rect 42156 755148 42208 755200
rect 672908 754944 672960 754996
rect 676036 754944 676088 754996
rect 42156 754876 42208 754928
rect 674472 754332 674524 754384
rect 676220 754332 676272 754384
rect 42064 754060 42116 754112
rect 43260 754060 43312 754112
rect 673184 753584 673236 753636
rect 676036 753584 676088 753636
rect 44916 753516 44968 753568
rect 62120 753516 62172 753568
rect 674380 753108 674432 753160
rect 676220 753108 676272 753160
rect 674564 752700 674616 752752
rect 676220 752700 676272 752752
rect 673000 752224 673052 752276
rect 676220 752224 676272 752276
rect 43076 752088 43128 752140
rect 44456 752088 44508 752140
rect 42156 751068 42208 751120
rect 42984 751068 43036 751120
rect 673092 750864 673144 750916
rect 676220 750864 676272 750916
rect 42156 749776 42208 749828
rect 43076 749776 43128 749828
rect 651564 749436 651616 749488
rect 672816 749436 672868 749488
rect 42984 749368 43036 749420
rect 44548 749368 44600 749420
rect 670056 749368 670108 749420
rect 683120 749368 683172 749420
rect 42984 746988 43036 747040
rect 42064 746920 42116 746972
rect 42156 746920 42208 746972
rect 42708 746920 42760 746972
rect 42708 746784 42760 746836
rect 42892 746784 42944 746836
rect 42616 746648 42668 746700
rect 43076 746648 43128 746700
rect 42156 746036 42208 746088
rect 42708 746036 42760 746088
rect 42708 745900 42760 745952
rect 44364 745900 44416 745952
rect 42156 745424 42208 745476
rect 43076 745424 43128 745476
rect 42156 743724 42208 743776
rect 42708 743724 42760 743776
rect 42156 743248 42208 743300
rect 42616 743248 42668 743300
rect 671988 743180 672040 743232
rect 675392 743180 675444 743232
rect 672356 742500 672408 742552
rect 675392 742500 675444 742552
rect 50436 741072 50488 741124
rect 62120 741072 62172 741124
rect 673184 739100 673236 739152
rect 675392 739100 675444 739152
rect 673736 738216 673788 738268
rect 675392 738216 675444 738268
rect 674288 735632 674340 735684
rect 675392 735632 675444 735684
rect 651564 735564 651616 735616
rect 660304 735564 660356 735616
rect 673092 734952 673144 735004
rect 675392 734952 675444 735004
rect 658924 734816 658976 734868
rect 674564 734340 674616 734392
rect 674472 733592 674524 733644
rect 675392 733592 675444 733644
rect 674564 732028 674616 732080
rect 675392 732028 675444 732080
rect 31392 731348 31444 731400
rect 44732 731348 44784 731400
rect 31576 731280 31628 731332
rect 49056 731212 49108 731264
rect 31668 731144 31720 731196
rect 51724 731076 51776 731128
rect 31484 731008 31536 731060
rect 54484 730940 54536 730992
rect 674472 730464 674524 730516
rect 675392 730464 675444 730516
rect 673828 728628 673880 728680
rect 675484 728628 675536 728680
rect 47676 727268 47728 727320
rect 62120 727268 62172 727320
rect 652024 723120 652076 723172
rect 658924 723120 658976 723172
rect 41512 719652 41564 719704
rect 50344 719652 50396 719704
rect 42156 716864 42208 716916
rect 42524 716864 42576 716916
rect 664444 716252 664496 716304
rect 676036 716252 676088 716304
rect 40868 716184 40920 716236
rect 41880 716184 41932 716236
rect 671436 716116 671488 716168
rect 676036 716116 676088 716168
rect 34428 715504 34480 715556
rect 42156 715504 42208 715556
rect 673368 715300 673420 715352
rect 675944 715300 675996 715352
rect 663064 714960 663116 715012
rect 676036 714960 676088 715012
rect 44824 714824 44876 714876
rect 62120 714824 62172 714876
rect 672908 714824 672960 714876
rect 676036 714824 676088 714876
rect 40684 714756 40736 714808
rect 42432 714756 42484 714808
rect 672264 714484 672316 714536
rect 676036 714484 676088 714536
rect 672264 714008 672316 714060
rect 676036 714008 676088 714060
rect 41880 713804 41932 713856
rect 42156 713804 42208 713856
rect 41880 713532 41932 713584
rect 674656 713668 674708 713720
rect 676036 713668 676088 713720
rect 673460 713192 673512 713244
rect 676036 713192 676088 713244
rect 673552 712376 673604 712428
rect 676036 712376 676088 712428
rect 42524 712104 42576 712156
rect 672632 712036 672684 712088
rect 676036 712036 676088 712088
rect 670608 711220 670660 711272
rect 676036 711220 676088 711272
rect 42524 710948 42576 711000
rect 42984 710948 43036 711000
rect 42156 710880 42208 710932
rect 43536 710880 43588 710932
rect 672540 710404 672592 710456
rect 676036 710404 676088 710456
rect 672172 709996 672224 710048
rect 676036 709996 676088 710048
rect 674196 709588 674248 709640
rect 676036 709588 676088 709640
rect 43168 709316 43220 709368
rect 44548 709316 44600 709368
rect 651564 709316 651616 709368
rect 671436 709316 671488 709368
rect 674012 709180 674064 709232
rect 676036 709180 676088 709232
rect 42156 708568 42208 708620
rect 42524 708568 42576 708620
rect 672448 708364 672500 708416
rect 676036 708364 676088 708416
rect 676036 708228 676088 708280
rect 677324 708228 677376 708280
rect 42156 708024 42208 708076
rect 43168 708024 43220 708076
rect 673276 707548 673328 707600
rect 676036 707548 676088 707600
rect 42156 707208 42208 707260
rect 44364 707208 44416 707260
rect 673644 707140 673696 707192
rect 676036 707140 676088 707192
rect 42156 706732 42208 706784
rect 42524 706732 42576 706784
rect 673920 706732 673972 706784
rect 676036 706732 676088 706784
rect 42064 704216 42116 704268
rect 43076 704216 43128 704268
rect 670148 703808 670200 703860
rect 676036 703808 676088 703860
rect 42156 703536 42208 703588
rect 42984 703536 43036 703588
rect 42432 702992 42484 703044
rect 42064 702856 42116 702908
rect 42248 702516 42300 702568
rect 42064 702244 42116 702296
rect 42156 700408 42208 700460
rect 42432 700408 42484 700460
rect 42156 699864 42208 699916
rect 42892 699864 42944 699916
rect 671896 698164 671948 698216
rect 675392 698164 675444 698216
rect 674656 694152 674708 694204
rect 675484 694152 675536 694204
rect 673276 692928 673328 692980
rect 675484 692928 675536 692980
rect 35716 692044 35768 692096
rect 44916 692044 44968 692096
rect 672632 690412 672684 690464
rect 675392 690412 675444 690464
rect 673920 690004 673972 690056
rect 675392 690004 675444 690056
rect 674380 689324 674432 689376
rect 675484 689324 675536 689376
rect 658924 689256 658976 689308
rect 674748 689256 674800 689308
rect 49056 688644 49108 688696
rect 62120 688644 62172 688696
rect 673000 688644 673052 688696
rect 675392 688644 675444 688696
rect 35808 687896 35860 687948
rect 47676 687896 47728 687948
rect 35624 687760 35676 687812
rect 50436 687760 50488 687812
rect 673368 687284 673420 687336
rect 675392 687284 675444 687336
rect 674748 687012 674800 687064
rect 675484 687012 675536 687064
rect 670608 686060 670660 686112
rect 675392 686060 675444 686112
rect 672540 684224 672592 684276
rect 675392 684224 675444 684276
rect 651840 683136 651892 683188
rect 658924 683136 658976 683188
rect 40684 683000 40736 683052
rect 41696 683000 41748 683052
rect 40776 681776 40828 681828
rect 41696 681776 41748 681828
rect 30472 676812 30524 676864
rect 51724 676812 51776 676864
rect 47676 674840 47728 674892
rect 62120 674840 62172 674892
rect 35164 672800 35216 672852
rect 42432 672800 42484 672852
rect 31024 672732 31076 672784
rect 41880 672732 41932 672784
rect 40776 670964 40828 671016
rect 42064 670964 42116 671016
rect 40684 670896 40736 670948
rect 42708 670896 42760 670948
rect 672724 670896 672776 670948
rect 676220 670896 676272 670948
rect 665824 670760 665876 670812
rect 676036 670760 676088 670812
rect 41880 670556 41932 670608
rect 41972 670556 42024 670608
rect 42984 670556 43036 670608
rect 41880 670352 41932 670404
rect 672264 669672 672316 669724
rect 676220 669672 676272 669724
rect 672908 669536 672960 669588
rect 676128 669536 676180 669588
rect 661776 669400 661828 669452
rect 676312 669400 676364 669452
rect 42708 669332 42760 669384
rect 46204 669332 46256 669384
rect 651564 669332 651616 669384
rect 659016 669332 659068 669384
rect 674196 668856 674248 668908
rect 676036 668856 676088 668908
rect 42984 668720 43036 668772
rect 42892 668516 42944 668568
rect 673460 668652 673512 668704
rect 676220 668652 676272 668704
rect 42156 667836 42208 667888
rect 42708 667836 42760 667888
rect 42708 667700 42760 667752
rect 44456 667904 44508 667956
rect 672724 667904 672776 667956
rect 676036 667904 676088 667956
rect 673552 667836 673604 667888
rect 676220 667836 676272 667888
rect 42156 666680 42208 666732
rect 42708 666680 42760 666732
rect 672264 666544 672316 666596
rect 676220 666544 676272 666596
rect 42708 666476 42760 666528
rect 43076 666476 43128 666528
rect 674472 666476 674524 666528
rect 676036 666476 676088 666528
rect 671988 665320 672040 665372
rect 676220 665320 676272 665372
rect 674288 665252 674340 665304
rect 676036 665252 676088 665304
rect 673828 664980 673880 665032
rect 676220 664980 676272 665032
rect 42156 664164 42208 664216
rect 42708 664164 42760 664216
rect 672356 663960 672408 664012
rect 676220 663960 676272 664012
rect 673184 663756 673236 663808
rect 676220 663756 676272 663808
rect 43536 662396 43588 662448
rect 62120 662396 62172 662448
rect 673736 662328 673788 662380
rect 676036 662328 676088 662380
rect 674564 661580 674616 661632
rect 676036 661580 676088 661632
rect 673092 661104 673144 661156
rect 676220 661104 676272 661156
rect 42156 661036 42208 661088
rect 43076 661036 43128 661088
rect 42156 659676 42208 659728
rect 42892 659676 42944 659728
rect 42156 658996 42208 659048
rect 42708 658996 42760 659048
rect 42892 658248 42944 658300
rect 44364 658248 44416 658300
rect 42156 657228 42208 657280
rect 42524 657228 42576 657280
rect 651564 656888 651616 656940
rect 663064 656888 663116 656940
rect 42156 656820 42208 656872
rect 42892 656820 42944 656872
rect 42156 656140 42208 656192
rect 42340 656140 42392 656192
rect 671988 652740 672040 652792
rect 675392 652740 675444 652792
rect 54484 650020 54536 650072
rect 62120 650020 62172 650072
rect 674564 649816 674616 649868
rect 675392 649816 675444 649868
rect 673184 647708 673236 647760
rect 675484 647708 675536 647760
rect 672908 645532 672960 645584
rect 675392 645532 675444 645584
rect 674288 644784 674340 644836
rect 675392 644784 675444 644836
rect 35808 644580 35860 644632
rect 47676 644580 47728 644632
rect 35624 644512 35676 644564
rect 49056 644512 49108 644564
rect 659016 643696 659068 643748
rect 674472 643696 674524 643748
rect 673092 643356 673144 643408
rect 675392 643356 675444 643408
rect 651564 643084 651616 643136
rect 668676 643084 668728 643136
rect 674472 641860 674524 641912
rect 675392 641860 675444 641912
rect 674012 639072 674064 639124
rect 675392 639072 675444 639124
rect 47676 636216 47728 636268
rect 62120 636216 62172 636268
rect 32404 629892 32456 629944
rect 41788 629892 41840 629944
rect 651564 629280 651616 629332
rect 661776 629280 661828 629332
rect 33784 628532 33836 628584
rect 42524 628532 42576 628584
rect 41788 627376 41840 627428
rect 41788 627036 41840 627088
rect 42984 626560 43036 626612
rect 44824 626560 44876 626612
rect 672816 625472 672868 625524
rect 676128 625472 676180 625524
rect 664536 625336 664588 625388
rect 676220 625336 676272 625388
rect 42156 625268 42208 625320
rect 42524 625268 42576 625320
rect 660304 625132 660356 625184
rect 676220 625132 676272 625184
rect 42156 624656 42208 624708
rect 42984 624656 43036 624708
rect 674196 624316 674248 624368
rect 676036 624316 676088 624368
rect 42524 623840 42576 623892
rect 672356 623840 672408 623892
rect 676036 623840 676088 623892
rect 42156 623432 42208 623484
rect 43628 623772 43680 623824
rect 62120 623772 62172 623824
rect 672448 623772 672500 623824
rect 676220 623772 676272 623824
rect 672264 622684 672316 622736
rect 676036 622684 676088 622736
rect 672724 622548 672776 622600
rect 676128 622548 676180 622600
rect 672264 622412 672316 622464
rect 676220 622412 676272 622464
rect 673644 622208 673696 622260
rect 676036 622208 676088 622260
rect 42064 622140 42116 622192
rect 42524 622140 42576 622192
rect 42524 622004 42576 622056
rect 42800 622004 42852 622056
rect 671896 621256 671948 621308
rect 676220 621256 676272 621308
rect 670608 621120 670660 621172
rect 676036 621120 676088 621172
rect 42064 620780 42116 620832
rect 43076 620780 43128 620832
rect 42064 620304 42116 620356
rect 42524 620304 42576 620356
rect 42524 620168 42576 620220
rect 42892 620168 42944 620220
rect 672632 619896 672684 619948
rect 676220 619896 676272 619948
rect 672540 619760 672592 619812
rect 676036 619760 676088 619812
rect 674656 619148 674708 619200
rect 676220 619148 676272 619200
rect 42156 617856 42208 617908
rect 42524 617856 42576 617908
rect 42524 617720 42576 617772
rect 44456 618264 44508 618316
rect 674380 617788 674432 617840
rect 676036 617788 676088 617840
rect 42064 617108 42116 617160
rect 42524 617108 42576 617160
rect 673368 617040 673420 617092
rect 676128 617040 676180 617092
rect 673920 616972 673972 617024
rect 676036 616972 676088 617024
rect 652392 616836 652444 616888
rect 659016 616836 659068 616888
rect 673276 616836 673328 616888
rect 676220 616836 676272 616888
rect 673000 615476 673052 615528
rect 676220 615476 676272 615528
rect 672724 614116 672776 614168
rect 683120 614116 683172 614168
rect 42156 613436 42208 613488
rect 42524 613436 42576 613488
rect 675208 610648 675260 610700
rect 675668 610648 675720 610700
rect 44824 609968 44876 610020
rect 62120 609968 62172 610020
rect 673368 607588 673420 607640
rect 675392 607588 675444 607640
rect 674472 604732 674524 604784
rect 675392 604732 675444 604784
rect 674656 604324 674708 604376
rect 675392 604324 675444 604376
rect 673828 603440 673880 603492
rect 675484 603440 675536 603492
rect 651564 603100 651616 603152
rect 660304 603100 660356 603152
rect 673276 603032 673328 603084
rect 675392 603032 675444 603084
rect 35808 601672 35860 601724
rect 47676 601672 47728 601724
rect 43628 601604 43680 601656
rect 35808 601536 35860 601588
rect 35716 601468 35768 601520
rect 44364 601468 44416 601520
rect 35808 601332 35860 601384
rect 54484 601332 54536 601384
rect 674380 599768 674432 599820
rect 675484 599768 675536 599820
rect 659016 599564 659068 599616
rect 674748 599156 674800 599208
rect 674196 598408 674248 598460
rect 675484 598408 675536 598460
rect 46204 597524 46256 597576
rect 62120 597524 62172 597576
rect 674748 596844 674800 596896
rect 675392 596844 675444 596896
rect 672632 595280 672684 595332
rect 675392 595280 675444 595332
rect 672816 593376 672868 593428
rect 675484 593376 675536 593428
rect 651564 590656 651616 590708
rect 664444 590656 664496 590708
rect 41512 589908 41564 589960
rect 54484 589908 54536 589960
rect 33784 585828 33836 585880
rect 41880 585828 41932 585880
rect 32404 585760 32456 585812
rect 41788 585760 41840 585812
rect 40776 584604 40828 584656
rect 42432 584604 42484 584656
rect 40684 584536 40736 584588
rect 41972 584536 42024 584588
rect 41880 584196 41932 584248
rect 42064 584196 42116 584248
rect 42708 584196 42760 584248
rect 41880 583924 41932 583976
rect 47768 583720 47820 583772
rect 62120 583720 62172 583772
rect 42892 581612 42944 581664
rect 43076 581612 43128 581664
rect 42156 581272 42208 581324
rect 43536 581272 43588 581324
rect 652024 581000 652076 581052
rect 676036 581000 676088 581052
rect 672448 580048 672500 580100
rect 676220 580048 676272 580100
rect 671436 579912 671488 579964
rect 676128 579912 676180 579964
rect 658924 579776 658976 579828
rect 676036 579776 676088 579828
rect 42892 579640 42944 579692
rect 44456 579640 44508 579692
rect 673736 579232 673788 579284
rect 676220 579232 676272 579284
rect 673920 578552 673972 578604
rect 676036 578552 676088 578604
rect 42156 578416 42208 578468
rect 42892 578416 42944 578468
rect 43168 578212 43220 578264
rect 44364 578212 44416 578264
rect 672356 578212 672408 578264
rect 676220 578212 676272 578264
rect 673644 577396 673696 577448
rect 676036 577396 676088 577448
rect 672264 576988 672316 577040
rect 676220 576988 676272 577040
rect 42156 576920 42208 576972
rect 43168 576920 43220 576972
rect 672540 576920 672592 576972
rect 676036 576920 676088 576972
rect 651564 576852 651616 576904
rect 659016 576852 659068 576904
rect 672448 576852 672500 576904
rect 676128 576852 676180 576904
rect 42432 576308 42484 576360
rect 42984 576308 43036 576360
rect 671988 575560 672040 575612
rect 676220 575560 676272 575612
rect 674564 575356 674616 575408
rect 676036 575356 676088 575408
rect 42156 574540 42208 574592
rect 42432 574540 42484 574592
rect 674012 574540 674064 574592
rect 676036 574540 676088 574592
rect 672908 574200 672960 574252
rect 676220 574200 676272 574252
rect 42156 574064 42208 574116
rect 42340 574064 42392 574116
rect 42156 573452 42208 573504
rect 43076 573452 43128 573504
rect 674288 571684 674340 571736
rect 676036 571684 676088 571736
rect 42340 571480 42392 571532
rect 673184 571480 673236 571532
rect 676220 571480 676272 571532
rect 42064 570868 42116 570920
rect 43536 571344 43588 571396
rect 62120 571344 62172 571396
rect 673092 569916 673144 569968
rect 676220 569916 676272 569968
rect 42064 569576 42116 569628
rect 42708 569576 42760 569628
rect 668584 568556 668636 568608
rect 683120 568556 683172 568608
rect 652116 563048 652168 563100
rect 658924 563048 658976 563100
rect 35624 562300 35676 562352
rect 43536 562300 43588 562352
rect 671988 561892 672040 561944
rect 675392 561892 675444 561944
rect 673092 560192 673144 560244
rect 675208 560192 675260 560244
rect 675208 559648 675260 559700
rect 675392 559648 675444 559700
rect 35716 558288 35768 558340
rect 46204 558288 46256 558340
rect 35808 558152 35860 558204
rect 47768 558152 47820 558204
rect 47676 557540 47728 557592
rect 62120 557540 62172 557592
rect 673184 557540 673236 557592
rect 675484 557540 675536 557592
rect 674288 555228 674340 555280
rect 675392 555228 675444 555280
rect 673000 554752 673052 554804
rect 675300 554752 675352 554804
rect 674564 554140 674616 554192
rect 675300 554140 675352 554192
rect 658924 554004 658976 554056
rect 675300 554004 675352 554056
rect 672908 553460 672960 553512
rect 675392 553460 675444 553512
rect 651564 550604 651616 550656
rect 661684 550604 661736 550656
rect 674932 549176 674984 549228
rect 675300 549176 675352 549228
rect 674748 548292 674800 548344
rect 675300 548292 675352 548344
rect 31668 547136 31720 547188
rect 35808 547136 35860 547188
rect 55864 547136 55916 547188
rect 31024 542988 31076 543040
rect 41788 542988 41840 543040
rect 40684 542308 40736 542360
rect 42708 542308 42760 542360
rect 41788 541016 41840 541068
rect 41788 540744 41840 540796
rect 43168 539588 43220 539640
rect 44824 539588 44876 539640
rect 42064 538908 42116 538960
rect 42708 538908 42760 538960
rect 44548 538228 44600 538280
rect 42156 538160 42208 538212
rect 43168 538160 43220 538212
rect 42064 537072 42116 537124
rect 42616 536800 42668 536852
rect 44456 536800 44508 536852
rect 651564 536800 651616 536852
rect 664536 536800 664588 536852
rect 42616 535984 42668 536036
rect 42156 535780 42208 535832
rect 668676 535712 668728 535764
rect 676220 535712 676272 535764
rect 663064 535576 663116 535628
rect 676036 535576 676088 535628
rect 42064 535236 42116 535288
rect 43076 535236 43128 535288
rect 673736 534896 673788 534948
rect 676036 534896 676088 534948
rect 661776 534216 661828 534268
rect 676220 534216 676272 534268
rect 673920 534080 673972 534132
rect 676036 534080 676088 534132
rect 42156 533944 42208 533996
rect 42616 533944 42668 533996
rect 672448 532856 672500 532908
rect 676220 532856 676272 532908
rect 51816 532720 51868 532772
rect 62120 532720 62172 532772
rect 42156 531428 42208 531480
rect 42616 531428 42668 531480
rect 42616 531292 42668 531344
rect 42984 531292 43036 531344
rect 672540 531292 672592 531344
rect 676220 531292 676272 531344
rect 674472 530408 674524 530460
rect 676036 530408 676088 530460
rect 42156 530068 42208 530120
rect 42616 530068 42668 530120
rect 672632 530000 672684 530052
rect 676220 530000 676272 530052
rect 42156 529456 42208 529508
rect 42340 529592 42392 529644
rect 674656 528844 674708 528896
rect 676036 528844 676088 528896
rect 673368 528776 673420 528828
rect 676220 528776 676272 528828
rect 672816 528640 672868 528692
rect 676128 528640 676180 528692
rect 42984 528572 43036 528624
rect 44364 528572 44416 528624
rect 673828 528368 673880 528420
rect 676036 528368 676088 528420
rect 42064 527212 42116 527264
rect 42340 527212 42392 527264
rect 42156 527144 42208 527196
rect 42984 527144 43036 527196
rect 674380 526736 674432 526788
rect 676036 526736 676088 526788
rect 42156 526600 42208 526652
rect 42616 526600 42668 526652
rect 674196 526328 674248 526380
rect 676036 526328 676088 526380
rect 673276 525920 673328 525972
rect 676220 525920 676272 525972
rect 668676 524424 668728 524476
rect 683120 524424 683172 524476
rect 651564 522996 651616 523048
rect 663156 522996 663208 523048
rect 676128 520956 676180 521008
rect 683304 520956 683356 521008
rect 676036 520888 676088 520940
rect 683672 520888 683724 520940
rect 40684 518916 40736 518968
rect 62120 518916 62172 518968
rect 651564 510620 651616 510672
rect 665824 510620 665876 510672
rect 49056 506472 49108 506524
rect 62120 506472 62172 506524
rect 40868 497428 40920 497480
rect 62764 497428 62816 497480
rect 651564 496816 651616 496868
rect 658924 496816 658976 496868
rect 53196 492668 53248 492720
rect 62120 492668 62172 492720
rect 664444 491648 664496 491700
rect 675944 491648 675996 491700
rect 660304 491512 660356 491564
rect 676036 491512 676088 491564
rect 659016 491376 659068 491428
rect 676036 491376 676088 491428
rect 675944 489268 675996 489320
rect 677324 489268 677376 489320
rect 675944 488588 675996 488640
rect 676128 488588 676180 488640
rect 675944 488452 675996 488504
rect 677508 488452 677560 488504
rect 674932 488316 674984 488368
rect 675944 488316 675996 488368
rect 675852 487976 675904 488028
rect 677232 487976 677284 488028
rect 674288 486004 674340 486056
rect 675944 486004 675996 486056
rect 673092 484576 673144 484628
rect 675944 484576 675996 484628
rect 651564 484372 651616 484424
rect 660396 484372 660448 484424
rect 671988 484372 672040 484424
rect 675852 484372 675904 484424
rect 674564 483556 674616 483608
rect 675944 483556 675996 483608
rect 673184 483080 673236 483132
rect 675944 483080 675996 483132
rect 673000 481856 673052 481908
rect 675852 481856 675904 481908
rect 672908 481720 672960 481772
rect 675944 481720 675996 481772
rect 50528 480224 50580 480276
rect 62120 480224 62172 480276
rect 674196 480224 674248 480276
rect 678980 480224 679032 480276
rect 651656 470568 651708 470620
rect 664444 470568 664496 470620
rect 55956 466420 56008 466472
rect 62120 466420 62172 466472
rect 651564 456764 651616 456816
rect 671528 456764 671580 456816
rect 50436 454044 50488 454096
rect 62120 454044 62172 454096
rect 651564 444388 651616 444440
rect 659016 444388 659068 444440
rect 44916 440240 44968 440292
rect 62120 440240 62172 440292
rect 40684 432556 40736 432608
rect 41788 432556 41840 432608
rect 43352 430584 43404 430636
rect 51816 430584 51868 430636
rect 651564 430584 651616 430636
rect 660304 430584 660356 430636
rect 40868 430108 40920 430160
rect 41788 430108 41840 430160
rect 54576 427796 54628 427848
rect 62120 427796 62172 427848
rect 40776 425688 40828 425740
rect 41788 425688 41840 425740
rect 41788 419432 41840 419484
rect 44824 419432 44876 419484
rect 651564 416780 651616 416832
rect 663064 416780 663116 416832
rect 51816 415420 51868 415472
rect 62120 415420 62172 415472
rect 32404 414808 32456 414860
rect 41880 414808 41932 414860
rect 31024 414672 31076 414724
rect 42524 414672 42576 414724
rect 41880 413380 41932 413432
rect 41880 413108 41932 413160
rect 42156 410660 42208 410712
rect 47676 410660 47728 410712
rect 42064 408144 42116 408196
rect 43076 408144 43128 408196
rect 42156 407600 42208 407652
rect 42524 407600 42576 407652
rect 42064 406784 42116 406836
rect 44456 406784 44508 406836
rect 652024 404336 652076 404388
rect 661776 404336 661828 404388
rect 42156 403860 42208 403912
rect 42800 403860 42852 403912
rect 664536 403384 664588 403436
rect 676220 403384 676272 403436
rect 663156 403248 663208 403300
rect 676220 403248 676272 403300
rect 661684 403112 661736 403164
rect 676404 403112 676456 403164
rect 42156 402908 42208 402960
rect 44364 402908 44416 402960
rect 43536 401616 43588 401668
rect 62120 401616 62172 401668
rect 673184 401616 673236 401668
rect 676220 401616 676272 401668
rect 673368 400256 673420 400308
rect 676220 400256 676272 400308
rect 673276 400188 673328 400240
rect 676128 400188 676180 400240
rect 674748 399576 674800 399628
rect 676220 399576 676272 399628
rect 675024 398216 675076 398268
rect 676036 398216 676088 398268
rect 674932 397468 674984 397520
rect 676036 397468 676088 397520
rect 674656 394000 674708 394052
rect 676036 394000 676088 394052
rect 673092 393320 673144 393372
rect 676220 393320 676272 393372
rect 670240 391960 670292 392012
rect 683120 391960 683172 392012
rect 651564 390532 651616 390584
rect 671436 390532 671488 390584
rect 43628 389172 43680 389224
rect 62120 389172 62172 389224
rect 35716 387744 35768 387796
rect 44272 387744 44324 387796
rect 675208 387744 675260 387796
rect 676956 387744 677008 387796
rect 675116 387676 675168 387728
rect 676496 387676 676548 387728
rect 35808 387608 35860 387660
rect 50528 387608 50580 387660
rect 675300 387608 675352 387660
rect 678244 387608 678296 387660
rect 35624 387472 35676 387524
rect 53196 387472 53248 387524
rect 35808 387336 35860 387388
rect 55956 387336 56008 387388
rect 675024 386112 675076 386164
rect 675392 386112 675444 386164
rect 675024 385976 675076 386028
rect 675300 385976 675352 386028
rect 675208 385772 675260 385824
rect 675392 385568 675444 385620
rect 675024 383868 675076 383920
rect 675300 383868 675352 383920
rect 674932 383052 674984 383104
rect 675392 383052 675444 383104
rect 675116 381080 675168 381132
rect 675392 381080 675444 381132
rect 651564 378156 651616 378208
rect 664536 378156 664588 378208
rect 673092 376728 673144 376780
rect 675300 376728 675352 376780
rect 674656 376660 674708 376712
rect 675484 376660 675536 376712
rect 35808 375980 35860 376032
rect 41512 375980 41564 376032
rect 53196 375980 53248 376032
rect 47676 375368 47728 375420
rect 62120 375368 62172 375420
rect 31024 371832 31076 371884
rect 42340 371832 42392 371884
rect 40868 371220 40920 371272
rect 42708 371220 42760 371272
rect 40684 370540 40736 370592
rect 41788 370540 41840 370592
rect 42156 369656 42208 369708
rect 42340 369656 42392 369708
rect 42156 368092 42208 368144
rect 42708 368092 42760 368144
rect 42156 366800 42208 366852
rect 42708 366800 42760 366852
rect 42156 364964 42208 365016
rect 43076 364964 43128 365016
rect 652024 364352 652076 364404
rect 674380 364352 674432 364404
rect 42156 364284 42208 364336
rect 44548 364284 44600 364336
rect 42708 364216 42760 364268
rect 49056 364216 49108 364268
rect 51908 362924 51960 362976
rect 62120 362924 62172 362976
rect 42064 360680 42116 360732
rect 42984 360680 43036 360732
rect 42156 359456 42208 359508
rect 42892 359456 42944 359508
rect 665824 357824 665876 357876
rect 675944 357824 675996 357876
rect 660396 357688 660448 357740
rect 676036 357688 676088 357740
rect 658924 357552 658976 357604
rect 675852 357552 675904 357604
rect 673184 357484 673236 357536
rect 676036 357484 676088 357536
rect 674656 357008 674708 357060
rect 676036 357008 676088 357060
rect 673276 356668 673328 356720
rect 676036 356668 676088 356720
rect 674472 356192 674524 356244
rect 676036 356192 676088 356244
rect 42156 355988 42208 356040
rect 44456 355988 44508 356040
rect 673368 355852 673420 355904
rect 676036 355852 676088 355904
rect 672908 355376 672960 355428
rect 676036 355376 676088 355428
rect 673276 354560 673328 354612
rect 676036 354560 676088 354612
rect 676036 351024 676088 351076
rect 676772 351024 676824 351076
rect 673368 350888 673420 350940
rect 676036 350888 676088 350940
rect 651564 350548 651616 350600
rect 674104 350548 674156 350600
rect 674564 350548 674616 350600
rect 676036 350548 676088 350600
rect 673184 349256 673236 349308
rect 676036 349256 676088 349308
rect 46204 349120 46256 349172
rect 62120 349120 62172 349172
rect 673092 348848 673144 348900
rect 676036 348848 676088 348900
rect 672816 346400 672868 346452
rect 676036 346400 676088 346452
rect 35716 344428 35768 344480
rect 44916 344428 44968 344480
rect 35808 344292 35860 344344
rect 51816 344292 51868 344344
rect 35624 344156 35676 344208
rect 54576 344156 54628 344208
rect 651656 338104 651708 338156
rect 673000 338104 673052 338156
rect 44916 336744 44968 336796
rect 62120 336744 62172 336796
rect 674840 336676 674892 336728
rect 675392 336676 675444 336728
rect 673368 336540 673420 336592
rect 675392 336540 675444 336592
rect 30380 333208 30432 333260
rect 49056 333208 49108 333260
rect 673184 332596 673236 332648
rect 675392 332596 675444 332648
rect 673092 331576 673144 331628
rect 675392 331576 675444 331628
rect 674564 330556 674616 330608
rect 675392 330556 675444 330608
rect 675116 327632 675168 327684
rect 675484 327632 675536 327684
rect 42064 326748 42116 326800
rect 43076 326748 43128 326800
rect 675760 325796 675812 325848
rect 675760 325592 675812 325644
rect 651564 324300 651616 324352
rect 671620 324300 671672 324352
rect 42156 323280 42208 323332
rect 42616 323280 42668 323332
rect 43720 322940 43772 322992
rect 62120 322940 62172 322992
rect 42064 322872 42116 322924
rect 42984 322872 43036 322924
rect 42616 321512 42668 321564
rect 50436 321512 50488 321564
rect 42156 321444 42208 321496
rect 42892 321444 42944 321496
rect 42156 319948 42208 320000
rect 44548 319948 44600 320000
rect 42156 316684 42208 316736
rect 44456 316684 44508 316736
rect 671528 313488 671580 313540
rect 676220 313488 676272 313540
rect 664444 313352 664496 313404
rect 676036 313352 676088 313404
rect 674656 312468 674708 312520
rect 676036 312468 676088 312520
rect 659016 311992 659068 312044
rect 676220 311992 676272 312044
rect 674748 311856 674800 311908
rect 676220 311856 676272 311908
rect 674472 311652 674524 311704
rect 676036 311652 676088 311704
rect 674656 311040 674708 311092
rect 676220 311040 676272 311092
rect 672908 310632 672960 310684
rect 676220 310632 676272 310684
rect 55956 310496 56008 310548
rect 62120 310496 62172 310548
rect 652392 310496 652444 310548
rect 672908 310496 672960 310548
rect 673276 309408 673328 309460
rect 676220 309408 676272 309460
rect 673368 309340 673420 309392
rect 676128 309340 676180 309392
rect 673368 309204 673420 309256
rect 676312 309204 676364 309256
rect 41972 307028 42024 307080
rect 51908 307028 51960 307080
rect 674564 304512 674616 304564
rect 676220 304512 676272 304564
rect 673184 303696 673236 303748
rect 676220 303696 676272 303748
rect 673092 303628 673144 303680
rect 676128 303628 676180 303680
rect 674288 302200 674340 302252
rect 683120 302200 683172 302252
rect 42064 300908 42116 300960
rect 47676 300908 47728 300960
rect 43628 298120 43680 298172
rect 62120 298120 62172 298172
rect 675116 298120 675168 298172
rect 676404 298120 676456 298172
rect 675760 298052 675812 298104
rect 679716 298052 679768 298104
rect 675208 297984 675260 298036
rect 676864 297984 676916 298036
rect 675760 296148 675812 296200
rect 675760 295944 675812 295996
rect 675208 295196 675260 295248
rect 675392 295196 675444 295248
rect 675116 294040 675168 294092
rect 675024 293972 675076 294024
rect 675024 291728 675076 291780
rect 675392 291728 675444 291780
rect 674564 291048 674616 291100
rect 675392 291048 675444 291100
rect 673092 287920 673144 287972
rect 675392 287920 675444 287972
rect 673184 286560 673236 286612
rect 675392 286560 675444 286612
rect 46296 284316 46348 284368
rect 62120 284316 62172 284368
rect 651564 284316 651616 284368
rect 671528 284316 671580 284368
rect 42156 283568 42208 283620
rect 42432 283568 42484 283620
rect 42156 281052 42208 281104
rect 43536 281052 43588 281104
rect 42156 279828 42208 279880
rect 42984 279828 43036 279880
rect 42064 278604 42116 278656
rect 44180 278604 44232 278656
rect 43444 278128 43496 278180
rect 647332 278128 647384 278180
rect 53196 278060 53248 278112
rect 659660 278060 659712 278112
rect 44824 277992 44876 278044
rect 658280 277992 658332 278044
rect 339408 277584 339460 277636
rect 454776 277584 454828 277636
rect 389088 277516 389140 277568
rect 587164 277516 587216 277568
rect 394424 277448 394476 277500
rect 601424 277448 601476 277500
rect 398380 277380 398432 277432
rect 612004 277380 612056 277432
rect 351828 277312 351880 277364
rect 489092 277312 489144 277364
rect 354588 277244 354640 277296
rect 496176 277244 496228 277296
rect 357348 277176 357400 277228
rect 503260 277176 503312 277228
rect 42156 277108 42208 277160
rect 42892 277108 42944 277160
rect 360108 277108 360160 277160
rect 510344 277108 510396 277160
rect 384948 277040 385000 277092
rect 574192 277040 574244 277092
rect 382004 276972 382056 277024
rect 567108 276972 567160 277024
rect 384580 276904 384632 276956
rect 575388 276904 575440 276956
rect 387248 276836 387300 276888
rect 582472 276836 582524 276888
rect 391756 276768 391808 276820
rect 593144 276768 593196 276820
rect 394608 276700 394660 276752
rect 600228 276700 600280 276752
rect 408408 276632 408460 276684
rect 638040 276632 638092 276684
rect 335268 276564 335320 276616
rect 444196 276564 444248 276616
rect 333888 276496 333940 276548
rect 439412 276496 439464 276548
rect 330760 276428 330812 276480
rect 432328 276428 432380 276480
rect 329748 276360 329800 276412
rect 428832 276360 428884 276412
rect 326988 276292 327040 276344
rect 421656 276292 421708 276344
rect 405648 276020 405700 276072
rect 142712 275952 142764 276004
rect 181168 275952 181220 276004
rect 185216 275952 185268 276004
rect 217324 275952 217376 276004
rect 346124 275952 346176 276004
rect 473728 275952 473780 276004
rect 629760 275952 629812 276004
rect 153292 275884 153344 275936
rect 204904 275884 204956 275936
rect 348792 275884 348844 275936
rect 480812 275884 480864 275936
rect 481180 275884 481232 275936
rect 581276 275884 581328 275936
rect 167552 275816 167604 275868
rect 223212 275816 223264 275868
rect 343364 275816 343416 275868
rect 466644 275816 466696 275868
rect 466736 275816 466788 275868
rect 603724 275816 603776 275868
rect 160468 275748 160520 275800
rect 220636 275748 220688 275800
rect 250260 275748 250312 275800
rect 251180 275748 251232 275800
rect 258540 275748 258592 275800
rect 264612 275748 264664 275800
rect 354496 275748 354548 275800
rect 494980 275748 495032 275800
rect 495072 275748 495124 275800
rect 588360 275748 588412 275800
rect 107200 275680 107252 275732
rect 208400 275680 208452 275732
rect 213644 275680 213696 275732
rect 223028 275680 223080 275732
rect 251456 275680 251508 275732
rect 252376 275680 252428 275732
rect 357256 275680 357308 275732
rect 502064 275680 502116 275732
rect 507860 275680 507912 275732
rect 100116 275612 100168 275664
rect 205824 275612 205876 275664
rect 212448 275612 212500 275664
rect 224960 275612 225012 275664
rect 360016 275612 360068 275664
rect 509148 275612 509200 275664
rect 577688 275680 577740 275732
rect 599032 275680 599084 275732
rect 591948 275612 592000 275664
rect 592040 275612 592092 275664
rect 614396 275612 614448 275664
rect 93032 275544 93084 275596
rect 201408 275544 201460 275596
rect 210056 275544 210108 275596
rect 231768 275544 231820 275596
rect 234896 275544 234948 275596
rect 245660 275544 245712 275596
rect 362316 275544 362368 275596
rect 516232 275544 516284 275596
rect 581644 275544 581696 275596
rect 607312 275544 607364 275596
rect 90640 275476 90692 275528
rect 201684 275476 201736 275528
rect 223120 275476 223172 275528
rect 244280 275476 244332 275528
rect 365444 275476 365496 275528
rect 523408 275476 523460 275528
rect 523592 275476 523644 275528
rect 594708 275476 594760 275528
rect 594800 275476 594852 275528
rect 617984 275476 618036 275528
rect 81256 275408 81308 275460
rect 197820 275408 197872 275460
rect 215944 275408 215996 275460
rect 240048 275408 240100 275460
rect 333796 275408 333848 275460
rect 438216 275408 438268 275460
rect 438860 275408 438912 275460
rect 622676 275408 622728 275460
rect 66996 275340 67048 275392
rect 185584 275340 185636 275392
rect 188804 275340 188856 275392
rect 215852 275340 215904 275392
rect 220728 275340 220780 275392
rect 243360 275340 243412 275392
rect 244372 275340 244424 275392
rect 259368 275340 259420 275392
rect 398840 275340 398892 275392
rect 413376 275340 413428 275392
rect 419540 275340 419592 275392
rect 643928 275340 643980 275392
rect 71780 275272 71832 275324
rect 193864 275272 193916 275324
rect 208860 275272 208912 275324
rect 234620 275272 234672 275324
rect 239588 275272 239640 275324
rect 252928 275272 252980 275324
rect 259736 275272 259788 275324
rect 265072 275272 265124 275324
rect 389272 275272 389324 275324
rect 409880 275272 409932 275324
rect 411168 275272 411220 275324
rect 646320 275272 646372 275324
rect 174636 275204 174688 275256
rect 207020 275204 207072 275256
rect 340604 275204 340656 275256
rect 459560 275204 459612 275256
rect 459744 275204 459796 275256
rect 577780 275204 577832 275256
rect 181720 275136 181772 275188
rect 213184 275136 213236 275188
rect 337844 275136 337896 275188
rect 452476 275136 452528 275188
rect 178132 275068 178184 275120
rect 195980 275068 196032 275120
rect 375932 275068 375984 275120
rect 487896 275068 487948 275120
rect 335176 275000 335228 275052
rect 445300 275000 445352 275052
rect 88340 274932 88392 274984
rect 90364 274932 90416 274984
rect 262128 274932 262180 274984
rect 264980 274932 265032 274984
rect 330668 274932 330720 274984
rect 431132 274932 431184 274984
rect 74080 274864 74132 274916
rect 77208 274864 77260 274916
rect 252652 274864 252704 274916
rect 96620 274796 96672 274848
rect 100024 274796 100076 274848
rect 70584 274660 70636 274712
rect 73804 274660 73856 274712
rect 103704 274660 103756 274712
rect 106924 274660 106976 274712
rect 207756 274660 207808 274712
rect 210608 274660 210660 274712
rect 227812 274660 227864 274712
rect 229928 274660 229980 274712
rect 159272 274592 159324 274644
rect 226892 274592 226944 274644
rect 260932 274864 260984 274916
rect 265440 274864 265492 274916
rect 403440 274864 403492 274916
rect 424048 274864 424100 274916
rect 409144 274796 409196 274848
rect 420552 274796 420604 274848
rect 264428 274728 264480 274780
rect 266728 274728 266780 274780
rect 263232 274660 263284 274712
rect 266452 274660 266504 274712
rect 266820 274660 266872 274712
rect 267740 274660 267792 274712
rect 262404 274592 262456 274644
rect 311164 274592 311216 274644
rect 333060 274592 333112 274644
rect 350448 274592 350500 274644
rect 483204 274592 483256 274644
rect 128544 274524 128596 274576
rect 196716 274524 196768 274576
rect 199476 274524 199528 274576
rect 242072 274524 242124 274576
rect 312452 274524 312504 274576
rect 336556 274524 336608 274576
rect 351736 274524 351788 274576
rect 486700 274524 486752 274576
rect 150992 274456 151044 274508
rect 223764 274456 223816 274508
rect 320824 274456 320876 274508
rect 349620 274456 349672 274508
rect 353208 274456 353260 274508
rect 490288 274456 490340 274508
rect 493324 274456 493376 274508
rect 505652 274456 505704 274508
rect 148600 274388 148652 274440
rect 222752 274388 222804 274440
rect 295984 274388 296036 274440
rect 329472 274388 329524 274440
rect 354404 274388 354456 274440
rect 493784 274388 493836 274440
rect 121368 274320 121420 274372
rect 196624 274320 196676 274372
rect 198280 274320 198332 274372
rect 241612 274320 241664 274372
rect 291016 274320 291068 274372
rect 324780 274320 324832 274372
rect 355968 274320 356020 274372
rect 497372 274320 497424 274372
rect 42156 274252 42208 274304
rect 44548 274252 44600 274304
rect 137928 274252 137980 274304
rect 219624 274252 219676 274304
rect 289084 274252 289136 274304
rect 318800 274252 318852 274304
rect 322204 274252 322256 274304
rect 356704 274252 356756 274304
rect 357164 274252 357216 274304
rect 500868 274252 500920 274304
rect 123760 274184 123812 274236
rect 214104 274184 214156 274236
rect 291108 274184 291160 274236
rect 325976 274184 326028 274236
rect 362776 274184 362828 274236
rect 518624 274184 518676 274236
rect 523684 274184 523736 274236
rect 533988 274184 534040 274236
rect 113180 274116 113232 274168
rect 209964 274116 210016 274168
rect 243176 274116 243228 274168
rect 258632 274116 258684 274168
rect 273168 274116 273220 274168
rect 279792 274116 279844 274168
rect 292488 274116 292540 274168
rect 328276 274116 328328 274168
rect 348976 274116 349028 274168
rect 479340 274116 479392 274168
rect 479524 274116 479576 274168
rect 640432 274116 640484 274168
rect 111984 274048 112036 274100
rect 208952 274048 209004 274100
rect 231400 274048 231452 274100
rect 254308 274048 254360 274100
rect 296444 274048 296496 274100
rect 342444 274048 342496 274100
rect 371056 274048 371108 274100
rect 539876 274048 539928 274100
rect 97724 273980 97776 274032
rect 203616 273980 203668 274032
rect 223028 273980 223080 274032
rect 247224 273980 247276 274032
rect 277308 273980 277360 274032
rect 289268 273980 289320 274032
rect 300768 273980 300820 274032
rect 353116 273980 353168 274032
rect 375656 273980 375708 274032
rect 551744 273980 551796 274032
rect 89536 273912 89588 273964
rect 200488 273912 200540 273964
rect 205364 273912 205416 273964
rect 244556 273912 244608 273964
rect 251180 273912 251232 273964
rect 261484 273912 261536 273964
rect 287704 273912 287756 273964
rect 304632 273912 304684 273964
rect 304724 273912 304776 273964
rect 363788 273912 363840 273964
rect 379428 273912 379480 273964
rect 562416 273912 562468 273964
rect 172244 273844 172296 273896
rect 232044 273844 232096 273896
rect 244280 273844 244332 273896
rect 251364 273844 251416 273896
rect 304264 273844 304316 273896
rect 323584 273844 323636 273896
rect 347688 273844 347740 273896
rect 476120 273844 476172 273896
rect 169852 273776 169904 273828
rect 231032 273776 231084 273828
rect 319444 273776 319496 273828
rect 338948 273776 339000 273828
rect 346216 273776 346268 273828
rect 472532 273776 472584 273828
rect 194692 273708 194744 273760
rect 240140 273708 240192 273760
rect 316684 273708 316736 273760
rect 331864 273708 331916 273760
rect 344560 273708 344612 273760
rect 468944 273708 468996 273760
rect 197084 273640 197136 273692
rect 238024 273640 238076 273692
rect 309784 273640 309836 273692
rect 322388 273640 322440 273692
rect 343456 273640 343508 273692
rect 465448 273640 465500 273692
rect 341892 273572 341944 273624
rect 461860 273572 461912 273624
rect 185584 273504 185636 273556
rect 192484 273504 192536 273556
rect 340696 273504 340748 273556
rect 458364 273504 458416 273556
rect 324964 273436 325016 273488
rect 402796 273436 402848 273488
rect 402888 273436 402940 273488
rect 438860 273436 438912 273488
rect 42064 273300 42116 273352
rect 44456 273300 44508 273352
rect 279424 273232 279476 273284
rect 285772 273232 285824 273284
rect 307024 273232 307076 273284
rect 315304 273232 315356 273284
rect 158076 273164 158128 273216
rect 226340 273164 226392 273216
rect 300124 273164 300176 273216
rect 319996 273164 320048 273216
rect 364248 273164 364300 273216
rect 522212 273164 522264 273216
rect 152188 273096 152240 273148
rect 223672 273096 223724 273148
rect 301504 273096 301556 273148
rect 321192 273096 321244 273148
rect 369768 273096 369820 273148
rect 536380 273096 536432 273148
rect 42156 273028 42208 273080
rect 42708 273028 42760 273080
rect 141516 273028 141568 273080
rect 220820 273028 220872 273080
rect 314476 273028 314528 273080
rect 387432 273028 387484 273080
rect 388444 273028 388496 273080
rect 565912 273028 565964 273080
rect 120264 272960 120316 273012
rect 212724 272960 212776 273012
rect 219532 272960 219584 273012
rect 117872 272892 117924 272944
rect 211988 272892 212040 272944
rect 101312 272824 101364 272876
rect 204812 272824 204864 272876
rect 94228 272756 94280 272808
rect 201592 272756 201644 272808
rect 204168 272756 204220 272808
rect 236736 272892 236788 272944
rect 314292 272960 314344 273012
rect 388628 272960 388680 273012
rect 397276 272960 397328 273012
rect 581644 272960 581696 273012
rect 315856 272892 315908 272944
rect 390928 272892 390980 272944
rect 398932 272892 398984 272944
rect 591948 272892 592000 272944
rect 249984 272824 250036 272876
rect 289176 272824 289228 272876
rect 301136 272824 301188 272876
rect 317236 272824 317288 272876
rect 394516 272824 394568 272876
rect 400312 272824 400364 272876
rect 594800 272824 594852 272876
rect 78864 272688 78916 272740
rect 191104 272688 191156 272740
rect 191196 272688 191248 272740
rect 239220 272756 239272 272808
rect 291844 272756 291896 272808
rect 311716 272756 311768 272808
rect 322664 272756 322716 272808
rect 411812 272756 411864 272808
rect 411904 272756 411956 272808
rect 610808 272756 610860 272808
rect 240048 272688 240100 272740
rect 248604 272688 248656 272740
rect 282828 272688 282880 272740
rect 305828 272688 305880 272740
rect 318616 272688 318668 272740
rect 398012 272688 398064 272740
rect 401968 272688 402020 272740
rect 621480 272688 621532 272740
rect 84752 272620 84804 272672
rect 198924 272620 198976 272672
rect 206560 272620 206612 272672
rect 244372 272620 244424 272672
rect 285588 272620 285640 272672
rect 312912 272620 312964 272672
rect 319996 272620 320048 272672
rect 401600 272620 401652 272672
rect 403256 272620 403308 272672
rect 625068 272620 625120 272672
rect 77208 272552 77260 272604
rect 194692 272552 194744 272604
rect 201776 272552 201828 272604
rect 243176 272552 243228 272604
rect 246764 272552 246816 272604
rect 259644 272552 259696 272604
rect 288348 272552 288400 272604
rect 317696 272552 317748 272604
rect 321376 272552 321428 272604
rect 405188 272552 405240 272604
rect 405556 272552 405608 272604
rect 632152 272552 632204 272604
rect 72976 272484 73028 272536
rect 194784 272484 194836 272536
rect 195888 272484 195940 272536
rect 240968 272484 241020 272536
rect 245568 272484 245620 272536
rect 259736 272484 259788 272536
rect 274180 272484 274232 272536
rect 282184 272484 282236 272536
rect 286876 272484 286928 272536
rect 316500 272484 316552 272536
rect 321468 272484 321520 272536
rect 408684 272484 408736 272536
rect 409788 272484 409840 272536
rect 642732 272484 642784 272536
rect 162768 272416 162820 272468
rect 228824 272416 228876 272468
rect 362684 272416 362736 272468
rect 515128 272416 515180 272468
rect 187608 272348 187660 272400
rect 235264 272348 235316 272400
rect 359924 272348 359976 272400
rect 507952 272348 508004 272400
rect 193496 272280 193548 272332
rect 240232 272280 240284 272332
rect 332508 272280 332560 272332
rect 182916 272212 182968 272264
rect 225604 272212 225656 272264
rect 329104 272212 329156 272264
rect 426440 272212 426492 272264
rect 435364 272280 435416 272332
rect 441804 272280 441856 272332
rect 491300 272280 491352 272332
rect 492220 272280 492272 272332
rect 437020 272212 437072 272264
rect 325608 272144 325660 272196
rect 419356 272144 419408 272196
rect 420184 272144 420236 272196
rect 434720 272144 434772 272196
rect 324136 272076 324188 272128
rect 415768 272076 415820 272128
rect 328368 272008 328420 272060
rect 403440 272008 403492 272060
rect 395804 271940 395856 271992
rect 466736 271940 466788 271992
rect 387064 271872 387116 271924
rect 399208 271872 399260 271924
rect 161572 271804 161624 271856
rect 227996 271804 228048 271856
rect 296536 271804 296588 271856
rect 340144 271804 340196 271856
rect 368112 271804 368164 271856
rect 531596 271804 531648 271856
rect 155684 271736 155736 271788
rect 226156 271736 226208 271788
rect 287796 271736 287848 271788
rect 294052 271736 294104 271788
rect 297824 271736 297876 271788
rect 343640 271736 343692 271788
rect 369492 271736 369544 271788
rect 535184 271736 535236 271788
rect 145012 271668 145064 271720
rect 222292 271668 222344 271720
rect 302148 271668 302200 271720
rect 354312 271668 354364 271720
rect 370780 271668 370832 271720
rect 538772 271668 538824 271720
rect 136824 271600 136876 271652
rect 218244 271600 218296 271652
rect 252928 271600 252980 271652
rect 257436 271600 257488 271652
rect 304816 271600 304868 271652
rect 362592 271600 362644 271652
rect 372160 271600 372212 271652
rect 542268 271600 542320 271652
rect 83556 271532 83608 271584
rect 164884 271532 164936 271584
rect 165160 271532 165212 271584
rect 229284 271532 229336 271584
rect 306288 271532 306340 271584
rect 366088 271532 366140 271584
rect 373816 271532 373868 271584
rect 547052 271532 547104 271584
rect 135628 271464 135680 271516
rect 218704 271464 218756 271516
rect 224960 271464 225012 271516
rect 247316 271464 247368 271516
rect 307576 271464 307628 271516
rect 369308 271464 369360 271516
rect 375288 271464 375340 271516
rect 550548 271464 550600 271516
rect 114284 271396 114336 271448
rect 200856 271396 200908 271448
rect 202972 271396 203024 271448
rect 242992 271396 243044 271448
rect 307484 271396 307536 271448
rect 370872 271396 370924 271448
rect 376576 271396 376628 271448
rect 554136 271396 554188 271448
rect 127348 271328 127400 271380
rect 215484 271328 215536 271380
rect 230204 271328 230256 271380
rect 254032 271328 254084 271380
rect 308956 271328 309008 271380
rect 373264 271328 373316 271380
rect 376484 271328 376536 271380
rect 555240 271328 555292 271380
rect 116676 271260 116728 271312
rect 211252 271260 211304 271312
rect 226616 271260 226668 271312
rect 252744 271260 252796 271312
rect 279976 271260 280028 271312
rect 297548 271260 297600 271312
rect 310336 271260 310388 271312
rect 376760 271260 376812 271312
rect 377956 271260 378008 271312
rect 557632 271260 557684 271312
rect 104900 271192 104952 271244
rect 206284 271192 206336 271244
rect 224224 271192 224276 271244
rect 251272 271192 251324 271244
rect 253848 271192 253900 271244
rect 262312 271192 262364 271244
rect 281356 271192 281408 271244
rect 299940 271192 299992 271244
rect 311716 271192 311768 271244
rect 380348 271192 380400 271244
rect 380624 271192 380676 271244
rect 564716 271192 564768 271244
rect 68192 271124 68244 271176
rect 193220 271124 193272 271176
rect 200580 271124 200632 271176
rect 242164 271124 242216 271176
rect 242256 271124 242308 271176
rect 258264 271124 258316 271176
rect 284024 271124 284076 271176
rect 308220 271124 308272 271176
rect 315304 271124 315356 271176
rect 383844 271124 383896 271176
rect 392584 271124 392636 271176
rect 594340 271124 594392 271176
rect 166356 271056 166408 271108
rect 230204 271056 230256 271108
rect 336004 271056 336056 271108
rect 364984 271056 365036 271108
rect 366824 271056 366876 271108
rect 528100 271056 528152 271108
rect 168656 270988 168708 271040
rect 230664 270988 230716 271040
rect 326344 270988 326396 271040
rect 350724 270988 350776 271040
rect 365536 270988 365588 271040
rect 524512 270988 524564 271040
rect 175832 270920 175884 270972
rect 233332 270920 233384 270972
rect 322296 270920 322348 270972
rect 347228 270920 347280 270972
rect 364156 270920 364208 270972
rect 521016 270920 521068 270972
rect 192300 270852 192352 270904
rect 238852 270852 238904 270904
rect 362868 270852 362920 270904
rect 517428 270852 517480 270904
rect 186412 270784 186464 270836
rect 227628 270784 227680 270836
rect 337936 270784 337988 270836
rect 451280 270784 451332 270836
rect 329656 270716 329708 270768
rect 429936 270716 429988 270768
rect 326896 270648 326948 270700
rect 422852 270648 422904 270700
rect 344284 270580 344336 270632
rect 374368 270580 374420 270632
rect 351644 270512 351696 270564
rect 375932 270512 375984 270564
rect 154488 270444 154540 270496
rect 225328 270444 225380 270496
rect 293868 270444 293920 270496
rect 335360 270444 335412 270496
rect 346768 270444 346820 270496
rect 474740 270444 474792 270496
rect 147588 270376 147640 270428
rect 222660 270376 222712 270428
rect 296076 270376 296128 270428
rect 340880 270376 340932 270428
rect 348056 270376 348108 270428
rect 477500 270376 477552 270428
rect 110788 270308 110840 270360
rect 140780 270308 140832 270360
rect 143908 270308 143960 270360
rect 221280 270308 221332 270360
rect 297916 270308 297968 270360
rect 345020 270308 345072 270360
rect 349068 270308 349120 270360
rect 481640 270308 481692 270360
rect 140688 270240 140740 270292
rect 219992 270240 220044 270292
rect 220636 270240 220688 270292
rect 228456 270240 228508 270292
rect 298744 270240 298796 270292
rect 347780 270240 347832 270292
rect 357532 270240 357584 270292
rect 503720 270240 503772 270292
rect 133788 270172 133840 270224
rect 216956 270172 217008 270224
rect 234620 270172 234672 270224
rect 246212 270172 246264 270224
rect 300400 270172 300452 270224
rect 351920 270172 351972 270224
rect 360200 270172 360252 270224
rect 510620 270172 510672 270224
rect 129556 270104 129608 270156
rect 215668 270104 215720 270156
rect 231768 270104 231820 270156
rect 246672 270104 246724 270156
rect 297456 270104 297508 270156
rect 343824 270104 343876 270156
rect 344008 270104 344060 270156
rect 467840 270104 467892 270156
rect 469312 270104 469364 270156
rect 625160 270104 625212 270156
rect 126888 270036 126940 270088
rect 214656 270036 214708 270088
rect 241428 270036 241480 270088
rect 258080 270036 258132 270088
rect 273352 270036 273404 270088
rect 280160 270036 280212 270088
rect 282736 270036 282788 270088
rect 289820 270036 289872 270088
rect 301412 270036 301464 270088
rect 354680 270036 354732 270088
rect 365628 270036 365680 270088
rect 524604 270036 524656 270088
rect 77116 269968 77168 270020
rect 124220 269968 124272 270020
rect 125508 269968 125560 270020
rect 215024 269968 215076 270020
rect 236092 269968 236144 270020
rect 256424 269968 256476 270020
rect 274732 269968 274784 270020
rect 284300 269968 284352 270020
rect 306012 269968 306064 270020
rect 358820 269968 358872 270020
rect 372252 269968 372304 270020
rect 542360 269968 542412 270020
rect 122748 269900 122800 269952
rect 213276 269900 213328 269952
rect 237196 269900 237248 269952
rect 256884 269900 256936 269952
rect 276020 269900 276072 269952
rect 287060 269900 287112 269952
rect 303252 269900 303304 269952
rect 360292 269900 360344 269952
rect 374368 269900 374420 269952
rect 547880 269900 547932 269952
rect 85948 269832 86000 269884
rect 116492 269832 116544 269884
rect 119068 269832 119120 269884
rect 211896 269832 211948 269884
rect 233700 269832 233752 269884
rect 255596 269832 255648 269884
rect 277860 269832 277912 269884
rect 292580 269832 292632 269884
rect 305920 269832 305972 269884
rect 367100 269832 367152 269884
rect 378048 269832 378100 269884
rect 557724 269832 557776 269884
rect 108948 269764 109000 269816
rect 207940 269764 207992 269816
rect 229928 269764 229980 269816
rect 253388 269764 253440 269816
rect 279148 269764 279200 269816
rect 295340 269764 295392 269816
rect 321928 269764 321980 269816
rect 389272 269764 389324 269816
rect 390008 269764 390060 269816
rect 590660 269764 590712 269816
rect 146208 269628 146260 269680
rect 177580 269628 177632 269680
rect 173808 269560 173860 269612
rect 232872 269696 232924 269748
rect 294788 269696 294840 269748
rect 336740 269696 336792 269748
rect 345112 269696 345164 269748
rect 470600 269696 470652 269748
rect 176936 269492 176988 269544
rect 234160 269628 234212 269680
rect 293408 269628 293460 269680
rect 333980 269628 334032 269680
rect 342444 269628 342496 269680
rect 463700 269628 463752 269680
rect 179328 269560 179380 269612
rect 234620 269560 234672 269612
rect 292120 269560 292172 269612
rect 329840 269560 329892 269612
rect 341064 269560 341116 269612
rect 459652 269560 459704 269612
rect 464712 269560 464764 269612
rect 469220 269560 469272 269612
rect 180708 269492 180760 269544
rect 235540 269492 235592 269544
rect 307760 269492 307812 269544
rect 327080 269492 327132 269544
rect 339776 269492 339828 269544
rect 456800 269492 456852 269544
rect 184848 269424 184900 269476
rect 236920 269424 236972 269476
rect 338396 269424 338448 269476
rect 452660 269424 452712 269476
rect 337108 269356 337160 269408
rect 449900 269356 449952 269408
rect 335728 269288 335780 269340
rect 445760 269288 445812 269340
rect 518992 269288 519044 269340
rect 525800 269288 525852 269340
rect 323584 269220 323636 269272
rect 376944 269220 376996 269272
rect 223212 269084 223264 269136
rect 231124 269084 231176 269136
rect 516140 269084 516192 269136
rect 518900 269084 518952 269136
rect 102508 269016 102560 269068
rect 206192 269016 206244 269068
rect 323216 269016 323268 269068
rect 398840 269016 398892 269068
rect 408684 269016 408736 269068
rect 583760 269016 583812 269068
rect 99288 268948 99340 269000
rect 204444 268948 204496 269000
rect 222108 268948 222160 269000
rect 236644 268948 236696 269000
rect 309048 268948 309100 269000
rect 375380 268948 375432 269000
rect 393136 268948 393188 269000
rect 577688 268948 577740 269000
rect 95424 268880 95476 268932
rect 203524 268880 203576 268932
rect 225420 268880 225472 268932
rect 245292 268880 245344 268932
rect 310428 268880 310480 268932
rect 378140 268880 378192 268932
rect 382188 268880 382240 268932
rect 568580 268880 568632 268932
rect 92388 268812 92440 268864
rect 202144 268812 202196 268864
rect 218336 268812 218388 268864
rect 239312 268812 239364 268864
rect 284852 268812 284904 268864
rect 298100 268812 298152 268864
rect 311808 268812 311860 268864
rect 382280 268812 382332 268864
rect 394608 268812 394660 268864
rect 601700 268812 601752 268864
rect 87144 268744 87196 268796
rect 200396 268744 200448 268796
rect 201408 268744 201460 268796
rect 203064 268744 203116 268796
rect 204904 268744 204956 268796
rect 225788 268744 225840 268796
rect 229008 268744 229060 268796
rect 253756 268744 253808 268796
rect 278688 268744 278740 268796
rect 294144 268744 294196 268796
rect 313004 268744 313056 268796
rect 385224 268744 385276 268796
rect 395436 268744 395488 268796
rect 604460 268744 604512 268796
rect 82728 268676 82780 268728
rect 198556 268676 198608 268728
rect 207020 268676 207072 268728
rect 233792 268676 233844 268728
rect 290924 268676 290976 268728
rect 306380 268676 306432 268728
rect 314384 268676 314436 268728
rect 389180 268676 389232 268728
rect 395896 268676 395948 268728
rect 605840 268676 605892 268728
rect 80060 268608 80112 268660
rect 197268 268608 197320 268660
rect 215208 268608 215260 268660
rect 244188 268608 244240 268660
rect 245660 268608 245712 268660
rect 256056 268608 256108 268660
rect 280528 268608 280580 268660
rect 291200 268608 291252 268660
rect 291476 268608 291528 268660
rect 310520 268608 310572 268660
rect 315672 268608 315724 268660
rect 393320 268608 393372 268660
rect 397184 268608 397236 268660
rect 608600 268608 608652 268660
rect 77668 268540 77720 268592
rect 196532 268540 196584 268592
rect 217140 268540 217192 268592
rect 249340 268540 249392 268592
rect 283012 268540 283064 268592
rect 302424 268540 302476 268592
rect 317052 268540 317104 268592
rect 396080 268540 396132 268592
rect 399852 268540 399904 268592
rect 615684 268540 615736 268592
rect 75828 268472 75880 268524
rect 195428 268472 195480 268524
rect 211344 268472 211396 268524
rect 247132 268472 247184 268524
rect 281448 268472 281500 268524
rect 302240 268472 302292 268524
rect 318340 268472 318392 268524
rect 400220 268472 400272 268524
rect 401140 268472 401192 268524
rect 619640 268472 619692 268524
rect 69388 268404 69440 268456
rect 193680 268404 193732 268456
rect 210608 268404 210660 268456
rect 245752 268404 245804 268456
rect 249708 268404 249760 268456
rect 261392 268404 261444 268456
rect 274272 268404 274324 268456
rect 282920 268404 282972 268456
rect 286784 268404 286836 268456
rect 309140 268404 309192 268456
rect 319720 268404 319772 268456
rect 402980 268404 403032 268456
rect 403900 268404 403952 268456
rect 626540 268404 626592 268456
rect 66168 268336 66220 268388
rect 192392 268336 192444 268388
rect 195980 268336 196032 268388
rect 235080 268336 235132 268388
rect 248328 268336 248380 268388
rect 260932 268336 260984 268388
rect 275652 268336 275704 268388
rect 285864 268336 285916 268388
rect 286232 268336 286284 268388
rect 313280 268336 313332 268388
rect 322388 268336 322440 268388
rect 409972 268336 410024 268388
rect 410432 268336 410484 268388
rect 636200 268336 636252 268388
rect 106188 268268 106240 268320
rect 207480 268268 207532 268320
rect 307668 268268 307720 268320
rect 371240 268268 371292 268320
rect 371884 268268 371936 268320
rect 394700 268268 394752 268320
rect 110328 268200 110380 268252
rect 208860 268200 208912 268252
rect 303712 268200 303764 268252
rect 360384 268200 360436 268252
rect 362960 268200 363012 268252
rect 385132 268200 385184 268252
rect 390468 268200 390520 268252
rect 507860 268200 507912 268252
rect 115848 268132 115900 268184
rect 210608 268132 210660 268184
rect 302332 268132 302384 268184
rect 357440 268132 357492 268184
rect 361488 268132 361540 268184
rect 380900 268132 380952 268184
rect 389180 268132 389232 268184
rect 495072 268132 495124 268184
rect 131028 268064 131080 268116
rect 216864 268064 216916 268116
rect 335360 268064 335412 268116
rect 368480 268064 368532 268116
rect 386512 268064 386564 268116
rect 481180 268064 481232 268116
rect 663064 268064 663116 268116
rect 676220 268064 676272 268116
rect 135168 267996 135220 268048
rect 218152 267996 218204 268048
rect 331128 267996 331180 268048
rect 413928 267996 413980 268048
rect 414020 267996 414072 268048
rect 426624 267996 426676 268048
rect 190368 267928 190420 267980
rect 230480 267928 230532 267980
rect 385132 267928 385184 267980
rect 459744 267928 459796 267980
rect 661776 267928 661828 267980
rect 676220 267928 676272 267980
rect 181168 267860 181220 267912
rect 221740 267860 221792 267912
rect 342168 267860 342220 267912
rect 407120 267860 407172 267912
rect 354680 267792 354732 267844
rect 416780 267792 416832 267844
rect 243360 267724 243412 267776
rect 250720 267724 250772 267776
rect 369676 267724 369728 267776
rect 391940 267724 391992 267776
rect 392032 267724 392084 267776
rect 523592 267724 523644 267776
rect 660304 267724 660356 267776
rect 676128 267724 676180 267776
rect 140780 267656 140832 267708
rect 209688 267656 209740 267708
rect 284944 267656 284996 267708
rect 291844 267656 291896 267708
rect 299204 267656 299256 267708
rect 320824 267656 320876 267708
rect 341984 267656 342036 267708
rect 462320 267656 462372 267708
rect 157248 267588 157300 267640
rect 227076 267588 227128 267640
rect 283196 267588 283248 267640
rect 290924 267588 290976 267640
rect 298284 267588 298336 267640
rect 322296 267588 322348 267640
rect 323676 267588 323728 267640
rect 331128 267588 331180 267640
rect 347320 267588 347372 267640
rect 476304 267588 476356 267640
rect 124220 267520 124272 267572
rect 196348 267520 196400 267572
rect 196716 267520 196768 267572
rect 216404 267520 216456 267572
rect 284484 267520 284536 267572
rect 291476 267520 291528 267572
rect 299664 267520 299716 267572
rect 326344 267520 326396 267572
rect 330852 267520 330904 267572
rect 350356 267520 350408 267572
rect 150348 267452 150400 267504
rect 224408 267452 224460 267504
rect 236736 267452 236788 267504
rect 244464 267452 244516 267504
rect 272064 267452 272116 267504
rect 277400 267452 277452 267504
rect 288532 267452 288584 267504
rect 301504 267452 301556 267504
rect 306380 267452 306432 267504
rect 335360 267452 335412 267504
rect 349988 267452 350040 267504
rect 483388 267520 483440 267572
rect 352656 267452 352708 267504
rect 491392 267452 491444 267504
rect 139308 267384 139360 267436
rect 220360 267384 220412 267436
rect 288072 267384 288124 267436
rect 300124 267384 300176 267436
rect 305000 267384 305052 267436
rect 336004 267384 336056 267436
rect 339316 267384 339368 267436
rect 116492 267316 116544 267368
rect 199936 267316 199988 267368
rect 132408 267248 132460 267300
rect 227628 267316 227680 267368
rect 237288 267316 237340 267368
rect 289452 267316 289504 267368
rect 304264 267316 304316 267368
rect 308588 267316 308640 267368
rect 344284 267316 344336 267368
rect 355324 267384 355376 267436
rect 498200 267384 498252 267436
rect 346400 267316 346452 267368
rect 346860 267316 346912 267368
rect 347688 267316 347740 267368
rect 348240 267316 348292 267368
rect 348976 267316 349028 267368
rect 349528 267316 349580 267368
rect 350448 267316 350500 267368
rect 350908 267316 350960 267368
rect 351736 267316 351788 267368
rect 352196 267316 352248 267368
rect 353208 267316 353260 267368
rect 353576 267316 353628 267368
rect 354404 267316 354456 267368
rect 360660 267316 360712 267368
rect 512000 267316 512052 267368
rect 217692 267248 217744 267300
rect 225604 267248 225656 267300
rect 236000 267248 236052 267300
rect 236644 267248 236696 267300
rect 251088 267248 251140 267300
rect 276940 267248 276992 267300
rect 282736 267248 282788 267300
rect 290740 267248 290792 267300
rect 307760 267248 307812 267300
rect 311256 267248 311308 267300
rect 361488 267248 361540 267300
rect 106924 267180 106976 267232
rect 200764 267180 200816 267232
rect 200856 267180 200908 267232
rect 100024 267112 100076 267164
rect 204352 267112 204404 267164
rect 90364 267044 90416 267096
rect 201224 267044 201276 267096
rect 217324 267180 217376 267232
rect 237748 267180 237800 267232
rect 238024 267180 238076 267232
rect 241796 267180 241848 267232
rect 245292 267180 245344 267232
rect 252468 267180 252520 267232
rect 256608 267180 256660 267232
rect 264060 267180 264112 267232
rect 288992 267180 289044 267232
rect 309784 267180 309836 267232
rect 312544 267180 312596 267232
rect 362960 267248 363012 267300
rect 363328 267248 363380 267300
rect 516140 267248 516192 267300
rect 361856 267180 361908 267232
rect 362684 267180 362736 267232
rect 368020 267180 368072 267232
rect 233148 267112 233200 267164
rect 255136 267112 255188 267164
rect 255228 267112 255280 267164
rect 263600 267112 263652 267164
rect 286324 267112 286376 267164
rect 307024 267112 307076 267164
rect 315212 267112 315264 267164
rect 369676 267112 369728 267164
rect 371332 267180 371384 267232
rect 371884 267112 371936 267164
rect 378784 267180 378836 267232
rect 523684 267180 523736 267232
rect 540980 267112 541032 267164
rect 211068 267044 211120 267096
rect 213184 267044 213236 267096
rect 73804 266976 73856 267028
rect 194140 266976 194192 267028
rect 202420 266976 202472 267028
rect 213736 266976 213788 267028
rect 215852 267044 215904 267096
rect 239128 267044 239180 267096
rect 239312 267044 239364 267096
rect 249800 267044 249852 267096
rect 252376 267044 252428 267096
rect 262220 267044 262272 267096
rect 292580 267044 292632 267096
rect 316684 267044 316736 267096
rect 317880 267044 317932 267096
rect 387064 267044 387116 267096
rect 236460 266976 236512 267028
rect 238668 266976 238720 267028
rect 257344 266976 257396 267028
rect 257988 266976 258040 267028
rect 264520 266976 264572 267028
rect 278320 266976 278372 267028
rect 287796 266976 287848 267028
rect 295248 266976 295300 267028
rect 319444 266976 319496 267028
rect 320548 266976 320600 267028
rect 400772 266976 400824 267028
rect 401508 266976 401560 267028
rect 402060 267044 402112 267096
rect 402888 267044 402940 267096
rect 404728 267044 404780 267096
rect 405648 267044 405700 267096
rect 410524 267044 410576 267096
rect 414756 267044 414808 267096
rect 405924 266976 405976 267028
rect 406108 266976 406160 267028
rect 632244 267044 632296 267096
rect 414940 266976 414992 267028
rect 644480 266976 644532 267028
rect 164148 266908 164200 266960
rect 170956 266840 171008 266892
rect 177580 266772 177632 266824
rect 223028 266772 223080 266824
rect 164884 266704 164936 266756
rect 199476 266704 199528 266756
rect 200764 266704 200816 266756
rect 207020 266704 207072 266756
rect 272524 266840 272576 266892
rect 277768 266840 277820 266892
rect 294328 266840 294380 266892
rect 312452 266908 312504 266960
rect 321008 266908 321060 266960
rect 342168 266908 342220 266960
rect 345480 266908 345532 266960
rect 346216 266908 346268 266960
rect 229744 266772 229796 266824
rect 311164 266840 311216 266892
rect 331312 266840 331364 266892
rect 232412 266704 232464 266756
rect 292948 266704 293000 266756
rect 301872 266704 301924 266756
rect 322204 266772 322256 266824
rect 325976 266772 326028 266824
rect 334072 266772 334124 266824
rect 328644 266704 328696 266756
rect 282276 266636 282328 266688
rect 287704 266636 287756 266688
rect 309876 266636 309928 266688
rect 323584 266636 323636 266688
rect 196624 266568 196676 266620
rect 202420 266568 202472 266620
rect 271604 266568 271656 266620
rect 276296 266568 276348 266620
rect 277400 266568 277452 266620
rect 280528 266568 280580 266620
rect 280988 266568 281040 266620
rect 289176 266568 289228 266620
rect 328184 266568 328236 266620
rect 329104 266568 329156 266620
rect 332600 266568 332652 266620
rect 333796 266568 333848 266620
rect 336648 266840 336700 266892
rect 334808 266772 334860 266824
rect 335268 266772 335320 266824
rect 337476 266772 337528 266824
rect 337936 266772 337988 266824
rect 340144 266772 340196 266824
rect 340696 266772 340748 266824
rect 342812 266772 342864 266824
rect 343456 266772 343508 266824
rect 344652 266840 344704 266892
rect 464712 266908 464764 266960
rect 346400 266840 346452 266892
rect 455420 266840 455472 266892
rect 674748 266840 674800 266892
rect 676220 266840 676272 266892
rect 448520 266772 448572 266824
rect 334256 266704 334308 266756
rect 435364 266704 435416 266756
rect 420184 266636 420236 266688
rect 674656 266636 674708 266688
rect 676036 266636 676088 266688
rect 414020 266568 414072 266620
rect 271144 266500 271196 266552
rect 274640 266500 274692 266552
rect 275192 266500 275244 266552
rect 279424 266500 279476 266552
rect 319260 266500 319312 266552
rect 324964 266500 325016 266552
rect 326344 266500 326396 266552
rect 326988 266500 327040 266552
rect 327264 266500 327316 266552
rect 328368 266500 328420 266552
rect 329012 266500 329064 266552
rect 329748 266500 329800 266552
rect 329932 266500 329984 266552
rect 330668 266500 330720 266552
rect 333060 266500 333112 266552
rect 333888 266500 333940 266552
rect 334072 266500 334124 266552
rect 409144 266500 409196 266552
rect 191104 266432 191156 266484
rect 197728 266432 197780 266484
rect 230480 266432 230532 266484
rect 238668 266432 238720 266484
rect 270684 266432 270736 266484
rect 273260 266432 273312 266484
rect 280068 266432 280120 266484
rect 284852 266432 284904 266484
rect 287612 266432 287664 266484
rect 289084 266432 289136 266484
rect 289820 266432 289872 266484
rect 291016 266432 291068 266484
rect 291660 266432 291712 266484
rect 295984 266432 296036 266484
rect 302792 266432 302844 266484
rect 306012 266432 306064 266484
rect 312084 266432 312136 266484
rect 315304 266432 315356 266484
rect 316592 266432 316644 266484
rect 368020 266432 368072 266484
rect 368664 266432 368716 266484
rect 378784 266432 378836 266484
rect 387800 266432 387852 266484
rect 193864 266364 193916 266416
rect 194600 266364 194652 266416
rect 235264 266364 235316 266416
rect 238208 266364 238260 266416
rect 242164 266364 242216 266416
rect 243084 266364 243136 266416
rect 244188 266364 244240 266416
rect 248420 266364 248472 266416
rect 270316 266364 270368 266416
rect 272156 266364 272208 266416
rect 276480 266364 276532 266416
rect 277308 266364 277360 266416
rect 280528 266364 280580 266416
rect 281356 266364 281408 266416
rect 281816 266364 281868 266416
rect 283012 266364 283064 266416
rect 284116 266364 284168 266416
rect 286784 266364 286836 266416
rect 287152 266364 287204 266416
rect 288348 266364 288400 266416
rect 290280 266364 290332 266416
rect 291108 266364 291160 266416
rect 291200 266364 291252 266416
rect 292488 266364 292540 266416
rect 295616 266364 295668 266416
rect 296536 266364 296588 266416
rect 296996 266364 297048 266416
rect 297824 266364 297876 266416
rect 300952 266364 301004 266416
rect 302148 266364 302200 266416
rect 304080 266364 304132 266416
rect 304816 266364 304868 266416
rect 305460 266364 305512 266416
rect 306288 266364 306340 266416
rect 306748 266364 306800 266416
rect 307576 266364 307628 266416
rect 308128 266364 308180 266416
rect 308956 266364 309008 266416
rect 309416 266364 309468 266416
rect 310336 266364 310388 266416
rect 310796 266364 310848 266416
rect 311716 266364 311768 266416
rect 313464 266364 313516 266416
rect 314476 266364 314528 266416
rect 314844 266364 314896 266416
rect 315856 266364 315908 266416
rect 316132 266364 316184 266416
rect 317236 266364 317288 266416
rect 317512 266364 317564 266416
rect 318616 266364 318668 266416
rect 318800 266364 318852 266416
rect 319996 266364 320048 266416
rect 320180 266364 320232 266416
rect 321376 266364 321428 266416
rect 324596 266364 324648 266416
rect 354680 266364 354732 266416
rect 354864 266364 354916 266416
rect 355968 266364 356020 266416
rect 356244 266364 356296 266416
rect 357164 266364 357216 266416
rect 358912 266364 358964 266416
rect 359924 266364 359976 266416
rect 362408 266364 362460 266416
rect 362868 266364 362920 266416
rect 364708 266364 364760 266416
rect 365444 266364 365496 266416
rect 367376 266364 367428 266416
rect 368388 266364 368440 266416
rect 370044 266364 370096 266416
rect 371148 266364 371200 266416
rect 372712 266364 372764 266416
rect 373908 266364 373960 266416
rect 376208 266364 376260 266416
rect 376576 266364 376628 266416
rect 381176 266364 381228 266416
rect 382004 266364 382056 266416
rect 383844 266364 383896 266416
rect 384948 266364 385000 266416
rect 390928 266364 390980 266416
rect 391756 266364 391808 266416
rect 393596 266432 393648 266484
rect 394516 266432 394568 266484
rect 394976 266432 395028 266484
rect 395804 266432 395856 266484
rect 396264 266432 396316 266484
rect 397276 266432 397328 266484
rect 408684 266432 408736 266484
rect 408776 266432 408828 266484
rect 479524 266432 479576 266484
rect 410064 266364 410116 266416
rect 411076 266364 411128 266416
rect 355784 266296 355836 266348
rect 499580 266296 499632 266348
rect 358452 266228 358504 266280
rect 506480 266228 506532 266280
rect 361120 266160 361172 266212
rect 513380 266160 513432 266212
rect 373172 266092 373224 266144
rect 545120 266092 545172 266144
rect 374460 266024 374512 266076
rect 549260 266024 549312 266076
rect 674656 266024 674708 266076
rect 676220 266024 676272 266076
rect 375840 265956 375892 266008
rect 552020 265956 552072 266008
rect 377128 265888 377180 265940
rect 556160 265888 556212 265940
rect 378508 265820 378560 265872
rect 558920 265820 558972 265872
rect 379796 265752 379848 265804
rect 563060 265752 563112 265804
rect 382464 265684 382516 265736
rect 569960 265684 570012 265736
rect 385592 265616 385644 265668
rect 578240 265616 578292 265668
rect 194692 265548 194744 265600
rect 195612 265548 195664 265600
rect 201592 265548 201644 265600
rect 202236 265548 202288 265600
rect 223672 265548 223724 265600
rect 224500 265548 224552 265600
rect 238852 265548 238904 265600
rect 239680 265548 239732 265600
rect 240140 265548 240192 265600
rect 240508 265548 240560 265600
rect 242992 265548 243044 265600
rect 243636 265548 243688 265600
rect 244372 265548 244424 265600
rect 245016 265548 245068 265600
rect 247224 265548 247276 265600
rect 247684 265548 247736 265600
rect 251272 265548 251324 265600
rect 251732 265548 251784 265600
rect 259644 265548 259696 265600
rect 260196 265548 260248 265600
rect 262312 265548 262364 265600
rect 262772 265548 262824 265600
rect 264980 265548 265032 265600
rect 265900 265548 265952 265600
rect 266360 265548 266412 265600
rect 267280 265548 267332 265600
rect 353116 265548 353168 265600
rect 491300 265548 491352 265600
rect 336188 265480 336240 265532
rect 447140 265480 447192 265532
rect 334348 265412 334400 265464
rect 443000 265412 443052 265464
rect 333520 265344 333572 265396
rect 440240 265344 440292 265396
rect 331680 265276 331732 265328
rect 434904 265276 434956 265328
rect 327724 265208 327776 265260
rect 425060 265208 425112 265260
rect 673368 265208 673420 265260
rect 676220 265208 676272 265260
rect 325056 265140 325108 265192
rect 418160 265140 418212 265192
rect 673276 265072 673328 265124
rect 676036 265072 676088 265124
rect 673368 264936 673420 264988
rect 676128 264936 676180 264988
rect 367008 264460 367060 264512
rect 528560 264460 528612 264512
rect 384948 264392 385000 264444
rect 575480 264392 575532 264444
rect 387616 264324 387668 264376
rect 582564 264324 582616 264376
rect 393044 264256 393096 264308
rect 597560 264256 597612 264308
rect 43996 264188 44048 264240
rect 662420 264188 662472 264240
rect 399760 264120 399812 264172
rect 401232 264120 401284 264172
rect 607404 264120 607456 264172
rect 615500 264052 615552 264104
rect 673276 263576 673328 263628
rect 676220 263576 676272 263628
rect 415308 262216 415360 262268
rect 572720 262216 572772 262268
rect 674564 259088 674616 259140
rect 676220 259088 676272 259140
rect 35808 258068 35860 258120
rect 44916 258068 44968 258120
rect 179420 258068 179472 258120
rect 189080 258068 189132 258120
rect 414204 258068 414256 258120
rect 571524 258068 571576 258120
rect 673184 258068 673236 258120
rect 676220 258068 676272 258120
rect 31668 258000 31720 258052
rect 43720 258000 43772 258052
rect 31576 257864 31628 257916
rect 44732 257864 44784 257916
rect 31668 257728 31720 257780
rect 46204 257728 46256 257780
rect 673092 256708 673144 256760
rect 683120 256708 683172 256760
rect 415308 255280 415360 255332
rect 571432 255280 571484 255332
rect 414388 252560 414440 252612
rect 574744 252560 574796 252612
rect 675760 252560 675812 252612
rect 678244 252560 678296 252612
rect 675208 251608 675260 251660
rect 676496 251608 676548 251660
rect 675024 251540 675076 251592
rect 676864 251540 676916 251592
rect 676956 251540 677008 251592
rect 674012 251472 674064 251524
rect 173900 251336 173952 251388
rect 179420 251336 179472 251388
rect 675760 251200 675812 251252
rect 675760 250928 675812 250980
rect 674472 249976 674524 250028
rect 675208 249976 675260 250028
rect 673644 249840 673696 249892
rect 674564 249840 674616 249892
rect 674564 249704 674616 249756
rect 675024 249704 675076 249756
rect 171784 249296 171836 249348
rect 173900 249296 173952 249348
rect 675208 248480 675260 248532
rect 414204 248412 414256 248464
rect 574100 248412 574152 248464
rect 675208 248276 675260 248328
rect 675024 247868 675076 247920
rect 675484 247868 675536 247920
rect 674472 247256 674524 247308
rect 675116 247256 675168 247308
rect 674564 247052 674616 247104
rect 675392 247052 675444 247104
rect 674012 246508 674064 246560
rect 675392 246508 675444 246560
rect 675116 246032 675168 246084
rect 675392 246032 675444 246084
rect 42432 245760 42484 245812
rect 42708 245760 42760 245812
rect 35808 245624 35860 245676
rect 191104 245624 191156 245676
rect 415308 245624 415360 245676
rect 565084 245624 565136 245676
rect 673920 243584 673972 243636
rect 675300 243584 675352 243636
rect 414388 242904 414440 242956
rect 623044 242904 623096 242956
rect 673644 242836 673696 242888
rect 675300 242836 675352 242888
rect 171784 241544 171836 241596
rect 164884 241408 164936 241460
rect 673184 241204 673236 241256
rect 675300 241204 675352 241256
rect 42156 240320 42208 240372
rect 42432 240320 42484 240372
rect 42708 238756 42760 238808
rect 43168 238756 43220 238808
rect 185584 237396 185636 237448
rect 189080 237396 189132 237448
rect 42156 235356 42208 235408
rect 44548 235356 44600 235408
rect 182916 234948 182968 235000
rect 185584 234948 185636 235000
rect 42156 233996 42208 234048
rect 44456 233996 44508 234048
rect 178040 233452 178092 233504
rect 182916 233452 182968 233504
rect 414204 232500 414256 232552
rect 639144 232500 639196 232552
rect 414940 232432 414992 232484
rect 638224 232432 638276 232484
rect 414296 232364 414348 232416
rect 577504 232364 577556 232416
rect 190368 231684 190420 231736
rect 604460 231684 604512 231736
rect 67548 231616 67600 231668
rect 178040 231616 178092 231668
rect 191104 231616 191156 231668
rect 663984 231616 664036 231668
rect 85028 231548 85080 231600
rect 663800 231548 663852 231600
rect 84844 231480 84896 231532
rect 663892 231480 663944 231532
rect 50344 231412 50396 231464
rect 650644 231412 650696 231464
rect 48964 231344 49016 231396
rect 649356 231344 649408 231396
rect 54484 231276 54536 231328
rect 655520 231276 655572 231328
rect 51724 231208 51776 231260
rect 652760 231208 652812 231260
rect 49056 231140 49108 231192
rect 661040 231140 661092 231192
rect 43812 231072 43864 231124
rect 662512 231072 662564 231124
rect 350172 230596 350224 230648
rect 423680 230596 423732 230648
rect 385132 230528 385184 230580
rect 507860 230528 507912 230580
rect 333612 230460 333664 230512
rect 179328 230392 179380 230444
rect 246120 230392 246172 230444
rect 262864 230392 262916 230444
rect 269948 230392 270000 230444
rect 42064 230324 42116 230376
rect 42984 230324 43036 230376
rect 175188 230324 175240 230376
rect 244648 230324 244700 230376
rect 246948 230324 247000 230376
rect 274640 230392 274692 230444
rect 276664 230392 276716 230444
rect 277768 230392 277820 230444
rect 271144 230324 271196 230376
rect 272800 230324 272852 230376
rect 169668 230256 169720 230308
rect 241796 230256 241848 230308
rect 244188 230256 244240 230308
rect 274272 230256 274324 230308
rect 274548 230256 274600 230308
rect 285312 230392 285364 230444
rect 286968 230392 287020 230444
rect 279424 230324 279476 230376
rect 283196 230324 283248 230376
rect 278044 230256 278096 230308
rect 287428 230324 287480 230376
rect 288348 230392 288400 230444
rect 292764 230392 292816 230444
rect 297456 230392 297508 230444
rect 299940 230392 299992 230444
rect 300216 230392 300268 230444
rect 303988 230392 304040 230444
rect 311716 230392 311768 230444
rect 315304 230392 315356 230444
rect 323124 230392 323176 230444
rect 291752 230324 291804 230376
rect 292580 230324 292632 230376
rect 293868 230324 293920 230376
rect 298100 230324 298152 230376
rect 299296 230324 299348 230376
rect 299572 230324 299624 230376
rect 300492 230324 300544 230376
rect 304172 230324 304224 230376
rect 304908 230324 304960 230376
rect 305644 230324 305696 230376
rect 306196 230324 306248 230376
rect 307024 230324 307076 230376
rect 307576 230324 307628 230376
rect 312084 230324 312136 230376
rect 313188 230324 313240 230376
rect 314936 230324 314988 230376
rect 315948 230324 316000 230376
rect 316316 230324 316368 230376
rect 317328 230324 317380 230376
rect 319260 230324 319312 230376
rect 319904 230324 319956 230376
rect 323492 230324 323544 230376
rect 324228 230324 324280 230376
rect 328460 230392 328512 230444
rect 329564 230392 329616 230444
rect 329840 230392 329892 230444
rect 330852 230392 330904 230444
rect 331680 230392 331732 230444
rect 332416 230392 332468 230444
rect 333060 230392 333112 230444
rect 333796 230392 333848 230444
rect 386236 230460 386288 230512
rect 511264 230460 511316 230512
rect 604460 230460 604512 230512
rect 605748 230460 605800 230512
rect 636844 230460 636896 230512
rect 371884 230392 371936 230444
rect 382280 230392 382332 230444
rect 383568 230392 383620 230444
rect 386880 230392 386932 230444
rect 388444 230392 388496 230444
rect 393320 230392 393372 230444
rect 394608 230392 394660 230444
rect 401876 230392 401928 230444
rect 456156 230392 456208 230444
rect 340144 230324 340196 230376
rect 341984 230324 342036 230376
rect 380440 230324 380492 230376
rect 381176 230324 381228 230376
rect 382188 230324 382240 230376
rect 382648 230324 382700 230376
rect 383384 230324 383436 230376
rect 383660 230324 383712 230376
rect 384948 230324 385000 230376
rect 385500 230324 385552 230376
rect 386328 230324 386380 230376
rect 386512 230324 386564 230376
rect 387708 230324 387760 230376
rect 387800 230324 387852 230376
rect 400680 230324 400732 230376
rect 403348 230324 403400 230376
rect 404176 230324 404228 230376
rect 406200 230324 406252 230376
rect 407028 230324 407080 230376
rect 409052 230324 409104 230376
rect 411168 230324 411220 230376
rect 411352 230324 411404 230376
rect 461584 230324 461636 230376
rect 285588 230256 285640 230308
rect 290648 230256 290700 230308
rect 310612 230256 310664 230308
rect 314476 230256 314528 230308
rect 317420 230256 317472 230308
rect 136364 230188 136416 230240
rect 213276 230188 213328 230240
rect 219256 230188 219308 230240
rect 263232 230188 263284 230240
rect 276756 230188 276808 230240
rect 287060 230188 287112 230240
rect 298836 230188 298888 230240
rect 302424 230188 302476 230240
rect 314568 230188 314620 230240
rect 155868 230120 155920 230172
rect 236092 230120 236144 230172
rect 240048 230120 240100 230172
rect 271788 230120 271840 230172
rect 275376 230120 275428 230172
rect 277676 230120 277728 230172
rect 277768 230120 277820 230172
rect 286048 230120 286100 230172
rect 317788 230188 317840 230240
rect 318708 230188 318760 230240
rect 319352 230120 319404 230172
rect 320272 230256 320324 230308
rect 337384 230256 337436 230308
rect 339132 230256 339184 230308
rect 378968 230256 379020 230308
rect 385868 230256 385920 230308
rect 391112 230256 391164 230308
rect 398656 230256 398708 230308
rect 405740 230256 405792 230308
rect 405832 230256 405884 230308
rect 409604 230256 409656 230308
rect 409788 230256 409840 230308
rect 467104 230256 467156 230308
rect 321652 230188 321704 230240
rect 338764 230188 338816 230240
rect 347688 230188 347740 230240
rect 387616 230188 387668 230240
rect 389088 230188 389140 230240
rect 396724 230188 396776 230240
rect 398104 230188 398156 230240
rect 403072 230188 403124 230240
rect 403992 230188 404044 230240
rect 406660 230188 406712 230240
rect 406844 230188 406896 230240
rect 411076 230188 411128 230240
rect 411260 230188 411312 230240
rect 468484 230188 468536 230240
rect 330116 230120 330168 230172
rect 330208 230120 330260 230172
rect 331036 230120 331088 230172
rect 336648 230120 336700 230172
rect 376024 230120 376076 230172
rect 378324 230120 378376 230172
rect 443644 230120 443696 230172
rect 146208 230052 146260 230104
rect 231860 230052 231912 230104
rect 234528 230052 234580 230104
rect 262864 230052 262916 230104
rect 139308 229984 139360 230036
rect 229008 229984 229060 230036
rect 233148 229984 233200 230036
rect 268936 230052 268988 230104
rect 271328 230052 271380 230104
rect 277124 230052 277176 230104
rect 270316 229984 270368 230036
rect 283840 230052 283892 230104
rect 315856 230052 315908 230104
rect 322204 230052 322256 230104
rect 323768 230052 323820 230104
rect 364524 230052 364576 230104
rect 368020 230052 368072 230104
rect 387524 230052 387576 230104
rect 387984 230052 388036 230104
rect 515404 230052 515456 230104
rect 277308 229984 277360 230036
rect 282460 229984 282512 230036
rect 284208 229984 284260 230036
rect 290280 229984 290332 230036
rect 312360 229984 312412 230036
rect 336924 229984 336976 230036
rect 343732 229984 343784 230036
rect 385684 229984 385736 230036
rect 399024 229984 399076 230036
rect 400128 229984 400180 230036
rect 401140 229984 401192 230036
rect 406752 229984 406804 230036
rect 407028 229984 407080 230036
rect 409788 229984 409840 230036
rect 132408 229916 132460 229968
rect 226156 229916 226208 229968
rect 226248 229916 226300 229968
rect 266084 229916 266136 229968
rect 270408 229916 270460 229968
rect 284576 229916 284628 229968
rect 285496 229916 285548 229968
rect 291384 229916 291436 229968
rect 303528 229916 303580 229968
rect 312544 229916 312596 229968
rect 313832 229916 313884 229968
rect 341248 229916 341300 229968
rect 356244 229916 356296 229968
rect 357072 229916 357124 229968
rect 359096 229916 359148 229968
rect 360108 229916 360160 229968
rect 360568 229916 360620 229968
rect 361304 229916 361356 229968
rect 361948 229916 362000 229968
rect 362684 229916 362736 229968
rect 362776 229916 362828 229968
rect 406476 229916 406528 229968
rect 407212 229916 407264 229968
rect 91744 229848 91796 229900
rect 203340 229848 203392 229900
rect 212448 229848 212500 229900
rect 260380 229848 260432 229900
rect 263508 229848 263560 229900
rect 281724 229848 281776 229900
rect 296720 229848 296772 229900
rect 299572 229848 299624 229900
rect 305000 229848 305052 229900
rect 311440 229848 311492 229900
rect 316684 229848 316736 229900
rect 346492 229848 346544 229900
rect 352012 229848 352064 229900
rect 398104 229848 398156 229900
rect 399760 229848 399812 229900
rect 407764 229848 407816 229900
rect 539600 229984 539652 230036
rect 85396 229780 85448 229832
rect 206192 229780 206244 229832
rect 206744 229780 206796 229832
rect 257528 229780 257580 229832
rect 259368 229780 259420 229832
rect 280344 229780 280396 229832
rect 281356 229780 281408 229832
rect 289912 229780 289964 229832
rect 302056 229780 302108 229832
rect 311164 229780 311216 229832
rect 318064 229780 318116 229832
rect 350908 229780 350960 229832
rect 354864 229780 354916 229832
rect 407120 229780 407172 229832
rect 411352 229916 411404 229968
rect 547144 229916 547196 229968
rect 71688 229712 71740 229764
rect 200488 229712 200540 229764
rect 200672 229712 200724 229764
rect 254676 229712 254728 229764
rect 255228 229712 255280 229764
rect 278504 229712 278556 229764
rect 278688 229712 278740 229764
rect 288532 229712 288584 229764
rect 315212 229712 315264 229764
rect 343732 229712 343784 229764
rect 344836 229712 344888 229764
rect 406384 229712 406436 229764
rect 406660 229712 406712 229764
rect 408316 229712 408368 229764
rect 410432 229780 410484 229832
rect 563704 229780 563756 229832
rect 411536 229712 411588 229764
rect 570604 229712 570656 229764
rect 140044 229644 140096 229696
rect 205824 229644 205876 229696
rect 227536 229644 227588 229696
rect 267096 229644 267148 229696
rect 268384 229644 268436 229696
rect 277216 229644 277268 229696
rect 277308 229644 277360 229696
rect 277492 229644 277544 229696
rect 277676 229644 277728 229696
rect 285680 229644 285732 229696
rect 318800 229644 318852 229696
rect 334716 229644 334768 229696
rect 340880 229644 340932 229696
rect 380256 229644 380308 229696
rect 391204 229644 391256 229696
rect 392584 229644 392636 229696
rect 400772 229644 400824 229696
rect 453304 229644 453356 229696
rect 151820 229576 151872 229628
rect 218980 229576 219032 229628
rect 248328 229576 248380 229628
rect 149704 229508 149756 229560
rect 216128 229508 216180 229560
rect 244924 229508 244976 229560
rect 254308 229508 254360 229560
rect 260104 229576 260156 229628
rect 262588 229576 262640 229628
rect 270132 229576 270184 229628
rect 271420 229576 271472 229628
rect 275652 229576 275704 229628
rect 280068 229576 280120 229628
rect 288900 229576 288952 229628
rect 313464 229576 313516 229628
rect 314568 229576 314620 229628
rect 328828 229576 328880 229628
rect 329656 229576 329708 229628
rect 330116 229576 330168 229628
rect 334624 229576 334676 229628
rect 338028 229576 338080 229628
rect 272984 229508 273036 229560
rect 281080 229508 281132 229560
rect 300676 229508 300728 229560
rect 305552 229508 305604 229560
rect 327356 229508 327408 229560
rect 341524 229508 341576 229560
rect 350540 229576 350592 229628
rect 388076 229576 388128 229628
rect 397644 229576 397696 229628
rect 398564 229576 398616 229628
rect 398656 229576 398708 229628
rect 404360 229576 404412 229628
rect 407120 229576 407172 229628
rect 407672 229576 407724 229628
rect 407764 229576 407816 229628
rect 449164 229576 449216 229628
rect 352564 229508 352616 229560
rect 366548 229508 366600 229560
rect 416688 229508 416740 229560
rect 146392 229440 146444 229492
rect 209044 229440 209096 229492
rect 275284 229440 275336 229492
rect 283932 229440 283984 229492
rect 339500 229440 339552 229492
rect 353944 229440 353996 229492
rect 355508 229440 355560 229492
rect 386972 229440 387024 229492
rect 393688 229440 393740 229492
rect 400956 229440 401008 229492
rect 401508 229440 401560 229492
rect 405004 229440 405056 229492
rect 405740 229440 405792 229492
rect 441712 229440 441764 229492
rect 186964 229372 187016 229424
rect 248972 229372 249024 229424
rect 273904 229372 273956 229424
rect 282828 229372 282880 229424
rect 298468 229372 298520 229424
rect 301136 229372 301188 229424
rect 332692 229372 332744 229424
rect 333888 229372 333940 229424
rect 334532 229372 334584 229424
rect 342904 229372 342956 229424
rect 361212 229372 361264 229424
rect 383108 229372 383160 229424
rect 392216 229372 392268 229424
rect 430764 229372 430816 229424
rect 162860 229304 162912 229356
rect 223304 229304 223356 229356
rect 277492 229304 277544 229356
rect 286692 229304 286744 229356
rect 295248 229304 295300 229356
rect 296904 229304 296956 229356
rect 331312 229304 331364 229356
rect 332232 229304 332284 229356
rect 342352 229304 342404 229356
rect 343272 229304 343324 229356
rect 371976 229304 372028 229356
rect 398656 229304 398708 229356
rect 402980 229304 403032 229356
rect 404268 229304 404320 229356
rect 404728 229304 404780 229356
rect 409788 229304 409840 229356
rect 410064 229304 410116 229356
rect 435548 229304 435600 229356
rect 180800 229236 180852 229288
rect 238944 229236 238996 229288
rect 271236 229236 271288 229288
rect 279976 229236 280028 229288
rect 281448 229236 281500 229288
rect 288164 229236 288216 229288
rect 313096 229236 313148 229288
rect 318064 229236 318116 229288
rect 357716 229236 357768 229288
rect 376116 229236 376168 229288
rect 384396 229236 384448 229288
rect 411352 229236 411404 229288
rect 255964 229168 256016 229220
rect 260012 229168 260064 229220
rect 282828 229168 282880 229220
rect 289268 229168 289320 229220
rect 296352 229168 296404 229220
rect 298468 229168 298520 229220
rect 369400 229168 369452 229220
rect 378600 229168 378652 229220
rect 395068 229168 395120 229220
rect 408408 229168 408460 229220
rect 409328 229168 409380 229220
rect 62120 229032 62172 229084
rect 67548 229100 67600 229152
rect 257344 229100 257396 229152
rect 258908 229100 258960 229152
rect 284116 229100 284168 229152
rect 289544 229100 289596 229152
rect 405096 229100 405148 229152
rect 411260 229100 411312 229152
rect 411904 229168 411956 229220
rect 420184 229168 420236 229220
rect 551284 229100 551336 229152
rect 120816 229032 120868 229084
rect 220820 229032 220872 229084
rect 365168 229032 365220 229084
rect 460940 229032 460992 229084
rect 117228 228964 117280 229016
rect 219348 228964 219400 229016
rect 332048 228964 332100 229016
rect 370228 228964 370280 229016
rect 373356 228964 373408 229016
rect 480260 228964 480312 229016
rect 114192 228896 114244 228948
rect 217968 228896 218020 228948
rect 224040 228896 224092 228948
rect 234712 228896 234764 228948
rect 329196 228896 329248 228948
rect 371332 228896 371384 228948
rect 375104 228896 375156 228948
rect 483480 228896 483532 228948
rect 110696 228828 110748 228880
rect 216496 228828 216548 228880
rect 227720 228828 227772 228880
rect 240416 228828 240468 228880
rect 327724 228828 327776 228880
rect 372712 228828 372764 228880
rect 376576 228828 376628 228880
rect 487712 228828 487764 228880
rect 107476 228760 107528 228812
rect 215116 228760 215168 228812
rect 216680 228760 216732 228812
rect 224684 228760 224736 228812
rect 230296 228760 230348 228812
rect 103980 228692 104032 228744
rect 213644 228692 213696 228744
rect 222108 228692 222160 228744
rect 230388 228692 230440 228744
rect 233516 228760 233568 228812
rect 268200 228760 268252 228812
rect 330576 228760 330628 228812
rect 375288 228760 375340 228812
rect 377956 228760 378008 228812
rect 491300 228760 491352 228812
rect 266728 228692 266780 228744
rect 328092 228692 328144 228744
rect 374000 228692 374052 228744
rect 391940 228692 391992 228744
rect 523040 228692 523092 228744
rect 100668 228624 100720 228676
rect 212264 228624 212316 228676
rect 215116 228624 215168 228676
rect 260748 228624 260800 228676
rect 334900 228624 334952 228676
rect 389272 228624 389324 228676
rect 392952 228624 393004 228676
rect 526352 228624 526404 228676
rect 97264 228556 97316 228608
rect 210792 228556 210844 228608
rect 213828 228556 213880 228608
rect 258540 228556 258592 228608
rect 336280 228556 336332 228608
rect 392492 228556 392544 228608
rect 398288 228556 398340 228608
rect 538220 228556 538272 228608
rect 77944 228488 77996 228540
rect 91744 228488 91796 228540
rect 93768 228488 93820 228540
rect 209412 228488 209464 228540
rect 209872 228488 209924 228540
rect 257160 228488 257212 228540
rect 306656 228488 306708 228540
rect 323676 228488 323728 228540
rect 337752 228488 337804 228540
rect 396172 228488 396224 228540
rect 397276 228488 397328 228540
rect 536840 228488 536892 228540
rect 54392 228420 54444 228472
rect 193312 228420 193364 228472
rect 194968 228420 195020 228472
rect 252192 228420 252244 228472
rect 53656 228352 53708 228404
rect 192300 228352 192352 228404
rect 194140 228352 194192 228404
rect 252836 228352 252888 228404
rect 127532 228284 127584 228336
rect 223672 228284 223724 228336
rect 252008 228284 252060 228336
rect 276388 228420 276440 228472
rect 309876 228420 309928 228472
rect 327816 228420 327868 228472
rect 340604 228420 340656 228472
rect 402980 228420 403032 228472
rect 409788 228420 409840 228472
rect 553952 228420 554004 228472
rect 260564 228352 260616 228404
rect 279608 228352 279660 228404
rect 308128 228352 308180 228404
rect 327080 228352 327132 228404
rect 345204 228352 345256 228404
rect 408500 228352 408552 228404
rect 410800 228352 410852 228404
rect 569132 228352 569184 228404
rect 353392 228284 353444 228336
rect 433340 228284 433392 228336
rect 131028 228216 131080 228268
rect 225052 228216 225104 228268
rect 349160 228216 349212 228268
rect 423036 228216 423088 228268
rect 137744 228148 137796 228200
rect 227904 228148 227956 228200
rect 334164 228148 334216 228200
rect 378508 228148 378560 228200
rect 378968 228148 379020 228200
rect 399392 228148 399444 228200
rect 404360 228148 404412 228200
rect 476120 228148 476172 228200
rect 144368 228080 144420 228132
rect 230756 228080 230808 228132
rect 346308 228080 346360 228132
rect 409972 228080 410024 228132
rect 420184 228080 420236 228132
rect 485136 228080 485188 228132
rect 154488 228012 154540 228064
rect 235080 228012 235132 228064
rect 343456 228012 343508 228064
rect 387248 228012 387300 228064
rect 406476 228012 406528 228064
rect 454040 228012 454092 228064
rect 161296 227944 161348 227996
rect 237932 227944 237984 227996
rect 388076 227944 388128 227996
rect 426440 227944 426492 227996
rect 171048 227876 171100 227928
rect 242164 227876 242216 227928
rect 387616 227876 387668 227928
rect 419540 227876 419592 227928
rect 403072 227808 403124 227860
rect 429660 227808 429712 227860
rect 375472 227740 375524 227792
rect 379704 227740 379756 227792
rect 380440 227740 380492 227792
rect 406108 227740 406160 227792
rect 160376 227672 160428 227724
rect 238576 227672 238628 227724
rect 364432 227672 364484 227724
rect 457352 227672 457404 227724
rect 157064 227604 157116 227656
rect 237196 227604 237248 227656
rect 360200 227604 360252 227656
rect 447324 227604 447376 227656
rect 449164 227604 449216 227656
rect 543004 227604 543056 227656
rect 153660 227536 153712 227588
rect 235724 227536 235776 227588
rect 365904 227536 365956 227588
rect 461216 227536 461268 227588
rect 461584 227536 461636 227588
rect 552664 227536 552716 227588
rect 108212 227468 108264 227520
rect 149704 227468 149756 227520
rect 150348 227468 150400 227520
rect 234344 227468 234396 227520
rect 367284 227468 367336 227520
rect 464160 227468 464212 227520
rect 147496 227400 147548 227452
rect 232228 227400 232280 227452
rect 309508 227400 309560 227452
rect 330392 227400 330444 227452
rect 368756 227400 368808 227452
rect 467840 227400 467892 227452
rect 468484 227400 468536 227452
rect 554964 227400 555016 227452
rect 91376 227332 91428 227384
rect 146392 227332 146444 227384
rect 146944 227332 146996 227384
rect 232872 227332 232924 227384
rect 315580 227332 315632 227384
rect 341340 227332 341392 227384
rect 370136 227332 370188 227384
rect 470876 227332 470928 227384
rect 141056 227264 141108 227316
rect 229376 227264 229428 227316
rect 312728 227264 312780 227316
rect 333980 227264 334032 227316
rect 335176 227264 335228 227316
rect 363144 227264 363196 227316
rect 371608 227264 371660 227316
rect 474188 227264 474240 227316
rect 143448 227196 143500 227248
rect 231492 227196 231544 227248
rect 232780 227196 232832 227248
rect 247500 227196 247552 227248
rect 318432 227196 318484 227248
rect 348056 227196 348108 227248
rect 372988 227196 373040 227248
rect 477592 227196 477644 227248
rect 478144 227196 478196 227248
rect 489368 227196 489420 227248
rect 82728 227128 82780 227180
rect 140044 227128 140096 227180
rect 140136 227128 140188 227180
rect 230020 227128 230072 227180
rect 237380 227128 237432 227180
rect 256056 227128 256108 227180
rect 258816 227128 258868 227180
rect 279240 227128 279292 227180
rect 321284 227128 321336 227180
rect 354772 227128 354824 227180
rect 374460 227128 374512 227180
rect 480904 227128 480956 227180
rect 134248 227060 134300 227112
rect 226524 227060 226576 227112
rect 234712 227060 234764 227112
rect 253204 227060 253256 227112
rect 255136 227060 255188 227112
rect 277860 227060 277912 227112
rect 325608 227060 325660 227112
rect 360292 227060 360344 227112
rect 374828 227060 374880 227112
rect 483112 227060 483164 227112
rect 124128 226992 124180 227044
rect 222200 226992 222252 227044
rect 237012 226992 237064 227044
rect 269580 226992 269632 227044
rect 305276 226992 305328 227044
rect 320272 226992 320324 227044
rect 329472 226992 329524 227044
rect 365352 226992 365404 227044
rect 409696 226992 409748 227044
rect 565912 226992 565964 227044
rect 125048 226924 125100 226976
rect 162860 226924 162912 226976
rect 163688 226924 163740 226976
rect 239772 226924 239824 226976
rect 363052 226924 363104 226976
rect 454132 226924 454184 226976
rect 166908 226856 166960 226908
rect 241428 226856 241480 226908
rect 361580 226856 361632 226908
rect 450636 226856 450688 226908
rect 164608 226788 164660 226840
rect 239312 226788 239364 226840
rect 358728 226788 358780 226840
rect 444380 226788 444432 226840
rect 173808 226720 173860 226772
rect 244280 226720 244332 226772
rect 357348 226720 357400 226772
rect 440608 226720 440660 226772
rect 42156 226652 42208 226704
rect 44364 226652 44416 226704
rect 174636 226652 174688 226704
rect 243636 226652 243688 226704
rect 355876 226652 355928 226704
rect 437480 226652 437532 226704
rect 177212 226584 177264 226636
rect 245752 226584 245804 226636
rect 354496 226584 354548 226636
rect 433800 226584 433852 226636
rect 190276 226516 190328 226568
rect 251456 226516 251508 226568
rect 351644 226516 351696 226568
rect 427084 226516 427136 226568
rect 57612 226312 57664 226364
rect 62120 226312 62172 226364
rect 116584 226244 116636 226296
rect 220084 226244 220136 226296
rect 364248 226244 364300 226296
rect 455696 226244 455748 226296
rect 456156 226244 456208 226296
rect 548156 226244 548208 226296
rect 112996 226176 113048 226228
rect 218612 226176 218664 226228
rect 223120 226176 223172 226228
rect 233240 226176 233292 226228
rect 365536 226176 365588 226228
rect 459560 226176 459612 226228
rect 109868 226108 109920 226160
rect 217232 226108 217284 226160
rect 218060 226108 218112 226160
rect 227260 226108 227312 226160
rect 227352 226108 227404 226160
rect 237564 226108 237616 226160
rect 366916 226108 366968 226160
rect 462412 226108 462464 226160
rect 106556 226040 106608 226092
rect 215760 226040 215812 226092
rect 224960 226040 225012 226092
rect 251824 226040 251876 226092
rect 253848 226040 253900 226092
rect 276480 226040 276532 226092
rect 335912 226040 335964 226092
rect 367744 226040 367796 226092
rect 368388 226040 368440 226092
rect 465080 226040 465132 226092
rect 103244 225972 103296 226024
rect 214380 225972 214432 226024
rect 220636 225972 220688 226024
rect 264244 225972 264296 226024
rect 358360 225972 358412 226024
rect 441620 225972 441672 226024
rect 441712 225972 441764 226024
rect 540428 225972 540480 226024
rect 99840 225904 99892 225956
rect 212908 225904 212960 225956
rect 215300 225904 215352 225956
rect 261392 225904 261444 225956
rect 322756 225904 322808 225956
rect 358176 225904 358228 225956
rect 369768 225904 369820 225956
rect 469220 225904 469272 225956
rect 96528 225836 96580 225888
rect 211528 225836 211580 225888
rect 211712 225836 211764 225888
rect 259000 225836 259052 225888
rect 326988 225836 327040 225888
rect 362960 225836 363012 225888
rect 371240 225836 371292 225888
rect 471980 225836 472032 225888
rect 86316 225768 86368 225820
rect 207204 225768 207256 225820
rect 208308 225768 208360 225820
rect 257896 225768 257948 225820
rect 324136 225768 324188 225820
rect 361580 225768 361632 225820
rect 372620 225768 372672 225820
rect 476212 225768 476264 225820
rect 76288 225700 76340 225752
rect 202972 225700 203024 225752
rect 206836 225700 206888 225752
rect 256792 225700 256844 225752
rect 303804 225700 303856 225752
rect 317420 225700 317472 225752
rect 343088 225700 343140 225752
rect 407120 225700 407172 225752
rect 408408 225700 408460 225752
rect 531412 225700 531464 225752
rect 539600 225700 539652 225752
rect 560300 225700 560352 225752
rect 56048 225632 56100 225684
rect 194416 225632 194468 225684
rect 199016 225632 199068 225684
rect 200672 225632 200724 225684
rect 203248 225632 203300 225684
rect 255320 225632 255372 225684
rect 263416 225632 263468 225684
rect 280988 225632 281040 225684
rect 302700 225632 302752 225684
rect 313556 225632 313608 225684
rect 314476 225632 314528 225684
rect 331220 225632 331272 225684
rect 341616 225632 341668 225684
rect 403532 225632 403584 225684
rect 403624 225632 403676 225684
rect 552020 225632 552072 225684
rect 52736 225564 52788 225616
rect 192668 225564 192720 225616
rect 201408 225564 201460 225616
rect 255044 225564 255096 225616
rect 257068 225564 257120 225616
rect 278136 225564 278188 225616
rect 310980 225564 311032 225616
rect 334072 225564 334124 225616
rect 344468 225564 344520 225616
rect 410248 225564 410300 225616
rect 411076 225564 411128 225616
rect 559196 225564 559248 225616
rect 119896 225496 119948 225548
rect 221188 225496 221240 225548
rect 362868 225496 362920 225548
rect 452660 225496 452712 225548
rect 123392 225428 123444 225480
rect 222936 225428 222988 225480
rect 359832 225428 359884 225480
rect 445760 225428 445812 225480
rect 126796 225360 126848 225412
rect 224316 225360 224368 225412
rect 356980 225360 357032 225412
rect 438860 225360 438912 225412
rect 130108 225292 130160 225344
rect 225788 225292 225840 225344
rect 348792 225292 348844 225344
rect 420368 225292 420420 225344
rect 133512 225224 133564 225276
rect 227168 225224 227220 225276
rect 345940 225224 345992 225276
rect 414020 225224 414072 225276
rect 170496 225156 170548 225208
rect 242900 225156 242952 225208
rect 339040 225156 339092 225208
rect 382280 225156 382332 225208
rect 383108 225156 383160 225208
rect 448980 225156 449032 225208
rect 180616 225088 180668 225140
rect 247132 225088 247184 225140
rect 340236 225088 340288 225140
rect 385684 225088 385736 225140
rect 386972 225088 387024 225140
rect 434720 225088 434772 225140
rect 192852 224952 192904 225004
rect 197636 224952 197688 225004
rect 162768 224884 162820 224936
rect 238208 224884 238260 224936
rect 374092 224884 374144 224936
rect 479248 224884 479300 224936
rect 159548 224816 159600 224868
rect 236828 224816 236880 224868
rect 370872 224816 370924 224868
rect 475016 224816 475068 224868
rect 155776 224748 155828 224800
rect 235356 224748 235408 224800
rect 372252 224748 372304 224800
rect 478972 224748 479024 224800
rect 114928 224680 114980 224732
rect 151820 224680 151872 224732
rect 152924 224680 152976 224732
rect 233976 224680 234028 224732
rect 332324 224680 332376 224732
rect 372620 224680 372672 224732
rect 373724 224680 373776 224732
rect 481824 224680 481876 224732
rect 149428 224612 149480 224664
rect 232320 224612 232372 224664
rect 338396 224612 338448 224664
rect 380164 224612 380216 224664
rect 388720 224612 388772 224664
rect 516232 224612 516284 224664
rect 146116 224544 146168 224596
rect 231124 224544 231176 224596
rect 337016 224544 337068 224596
rect 378692 224544 378744 224596
rect 389732 224544 389784 224596
rect 518900 224544 518952 224596
rect 142712 224476 142764 224528
rect 229652 224476 229704 224528
rect 342720 224476 342772 224528
rect 405924 224476 405976 224528
rect 406752 224476 406804 224528
rect 545764 224476 545816 224528
rect 139216 224408 139268 224460
rect 228272 224408 228324 224460
rect 234620 224408 234672 224460
rect 250352 224408 250404 224460
rect 268936 224408 268988 224460
rect 283564 224408 283616 224460
rect 333704 224408 333756 224460
rect 378048 224408 378100 224460
rect 400036 224408 400088 224460
rect 543188 224408 543240 224460
rect 135996 224340 136048 224392
rect 226800 224340 226852 224392
rect 246856 224340 246908 224392
rect 273628 224340 273680 224392
rect 307760 224340 307812 224392
rect 325700 224340 325752 224392
rect 339868 224340 339920 224392
rect 386972 224340 387024 224392
rect 402244 224340 402296 224392
rect 548248 224340 548300 224392
rect 101496 224272 101548 224324
rect 136364 224272 136416 224324
rect 136456 224272 136508 224324
rect 228640 224272 228692 224324
rect 232412 224272 232464 224324
rect 243268 224272 243320 224324
rect 243636 224272 243688 224324
rect 272248 224272 272300 224324
rect 309232 224272 309284 224324
rect 328736 224272 328788 224324
rect 341432 224272 341484 224324
rect 401876 224272 401928 224324
rect 408684 224272 408736 224324
rect 88156 224204 88208 224256
rect 207572 224204 207624 224256
rect 239956 224204 240008 224256
rect 271052 224204 271104 224256
rect 292580 224204 292632 224256
rect 293500 224204 293552 224256
rect 311348 224204 311400 224256
rect 331312 224204 331364 224256
rect 344100 224204 344152 224256
rect 408592 224204 408644 224256
rect 411352 224204 411404 224256
rect 412272 224272 412324 224324
rect 556160 224272 556212 224324
rect 166264 224136 166316 224188
rect 239680 224136 239732 224188
rect 345572 224136 345624 224188
rect 411996 224136 412048 224188
rect 563612 224204 563664 224256
rect 506480 224136 506532 224188
rect 169576 224068 169628 224120
rect 241060 224068 241112 224120
rect 335544 224068 335596 224120
rect 377312 224068 377364 224120
rect 378600 224068 378652 224120
rect 472072 224068 472124 224120
rect 172980 224000 173032 224052
rect 242532 224000 242584 224052
rect 387524 224000 387576 224052
rect 468300 224000 468352 224052
rect 176476 223932 176528 223984
rect 243912 223932 243964 223984
rect 349804 223932 349856 223984
rect 422392 223932 422444 223984
rect 179696 223864 179748 223916
rect 245384 223864 245436 223916
rect 347320 223864 347372 223916
rect 417056 223864 417108 223916
rect 183192 223796 183244 223848
rect 246764 223796 246816 223848
rect 348424 223796 348476 223848
rect 418712 223796 418764 223848
rect 186228 223728 186280 223780
rect 248236 223728 248288 223780
rect 346952 223728 347004 223780
rect 415492 223728 415544 223780
rect 416688 223728 416740 223780
rect 465172 223728 465224 223780
rect 405464 223660 405516 223712
rect 412272 223660 412324 223712
rect 125876 223524 125928 223576
rect 222568 223524 222620 223576
rect 357992 223524 358044 223576
rect 444748 223524 444800 223576
rect 115756 223456 115808 223508
rect 210424 223456 210476 223508
rect 213920 223456 213972 223508
rect 221832 223456 221884 223508
rect 359464 223456 359516 223508
rect 448612 223456 448664 223508
rect 108856 223388 108908 223440
rect 215392 223388 215444 223440
rect 361120 223388 361172 223440
rect 451464 223388 451516 223440
rect 105728 223320 105780 223372
rect 214012 223320 214064 223372
rect 352288 223320 352340 223372
rect 431316 223320 431368 223372
rect 431408 223320 431460 223372
rect 525064 223320 525116 223372
rect 101956 223252 102008 223304
rect 95608 223184 95660 223236
rect 210424 223252 210476 223304
rect 218244 223252 218296 223304
rect 390100 223252 390152 223304
rect 395712 223252 395764 223304
rect 396356 223252 396408 223304
rect 523132 223252 523184 223304
rect 82176 223116 82228 223168
rect 203984 223116 204036 223168
rect 212540 223184 212592 223236
rect 314200 223184 314252 223236
rect 338120 223184 338172 223236
rect 353760 223184 353812 223236
rect 434812 223184 434864 223236
rect 435548 223184 435600 223236
rect 567200 223184 567252 223236
rect 209688 223116 209740 223168
rect 250352 223116 250404 223168
rect 275100 223116 275152 223168
rect 317052 223116 317104 223168
rect 345020 223116 345072 223168
rect 395804 223116 395856 223168
rect 75368 223048 75420 223100
rect 201132 223048 201184 223100
rect 204904 223048 204956 223100
rect 256424 223048 256476 223100
rect 319260 223048 319312 223100
rect 350632 223048 350684 223100
rect 391572 223048 391624 223100
rect 396356 223048 396408 223100
rect 398840 223116 398892 223168
rect 530584 223116 530636 223168
rect 671436 223116 671488 223168
rect 675944 223116 675996 223168
rect 533068 223048 533120 223100
rect 68744 222980 68796 223032
rect 65340 222912 65392 222964
rect 196900 222912 196952 222964
rect 198188 222980 198240 223032
rect 253572 222980 253624 223032
rect 311440 222980 311492 223032
rect 318892 222980 318944 223032
rect 330944 222980 330996 223032
rect 365996 222980 366048 223032
rect 397920 222980 397972 223032
rect 538312 222980 538364 223032
rect 198280 222912 198332 222964
rect 199936 222912 199988 222964
rect 253940 222912 253992 222964
rect 265532 222912 265584 222964
rect 282092 222912 282144 222964
rect 306380 222912 306432 222964
rect 321928 222912 321980 222964
rect 326620 222912 326672 222964
rect 371240 222912 371292 222964
rect 379796 222912 379848 222964
rect 389180 222912 389232 222964
rect 394792 222912 394844 222964
rect 398840 222912 398892 222964
rect 404636 222912 404688 222964
rect 553676 222912 553728 222964
rect 66076 222844 66128 222896
rect 198372 222844 198424 222896
rect 200764 222844 200816 222896
rect 255688 222844 255740 222896
rect 262128 222844 262180 222896
rect 280712 222844 280764 222896
rect 308496 222844 308548 222896
rect 324504 222844 324556 222896
rect 337660 222844 337712 222896
rect 390652 222844 390704 222896
rect 407580 222844 407632 222896
rect 560944 222844 560996 222896
rect 132316 222776 132368 222828
rect 225420 222776 225472 222828
rect 356612 222776 356664 222828
rect 441712 222776 441764 222828
rect 177856 222708 177908 222760
rect 245016 222708 245068 222760
rect 355140 222708 355192 222760
rect 438032 222708 438084 222760
rect 674380 222708 674432 222760
rect 675944 222708 675996 222760
rect 162032 222640 162084 222692
rect 180800 222640 180852 222692
rect 181352 222640 181404 222692
rect 246488 222640 246540 222692
rect 352656 222640 352708 222692
rect 429292 222640 429344 222692
rect 187332 222572 187384 222624
rect 249984 222572 250036 222624
rect 351184 222572 351236 222624
rect 427912 222572 427964 222624
rect 428648 222572 428700 222624
rect 488540 222572 488592 222624
rect 184756 222504 184808 222556
rect 247868 222504 247920 222556
rect 349436 222504 349488 222556
rect 425060 222504 425112 222556
rect 188160 222436 188212 222488
rect 249340 222436 249392 222488
rect 348148 222436 348200 222488
rect 421196 222436 421248 222488
rect 191564 222368 191616 222420
rect 250720 222368 250772 222420
rect 346676 222368 346728 222420
rect 415308 222368 415360 222420
rect 196532 222300 196584 222352
rect 252284 222300 252336 222352
rect 664536 222164 664588 222216
rect 676036 222164 676088 222216
rect 122472 222096 122524 222148
rect 221004 222096 221056 222148
rect 228456 222096 228508 222148
rect 266452 222096 266504 222148
rect 311164 222096 311216 222148
rect 311992 222096 312044 222148
rect 312544 222096 312596 222148
rect 315304 222096 315356 222148
rect 318708 222096 318760 222148
rect 349160 222096 349212 222148
rect 362684 222096 362736 222148
rect 453212 222096 453264 222148
rect 453304 222096 453356 222148
rect 545212 222096 545264 222148
rect 119160 222028 119212 222080
rect 219532 222028 219584 222080
rect 226800 222028 226852 222080
rect 265164 222028 265216 222080
rect 320824 222028 320876 222080
rect 356060 222028 356112 222080
rect 363604 222028 363656 222080
rect 456800 222028 456852 222080
rect 100760 221960 100812 222012
rect 204444 221960 204496 222012
rect 224868 221960 224920 222012
rect 265072 221960 265124 222012
rect 322296 221960 322348 222012
rect 359096 221960 359148 222012
rect 365076 221960 365128 222012
rect 460020 221960 460072 222012
rect 112444 221892 112496 221944
rect 216772 221892 216824 221944
rect 223488 221892 223540 221944
rect 263784 221892 263836 221944
rect 321192 221892 321244 221944
rect 357532 221892 357584 221944
rect 363972 221892 364024 221944
rect 458364 221892 458416 221944
rect 88892 221824 88944 221876
rect 85488 221756 85540 221808
rect 205180 221756 205232 221808
rect 205548 221824 205600 221876
rect 206744 221824 206796 221876
rect 220084 221824 220136 221876
rect 262312 221824 262364 221876
rect 322664 221824 322716 221876
rect 360752 221824 360804 221876
rect 366456 221824 366508 221876
rect 463700 221824 463752 221876
rect 672632 221824 672684 221876
rect 676036 221824 676088 221876
rect 206652 221756 206704 221808
rect 208216 221756 208268 221808
rect 220176 221756 220228 221808
rect 221740 221756 221792 221808
rect 263692 221756 263744 221808
rect 324228 221756 324280 221808
rect 362408 221756 362460 221808
rect 367928 221756 367980 221808
rect 466736 221756 466788 221808
rect 467104 221756 467156 221808
rect 557816 221756 557868 221808
rect 83832 221688 83884 221740
rect 204812 221688 204864 221740
rect 206928 221688 206980 221740
rect 217324 221688 217376 221740
rect 218428 221688 218480 221740
rect 261852 221688 261904 221740
rect 325148 221688 325200 221740
rect 365812 221688 365864 221740
rect 369308 221688 369360 221740
rect 470140 221688 470192 221740
rect 80428 221620 80480 221672
rect 203432 221620 203484 221672
rect 203708 221620 203760 221672
rect 214472 221620 214524 221672
rect 216588 221620 216640 221672
rect 261024 221620 261076 221672
rect 326528 221620 326580 221672
rect 369124 221620 369176 221672
rect 370780 221620 370832 221672
rect 473544 221620 473596 221672
rect 551284 221620 551336 221672
rect 565452 221620 565504 221672
rect 77024 221552 77076 221604
rect 201960 221552 202012 221604
rect 202420 221552 202472 221604
rect 210148 221552 210200 221604
rect 213368 221552 213420 221604
rect 259644 221552 259696 221604
rect 325516 221552 325568 221604
rect 367468 221552 367520 221604
rect 400128 221552 400180 221604
rect 541440 221552 541492 221604
rect 547144 221552 547196 221604
rect 561772 221552 561824 221604
rect 63408 221484 63460 221536
rect 196256 221484 196308 221536
rect 197268 221484 197320 221536
rect 244924 221484 244976 221536
rect 245292 221484 245344 221536
rect 273444 221484 273496 221536
rect 275560 221484 275612 221536
rect 286140 221484 286192 221536
rect 319444 221484 319496 221536
rect 352380 221484 352432 221536
rect 352564 221484 352616 221536
rect 397736 221484 397788 221536
rect 404176 221484 404228 221536
rect 551284 221484 551336 221536
rect 674656 221484 674708 221536
rect 676036 221484 676088 221536
rect 60280 221416 60332 221468
rect 194876 221416 194928 221468
rect 209688 221416 209740 221468
rect 258264 221416 258316 221468
rect 272248 221416 272300 221468
rect 284668 221416 284720 221468
rect 301228 221416 301280 221468
rect 310520 221416 310572 221468
rect 319812 221416 319864 221468
rect 354036 221416 354088 221468
rect 129280 221348 129332 221400
rect 223764 221348 223816 221400
rect 231676 221348 231728 221400
rect 267832 221348 267884 221400
rect 317328 221348 317380 221400
rect 345572 221348 345624 221400
rect 151084 221280 151136 221332
rect 233424 221280 233476 221332
rect 235264 221280 235316 221332
rect 269212 221280 269264 221332
rect 315948 221280 316000 221332
rect 342260 221280 342312 221332
rect 353944 221280 353996 221332
rect 401140 221416 401192 221468
rect 406292 221416 406344 221468
rect 558460 221416 558512 221468
rect 565084 221416 565136 221468
rect 573548 221416 573600 221468
rect 361304 221348 361356 221400
rect 449900 221348 449952 221400
rect 360108 221280 360160 221332
rect 446588 221280 446640 221332
rect 157800 221212 157852 221264
rect 236184 221212 236236 221264
rect 238576 221212 238628 221264
rect 270684 221212 270736 221264
rect 314568 221212 314620 221264
rect 338856 221212 338908 221264
rect 357072 221212 357124 221264
rect 439780 221212 439832 221264
rect 443644 221212 443696 221264
rect 491392 221212 491444 221264
rect 167920 221144 167972 221196
rect 240508 221144 240560 221196
rect 241980 221144 242032 221196
rect 271972 221144 272024 221196
rect 313188 221144 313240 221196
rect 335544 221144 335596 221196
rect 351552 221144 351604 221196
rect 425520 221144 425572 221196
rect 183928 221076 183980 221128
rect 248512 221076 248564 221128
rect 248696 221076 248748 221128
rect 274824 221076 274876 221128
rect 376116 221076 376168 221128
rect 443184 221076 443236 221128
rect 189816 221008 189868 221060
rect 249432 221008 249484 221060
rect 343272 221008 343324 221060
rect 407856 221008 407908 221060
rect 192944 220940 192996 220992
rect 250812 220940 250864 220992
rect 385776 220940 385828 220992
rect 411260 220940 411312 220992
rect 195152 220872 195204 220924
rect 211620 220872 211672 220924
rect 380256 220872 380308 220924
rect 404452 220872 404504 220924
rect 407672 220872 407724 220924
rect 436468 221008 436520 221060
rect 672540 221008 672592 221060
rect 676036 221008 676088 221060
rect 563612 220940 563664 220992
rect 563704 220872 563756 220924
rect 567936 220872 567988 220924
rect 569132 220940 569184 220992
rect 621204 220940 621256 220992
rect 619824 220872 619876 220924
rect 52460 220736 52512 220788
rect 57612 220804 57664 220856
rect 71228 220736 71280 220788
rect 71688 220736 71740 220788
rect 84660 220736 84712 220788
rect 85396 220736 85448 220788
rect 131764 220736 131816 220788
rect 132408 220736 132460 220788
rect 138480 220736 138532 220788
rect 139308 220736 139360 220788
rect 141884 220736 141936 220788
rect 222108 220736 222160 220788
rect 232688 220736 232740 220788
rect 233148 220736 233200 220788
rect 239404 220736 239456 220788
rect 240048 220736 240100 220788
rect 241152 220736 241204 220788
rect 269672 220736 269724 220788
rect 270408 220736 270460 220788
rect 305552 220804 305604 220856
rect 308588 220804 308640 220856
rect 558460 220804 558512 220856
rect 618812 220804 618864 220856
rect 271144 220736 271196 220788
rect 273904 220736 273956 220788
rect 274548 220736 274600 220788
rect 278136 220736 278188 220788
rect 278688 220736 278740 220788
rect 282368 220736 282420 220788
rect 282828 220736 282880 220788
rect 286508 220736 286560 220788
rect 286968 220736 287020 220788
rect 287336 220736 287388 220788
rect 290648 220736 290700 220788
rect 290740 220736 290792 220788
rect 292212 220736 292264 220788
rect 292488 220736 292540 220788
rect 293224 220736 293276 220788
rect 294972 220736 295024 220788
rect 295524 220736 295576 220788
rect 298008 220736 298060 220788
rect 302240 220736 302292 220788
rect 324780 220736 324832 220788
rect 363236 220736 363288 220788
rect 365996 220736 366048 220788
rect 380900 220736 380952 220788
rect 383384 220736 383436 220788
rect 502432 220736 502484 220788
rect 505008 220736 505060 220788
rect 623872 220736 623924 220788
rect 134984 220668 135036 220720
rect 57612 220600 57664 220652
rect 58624 220600 58676 220652
rect 128176 220600 128228 220652
rect 214196 220668 214248 220720
rect 215300 220668 215352 220720
rect 237748 220668 237800 220720
rect 270132 220668 270184 220720
rect 274456 220668 274508 220720
rect 276756 220668 276808 220720
rect 289084 220668 289136 220720
rect 291844 220668 291896 220720
rect 303068 220668 303120 220720
rect 311164 220668 311216 220720
rect 326252 220668 326304 220720
rect 366640 220668 366692 220720
rect 367744 220668 367796 220720
rect 390560 220668 390612 220720
rect 396724 220668 396776 220720
rect 517520 220668 517572 220720
rect 525064 220668 525116 220720
rect 577228 220668 577280 220720
rect 673368 220668 673420 220720
rect 676036 220668 676088 220720
rect 118332 220532 118384 220584
rect 218060 220600 218112 220652
rect 235908 220600 235960 220652
rect 270040 220600 270092 220652
rect 271420 220600 271472 220652
rect 275376 220600 275428 220652
rect 303436 220600 303488 220652
rect 312820 220600 312872 220652
rect 329564 220600 329616 220652
rect 371700 220600 371752 220652
rect 371884 220600 371936 220652
rect 385960 220600 386012 220652
rect 388444 220600 388496 220652
rect 512828 220600 512880 220652
rect 552664 220600 552716 220652
rect 632336 220600 632388 220652
rect 121276 220464 121328 220516
rect 206192 220464 206244 220516
rect 216680 220532 216732 220584
rect 231032 220532 231084 220584
rect 268292 220532 268344 220584
rect 273076 220532 273128 220584
rect 276664 220532 276716 220584
rect 293224 220532 293276 220584
rect 294328 220532 294380 220584
rect 299296 220532 299348 220584
rect 303620 220532 303672 220584
rect 306196 220532 306248 220584
rect 317880 220532 317932 220584
rect 329656 220532 329708 220584
rect 373356 220532 373408 220584
rect 375288 220532 375340 220584
rect 379520 220532 379572 220584
rect 379612 220532 379664 220584
rect 394700 220532 394752 220584
rect 395712 220532 395764 220584
rect 520004 220532 520056 220584
rect 208216 220464 208268 220516
rect 111616 220396 111668 220448
rect 206928 220396 206980 220448
rect 145196 220328 145248 220380
rect 146208 220328 146260 220380
rect 155316 220328 155368 220380
rect 155868 220328 155920 220380
rect 168748 220328 168800 220380
rect 169668 220328 169720 220380
rect 178868 220328 178920 220380
rect 179328 220328 179380 220380
rect 192300 220328 192352 220380
rect 224960 220464 225012 220516
rect 229376 220464 229428 220516
rect 262588 220464 262640 220516
rect 262956 220464 263008 220516
rect 263508 220464 263560 220516
rect 304816 220464 304868 220516
rect 316132 220464 316184 220516
rect 322204 220464 322256 220516
rect 342996 220464 343048 220516
rect 343088 220464 343140 220516
rect 386788 220464 386840 220516
rect 392584 220464 392636 220516
rect 522580 220464 522632 220516
rect 560576 220464 560628 220516
rect 574744 220532 574796 220584
rect 575480 220532 575532 220584
rect 576400 220464 576452 220516
rect 222568 220396 222620 220448
rect 264336 220396 264388 220448
rect 299388 220396 299440 220448
rect 305276 220396 305328 220448
rect 306104 220396 306156 220448
rect 319536 220396 319588 220448
rect 330852 220396 330904 220448
rect 375380 220396 375432 220448
rect 376024 220396 376076 220448
rect 224316 220328 224368 220380
rect 265440 220328 265492 220380
rect 307576 220328 307628 220380
rect 321560 220328 321612 220380
rect 332232 220328 332284 220380
rect 376208 220328 376260 220380
rect 377312 220396 377364 220448
rect 388536 220396 388588 220448
rect 394608 220396 394660 220448
rect 527272 220396 527324 220448
rect 379612 220328 379664 220380
rect 395620 220328 395672 220380
rect 79600 220260 79652 220312
rect 100760 220260 100812 220312
rect 104716 220260 104768 220312
rect 203708 220260 203760 220312
rect 206192 220260 206244 220312
rect 213920 220260 213972 220312
rect 217600 220260 217652 220312
rect 260104 220260 260156 220312
rect 264704 220260 264756 220312
rect 273812 220260 273864 220312
rect 283196 220260 283248 220312
rect 284208 220260 284260 220312
rect 291568 220260 291620 220312
rect 293960 220260 294012 220312
rect 307392 220260 307444 220312
rect 322940 220260 322992 220312
rect 331036 220260 331088 220312
rect 376944 220260 376996 220312
rect 378692 220260 378744 220312
rect 391940 220260 391992 220312
rect 396816 220260 396868 220312
rect 415308 220328 415360 220380
rect 418160 220328 418212 220380
rect 574192 220328 574244 220380
rect 94780 220192 94832 220244
rect 202420 220192 202472 220244
rect 81256 220124 81308 220176
rect 204536 220192 204588 220244
rect 207480 220192 207532 220244
rect 213828 220192 213880 220244
rect 215852 220192 215904 220244
rect 261484 220192 261536 220244
rect 262588 220192 262640 220244
rect 267188 220192 267240 220244
rect 304908 220192 304960 220244
rect 314660 220192 314712 220244
rect 315396 220192 315448 220244
rect 332968 220192 333020 220244
rect 333888 220192 333940 220244
rect 381820 220192 381872 220244
rect 382280 220192 382332 220244
rect 396908 220192 396960 220244
rect 532700 220260 532752 220312
rect 560576 220260 560628 220312
rect 577136 220464 577188 220516
rect 535368 220192 535420 220244
rect 605932 220192 605984 220244
rect 674656 220192 674708 220244
rect 676036 220192 676088 220244
rect 204076 220124 204128 220176
rect 209872 220124 209924 220176
rect 210792 220124 210844 220176
rect 64512 220056 64564 220108
rect 192852 220056 192904 220108
rect 209136 220056 209188 220108
rect 252100 220056 252152 220108
rect 254584 220124 254636 220176
rect 255228 220124 255280 220176
rect 257896 220124 257948 220176
rect 271236 220124 271288 220176
rect 255964 220056 256016 220108
rect 266176 220056 266228 220108
rect 279424 220124 279476 220176
rect 280620 220124 280672 220176
rect 281448 220124 281500 220176
rect 278596 220056 278648 220108
rect 287520 220124 287572 220176
rect 308772 220124 308824 220176
rect 326252 220124 326304 220176
rect 332416 220124 332468 220176
rect 380072 220124 380124 220176
rect 380164 220124 380216 220176
rect 395252 220124 395304 220176
rect 398564 220124 398616 220176
rect 537392 220124 537444 220176
rect 548156 220124 548208 220176
rect 615500 220124 615552 220176
rect 284852 220056 284904 220108
rect 285496 220056 285548 220108
rect 301964 220056 302016 220108
rect 309416 220056 309468 220108
rect 310244 220056 310296 220108
rect 329840 220056 329892 220108
rect 333796 220056 333848 220108
rect 383660 220056 383712 220108
rect 385684 220056 385736 220108
rect 400312 220056 400364 220108
rect 404268 220056 404320 220108
rect 549996 220056 550048 220108
rect 551284 220056 551336 220108
rect 609612 220056 609664 220108
rect 148600 219988 148652 220040
rect 223120 219988 223172 220040
rect 247868 219988 247920 220040
rect 248328 219988 248380 220040
rect 151728 219920 151780 219972
rect 224040 219920 224092 219972
rect 246120 219920 246172 219972
rect 246948 219920 247000 219972
rect 272892 219988 272944 220040
rect 289636 219988 289688 220040
rect 292856 219988 292908 220040
rect 319352 219988 319404 220040
rect 339684 219988 339736 220040
rect 341524 219988 341576 220040
rect 370044 219988 370096 220040
rect 370228 219988 370280 220040
rect 382648 219988 382700 220040
rect 384948 219988 385000 220040
rect 505008 219988 505060 220040
rect 543004 219988 543056 220040
rect 614120 219988 614172 220040
rect 158628 219852 158680 219904
rect 227352 219852 227404 219904
rect 242808 219852 242860 219904
rect 249524 219852 249576 219904
rect 276204 219920 276256 219972
rect 318064 219920 318116 219972
rect 336740 219920 336792 219972
rect 340144 219920 340196 219972
rect 360200 219920 360252 219972
rect 363144 219920 363196 219972
rect 391020 219920 391072 219972
rect 391112 219920 391164 219972
rect 509884 219920 509936 219972
rect 540428 219920 540480 219972
rect 613384 219920 613436 219972
rect 252928 219852 252980 219904
rect 277584 219852 277636 219904
rect 338764 219852 338816 219904
rect 356520 219852 356572 219904
rect 365352 219852 365404 219904
rect 377588 219852 377640 219904
rect 386972 219852 387024 219904
rect 398840 219852 398892 219904
rect 400680 219852 400732 219904
rect 513840 219852 513892 219904
rect 517520 219852 517572 219904
rect 574836 219852 574888 219904
rect 673276 219852 673328 219904
rect 676036 219852 676088 219904
rect 165436 219784 165488 219836
rect 227720 219784 227772 219836
rect 256240 219784 256292 219836
rect 278964 219784 279016 219836
rect 337384 219784 337436 219836
rect 353300 219784 353352 219836
rect 362960 219784 363012 219836
rect 368480 219784 368532 219836
rect 376208 219784 376260 219836
rect 378416 219784 378468 219836
rect 379704 219784 379756 219836
rect 484400 219784 484452 219836
rect 529940 219784 529992 219836
rect 612004 219784 612056 219836
rect 172152 219716 172204 219768
rect 232412 219716 232464 219768
rect 250996 219716 251048 219768
rect 271328 219716 271380 219768
rect 334716 219716 334768 219768
rect 349804 219716 349856 219768
rect 372620 219716 372672 219768
rect 384304 219716 384356 219768
rect 387248 219716 387300 219768
rect 409880 219716 409932 219768
rect 409972 219716 410024 219768
rect 416228 219716 416280 219768
rect 515404 219716 515456 219768
rect 625252 219716 625304 219768
rect 185584 219648 185636 219700
rect 186964 219648 187016 219700
rect 181996 219580 182048 219632
rect 232780 219648 232832 219700
rect 252100 219648 252152 219700
rect 257344 219648 257396 219700
rect 268016 219648 268068 219700
rect 275284 219648 275336 219700
rect 334624 219648 334676 219700
rect 346492 219648 346544 219700
rect 378048 219648 378100 219700
rect 387800 219648 387852 219700
rect 512828 219648 512880 219700
rect 625528 219648 625580 219700
rect 188896 219580 188948 219632
rect 234620 219580 234672 219632
rect 261300 219580 261352 219632
rect 272984 219580 273036 219632
rect 300492 219580 300544 219632
rect 306932 219580 306984 219632
rect 406384 219580 406436 219632
rect 412916 219580 412968 219632
rect 509884 219580 509936 219632
rect 623780 219580 623832 219632
rect 61108 219512 61160 219564
rect 66904 219512 66956 219564
rect 97816 219512 97868 219564
rect 195704 219512 195756 219564
rect 234712 219512 234764 219564
rect 301596 219512 301648 219564
rect 307760 219512 307812 219564
rect 408500 219512 408552 219564
rect 414572 219512 414624 219564
rect 502432 219512 502484 219564
rect 622952 219512 623004 219564
rect 195152 219444 195204 219496
rect 202420 219444 202472 219496
rect 237380 219444 237432 219496
rect 267188 219444 267240 219496
rect 268384 219444 268436 219496
rect 276480 219444 276532 219496
rect 278044 219444 278096 219496
rect 300584 219444 300636 219496
rect 306380 219444 306432 219496
rect 360292 219444 360344 219496
rect 364984 219444 365036 219496
rect 371332 219444 371384 219496
rect 375932 219444 375984 219496
rect 378508 219444 378560 219496
rect 385132 219444 385184 219496
rect 390652 219444 390704 219496
rect 393596 219444 393648 219496
rect 394516 219444 394568 219496
rect 529940 219444 529992 219496
rect 565452 219444 565504 219496
rect 354404 219376 354456 219428
rect 432236 219376 432288 219428
rect 577044 219444 577096 219496
rect 353208 219308 353260 219360
rect 430580 219308 430632 219360
rect 379428 219240 379480 219292
rect 494520 219240 494572 219292
rect 380808 219172 380860 219224
rect 498200 219172 498252 219224
rect 567936 219172 567988 219224
rect 616788 219172 616840 219224
rect 383568 219104 383620 219156
rect 501236 219104 501288 219156
rect 545764 219104 545816 219156
rect 576308 219104 576360 219156
rect 383476 219036 383528 219088
rect 503720 219036 503772 219088
rect 543188 219036 543240 219088
rect 543648 219036 543700 219088
rect 576216 219036 576268 219088
rect 386328 218968 386380 219020
rect 508780 218968 508832 219020
rect 541440 218968 541492 219020
rect 576124 218968 576176 219020
rect 35716 218900 35768 218952
rect 55956 218900 56008 218952
rect 387708 218900 387760 218952
rect 511356 218900 511408 218952
rect 570604 218900 570656 218952
rect 617524 218900 617576 218952
rect 47584 218832 47636 218884
rect 647148 218832 647200 218884
rect 55864 218764 55916 218816
rect 656900 218764 656952 218816
rect 45008 218696 45060 218748
rect 662512 218696 662564 218748
rect 553676 218628 553728 218680
rect 576032 218628 576084 218680
rect 518164 218560 518216 218612
rect 518440 218560 518492 218612
rect 575940 218560 575992 218612
rect 515496 218492 515548 218544
rect 516048 218492 516100 218544
rect 608416 218492 608468 218544
rect 511264 218424 511316 218476
rect 609888 218424 609940 218476
rect 487804 218356 487856 218408
rect 606668 218356 606720 218408
rect 489368 218288 489420 218340
rect 489828 218288 489880 218340
rect 620284 218288 620336 218340
rect 499672 218220 499724 218272
rect 500224 218220 500276 218272
rect 636016 218220 636068 218272
rect 493416 218152 493468 218204
rect 629944 218152 629996 218204
rect 486424 218084 486476 218136
rect 487528 218016 487580 218068
rect 487804 218016 487856 218068
rect 496084 218084 496136 218136
rect 636108 218084 636160 218136
rect 638316 218016 638368 218068
rect 523040 217880 523092 217932
rect 523960 217880 524012 217932
rect 538220 217880 538272 217932
rect 539048 217880 539100 217932
rect 296720 217812 296772 217864
rect 297640 217812 297692 217864
rect 299572 217812 299624 217864
rect 300216 217812 300268 217864
rect 331220 217812 331272 217864
rect 332140 217812 332192 217864
rect 333980 217812 334032 217864
rect 334716 217812 334768 217864
rect 350632 217812 350684 217864
rect 351460 217812 351512 217864
rect 434720 217812 434772 217864
rect 435640 217812 435692 217864
rect 441620 217812 441672 217864
rect 442356 217812 442408 217864
rect 454040 217812 454092 217864
rect 454960 217812 455012 217864
rect 460940 217812 460992 217864
rect 461676 217812 461728 217864
rect 465080 217812 465132 217864
rect 465908 217812 465960 217864
rect 471980 217812 472032 217864
rect 472624 217812 472676 217864
rect 476120 217812 476172 217864
rect 476856 217812 476908 217864
rect 491392 217812 491444 217864
rect 492588 217812 492640 217864
rect 619916 217812 619968 217864
rect 508412 217744 508464 217796
rect 575848 217744 575900 217796
rect 561772 217676 561824 217728
rect 562876 217676 562928 217728
rect 634544 217676 634596 217728
rect 560300 217608 560352 217660
rect 634084 217608 634136 217660
rect 557816 217540 557868 217592
rect 633624 217540 633676 217592
rect 545212 217472 545264 217524
rect 621020 217472 621072 217524
rect 555700 217404 555752 217456
rect 633164 217404 633216 217456
rect 499580 217336 499632 217388
rect 500868 217336 500920 217388
rect 576952 217336 577004 217388
rect 35624 217268 35676 217320
rect 46296 217268 46348 217320
rect 52184 217268 52236 217320
rect 164884 217268 164936 217320
rect 550548 217268 550600 217320
rect 629208 217268 629260 217320
rect 497648 217200 497700 217252
rect 575756 217200 575808 217252
rect 537852 217132 537904 217184
rect 618996 217132 619048 217184
rect 532976 217064 533028 217116
rect 618168 217064 618220 217116
rect 513656 216996 513708 217048
rect 610808 216996 610860 217048
rect 506112 216928 506164 216980
rect 607496 216928 607548 216980
rect 502524 216860 502576 216912
rect 503536 216860 503588 216912
rect 608508 216860 608560 216912
rect 494336 216792 494388 216844
rect 607588 216792 607640 216844
rect 499120 216724 499172 216776
rect 622584 216724 622636 216776
rect 566648 216656 566700 216708
rect 575664 216656 575716 216708
rect 490932 216384 490984 216436
rect 521200 216384 521252 216436
rect 523776 216384 523828 216436
rect 526260 216384 526312 216436
rect 528560 216384 528612 216436
rect 531228 216384 531280 216436
rect 533804 216384 533856 216436
rect 536380 216384 536432 216436
rect 538864 216384 538916 216436
rect 548984 216384 549036 216436
rect 556528 216384 556580 216436
rect 561588 216384 561640 216436
rect 615500 216452 615552 216504
rect 631784 216452 631836 216504
rect 574192 216384 574244 216436
rect 574836 216384 574888 216436
rect 613384 216384 613436 216436
rect 630404 216384 630456 216436
rect 612004 216316 612056 216368
rect 628472 216316 628524 216368
rect 614120 216248 614172 216300
rect 630864 216248 630916 216300
rect 626172 216180 626224 216232
rect 628012 216112 628064 216164
rect 674380 216112 674432 216164
rect 676036 216112 676088 216164
rect 577872 216044 577924 216096
rect 605932 216044 605984 216096
rect 629484 216044 629536 216096
rect 619640 215976 619692 216028
rect 618720 215908 618772 215960
rect 676220 215908 676272 215960
rect 676864 215908 676916 215960
rect 615500 215840 615552 215892
rect 615040 215772 615092 215824
rect 614580 215704 614632 215756
rect 674472 215704 674524 215756
rect 676036 215704 676088 215756
rect 614028 215636 614080 215688
rect 613568 215568 613620 215620
rect 613108 215500 613160 215552
rect 612648 215432 612700 215484
rect 612188 215364 612240 215416
rect 607128 215296 607180 215348
rect 577136 214820 577188 214872
rect 627092 214820 627144 214872
rect 577228 214684 577280 214736
rect 627552 214684 627604 214736
rect 576400 214616 576452 214668
rect 626632 214616 626684 214668
rect 35808 214548 35860 214600
rect 43628 214548 43680 214600
rect 577044 214548 577096 214600
rect 635004 214548 635056 214600
rect 48964 214344 49016 214396
rect 665272 214344 665324 214396
rect 46572 214276 46624 214328
rect 668952 214276 669004 214328
rect 40868 214208 40920 214260
rect 666192 214208 666244 214260
rect 42800 214140 42852 214192
rect 668124 214140 668176 214192
rect 40684 214072 40736 214124
rect 665732 214072 665784 214124
rect 673184 214072 673236 214124
rect 676036 214072 676088 214124
rect 41788 214004 41840 214056
rect 668860 214004 668912 214056
rect 41328 213936 41380 213988
rect 668768 213936 668820 213988
rect 576952 213868 577004 213920
rect 608508 213868 608560 213920
rect 636108 213868 636160 213920
rect 637396 213868 637448 213920
rect 638224 213868 638276 213920
rect 640616 213868 640668 213920
rect 575756 213800 575808 213852
rect 608048 213800 608100 213852
rect 609612 213800 609664 213852
rect 617800 213800 617852 213852
rect 619916 213800 619968 213852
rect 622032 213800 622084 213852
rect 629944 213800 629996 213852
rect 636568 213800 636620 213852
rect 636844 213800 636896 213852
rect 639236 213800 639288 213852
rect 575848 213732 575900 213784
rect 609888 213732 609940 213784
rect 610348 213732 610400 213784
rect 621480 213732 621532 213784
rect 636016 213732 636068 213784
rect 637856 213732 637908 213784
rect 575940 213664 575992 213716
rect 611728 213664 611780 213716
rect 621020 213664 621072 213716
rect 631324 213664 631376 213716
rect 674564 213664 674616 213716
rect 676036 213664 676088 213716
rect 577872 213596 577924 213648
rect 617340 213596 617392 213648
rect 618168 213596 618220 213648
rect 628932 213596 628984 213648
rect 629208 213596 629260 213648
rect 632244 213596 632296 213648
rect 576124 213528 576176 213580
rect 615960 213528 616012 213580
rect 618996 213528 619048 213580
rect 629944 213528 629996 213580
rect 576216 213460 576268 213512
rect 616420 213460 616472 213512
rect 616788 213460 616840 213512
rect 635464 213460 635516 213512
rect 576308 213392 576360 213444
rect 616880 213392 616932 213444
rect 617524 213392 617576 213444
rect 635924 213392 635976 213444
rect 576032 213324 576084 213376
rect 618260 213324 618312 213376
rect 620284 213324 620336 213376
rect 636384 213324 636436 213376
rect 575664 213256 575716 213308
rect 620560 213256 620612 213308
rect 623044 213256 623096 213308
rect 641076 213256 641128 213308
rect 642732 213256 642784 213308
rect 650000 213256 650052 213308
rect 577504 213188 577556 213240
rect 640156 213188 640208 213240
rect 643836 213188 643888 213240
rect 651380 213188 651432 213240
rect 607496 213120 607548 213172
rect 609428 213120 609480 213172
rect 608416 213052 608468 213104
rect 611268 213052 611320 213104
rect 646964 212984 647016 213036
rect 651472 212984 651524 213036
rect 645584 212576 645636 212628
rect 650092 212576 650144 212628
rect 623780 212372 623832 212424
rect 624424 212372 624476 212424
rect 625252 212372 625304 212424
rect 625712 212372 625764 212424
rect 663800 212372 663852 212424
rect 664444 212372 664496 212424
rect 663892 212304 663944 212356
rect 664352 212304 664404 212356
rect 671436 211148 671488 211200
rect 676036 211148 676088 211200
rect 662420 210536 662472 210588
rect 663064 210536 663116 210588
rect 652024 210400 652076 210452
rect 667204 210400 667256 210452
rect 580264 209788 580316 209840
rect 638408 209788 638460 209840
rect 579068 209720 579120 209772
rect 603172 209720 603224 209772
rect 578884 209652 578936 209704
rect 603080 209652 603132 209704
rect 665456 209652 665508 209704
rect 666928 209652 666980 209704
rect 578976 208292 579028 208344
rect 603080 208292 603132 208344
rect 578424 206932 578476 206984
rect 603080 206932 603132 206984
rect 578516 205572 578568 205624
rect 603080 205572 603132 205624
rect 579528 205504 579580 205556
rect 603172 205504 603224 205556
rect 578792 204212 578844 204264
rect 603080 204212 603132 204264
rect 35808 202852 35860 202904
rect 48964 202852 49016 202904
rect 579436 202784 579488 202836
rect 603080 202784 603132 202836
rect 674380 201832 674432 201884
rect 675392 201832 675444 201884
rect 579252 201424 579304 201476
rect 603172 201424 603224 201476
rect 674472 201424 674524 201476
rect 675392 201424 675444 201476
rect 578884 201356 578936 201408
rect 603080 201356 603132 201408
rect 675116 200676 675168 200728
rect 675392 200676 675444 200728
rect 578240 200064 578292 200116
rect 603080 200064 603132 200116
rect 578424 198636 578476 198688
rect 603080 198636 603132 198688
rect 673184 197412 673236 197464
rect 675484 197412 675536 197464
rect 579068 197276 579120 197328
rect 603172 197276 603224 197328
rect 674840 197004 674892 197056
rect 675392 197004 675444 197056
rect 579528 196596 579580 196648
rect 603080 196596 603132 196648
rect 674564 196528 674616 196580
rect 675392 196528 675444 196580
rect 579528 195236 579580 195288
rect 603080 195236 603132 195288
rect 579528 193808 579580 193860
rect 603080 193808 603132 193860
rect 42064 193128 42116 193180
rect 44456 193128 44508 193180
rect 579528 192448 579580 192500
rect 603080 192448 603132 192500
rect 674840 192448 674892 192500
rect 675392 192448 675444 192500
rect 579252 191836 579304 191888
rect 603080 191836 603132 191888
rect 42064 191632 42116 191684
rect 42984 191632 43036 191684
rect 42156 191564 42208 191616
rect 44364 191564 44416 191616
rect 42156 190816 42208 190868
rect 43076 190816 43128 190868
rect 675760 190612 675812 190664
rect 578240 190476 578292 190528
rect 603080 190476 603132 190528
rect 675760 190340 675812 190392
rect 579528 189116 579580 189168
rect 603080 189116 603132 189168
rect 579252 189048 579304 189100
rect 603172 189048 603224 189100
rect 578792 187688 578844 187740
rect 603080 187688 603132 187740
rect 42156 187620 42208 187672
rect 44272 187620 44324 187672
rect 579344 186328 579396 186380
rect 603080 186328 603132 186380
rect 42064 186260 42116 186312
rect 42892 186260 42944 186312
rect 42156 185852 42208 185904
rect 42800 185852 42852 185904
rect 578976 184968 579028 185020
rect 603080 184968 603132 185020
rect 579068 184900 579120 184952
rect 603172 184900 603224 184952
rect 668308 184152 668360 184204
rect 671344 184152 671396 184204
rect 579252 183540 579304 183592
rect 603080 183540 603132 183592
rect 42156 183404 42208 183456
rect 44180 183404 44232 183456
rect 578240 182180 578292 182232
rect 603080 182180 603132 182232
rect 578332 180888 578384 180940
rect 603172 180888 603224 180940
rect 578424 180820 578476 180872
rect 603080 180820 603132 180872
rect 578792 179392 578844 179444
rect 603080 179392 603132 179444
rect 667940 178780 667992 178832
rect 670056 178780 670108 178832
rect 673000 178168 673052 178220
rect 676036 178168 676088 178220
rect 578700 178032 578752 178084
rect 603080 178032 603132 178084
rect 674104 178032 674156 178084
rect 676036 178032 676088 178084
rect 672632 176944 672684 176996
rect 676036 176944 676088 176996
rect 671620 176808 671672 176860
rect 675944 176808 675996 176860
rect 579436 176740 579488 176792
rect 603172 176740 603224 176792
rect 674012 176740 674064 176792
rect 676036 176740 676088 176792
rect 579252 176672 579304 176724
rect 603080 176672 603132 176724
rect 672540 176468 672592 176520
rect 676036 176468 676088 176520
rect 674564 175992 674616 176044
rect 676036 175992 676088 176044
rect 674656 175652 674708 175704
rect 676036 175652 676088 175704
rect 581644 175244 581696 175296
rect 603080 175244 603132 175296
rect 674564 175176 674616 175228
rect 676036 175176 676088 175228
rect 673368 174360 673420 174412
rect 676036 174360 676088 174412
rect 580356 173884 580408 173936
rect 603080 173884 603132 173936
rect 667940 173612 667992 173664
rect 670148 173612 670200 173664
rect 579160 172524 579212 172576
rect 603080 172524 603132 172576
rect 674840 172524 674892 172576
rect 676036 172524 676088 172576
rect 579344 171096 579396 171148
rect 603080 171096 603132 171148
rect 674472 170280 674524 170332
rect 676036 170280 676088 170332
rect 578976 169804 579028 169856
rect 603080 169804 603132 169856
rect 579068 169736 579120 169788
rect 603172 169736 603224 169788
rect 673184 169464 673236 169516
rect 676036 169464 676088 169516
rect 674380 169056 674432 169108
rect 676036 169056 676088 169108
rect 673276 168648 673328 168700
rect 676036 168648 676088 168700
rect 578884 168376 578936 168428
rect 603080 168376 603132 168428
rect 674104 168240 674156 168292
rect 676036 168240 676088 168292
rect 673000 167832 673052 167884
rect 676036 167832 676088 167884
rect 583116 167016 583168 167068
rect 603080 167016 603132 167068
rect 671344 167016 671396 167068
rect 676036 167016 676088 167068
rect 578700 166676 578752 166728
rect 581644 166676 581696 166728
rect 581736 165588 581788 165640
rect 603080 165588 603132 165640
rect 578240 164568 578292 164620
rect 580356 164568 580408 164620
rect 581644 164228 581696 164280
rect 603080 164228 603132 164280
rect 579528 164160 579580 164212
rect 603724 164160 603776 164212
rect 668400 163956 668452 164008
rect 672724 163956 672776 164008
rect 580356 162868 580408 162920
rect 603080 162868 603132 162920
rect 583024 161440 583076 161492
rect 603080 161440 603132 161492
rect 674840 160760 674892 160812
rect 675484 160760 675536 160812
rect 579436 160080 579488 160132
rect 603080 160080 603132 160132
rect 579344 158720 579396 158772
rect 603080 158720 603132 158772
rect 585876 157428 585928 157480
rect 603080 157428 603132 157480
rect 584404 157360 584456 157412
rect 603172 157360 603224 157412
rect 587256 155932 587308 155984
rect 603080 155932 603132 155984
rect 673184 155456 673236 155508
rect 675484 155456 675536 155508
rect 578516 154640 578568 154692
rect 583116 154640 583168 154692
rect 579160 154572 579212 154624
rect 603080 154572 603132 154624
rect 579068 153280 579120 153332
rect 603172 153280 603224 153332
rect 578976 153212 579028 153264
rect 603080 153212 603132 153264
rect 579252 153076 579304 153128
rect 581736 153076 581788 153128
rect 579252 152940 579304 152992
rect 579436 152940 579488 152992
rect 674380 152532 674432 152584
rect 675392 152532 675444 152584
rect 587164 151784 587216 151836
rect 603080 151784 603132 151836
rect 579528 151716 579580 151768
rect 603816 151716 603868 151768
rect 673276 151376 673328 151428
rect 675392 151376 675444 151428
rect 578884 150424 578936 150476
rect 603080 150424 603132 150476
rect 674472 150356 674524 150408
rect 675392 150356 675444 150408
rect 579436 150220 579488 150272
rect 581644 150220 581696 150272
rect 592776 149132 592828 149184
rect 603080 149132 603132 149184
rect 589924 149064 589976 149116
rect 603172 149064 603224 149116
rect 578516 148656 578568 148708
rect 580356 148656 580408 148708
rect 668308 148520 668360 148572
rect 674196 148520 674248 148572
rect 584588 147636 584640 147688
rect 603080 147636 603132 147688
rect 578516 147296 578568 147348
rect 580264 147296 580316 147348
rect 588544 146276 588596 146328
rect 603080 146276 603132 146328
rect 579528 146072 579580 146124
rect 583024 146072 583076 146124
rect 583116 144916 583168 144968
rect 603172 144916 603224 144968
rect 578608 144848 578660 144900
rect 603724 144848 603776 144900
rect 580356 143556 580408 143608
rect 603080 143556 603132 143608
rect 667940 143284 667992 143336
rect 670240 143284 670292 143336
rect 579528 142604 579580 142656
rect 584404 142604 584456 142656
rect 585784 142128 585836 142180
rect 603080 142128 603132 142180
rect 591304 140768 591356 140820
rect 603080 140768 603132 140820
rect 584404 139408 584456 139460
rect 603080 139408 603132 139460
rect 668032 138184 668084 138236
rect 672816 138184 672868 138236
rect 598296 138048 598348 138100
rect 603172 138048 603224 138100
rect 583024 137980 583076 138032
rect 603080 137980 603132 138032
rect 579528 137912 579580 137964
rect 587256 137912 587308 137964
rect 581644 136620 581696 136672
rect 603080 136620 603132 136672
rect 579528 136484 579580 136536
rect 585876 136484 585928 136536
rect 587348 135260 587400 135312
rect 603080 135260 603132 135312
rect 580264 133900 580316 133952
rect 603080 133900 603132 133952
rect 668584 132948 668636 133000
rect 674288 132948 674340 133000
rect 672908 132880 672960 132932
rect 676036 132880 676088 132932
rect 671528 132744 671580 132796
rect 676220 132744 676272 132796
rect 667204 132608 667256 132660
rect 676128 132608 676180 132660
rect 590016 132472 590068 132524
rect 603080 132472 603132 132524
rect 674012 132268 674064 132320
rect 676220 132268 676272 132320
rect 588636 131724 588688 131776
rect 603172 131724 603224 131776
rect 674656 131316 674708 131368
rect 676036 131316 676088 131368
rect 596916 131112 596968 131164
rect 603080 131112 603132 131164
rect 668676 131112 668728 131164
rect 668952 131112 669004 131164
rect 676220 131112 676272 131164
rect 579252 131044 579304 131096
rect 587164 131044 587216 131096
rect 674564 130500 674616 130552
rect 676036 130500 676088 130552
rect 672724 129888 672776 129940
rect 676220 129888 676272 129940
rect 585876 129752 585928 129804
rect 603080 129752 603132 129804
rect 668584 129752 668636 129804
rect 668860 129752 668912 129804
rect 676220 129752 676272 129804
rect 581736 129004 581788 129056
rect 603908 129004 603960 129056
rect 673368 128528 673420 128580
rect 676128 128528 676180 128580
rect 594064 128324 594116 128376
rect 603080 128324 603132 128376
rect 668768 128324 668820 128376
rect 676220 128324 676272 128376
rect 578884 128256 578936 128308
rect 584588 128256 584640 128308
rect 668032 128120 668084 128172
rect 673092 128120 673144 128172
rect 584496 126964 584548 127016
rect 603080 126964 603132 127016
rect 675116 126964 675168 127016
rect 676036 126964 676088 127016
rect 579068 126896 579120 126948
rect 592776 126896 592828 126948
rect 601056 125672 601108 125724
rect 603080 125672 603132 125724
rect 592684 125604 592736 125656
rect 603172 125604 603224 125656
rect 578424 125536 578476 125588
rect 589924 125536 589976 125588
rect 591396 124176 591448 124228
rect 603080 124176 603132 124228
rect 579252 124108 579304 124160
rect 588544 124108 588596 124160
rect 667940 123836 667992 123888
rect 671436 123836 671488 123888
rect 673368 122952 673420 123004
rect 676220 122952 676272 123004
rect 589924 122816 589976 122868
rect 603080 122816 603132 122868
rect 668860 122816 668912 122868
rect 676220 122816 676272 122868
rect 587256 121456 587308 121508
rect 603080 121456 603132 121508
rect 670148 121456 670200 121508
rect 676128 121456 676180 121508
rect 579528 121388 579580 121440
rect 583116 121388 583168 121440
rect 670056 120708 670108 120760
rect 676220 120708 676272 120760
rect 588544 120096 588596 120148
rect 603080 120096 603132 120148
rect 579252 120028 579304 120080
rect 581736 120028 581788 120080
rect 579160 118668 579212 118720
rect 603080 118668 603132 118720
rect 578608 118396 578660 118448
rect 580356 118396 580408 118448
rect 669228 117784 669280 117836
rect 674104 117784 674156 117836
rect 579068 117308 579120 117360
rect 603080 117308 603132 117360
rect 579528 117240 579580 117292
rect 603724 117240 603776 117292
rect 668492 117240 668544 117292
rect 673000 117240 673052 117292
rect 675208 116560 675260 116612
rect 683304 116560 683356 116612
rect 674656 116220 674708 116272
rect 677600 116220 677652 116272
rect 600964 115948 601016 116000
rect 603448 115948 603500 116000
rect 579528 115540 579580 115592
rect 585784 115540 585836 115592
rect 678244 116152 678296 116204
rect 675116 115540 675168 115592
rect 675392 115540 675444 115592
rect 675116 115404 675168 115456
rect 675208 114792 675260 114844
rect 675392 114792 675444 114844
rect 599584 114588 599636 114640
rect 603172 114588 603224 114640
rect 674656 114588 674708 114640
rect 675116 114588 675168 114640
rect 578976 114520 579028 114572
rect 603080 114520 603132 114572
rect 579252 114452 579304 114504
rect 591304 114452 591356 114504
rect 668492 114316 668544 114368
rect 671344 114316 671396 114368
rect 578884 113160 578936 113212
rect 603080 113160 603132 113212
rect 578424 112616 578476 112668
rect 584404 112616 584456 112668
rect 583116 112412 583168 112464
rect 603816 112412 603868 112464
rect 598204 111800 598256 111852
rect 603080 111800 603132 111852
rect 578700 111732 578752 111784
rect 598296 111732 598348 111784
rect 667940 111256 667992 111308
rect 670148 111256 670200 111308
rect 675208 111120 675260 111172
rect 675392 111120 675444 111172
rect 675116 110644 675168 110696
rect 675392 110644 675444 110696
rect 595444 110440 595496 110492
rect 603080 110440 603132 110492
rect 667940 110304 667992 110356
rect 670056 110304 670108 110356
rect 579436 109556 579488 109608
rect 583024 109556 583076 109608
rect 587164 109012 587216 109064
rect 603080 109012 603132 109064
rect 579252 108740 579304 108792
rect 581644 108740 581696 108792
rect 581736 107652 581788 107704
rect 603080 107652 603132 107704
rect 579528 107584 579580 107636
rect 587348 107584 587400 107636
rect 675116 106972 675168 107024
rect 675392 106972 675444 107024
rect 675484 106564 675536 106616
rect 585784 106292 585836 106344
rect 603080 106292 603132 106344
rect 673368 106292 673420 106344
rect 579528 106224 579580 106276
rect 588636 106224 588688 106276
rect 674748 106224 674800 106276
rect 675392 106224 675444 106276
rect 669228 106088 669280 106140
rect 672724 106088 672776 106140
rect 584404 104864 584456 104916
rect 603080 104864 603132 104916
rect 596824 103912 596876 103964
rect 603172 103912 603224 103964
rect 578516 103436 578568 103488
rect 580264 103436 580316 103488
rect 583024 102212 583076 102264
rect 603172 102212 603224 102264
rect 581644 102144 581696 102196
rect 603080 102144 603132 102196
rect 578332 102076 578384 102128
rect 590016 102076 590068 102128
rect 580264 100716 580316 100768
rect 603080 100716 603132 100768
rect 578700 100648 578752 100700
rect 596916 100648 596968 100700
rect 591304 99356 591356 99408
rect 603080 99356 603132 99408
rect 579528 98880 579580 98932
rect 585876 98880 585928 98932
rect 580356 98608 580408 98660
rect 603816 98608 603868 98660
rect 625068 97928 625120 97980
rect 625988 97928 626040 97980
rect 634452 97928 634504 97980
rect 637580 97928 637632 97980
rect 638316 97928 638368 97980
rect 644664 97928 644716 97980
rect 663064 97928 663116 97980
rect 665364 97928 665416 97980
rect 624608 97860 624660 97912
rect 625804 97860 625856 97912
rect 633072 97860 633124 97912
rect 635280 97860 635332 97912
rect 633808 97792 633860 97844
rect 636384 97792 636436 97844
rect 647516 97792 647568 97844
rect 654784 97792 654836 97844
rect 637028 97724 637080 97776
rect 642180 97724 642232 97776
rect 632428 97656 632480 97708
rect 634084 97656 634136 97708
rect 635740 97656 635792 97708
rect 639880 97656 639932 97708
rect 579528 97588 579580 97640
rect 583116 97588 583168 97640
rect 631140 97588 631192 97640
rect 632152 97588 632204 97640
rect 637488 97588 637540 97640
rect 644572 97588 644624 97640
rect 635096 97520 635148 97572
rect 639052 97520 639104 97572
rect 614856 97452 614908 97504
rect 621664 97452 621716 97504
rect 643560 97452 643612 97504
rect 660396 97452 660448 97504
rect 620744 97384 620796 97436
rect 646044 97384 646096 97436
rect 649448 97384 649500 97436
rect 658832 97384 658884 97436
rect 648160 97316 648212 97368
rect 660120 97316 660172 97368
rect 622032 97248 622084 97300
rect 648804 97248 648856 97300
rect 652024 97248 652076 97300
rect 661960 97248 662012 97300
rect 621388 97180 621440 97232
rect 647424 97180 647476 97232
rect 654692 97180 654744 97232
rect 658372 97180 658424 97232
rect 659200 97180 659252 97232
rect 662512 97180 662564 97232
rect 623688 97112 623740 97164
rect 624424 97112 624476 97164
rect 657728 97112 657780 97164
rect 660672 97112 660724 97164
rect 662328 97112 662380 97164
rect 663984 97112 664036 97164
rect 610072 96908 610124 96960
rect 610900 96908 610952 96960
rect 616144 96908 616196 96960
rect 616788 96908 616840 96960
rect 617432 96908 617484 96960
rect 618168 96908 618220 96960
rect 622676 96908 622728 96960
rect 623596 96908 623648 96960
rect 625896 96908 625948 96960
rect 626448 96908 626500 96960
rect 644848 96908 644900 96960
rect 646504 96908 646556 96960
rect 650736 96908 650788 96960
rect 651196 96908 651248 96960
rect 655428 96908 655480 96960
rect 659292 96908 659344 96960
rect 618720 96840 618772 96892
rect 619548 96840 619600 96892
rect 620008 96840 620060 96892
rect 620928 96840 620980 96892
rect 640984 96840 641036 96892
rect 643284 96840 643336 96892
rect 660580 96840 660632 96892
rect 661408 96840 661460 96892
rect 655980 96772 656032 96824
rect 659568 96772 659620 96824
rect 631784 96704 631836 96756
rect 632980 96704 633032 96756
rect 636108 96704 636160 96756
rect 640984 96704 641036 96756
rect 661868 96704 661920 96756
rect 663064 96704 663116 96756
rect 578608 96568 578660 96620
rect 594064 96568 594116 96620
rect 640248 96568 640300 96620
rect 643192 96568 643244 96620
rect 656808 96568 656860 96620
rect 658280 96568 658332 96620
rect 638868 96500 638920 96552
rect 643100 96500 643152 96552
rect 656624 96160 656676 96212
rect 663892 96160 663944 96212
rect 646780 96024 646832 96076
rect 663800 96024 663852 96076
rect 653312 95956 653364 96008
rect 665272 95956 665324 96008
rect 639604 95888 639656 95940
rect 644480 95888 644532 95940
rect 646136 95888 646188 95940
rect 665180 95888 665232 95940
rect 641628 95820 641680 95872
rect 645860 95820 645912 95872
rect 607220 95480 607272 95532
rect 607680 95480 607732 95532
rect 657268 95208 657320 95260
rect 664076 95208 664128 95260
rect 578700 95140 578752 95192
rect 584496 95140 584548 95192
rect 579528 93780 579580 93832
rect 592684 93780 592736 93832
rect 646504 93100 646556 93152
rect 654876 93100 654928 93152
rect 579528 92420 579580 92472
rect 601056 92420 601108 92472
rect 644388 92420 644440 92472
rect 654324 92420 654376 92472
rect 579528 90992 579580 91044
rect 591396 90992 591448 91044
rect 579528 89632 579580 89684
rect 602436 89632 602488 89684
rect 616696 89632 616748 89684
rect 626448 89632 626500 89684
rect 656808 88816 656860 88868
rect 658096 88816 658148 88868
rect 662328 88816 662380 88868
rect 663984 88816 664036 88868
rect 616788 88272 616840 88324
rect 626448 88272 626500 88324
rect 659476 88272 659528 88324
rect 663156 88272 663208 88324
rect 620928 88204 620980 88256
rect 626356 88204 626408 88256
rect 579528 86912 579580 86964
rect 589924 86912 589976 86964
rect 651288 86844 651340 86896
rect 657176 86844 657228 86896
rect 649908 86776 649960 86828
rect 660672 86776 660724 86828
rect 651196 86708 651248 86760
rect 657728 86708 657780 86760
rect 652668 86640 652720 86692
rect 662512 86640 662564 86692
rect 645676 86572 645728 86624
rect 660120 86572 660172 86624
rect 648528 86504 648580 86556
rect 661408 86504 661460 86556
rect 653956 86436 654008 86488
rect 658832 86436 658884 86488
rect 619456 86232 619508 86284
rect 626448 86232 626500 86284
rect 579528 85484 579580 85536
rect 587256 85484 587308 85536
rect 619548 85484 619600 85536
rect 626448 85484 626500 85536
rect 579528 84124 579580 84176
rect 588544 84124 588596 84176
rect 618076 84124 618128 84176
rect 625620 84124 625672 84176
rect 618168 84056 618220 84108
rect 626448 84056 626500 84108
rect 578516 81336 578568 81388
rect 602344 81336 602396 81388
rect 579528 78616 579580 78668
rect 600964 78616 601016 78668
rect 626448 78140 626500 78192
rect 642456 78140 642508 78192
rect 631048 78072 631100 78124
rect 638960 78072 639012 78124
rect 629208 78004 629260 78056
rect 645308 78004 645360 78056
rect 605748 77936 605800 77988
rect 636752 77936 636804 77988
rect 628380 77596 628432 77648
rect 631508 77596 631560 77648
rect 579068 77324 579120 77376
rect 628380 77324 628432 77376
rect 576124 77256 576176 77308
rect 631048 77256 631100 77308
rect 623596 76576 623648 76628
rect 646320 76576 646372 76628
rect 624424 76508 624476 76560
rect 646964 76508 647016 76560
rect 579528 75828 579580 75880
rect 599584 75828 599636 75880
rect 623688 75216 623740 75268
rect 646136 75216 646188 75268
rect 615408 75148 615460 75200
rect 646872 75148 646924 75200
rect 646320 74468 646372 74520
rect 647240 74468 647292 74520
rect 579528 71680 579580 71732
rect 598204 71680 598256 71732
rect 623044 70388 623096 70440
rect 623780 70388 623832 70440
rect 579528 70320 579580 70372
rect 595444 70320 595496 70372
rect 578332 68892 578384 68944
rect 580356 68892 580408 68944
rect 579528 67532 579580 67584
rect 587164 67532 587216 67584
rect 579252 65764 579304 65816
rect 581736 65764 581788 65816
rect 579528 64268 579580 64320
rect 585784 64268 585836 64320
rect 579528 63452 579580 63504
rect 596824 63452 596876 63504
rect 578700 61344 578752 61396
rect 584404 61344 584456 61396
rect 578976 60664 579028 60716
rect 603724 60664 603776 60716
rect 618904 59848 618956 59900
rect 623044 59848 623096 59900
rect 578884 58760 578936 58812
rect 583024 58760 583076 58812
rect 621664 58624 621716 58676
rect 662420 58624 662472 58676
rect 578884 57876 578936 57928
rect 581644 57876 581696 57928
rect 578332 57196 578384 57248
rect 591304 57196 591356 57248
rect 578240 55632 578292 55684
rect 580264 55632 580316 55684
rect 616328 53796 616380 53848
rect 618904 53796 618956 53848
rect 52276 53116 52328 53168
rect 346308 53116 346360 53168
rect 145380 53048 145432 53100
rect 579068 53048 579120 53100
rect 347136 52368 347188 52420
rect 616328 52368 616380 52420
rect 52184 51688 52236 51740
rect 60740 51688 60792 51740
rect 60740 51008 60792 51060
rect 150348 51008 150400 51060
rect 189080 51008 189132 51060
rect 478144 49716 478196 49768
rect 478788 49716 478840 49768
rect 664444 49036 664496 49088
rect 669964 49036 670016 49088
rect 648157 46658 649617 47126
rect 241520 44956 241572 45008
rect 246120 44956 246172 45008
rect 251088 44888 251140 44940
rect 255872 44888 255924 44940
rect 241520 44820 241572 44872
rect 246120 44820 246172 44872
rect 405556 44820 405608 44872
rect 608784 44820 608836 44872
rect 251088 44752 251140 44804
rect 255872 44752 255924 44804
rect 473176 42476 473228 42528
<< metal2 >>
rect 110170 1029098 110262 1029126
rect 212934 1029098 213026 1029126
rect 264362 1029098 264454 1029126
rect 315974 1029098 316066 1029126
rect 366390 1029098 366482 1029126
rect 433734 1029098 433826 1029126
rect 510738 1029098 510830 1029126
rect 562166 1029098 562258 1029126
rect 110170 1028622 110262 1028650
rect 212934 1028622 213026 1028650
rect 264362 1028622 264454 1028650
rect 315974 1028622 316066 1028650
rect 366390 1028622 366482 1028650
rect 433734 1028622 433826 1028650
rect 510738 1028622 510830 1028650
rect 562166 1028622 562258 1028650
rect 110170 1028177 110262 1028205
rect 212934 1028177 213026 1028205
rect 264362 1028177 264454 1028205
rect 315974 1028177 316066 1028205
rect 366390 1028177 366482 1028205
rect 433734 1028177 433826 1028205
rect 510738 1028177 510830 1028205
rect 562166 1028177 562258 1028205
rect 366284 1027806 366496 1027834
rect 110170 1027738 110262 1027766
rect 212934 1027738 213026 1027766
rect 264362 1027738 264454 1027766
rect 315974 1027738 316066 1027766
rect 366284 1027752 366312 1027806
rect 366468 1027752 366496 1027806
rect 433734 1027738 433826 1027766
rect 510738 1027738 510830 1027766
rect 562166 1027738 562258 1027766
rect 110170 1027262 110262 1027290
rect 212934 1027262 213026 1027290
rect 264362 1027262 264454 1027290
rect 315974 1027262 316066 1027290
rect 366390 1027262 366482 1027290
rect 433734 1027262 433826 1027290
rect 510738 1027262 510830 1027290
rect 562166 1027262 562258 1027290
rect 110170 1026786 110262 1026814
rect 212934 1026786 213026 1026814
rect 264362 1026786 264454 1026814
rect 315974 1026786 316066 1026814
rect 366390 1026786 366482 1026814
rect 433734 1026786 433826 1026814
rect 510738 1026786 510830 1026814
rect 562166 1026786 562258 1026814
rect 110170 1026310 110262 1026338
rect 212934 1026310 213026 1026338
rect 264362 1026310 264454 1026338
rect 315974 1026310 316066 1026338
rect 366284 1026202 366312 1026324
rect 366468 1026202 366496 1026324
rect 433734 1026310 433826 1026338
rect 510738 1026310 510830 1026338
rect 562166 1026310 562258 1026338
rect 366284 1026174 366496 1026202
rect 366284 1026038 366496 1026066
rect 110170 1025902 110262 1025930
rect 212934 1025902 213026 1025930
rect 264362 1025902 264454 1025930
rect 315974 1025902 316066 1025930
rect 366284 1025916 366312 1026038
rect 366468 1025916 366496 1026038
rect 433734 1025902 433826 1025930
rect 510738 1025902 510830 1025930
rect 562166 1025902 562258 1025930
rect 110170 1025426 110262 1025454
rect 212934 1025426 213026 1025454
rect 264362 1025426 264454 1025454
rect 315974 1025426 316066 1025454
rect 366390 1025426 366482 1025454
rect 433734 1025426 433826 1025454
rect 510738 1025426 510830 1025454
rect 562166 1025426 562258 1025454
rect 110170 1024950 110262 1024978
rect 212934 1024950 213026 1024978
rect 264362 1024950 264454 1024978
rect 315974 1024950 316066 1024978
rect 366390 1024950 366482 1024978
rect 433734 1024950 433826 1024978
rect 510738 1024950 510830 1024978
rect 562166 1024950 562258 1024978
rect 110170 1024474 110262 1024502
rect 212934 1024474 213026 1024502
rect 264362 1024474 264454 1024502
rect 315974 1024474 316066 1024502
rect 366284 1024434 366312 1024488
rect 366468 1024434 366496 1024488
rect 433734 1024474 433826 1024502
rect 510738 1024474 510830 1024502
rect 562166 1024474 562258 1024502
rect 366284 1024406 366496 1024434
rect 110170 1024037 110262 1024065
rect 212934 1024037 213026 1024065
rect 264362 1024037 264454 1024065
rect 315974 1024037 316066 1024065
rect 366390 1024037 366482 1024065
rect 433734 1024037 433826 1024065
rect 510738 1024037 510830 1024065
rect 562166 1024037 562258 1024065
rect 110170 1023590 110262 1023618
rect 212934 1023590 213026 1023618
rect 264362 1023590 264454 1023618
rect 315974 1023590 316066 1023618
rect 366390 1023590 366482 1023618
rect 433734 1023590 433826 1023618
rect 510738 1023590 510830 1023618
rect 562166 1023590 562258 1023618
rect 154578 1007176 154634 1007185
rect 146944 1007140 146996 1007146
rect 154578 1007111 154580 1007120
rect 146944 1007082 146996 1007088
rect 154632 1007111 154634 1007120
rect 154580 1007082 154632 1007088
rect 95884 1006528 95936 1006534
rect 103612 1006528 103664 1006534
rect 95884 1006470 95936 1006476
rect 103150 1006496 103206 1006505
rect 94504 1006460 94556 1006466
rect 94504 1006402 94556 1006408
rect 93308 1006324 93360 1006330
rect 93308 1006266 93360 1006272
rect 93124 1006256 93176 1006262
rect 93124 1006198 93176 1006204
rect 92296 1001224 92348 1001230
rect 92296 1001166 92348 1001172
rect 92308 999274 92336 1001166
rect 92216 999246 92336 999274
rect 89628 995852 89680 995858
rect 89628 995794 89680 995800
rect 80978 995752 81034 995761
rect 80730 995710 80978 995738
rect 82358 995752 82414 995761
rect 82018 995710 82358 995738
rect 80978 995687 81034 995696
rect 89640 995738 89668 995794
rect 91560 995784 91612 995790
rect 86342 995722 86632 995738
rect 86342 995716 86644 995722
rect 86342 995710 86592 995716
rect 82358 995687 82414 995696
rect 89378 995710 89668 995738
rect 91218 995732 91560 995738
rect 91218 995726 91612 995732
rect 91218 995710 91600 995726
rect 92216 995722 92244 999246
rect 92296 999116 92348 999122
rect 92296 999058 92348 999064
rect 92308 995790 92336 999058
rect 92388 998436 92440 998442
rect 92388 998378 92440 998384
rect 92400 995858 92428 998378
rect 92664 997552 92716 997558
rect 92664 997494 92716 997500
rect 92480 997144 92532 997150
rect 92480 997086 92532 997092
rect 92388 995852 92440 995858
rect 92388 995794 92440 995800
rect 92296 995784 92348 995790
rect 92492 995761 92520 997086
rect 92572 997076 92624 997082
rect 92572 997018 92624 997024
rect 92296 995726 92348 995732
rect 92478 995752 92534 995761
rect 92204 995716 92256 995722
rect 86592 995658 86644 995664
rect 92478 995687 92534 995696
rect 92204 995658 92256 995664
rect 55864 995648 55916 995654
rect 84658 995616 84714 995625
rect 55864 995590 55916 995596
rect 46204 992928 46256 992934
rect 46204 992870 46256 992876
rect 44824 991500 44876 991506
rect 44824 991442 44876 991448
rect 42708 975724 42760 975730
rect 42708 975666 42760 975672
rect 41800 968833 41828 969272
rect 41786 968824 41842 968833
rect 41786 968759 41842 968768
rect 41800 967337 41828 967405
rect 41786 967328 41842 967337
rect 42720 967298 42748 975666
rect 41786 967263 41842 967272
rect 42156 967292 42208 967298
rect 42156 967234 42208 967240
rect 42708 967292 42760 967298
rect 42708 967234 42760 967240
rect 42168 966756 42196 967234
rect 41800 965161 41828 965565
rect 41786 965152 41842 965161
rect 41786 965087 41842 965096
rect 42168 964034 42196 964376
rect 42156 964028 42208 964034
rect 42156 963970 42208 963976
rect 42800 964028 42852 964034
rect 42800 963970 42852 963976
rect 41800 963529 41828 963725
rect 41786 963520 41842 963529
rect 41786 963455 41842 963464
rect 42168 962878 42196 963084
rect 42156 962872 42208 962878
rect 42156 962814 42208 962820
rect 41800 962169 41828 962540
rect 41786 962160 41842 962169
rect 41786 962095 41842 962104
rect 42076 959750 42104 960024
rect 42064 959744 42116 959750
rect 42064 959686 42116 959692
rect 42168 959138 42196 959412
rect 42156 959132 42208 959138
rect 42156 959074 42208 959080
rect 42076 958497 42104 958732
rect 42062 958488 42118 958497
rect 42062 958423 42118 958432
rect 41800 957817 41828 958188
rect 41786 957808 41842 957817
rect 41786 957743 41842 957752
rect 42182 956338 42288 956366
rect 42168 955398 42196 955740
rect 42156 955392 42208 955398
rect 42156 955334 42208 955340
rect 41800 954650 41828 955060
rect 41788 954644 41840 954650
rect 41788 954586 41840 954592
rect 41788 954440 41840 954446
rect 41788 954382 41840 954388
rect 31022 952912 31078 952921
rect 41800 952882 41828 954382
rect 42260 953578 42288 956338
rect 42340 955392 42392 955398
rect 42340 955334 42392 955340
rect 42168 953550 42288 953578
rect 31022 952847 31078 952856
rect 32404 952876 32456 952882
rect 27620 947368 27672 947374
rect 27620 947310 27672 947316
rect 8588 944180 8616 944316
rect 9048 944180 9076 944316
rect 9508 944180 9536 944316
rect 9968 944180 9996 944316
rect 10428 944180 10456 944316
rect 10888 944180 10916 944316
rect 11348 944180 11376 944316
rect 11808 944180 11836 944316
rect 12268 944180 12296 944316
rect 12728 944180 12756 944316
rect 13188 944180 13216 944316
rect 13648 944180 13676 944316
rect 14108 944180 14136 944316
rect 27632 943809 27660 947310
rect 27618 943800 27674 943809
rect 27618 943735 27674 943744
rect 31036 937417 31064 952847
rect 32404 952818 32456 952824
rect 41788 952876 41840 952882
rect 41788 952818 41840 952824
rect 32416 938233 32444 952818
rect 36726 952368 36782 952377
rect 36726 952303 36782 952312
rect 36542 952232 36598 952241
rect 36542 952167 36598 952176
rect 35808 943288 35860 943294
rect 35808 943230 35860 943236
rect 35716 943220 35768 943226
rect 35716 943162 35768 943168
rect 35728 942721 35756 943162
rect 35820 943129 35848 943230
rect 35806 943120 35862 943129
rect 35806 943055 35862 943064
rect 35714 942712 35770 942721
rect 35714 942647 35770 942656
rect 32402 938224 32458 938233
rect 32402 938159 32458 938168
rect 31022 937408 31078 937417
rect 31022 937343 31078 937352
rect 36556 935377 36584 952167
rect 36740 936193 36768 952303
rect 37924 952264 37976 952270
rect 37924 952206 37976 952212
rect 37936 936601 37964 952206
rect 41970 943800 42026 943809
rect 41970 943735 42026 943744
rect 41786 941896 41842 941905
rect 41786 941831 41842 941840
rect 41800 941746 41828 941831
rect 41524 941718 41828 941746
rect 37922 936592 37978 936601
rect 37922 936527 37978 936536
rect 36726 936184 36782 936193
rect 36726 936119 36782 936128
rect 36542 935368 36598 935377
rect 36542 935303 36598 935312
rect 39946 933328 40002 933337
rect 39946 933263 40002 933272
rect 39960 932414 39988 933263
rect 39948 932408 40000 932414
rect 39948 932350 40000 932356
rect 8588 818380 8616 818516
rect 9048 818380 9076 818516
rect 9508 818380 9536 818516
rect 9968 818380 9996 818516
rect 10428 818380 10456 818516
rect 10888 818380 10916 818516
rect 11348 818380 11376 818516
rect 11808 818380 11836 818516
rect 12268 818380 12296 818516
rect 12728 818380 12756 818516
rect 13188 818380 13216 818516
rect 13648 818380 13676 818516
rect 14108 818380 14136 818516
rect 41234 818000 41290 818009
rect 41234 817935 41290 817944
rect 41248 817426 41276 817935
rect 41328 817556 41380 817562
rect 41328 817498 41380 817504
rect 41236 817420 41288 817426
rect 41236 817362 41288 817368
rect 41340 817329 41368 817498
rect 41326 817320 41382 817329
rect 41326 817255 41382 817264
rect 41524 816626 41552 941718
rect 41786 941080 41842 941089
rect 41786 941015 41842 941024
rect 41694 939312 41750 939321
rect 41616 939270 41694 939298
rect 41616 821114 41644 939270
rect 41694 939247 41750 939256
rect 41696 932408 41748 932414
rect 41696 932350 41748 932356
rect 41708 932249 41736 932350
rect 41694 932240 41750 932249
rect 41694 932175 41696 932184
rect 41748 932175 41750 932184
rect 41696 932146 41748 932152
rect 41708 932115 41736 932146
rect 41800 923234 41828 941015
rect 41878 940264 41934 940273
rect 41878 940199 41934 940208
rect 41708 923206 41828 923234
rect 41708 828014 41736 923206
rect 41708 827986 41828 828014
rect 41616 821086 41736 821114
rect 41708 816762 41736 821086
rect 41800 819210 41828 827986
rect 41892 823874 41920 940199
rect 41984 938641 42012 943735
rect 42168 939049 42196 953550
rect 42352 952270 42380 955334
rect 42340 952264 42392 952270
rect 42340 952206 42392 952212
rect 42154 939040 42210 939049
rect 42154 938975 42210 938984
rect 41970 938632 42026 938641
rect 41970 938567 42026 938576
rect 42812 933745 42840 963970
rect 42892 962872 42944 962878
rect 42892 962814 42944 962820
rect 42904 934153 42932 962814
rect 44180 959744 44232 959750
rect 44180 959686 44232 959692
rect 42984 959132 43036 959138
rect 42984 959074 43036 959080
rect 42996 935785 43024 959074
rect 42982 935776 43038 935785
rect 42982 935711 43038 935720
rect 44192 934561 44220 959686
rect 44836 940681 44864 991442
rect 44916 961920 44968 961926
rect 44916 961862 44968 961868
rect 44928 943226 44956 961862
rect 45744 943288 45796 943294
rect 45744 943230 45796 943236
rect 44916 943220 44968 943226
rect 44916 943162 44968 943168
rect 44822 940672 44878 940681
rect 44822 940607 44878 940616
rect 45756 937038 45784 943230
rect 46216 942313 46244 992870
rect 47584 990140 47636 990146
rect 47584 990082 47636 990088
rect 46202 942304 46258 942313
rect 46202 942239 46258 942248
rect 47596 941497 47624 990082
rect 47582 941488 47638 941497
rect 47582 941423 47638 941432
rect 55876 939865 55904 995590
rect 84502 995574 84658 995602
rect 85210 995616 85266 995625
rect 85054 995574 85210 995602
rect 84658 995551 84714 995560
rect 86038 995616 86094 995625
rect 85698 995574 86038 995602
rect 85210 995551 85266 995560
rect 86038 995551 86094 995560
rect 88890 995480 88946 995489
rect 77036 995042 77064 995452
rect 77680 995178 77708 995452
rect 77668 995172 77720 995178
rect 77668 995114 77720 995120
rect 78324 995110 78352 995452
rect 78312 995104 78364 995110
rect 80164 995081 80192 995452
rect 81360 995246 81388 995452
rect 81348 995240 81400 995246
rect 87524 995217 87552 995452
rect 88734 995438 88890 995466
rect 88890 995415 88946 995424
rect 81348 995182 81400 995188
rect 87510 995208 87566 995217
rect 92584 995178 92612 997018
rect 92676 995246 92704 997494
rect 93136 995897 93164 1006198
rect 93122 995888 93178 995897
rect 93122 995823 93178 995832
rect 93320 995625 93348 1006266
rect 94516 996985 94544 1006402
rect 94596 1004692 94648 1004698
rect 94596 1004634 94648 1004640
rect 94608 999122 94636 1004634
rect 94780 999388 94832 999394
rect 94780 999330 94832 999336
rect 94596 999116 94648 999122
rect 94596 999058 94648 999064
rect 94792 997257 94820 999330
rect 94778 997248 94834 997257
rect 94778 997183 94834 997192
rect 94502 996976 94558 996985
rect 94502 996911 94558 996920
rect 93306 995616 93362 995625
rect 93306 995551 93362 995560
rect 92664 995240 92716 995246
rect 92664 995182 92716 995188
rect 87510 995143 87566 995152
rect 92572 995172 92624 995178
rect 92572 995114 92624 995120
rect 95896 995081 95924 1006470
rect 103150 1006431 103152 1006440
rect 103204 1006431 103206 1006440
rect 103610 1006496 103612 1006505
rect 145748 1006528 145800 1006534
rect 103664 1006496 103666 1006505
rect 145748 1006470 145800 1006476
rect 103610 1006431 103666 1006440
rect 144184 1006460 144236 1006466
rect 103152 1006402 103204 1006408
rect 144184 1006402 144236 1006408
rect 100116 1006392 100168 1006398
rect 104348 1006392 104400 1006398
rect 100116 1006334 100168 1006340
rect 100666 1006360 100722 1006369
rect 97264 1006188 97316 1006194
rect 97264 1006130 97316 1006136
rect 95976 1002176 96028 1002182
rect 95976 1002118 96028 1002124
rect 95988 1001230 96016 1002118
rect 95976 1001224 96028 1001230
rect 95976 1001166 96028 1001172
rect 95976 999728 96028 999734
rect 95976 999670 96028 999676
rect 95988 997558 96016 999670
rect 95976 997552 96028 997558
rect 95976 997494 96028 997500
rect 97276 995110 97304 1006130
rect 98276 1006120 98328 1006126
rect 98274 1006088 98276 1006097
rect 99104 1006120 99156 1006126
rect 98328 1006088 98330 1006097
rect 98274 1006023 98330 1006032
rect 99102 1006088 99104 1006097
rect 99156 1006088 99158 1006097
rect 99102 1006023 99158 1006032
rect 97356 1002244 97408 1002250
rect 97356 1002186 97408 1002192
rect 97368 997150 97396 1002186
rect 99472 1002176 99524 1002182
rect 99470 1002144 99472 1002153
rect 99524 1002144 99526 1002153
rect 98828 1002108 98880 1002114
rect 99470 1002079 99526 1002088
rect 98828 1002050 98880 1002056
rect 98644 1002040 98696 1002046
rect 98644 1001982 98696 1001988
rect 97540 1001972 97592 1001978
rect 97540 1001914 97592 1001920
rect 97552 999394 97580 1001914
rect 97540 999388 97592 999394
rect 97540 999330 97592 999336
rect 97356 997144 97408 997150
rect 97356 997086 97408 997092
rect 98656 995217 98684 1001982
rect 98840 999734 98868 1002050
rect 99930 1002008 99986 1002017
rect 99930 1001943 99932 1001952
rect 99984 1001943 99986 1001952
rect 100024 1001972 100076 1001978
rect 99932 1001914 99984 1001920
rect 100024 1001914 100076 1001920
rect 98828 999728 98880 999734
rect 98828 999670 98880 999676
rect 100036 997082 100064 1001914
rect 100128 998442 100156 1006334
rect 100666 1006295 100668 1006304
rect 100720 1006295 100722 1006304
rect 104346 1006360 104348 1006369
rect 104400 1006360 104402 1006369
rect 104346 1006295 104402 1006304
rect 108854 1006360 108910 1006369
rect 108854 1006295 108856 1006304
rect 100668 1006266 100720 1006272
rect 108908 1006295 108910 1006304
rect 108856 1006266 108908 1006272
rect 101956 1006256 102008 1006262
rect 101954 1006224 101956 1006233
rect 102784 1006256 102836 1006262
rect 102008 1006224 102010 1006233
rect 108488 1006256 108540 1006262
rect 102784 1006198 102836 1006204
rect 104806 1006224 104862 1006233
rect 101954 1006159 102010 1006168
rect 100298 1002280 100354 1002289
rect 100298 1002215 100300 1002224
rect 100352 1002215 100354 1002224
rect 100300 1002186 100352 1002192
rect 101494 1002144 101550 1002153
rect 101494 1002079 101496 1002088
rect 101548 1002079 101550 1002088
rect 101496 1002050 101548 1002056
rect 101128 1002040 101180 1002046
rect 101126 1002008 101128 1002017
rect 101180 1002008 101182 1002017
rect 101126 1001943 101182 1001952
rect 102322 1002008 102378 1002017
rect 102322 1001943 102324 1001952
rect 102376 1001943 102378 1001952
rect 102324 1001914 102376 1001920
rect 100116 998436 100168 998442
rect 100116 998378 100168 998384
rect 100024 997076 100076 997082
rect 100024 997018 100076 997024
rect 98642 995208 98698 995217
rect 98642 995143 98698 995152
rect 97264 995104 97316 995110
rect 78312 995046 78364 995052
rect 80150 995072 80206 995081
rect 77024 995036 77076 995042
rect 80150 995007 80206 995016
rect 95882 995072 95938 995081
rect 97264 995046 97316 995052
rect 95882 995007 95938 995016
rect 77024 994978 77076 994984
rect 88340 992996 88392 993002
rect 88340 992938 88392 992944
rect 88352 986678 88380 992938
rect 88340 986672 88392 986678
rect 88340 986614 88392 986620
rect 89628 986672 89680 986678
rect 89628 986614 89680 986620
rect 73436 985992 73488 985998
rect 73436 985934 73488 985940
rect 73448 983620 73476 985934
rect 89640 983620 89668 986614
rect 102796 985998 102824 1006198
rect 104806 1006159 104808 1006168
rect 104860 1006159 104862 1006168
rect 108486 1006224 108488 1006233
rect 113824 1006256 113876 1006262
rect 108540 1006224 108542 1006233
rect 113824 1006198 113876 1006204
rect 108486 1006159 108542 1006168
rect 104808 1006130 104860 1006136
rect 103150 1004728 103206 1004737
rect 103150 1004663 103152 1004672
rect 103204 1004663 103206 1004672
rect 103152 1004634 103204 1004640
rect 106830 1002416 106886 1002425
rect 106830 1002351 106832 1002360
rect 106884 1002351 106886 1002360
rect 109868 1002380 109920 1002386
rect 106832 1002322 106884 1002328
rect 109868 1002322 109920 1002328
rect 106188 1002312 106240 1002318
rect 106002 1002280 106058 1002289
rect 108488 1002312 108540 1002318
rect 106188 1002254 106240 1002260
rect 108486 1002280 108488 1002289
rect 108540 1002280 108542 1002289
rect 106002 1002215 106004 1002224
rect 106056 1002215 106058 1002224
rect 106004 1002186 106056 1002192
rect 105634 1002144 105690 1002153
rect 105634 1002079 105636 1002088
rect 105688 1002079 105690 1002088
rect 105636 1002050 105688 1002056
rect 104348 1002040 104400 1002046
rect 104346 1002008 104348 1002017
rect 104400 1002008 104402 1002017
rect 104346 1001943 104402 1001952
rect 102784 985992 102836 985998
rect 102784 985934 102836 985940
rect 106200 983634 106228 1002254
rect 108304 1002244 108356 1002250
rect 108486 1002215 108542 1002224
rect 108304 1002186 108356 1002192
rect 107660 1002176 107712 1002182
rect 107658 1002144 107660 1002153
rect 107712 1002144 107714 1002153
rect 107658 1002079 107714 1002088
rect 107752 1002108 107804 1002114
rect 107752 1002050 107804 1002056
rect 106648 1002040 106700 1002046
rect 106462 1002008 106518 1002017
rect 107200 1002040 107252 1002046
rect 106648 1001982 106700 1001988
rect 107198 1002008 107200 1002017
rect 107252 1002008 107254 1002017
rect 106462 1001943 106464 1001952
rect 106516 1001943 106518 1001952
rect 106464 1001914 106516 1001920
rect 106660 995042 106688 1001982
rect 107198 1001943 107254 1001952
rect 107764 995654 107792 1002050
rect 108026 1002008 108082 1002017
rect 107936 1001972 107988 1001978
rect 108026 1001943 108028 1001952
rect 107936 1001914 107988 1001920
rect 108080 1001943 108082 1001952
rect 108028 1001914 108080 1001920
rect 107752 995648 107804 995654
rect 107752 995590 107804 995596
rect 106648 995036 106700 995042
rect 106648 994978 106700 994984
rect 107948 991506 107976 1001914
rect 108316 996130 108344 1002186
rect 109684 1002176 109736 1002182
rect 109684 1002118 109736 1002124
rect 109040 1002040 109092 1002046
rect 109040 1001982 109092 1001988
rect 108304 996124 108356 996130
rect 108304 996066 108356 996072
rect 107936 991500 107988 991506
rect 107936 991442 107988 991448
rect 109052 990146 109080 1001982
rect 109696 996062 109724 1002118
rect 109880 997257 109908 1002322
rect 111798 1002008 111854 1002017
rect 110512 1001972 110564 1001978
rect 111798 1001943 111854 1001952
rect 110512 1001914 110564 1001920
rect 109866 997248 109922 997257
rect 109866 997183 109922 997192
rect 109684 996056 109736 996062
rect 109684 995998 109736 996004
rect 110524 992934 110552 1001914
rect 111812 993002 111840 1001943
rect 113836 997286 113864 1006198
rect 126244 1006052 126296 1006058
rect 126244 1005994 126296 1006000
rect 113824 997280 113876 997286
rect 112994 997248 113050 997257
rect 116124 997280 116176 997286
rect 113824 997222 113876 997228
rect 116122 997248 116124 997257
rect 116176 997248 116178 997257
rect 112994 997183 113050 997192
rect 116122 997183 116178 997192
rect 113008 997150 113036 997183
rect 112996 997144 113048 997150
rect 116124 997144 116176 997150
rect 112996 997086 113048 997092
rect 116122 997112 116124 997121
rect 116176 997112 116178 997121
rect 116122 997047 116178 997056
rect 111800 992996 111852 993002
rect 111800 992938 111852 992944
rect 110512 992928 110564 992934
rect 110512 992870 110564 992876
rect 122102 990992 122158 991001
rect 122102 990927 122158 990936
rect 109040 990140 109092 990146
rect 109040 990082 109092 990088
rect 105846 983606 106228 983634
rect 122116 983620 122144 990927
rect 126256 984638 126284 1005994
rect 143724 1005440 143776 1005446
rect 143724 1005382 143776 1005388
rect 143736 1001894 143764 1005382
rect 144092 1002108 144144 1002114
rect 144092 1002050 144144 1002056
rect 143644 1001866 143764 1001894
rect 137376 995852 137428 995858
rect 137376 995794 137428 995800
rect 137928 995852 137980 995858
rect 137928 995794 137980 995800
rect 139216 995852 139268 995858
rect 139216 995794 139268 995800
rect 142896 995852 142948 995858
rect 142896 995794 142948 995800
rect 129370 995752 129426 995761
rect 129122 995710 129370 995738
rect 133142 995752 133198 995761
rect 132802 995710 133142 995738
rect 129370 995687 129426 995696
rect 137388 995738 137416 995794
rect 137940 995738 137968 995794
rect 139228 995738 139256 995794
rect 141056 995784 141108 995790
rect 137126 995710 137416 995738
rect 137770 995710 137968 995738
rect 138966 995710 139256 995738
rect 140806 995732 141056 995738
rect 142908 995738 142936 995794
rect 143644 995790 143672 1001866
rect 143998 1000648 144054 1000657
rect 143998 1000583 144054 1000592
rect 143724 997824 143776 997830
rect 143724 997766 143776 997772
rect 143736 995858 143764 997766
rect 143816 997756 143868 997762
rect 143816 997698 143868 997704
rect 143828 997257 143856 997698
rect 143908 997688 143960 997694
rect 143908 997630 143960 997636
rect 143814 997248 143870 997257
rect 143814 997183 143870 997192
rect 143724 995852 143776 995858
rect 143724 995794 143776 995800
rect 140806 995726 141108 995732
rect 140806 995710 141096 995726
rect 142646 995710 142936 995738
rect 143632 995784 143684 995790
rect 143632 995726 143684 995732
rect 143920 995722 143948 997630
rect 144012 995926 144040 1000583
rect 144104 995994 144132 1002050
rect 144092 995988 144144 995994
rect 144092 995930 144144 995936
rect 144000 995920 144052 995926
rect 144000 995862 144052 995868
rect 143908 995716 143960 995722
rect 133142 995687 133198 995696
rect 143908 995658 143960 995664
rect 136546 995616 136602 995625
rect 136482 995574 136546 995602
rect 136546 995551 136602 995560
rect 130014 995480 130070 995489
rect 128464 995110 128492 995452
rect 129766 995438 130014 995466
rect 130014 995415 130070 995424
rect 131592 995217 131620 995452
rect 132144 995353 132172 995452
rect 132130 995344 132186 995353
rect 132130 995279 132186 995288
rect 131578 995208 131634 995217
rect 133432 995178 133460 995452
rect 135930 995438 136312 995466
rect 131578 995143 131634 995152
rect 133420 995172 133472 995178
rect 133420 995114 133472 995120
rect 128452 995104 128504 995110
rect 136284 995081 136312 995438
rect 140148 995081 140176 995452
rect 144196 995178 144224 1006402
rect 145564 1006188 145616 1006194
rect 145564 1006130 145616 1006136
rect 144828 996396 144880 996402
rect 144828 996338 144880 996344
rect 144840 995761 144868 996338
rect 144826 995752 144882 995761
rect 144826 995687 144882 995696
rect 145576 995489 145604 1006130
rect 145656 1006052 145708 1006058
rect 145656 1005994 145708 1006000
rect 145668 997121 145696 1005994
rect 145760 997830 145788 1006470
rect 145748 997824 145800 997830
rect 145748 997766 145800 997772
rect 145654 997112 145710 997121
rect 145654 997047 145710 997056
rect 146956 996169 146984 1007082
rect 203890 1007040 203946 1007049
rect 195428 1007004 195480 1007010
rect 308954 1007040 309010 1007049
rect 203890 1006975 203892 1006984
rect 195428 1006946 195480 1006952
rect 203944 1006975 203946 1006984
rect 300308 1007004 300360 1007010
rect 203892 1006946 203944 1006952
rect 308954 1006975 308956 1006984
rect 300308 1006946 300360 1006952
rect 309008 1006975 309010 1006984
rect 308956 1006946 309008 1006952
rect 154118 1006496 154174 1006505
rect 151636 1006460 151688 1006466
rect 154118 1006431 154120 1006440
rect 151636 1006402 151688 1006408
rect 154172 1006431 154174 1006440
rect 154120 1006402 154172 1006408
rect 150440 1006392 150492 1006398
rect 150440 1006334 150492 1006340
rect 150452 1006126 150480 1006334
rect 149704 1006120 149756 1006126
rect 149702 1006088 149704 1006097
rect 150440 1006120 150492 1006126
rect 149756 1006088 149758 1006097
rect 149702 1006023 149758 1006032
rect 150438 1006088 150440 1006097
rect 150492 1006088 150494 1006097
rect 151648 1006074 151676 1006402
rect 177304 1006392 177356 1006398
rect 177304 1006334 177356 1006340
rect 156142 1006224 156198 1006233
rect 156142 1006159 156144 1006168
rect 156196 1006159 156198 1006168
rect 156144 1006130 156196 1006136
rect 157432 1006120 157484 1006126
rect 151726 1006088 151782 1006097
rect 151648 1006046 151726 1006074
rect 150438 1006023 150494 1006032
rect 157430 1006088 157432 1006097
rect 159088 1006120 159140 1006126
rect 157484 1006088 157486 1006097
rect 151726 1006023 151782 1006032
rect 154488 1006052 154540 1006058
rect 157430 1006023 157486 1006032
rect 159086 1006088 159088 1006097
rect 166264 1006120 166316 1006126
rect 159140 1006088 159142 1006097
rect 159086 1006023 159142 1006032
rect 160650 1006088 160706 1006097
rect 166264 1006062 166316 1006068
rect 160650 1006023 160652 1006032
rect 154488 1005994 154540 1006000
rect 160704 1006023 160706 1006032
rect 160652 1005994 160704 1006000
rect 152556 1005440 152608 1005446
rect 152554 1005408 152556 1005417
rect 152608 1005408 152610 1005417
rect 152554 1005343 152610 1005352
rect 152922 1005000 152978 1005009
rect 149704 1004964 149756 1004970
rect 152922 1004935 152924 1004944
rect 149704 1004906 149756 1004912
rect 152976 1004935 152978 1004944
rect 152924 1004906 152976 1004912
rect 148324 1002040 148376 1002046
rect 148324 1001982 148376 1001988
rect 146942 996160 146998 996169
rect 146942 996095 146998 996104
rect 148336 995625 148364 1001982
rect 148508 1001972 148560 1001978
rect 148508 1001914 148560 1001920
rect 148520 1000657 148548 1001914
rect 148506 1000648 148562 1000657
rect 148506 1000583 148562 1000592
rect 149716 996402 149744 1004906
rect 153750 1004864 153806 1004873
rect 151084 1004828 151136 1004834
rect 153750 1004799 153752 1004808
rect 151084 1004770 151136 1004776
rect 153804 1004799 153806 1004808
rect 153752 1004770 153804 1004776
rect 150348 1004760 150400 1004766
rect 150348 1004702 150400 1004708
rect 150360 1002114 150388 1004702
rect 150348 1002108 150400 1002114
rect 150348 1002050 150400 1002056
rect 150898 1002008 150954 1002017
rect 150898 1001943 150900 1001952
rect 150952 1001943 150954 1001952
rect 150900 1001914 150952 1001920
rect 149704 996396 149756 996402
rect 149704 996338 149756 996344
rect 151096 995897 151124 1004770
rect 152096 1004760 152148 1004766
rect 152094 1004728 152096 1004737
rect 152148 1004728 152150 1004737
rect 151268 1004692 151320 1004698
rect 152094 1004663 152150 1004672
rect 153290 1004728 153346 1004737
rect 153290 1004663 153292 1004672
rect 151268 1004634 151320 1004640
rect 153344 1004663 153346 1004672
rect 153292 1004634 153344 1004640
rect 151082 995888 151138 995897
rect 151082 995823 151138 995832
rect 148322 995616 148378 995625
rect 148322 995551 148378 995560
rect 145562 995480 145618 995489
rect 145562 995415 145618 995424
rect 151280 995353 151308 1004634
rect 151728 1002040 151780 1002046
rect 151726 1002008 151728 1002017
rect 151780 1002008 151782 1002017
rect 151726 1001943 151782 1001952
rect 151266 995344 151322 995353
rect 151266 995279 151322 995288
rect 144184 995172 144236 995178
rect 144184 995114 144236 995120
rect 128452 995046 128504 995052
rect 136270 995072 136326 995081
rect 136270 995007 136326 995016
rect 140134 995072 140190 995081
rect 140134 995007 140190 995016
rect 138296 990140 138348 990146
rect 138296 990082 138348 990088
rect 126244 984632 126296 984638
rect 126244 984574 126296 984580
rect 138308 983620 138336 990082
rect 154500 983620 154528 1005994
rect 160650 1005000 160706 1005009
rect 160650 1004935 160652 1004944
rect 160704 1004935 160706 1004944
rect 162860 1004964 162912 1004970
rect 160652 1004906 160704 1004912
rect 162860 1004906 162912 1004912
rect 159454 1004864 159510 1004873
rect 159454 1004799 159456 1004808
rect 159508 1004799 159510 1004808
rect 161480 1004828 161532 1004834
rect 159456 1004770 159508 1004776
rect 161480 1004770 161532 1004776
rect 160284 1004760 160336 1004766
rect 159822 1004728 159878 1004737
rect 159822 1004663 159824 1004672
rect 159876 1004663 159878 1004672
rect 160282 1004728 160284 1004737
rect 160336 1004728 160338 1004737
rect 160282 1004663 160338 1004672
rect 159824 1004634 159876 1004640
rect 158260 1002176 158312 1002182
rect 155774 1002144 155830 1002153
rect 157430 1002144 157486 1002153
rect 155774 1002079 155776 1002088
rect 155828 1002079 155830 1002088
rect 157340 1002108 157392 1002114
rect 155776 1002050 155828 1002056
rect 157430 1002079 157432 1002088
rect 157340 1002050 157392 1002056
rect 157484 1002079 157486 1002088
rect 158258 1002144 158260 1002153
rect 161112 1002176 161164 1002182
rect 158312 1002144 158314 1002153
rect 161112 1002118 161164 1002124
rect 158258 1002079 158314 1002088
rect 159364 1002108 159416 1002114
rect 157432 1002050 157484 1002056
rect 159364 1002050 159416 1002056
rect 155774 1002008 155830 1002017
rect 155774 1001943 155830 1001952
rect 156970 1002008 157026 1002017
rect 156970 1001943 156972 1001952
rect 155788 997694 155816 1001943
rect 157024 1001943 157026 1001952
rect 156972 1001914 157024 1001920
rect 155776 997688 155828 997694
rect 155776 997630 155828 997636
rect 157352 997422 157380 1002050
rect 158628 1002040 158680 1002046
rect 158626 1002008 158628 1002017
rect 158680 1002008 158682 1002017
rect 158626 1001943 158682 1001952
rect 158720 1001972 158772 1001978
rect 158720 1001914 158772 1001920
rect 154580 997416 154632 997422
rect 154580 997358 154632 997364
rect 157340 997416 157392 997422
rect 157340 997358 157392 997364
rect 154592 995110 154620 997358
rect 158732 996130 158760 1001914
rect 159376 996198 159404 1002050
rect 160192 1002040 160244 1002046
rect 160192 1001982 160244 1001988
rect 159364 996192 159416 996198
rect 159364 996134 159416 996140
rect 158720 996124 158772 996130
rect 158720 996066 158772 996072
rect 160204 996062 160232 1001982
rect 161124 997121 161152 1002118
rect 161492 997762 161520 1004770
rect 162124 1004692 162176 1004698
rect 162124 1004634 162176 1004640
rect 161480 997756 161532 997762
rect 161480 997698 161532 997704
rect 162136 997393 162164 1004634
rect 162122 997384 162178 997393
rect 162122 997319 162178 997328
rect 161110 997112 161166 997121
rect 161110 997047 161166 997056
rect 160192 996056 160244 996062
rect 160192 995998 160244 996004
rect 154580 995104 154632 995110
rect 154580 995046 154632 995052
rect 162872 990146 162900 1004906
rect 163504 1004760 163556 1004766
rect 163504 1004702 163556 1004708
rect 162860 990140 162912 990146
rect 162860 990082 162912 990088
rect 163516 985930 163544 1004702
rect 164422 997384 164478 997393
rect 164422 997319 164478 997328
rect 164436 997286 164464 997319
rect 164424 997280 164476 997286
rect 164424 997222 164476 997228
rect 164424 997144 164476 997150
rect 164422 997112 164424 997121
rect 164476 997112 164478 997121
rect 164422 997047 164478 997056
rect 166276 996062 166304 1006062
rect 167552 997280 167604 997286
rect 167550 997248 167552 997257
rect 167604 997248 167606 997257
rect 167550 997183 167606 997192
rect 167552 997144 167604 997150
rect 167550 997112 167552 997121
rect 167604 997112 167606 997121
rect 167550 997047 167606 997056
rect 166264 996056 166316 996062
rect 166264 995998 166316 996004
rect 165986 995072 166042 995081
rect 165986 995007 165988 995016
rect 166040 995007 166042 995016
rect 167550 995072 167606 995081
rect 167550 995007 167552 995016
rect 165988 994978 166040 994984
rect 167604 995007 167606 995016
rect 167552 994978 167604 994984
rect 163504 985924 163556 985930
rect 163504 985866 163556 985872
rect 170772 985924 170824 985930
rect 170772 985866 170824 985872
rect 170784 983620 170812 985866
rect 177316 984706 177344 1006334
rect 195152 1006324 195204 1006330
rect 195152 1006266 195204 1006272
rect 195164 1001910 195192 1006266
rect 195244 1006120 195296 1006126
rect 195244 1006062 195296 1006068
rect 195152 1001904 195204 1001910
rect 195058 1001872 195114 1001881
rect 195256 1001881 195284 1006062
rect 195336 1001904 195388 1001910
rect 195152 1001846 195204 1001852
rect 195242 1001872 195298 1001881
rect 195058 1001807 195114 1001816
rect 195440 1001894 195468 1006946
rect 261022 1006904 261078 1006913
rect 261022 1006839 261024 1006848
rect 261076 1006839 261078 1006848
rect 268384 1006868 268436 1006874
rect 261024 1006810 261076 1006816
rect 268384 1006810 268436 1006816
rect 203522 1006632 203578 1006641
rect 198004 1006596 198056 1006602
rect 203522 1006567 203524 1006576
rect 198004 1006538 198056 1006544
rect 203576 1006567 203578 1006576
rect 203524 1006538 203576 1006544
rect 196624 1006188 196676 1006194
rect 196624 1006130 196676 1006136
rect 195440 1001866 195744 1001894
rect 195336 1001846 195388 1001852
rect 195242 1001807 195298 1001816
rect 189448 995852 189500 995858
rect 189448 995794 189500 995800
rect 194324 995852 194376 995858
rect 194324 995794 194376 995800
rect 184662 995752 184718 995761
rect 188158 995752 188214 995761
rect 184718 995710 184828 995738
rect 187864 995710 188158 995738
rect 184662 995687 184718 995696
rect 189460 995738 189488 995794
rect 192484 995784 192536 995790
rect 189152 995710 189488 995738
rect 190348 995722 190684 995738
rect 192188 995732 192484 995738
rect 194336 995738 194364 995794
rect 192188 995726 192536 995732
rect 190348 995716 190696 995722
rect 190348 995710 190644 995716
rect 188158 995687 188214 995696
rect 192188 995710 192524 995726
rect 194028 995710 194364 995738
rect 190644 995658 190696 995664
rect 188802 995616 188858 995625
rect 188508 995574 188802 995602
rect 188802 995551 188858 995560
rect 195072 995489 195100 1001807
rect 195152 1001632 195204 1001638
rect 195152 1001574 195204 1001580
rect 195164 995790 195192 1001574
rect 195348 998186 195376 1001846
rect 195348 998158 195560 998186
rect 195428 998028 195480 998034
rect 195428 997970 195480 997976
rect 195336 997824 195388 997830
rect 195336 997766 195388 997772
rect 195244 997756 195296 997762
rect 195244 997698 195296 997704
rect 195256 997257 195284 997698
rect 195242 997248 195298 997257
rect 195242 997183 195298 997192
rect 195244 997144 195296 997150
rect 195244 997086 195296 997092
rect 195152 995784 195204 995790
rect 195152 995726 195204 995732
rect 195256 995625 195284 997086
rect 195348 995858 195376 997766
rect 195440 995926 195468 997970
rect 195428 995920 195480 995926
rect 195428 995862 195480 995868
rect 195336 995852 195388 995858
rect 195336 995794 195388 995800
rect 195242 995616 195298 995625
rect 195242 995551 195298 995560
rect 184478 995480 184534 995489
rect 179860 995438 180196 995466
rect 180504 995438 180656 995466
rect 180168 995178 180196 995438
rect 180156 995172 180208 995178
rect 180156 995114 180208 995120
rect 180628 995110 180656 995438
rect 181134 995217 181162 995452
rect 182988 995438 183324 995466
rect 181120 995208 181176 995217
rect 181120 995143 181176 995152
rect 180616 995104 180668 995110
rect 180616 995046 180668 995052
rect 183296 995042 183324 995438
rect 183526 995246 183554 995452
rect 184184 995438 184478 995466
rect 195058 995480 195114 995489
rect 184478 995415 184534 995424
rect 187298 995353 187326 995452
rect 191544 995438 191788 995466
rect 187284 995344 187340 995353
rect 187284 995279 187340 995288
rect 183514 995240 183566 995246
rect 183514 995182 183566 995188
rect 191760 995081 191788 995438
rect 195058 995415 195114 995424
rect 195532 995246 195560 998158
rect 195716 995722 195744 1001866
rect 195980 998436 196032 998442
rect 195980 998378 196032 998384
rect 195704 995716 195756 995722
rect 195704 995658 195756 995664
rect 195520 995240 195572 995246
rect 195520 995182 195572 995188
rect 195992 995178 196020 998378
rect 196636 997830 196664 1006130
rect 197360 1000408 197412 1000414
rect 197360 1000350 197412 1000356
rect 196624 997824 196676 997830
rect 196624 997766 196676 997772
rect 197372 996305 197400 1000350
rect 198016 997150 198044 1006538
rect 204718 1006360 204774 1006369
rect 258170 1006360 258226 1006369
rect 204718 1006295 204720 1006304
rect 204772 1006295 204774 1006304
rect 228364 1006324 228416 1006330
rect 204720 1006266 204772 1006272
rect 228364 1006266 228416 1006272
rect 254676 1006324 254728 1006330
rect 258170 1006295 258172 1006304
rect 254676 1006266 254728 1006272
rect 258224 1006295 258226 1006304
rect 258172 1006266 258224 1006272
rect 205546 1006224 205602 1006233
rect 205546 1006159 205548 1006168
rect 205600 1006159 205602 1006168
rect 205548 1006130 205600 1006136
rect 204352 1006120 204404 1006126
rect 201038 1006088 201094 1006097
rect 201038 1006023 201040 1006032
rect 201092 1006023 201094 1006032
rect 201866 1006088 201922 1006097
rect 201866 1006023 201868 1006032
rect 201040 1005994 201092 1006000
rect 201920 1006023 201922 1006032
rect 204350 1006088 204352 1006097
rect 209596 1006120 209648 1006126
rect 204404 1006088 204406 1006097
rect 208766 1006088 208822 1006097
rect 204350 1006023 204406 1006032
rect 204904 1006052 204956 1006058
rect 201868 1005994 201920 1006000
rect 208766 1006023 208768 1006032
rect 204904 1005994 204956 1006000
rect 208820 1006023 208822 1006032
rect 209594 1006088 209596 1006097
rect 216036 1006120 216088 1006126
rect 209648 1006088 209650 1006097
rect 209594 1006023 209650 1006032
rect 215206 1006088 215262 1006097
rect 216036 1006062 216088 1006068
rect 215206 1006023 215262 1006032
rect 208768 1005994 208820 1006000
rect 202326 1004728 202382 1004737
rect 199384 1004692 199436 1004698
rect 202326 1004663 202328 1004672
rect 199384 1004634 199436 1004640
rect 202380 1004663 202382 1004672
rect 202328 1004634 202380 1004640
rect 199396 998034 199424 1004634
rect 202144 1002108 202196 1002114
rect 202144 1002050 202196 1002056
rect 200764 1002040 200816 1002046
rect 200764 1001982 200816 1001988
rect 199384 998028 199436 998034
rect 199384 997970 199436 997976
rect 198004 997144 198056 997150
rect 200212 997144 200264 997150
rect 198004 997086 198056 997092
rect 200210 997112 200212 997121
rect 200264 997112 200266 997121
rect 200210 997047 200266 997056
rect 197358 996296 197414 996305
rect 197358 996231 197414 996240
rect 200776 995761 200804 1001982
rect 200948 1001972 201000 1001978
rect 200948 1001914 201000 1001920
rect 200960 1000414 200988 1001914
rect 200948 1000408 201000 1000414
rect 200948 1000350 201000 1000356
rect 200762 995752 200818 995761
rect 200762 995687 200818 995696
rect 195980 995172 196032 995178
rect 195980 995114 196032 995120
rect 202156 995110 202184 1002050
rect 202696 1002040 202748 1002046
rect 202694 1002008 202696 1002017
rect 202748 1002008 202750 1002017
rect 202694 1001943 202750 1001952
rect 203062 1002008 203118 1002017
rect 203062 1001943 203064 1001952
rect 203116 1001943 203118 1001952
rect 203524 1001972 203576 1001978
rect 203064 1001914 203116 1001920
rect 203524 1001914 203576 1001920
rect 202420 998300 202472 998306
rect 202420 998242 202472 998248
rect 202432 995217 202460 998242
rect 203536 995353 203564 1001914
rect 204916 997150 204944 1005994
rect 215220 1005310 215248 1006023
rect 215208 1005304 215260 1005310
rect 215208 1005246 215260 1005252
rect 208400 1004896 208452 1004902
rect 208398 1004864 208400 1004873
rect 209780 1004896 209832 1004902
rect 208452 1004864 208454 1004873
rect 209780 1004838 209832 1004844
rect 208398 1004799 208454 1004808
rect 208768 1004760 208820 1004766
rect 208766 1004728 208768 1004737
rect 208820 1004728 208822 1004737
rect 208766 1004663 208822 1004672
rect 207204 1002584 207256 1002590
rect 207202 1002552 207204 1002561
rect 207256 1002552 207258 1002561
rect 207202 1002487 207258 1002496
rect 205178 1002144 205234 1002153
rect 205178 1002079 205180 1002088
rect 205232 1002079 205234 1002088
rect 206742 1002144 206798 1002153
rect 206742 1002079 206744 1002088
rect 205180 1002050 205232 1002056
rect 206796 1002079 206798 1002088
rect 208400 1002108 208452 1002114
rect 206744 1002050 206796 1002056
rect 208400 1002050 208452 1002056
rect 205914 1002008 205970 1002017
rect 206742 1002008 206798 1002017
rect 205914 1001943 205916 1001952
rect 205968 1001943 205970 1001952
rect 206296 1001966 206742 1001994
rect 205916 1001914 205968 1001920
rect 206296 998442 206324 1001966
rect 206742 1001943 206798 1001952
rect 207570 1002008 207626 1002017
rect 207570 1001943 207626 1001952
rect 207584 1001910 207612 1001943
rect 206928 1001904 206980 1001910
rect 206928 1001846 206980 1001852
rect 207572 1001904 207624 1001910
rect 207572 1001846 207624 1001852
rect 206284 998436 206336 998442
rect 206284 998378 206336 998384
rect 206940 998306 206968 1001846
rect 206928 998300 206980 998306
rect 206928 998242 206980 998248
rect 204904 997144 204956 997150
rect 204904 997086 204956 997092
rect 203522 995344 203578 995353
rect 203522 995279 203578 995288
rect 202418 995208 202474 995217
rect 202418 995143 202474 995152
rect 202144 995104 202196 995110
rect 186502 995072 186558 995081
rect 183284 995036 183336 995042
rect 186502 995007 186558 995016
rect 191746 995072 191802 995081
rect 202144 995046 202196 995052
rect 208412 995042 208440 1002050
rect 209792 996198 209820 1004838
rect 211804 1004760 211856 1004766
rect 211804 1004702 211856 1004708
rect 210422 1002280 210478 1002289
rect 210422 1002215 210424 1002224
rect 210476 1002215 210478 1002224
rect 210424 1002186 210476 1002192
rect 210056 1002176 210108 1002182
rect 210054 1002144 210056 1002153
rect 210108 1002144 210110 1002153
rect 210054 1002079 210110 1002088
rect 211250 1002144 211306 1002153
rect 211250 1002079 211252 1002088
rect 211304 1002079 211306 1002088
rect 211252 1002050 211304 1002056
rect 211712 1002040 211764 1002046
rect 210882 1002008 210938 1002017
rect 211710 1002008 211712 1002017
rect 211764 1002008 211766 1002017
rect 210938 1001966 211292 1001994
rect 210882 1001943 210938 1001952
rect 211264 997762 211292 1001966
rect 211710 1001943 211766 1001952
rect 211252 997756 211304 997762
rect 211252 997698 211304 997704
rect 209780 996192 209832 996198
rect 209780 996134 209832 996140
rect 211816 996130 211844 1004702
rect 213184 1002244 213236 1002250
rect 213184 1002186 213236 1002192
rect 212540 1002176 212592 1002182
rect 212540 1002118 212592 1002124
rect 212078 1002008 212134 1002017
rect 212078 1001943 212080 1001952
rect 212132 1001943 212134 1001952
rect 212080 1001914 212132 1001920
rect 211804 996124 211856 996130
rect 211804 996066 211856 996072
rect 212552 996062 212580 1002118
rect 213196 996198 213224 1002186
rect 213368 1002108 213420 1002114
rect 213368 1002050 213420 1002056
rect 213380 997393 213408 1002050
rect 215944 1002040 215996 1002046
rect 215944 1001982 215996 1001988
rect 213920 1001972 213972 1001978
rect 213920 1001914 213972 1001920
rect 213366 997384 213422 997393
rect 213366 997319 213422 997328
rect 213184 996192 213236 996198
rect 213184 996134 213236 996140
rect 212540 996056 212592 996062
rect 212540 995998 212592 996004
rect 191746 995007 191802 995016
rect 208400 995036 208452 995042
rect 183284 994978 183336 994984
rect 177304 984700 177356 984706
rect 177304 984642 177356 984648
rect 186516 983634 186544 995007
rect 208400 994978 208452 994984
rect 213932 991506 213960 1001914
rect 215758 997384 215814 997393
rect 215758 997319 215760 997328
rect 215812 997319 215814 997328
rect 215760 997290 215812 997296
rect 215956 991506 215984 1001982
rect 216048 996062 216076 1006062
rect 219440 1005304 219492 1005310
rect 219440 1005246 219492 1005252
rect 218888 997348 218940 997354
rect 218888 997290 218940 997296
rect 218900 997257 218928 997290
rect 218886 997248 218942 997257
rect 218886 997183 218942 997192
rect 216036 996056 216088 996062
rect 216036 995998 216088 996004
rect 217416 995104 217468 995110
rect 217414 995072 217416 995081
rect 218888 995104 218940 995110
rect 217468 995072 217470 995081
rect 217414 995007 217470 995016
rect 218886 995072 218888 995081
rect 218940 995072 218942 995081
rect 218886 995007 218942 995016
rect 203156 991500 203208 991506
rect 203156 991442 203208 991448
rect 213920 991500 213972 991506
rect 213920 991442 213972 991448
rect 215944 991500 215996 991506
rect 215944 991442 215996 991448
rect 186516 983606 186990 983634
rect 203168 983620 203196 991442
rect 219452 983620 219480 1005246
rect 228376 984774 228404 1006266
rect 252468 1006256 252520 1006262
rect 252466 1006224 252468 1006233
rect 253296 1006256 253348 1006262
rect 252520 1006224 252522 1006233
rect 250444 1006188 250496 1006194
rect 252466 1006159 252522 1006168
rect 253294 1006224 253296 1006233
rect 253348 1006224 253350 1006233
rect 253294 1006159 253350 1006168
rect 250444 1006130 250496 1006136
rect 247684 1006120 247736 1006126
rect 247684 1006062 247736 1006068
rect 246672 1002584 246724 1002590
rect 246672 1002526 246724 1002532
rect 246580 1001904 246632 1001910
rect 246580 1001846 246632 1001852
rect 246592 997914 246620 1001846
rect 246500 997886 246620 997914
rect 246500 995858 246528 997886
rect 246580 997756 246632 997762
rect 246580 997698 246632 997704
rect 246592 997257 246620 997698
rect 246578 997248 246634 997257
rect 246578 997183 246634 997192
rect 240876 995852 240928 995858
rect 240876 995794 240928 995800
rect 246488 995852 246540 995858
rect 246488 995794 246540 995800
rect 240048 995784 240100 995790
rect 235262 995752 235318 995761
rect 234968 995710 235262 995738
rect 239936 995732 240048 995738
rect 240888 995738 240916 995794
rect 246684 995790 246712 1002526
rect 247040 1001292 247092 1001298
rect 247040 1001234 247092 1001240
rect 246764 998436 246816 998442
rect 246764 998378 246816 998384
rect 246672 995784 246724 995790
rect 243818 995752 243874 995761
rect 239936 995726 240100 995732
rect 239936 995710 240088 995726
rect 240580 995710 240916 995738
rect 243616 995710 243818 995738
rect 235262 995687 235318 995696
rect 245456 995722 245608 995738
rect 246672 995726 246724 995732
rect 246776 995722 246804 998378
rect 246856 997824 246908 997830
rect 246856 997766 246908 997772
rect 245456 995716 245620 995722
rect 245456 995710 245568 995716
rect 243818 995687 243874 995696
rect 245568 995658 245620 995664
rect 246764 995716 246816 995722
rect 246764 995658 246816 995664
rect 246868 995654 246896 997766
rect 243268 995648 243320 995654
rect 232226 995616 232282 995625
rect 231932 995574 232226 995602
rect 242070 995616 242126 995625
rect 241776 995574 242070 995602
rect 232226 995551 232282 995560
rect 242972 995596 243268 995602
rect 242972 995590 243320 995596
rect 246856 995648 246908 995654
rect 246856 995590 246908 995596
rect 242972 995574 243308 995590
rect 242070 995551 242126 995560
rect 247052 995489 247080 1001234
rect 247132 1001224 247184 1001230
rect 247132 1001166 247184 1001172
rect 236550 995480 236606 995489
rect 231288 995438 231624 995466
rect 232576 995438 232912 995466
rect 234416 995438 234568 995466
rect 235612 995438 235948 995466
rect 236256 995438 236550 995466
rect 231596 995110 231624 995438
rect 231584 995104 231636 995110
rect 231584 995046 231636 995052
rect 232884 995042 232912 995438
rect 234540 995194 234568 995438
rect 234618 995208 234674 995217
rect 234540 995166 234618 995194
rect 235920 995178 235948 995438
rect 247038 995480 247094 995489
rect 236550 995415 236606 995424
rect 238726 995353 238754 995452
rect 238712 995344 238768 995353
rect 238712 995279 238768 995288
rect 239278 995246 239306 995452
rect 247038 995415 247094 995424
rect 239266 995240 239318 995246
rect 239266 995182 239318 995188
rect 247144 995178 247172 1001166
rect 247696 996441 247724 1006062
rect 249064 1006052 249116 1006058
rect 249064 1005994 249116 1006000
rect 247682 996432 247738 996441
rect 247682 996367 247738 996376
rect 249076 995625 249104 1005994
rect 249156 1001972 249208 1001978
rect 249156 1001914 249208 1001920
rect 249062 995616 249118 995625
rect 249062 995551 249118 995560
rect 249168 995246 249196 1001914
rect 250456 1001894 250484 1006130
rect 253662 1002688 253718 1002697
rect 253662 1002623 253664 1002632
rect 253716 1002623 253718 1002632
rect 253664 1002594 253716 1002600
rect 253204 1002176 253256 1002182
rect 253204 1002118 253256 1002124
rect 251916 1002040 251968 1002046
rect 251916 1001982 251968 1001988
rect 250364 1001866 250484 1001894
rect 250364 996033 250392 1001866
rect 251928 1001298 251956 1001982
rect 251916 1001292 251968 1001298
rect 251916 1001234 251968 1001240
rect 251548 1000612 251600 1000618
rect 251548 1000554 251600 1000560
rect 250444 1000544 250496 1000550
rect 250444 1000486 250496 1000492
rect 250456 996169 250484 1000486
rect 251364 999184 251416 999190
rect 251364 999126 251416 999132
rect 250442 996160 250498 996169
rect 250442 996095 250498 996104
rect 250350 996024 250406 996033
rect 250350 995959 250406 995968
rect 251376 995353 251404 999126
rect 251362 995344 251418 995353
rect 251362 995279 251418 995288
rect 249156 995240 249208 995246
rect 249156 995182 249208 995188
rect 234618 995143 234674 995152
rect 235908 995172 235960 995178
rect 235908 995114 235960 995120
rect 247132 995172 247184 995178
rect 247132 995114 247184 995120
rect 251560 995110 251588 1000554
rect 253216 1000550 253244 1002118
rect 253388 1002108 253440 1002114
rect 253388 1002050 253440 1002056
rect 253400 1001230 253428 1002050
rect 254492 1002040 254544 1002046
rect 254122 1002008 254178 1002017
rect 254122 1001943 254124 1001952
rect 254176 1001943 254178 1001952
rect 254490 1002008 254492 1002017
rect 254584 1002040 254636 1002046
rect 254544 1002008 254546 1002017
rect 254584 1001982 254636 1001988
rect 254490 1001943 254546 1001952
rect 254124 1001914 254176 1001920
rect 253388 1001224 253440 1001230
rect 253388 1001166 253440 1001172
rect 253204 1000544 253256 1000550
rect 253204 1000486 253256 1000492
rect 254596 998442 254624 1001982
rect 254688 1000618 254716 1006266
rect 256514 1006224 256570 1006233
rect 256514 1006159 256516 1006168
rect 256568 1006159 256570 1006168
rect 256516 1006130 256568 1006136
rect 258540 1006120 258592 1006126
rect 255318 1006088 255374 1006097
rect 258538 1006088 258540 1006097
rect 263048 1006120 263100 1006126
rect 258592 1006088 258594 1006097
rect 255318 1006023 255320 1006032
rect 255372 1006023 255374 1006032
rect 257344 1006052 257396 1006058
rect 255320 1005994 255372 1006000
rect 258538 1006023 258594 1006032
rect 258998 1006088 259054 1006097
rect 258998 1006023 259000 1006032
rect 257344 1005994 257396 1006000
rect 259052 1006023 259054 1006032
rect 262678 1006088 262734 1006097
rect 262678 1006023 262680 1006032
rect 259000 1005994 259052 1006000
rect 262732 1006023 262734 1006032
rect 263046 1006088 263048 1006097
rect 263100 1006088 263102 1006097
rect 263046 1006023 263102 1006032
rect 262680 1005994 262732 1006000
rect 254952 1002584 255004 1002590
rect 254950 1002552 254952 1002561
rect 255004 1002552 255006 1002561
rect 254950 1002487 255006 1002496
rect 256148 1002176 256200 1002182
rect 255686 1002144 255742 1002153
rect 255686 1002079 255688 1002088
rect 255740 1002079 255742 1002088
rect 256146 1002144 256148 1002153
rect 256200 1002144 256202 1002153
rect 256146 1002079 256202 1002088
rect 255688 1002050 255740 1002056
rect 256976 1002040 257028 1002046
rect 256974 1002008 256976 1002017
rect 257028 1002008 257030 1002017
rect 254768 1001972 254820 1001978
rect 256974 1001943 257030 1001952
rect 254768 1001914 254820 1001920
rect 254676 1000612 254728 1000618
rect 254676 1000554 254728 1000560
rect 254780 999190 254808 1001914
rect 254768 999184 254820 999190
rect 254768 999126 254820 999132
rect 254584 998436 254636 998442
rect 254584 998378 254636 998384
rect 251548 995104 251600 995110
rect 245658 995072 245714 995081
rect 232872 995036 232924 995042
rect 251548 995046 251600 995052
rect 257356 995042 257384 1005994
rect 260194 1002280 260250 1002289
rect 260194 1002215 260196 1002224
rect 260248 1002215 260250 1002224
rect 262864 1002244 262916 1002250
rect 260196 1002186 260248 1002192
rect 262864 1002186 262916 1002192
rect 261852 1002176 261904 1002182
rect 261482 1002144 261538 1002153
rect 261482 1002079 261484 1002088
rect 261536 1002079 261538 1002088
rect 261850 1002144 261852 1002153
rect 261904 1002144 261906 1002153
rect 261850 1002079 261906 1002088
rect 261484 1002050 261536 1002056
rect 260656 1002040 260708 1002046
rect 257802 1002008 257858 1002017
rect 257802 1001943 257804 1001952
rect 257856 1001943 257858 1001952
rect 259826 1002008 259882 1002017
rect 259826 1001943 259828 1001952
rect 257804 1001914 257856 1001920
rect 259880 1001943 259882 1001952
rect 260654 1002008 260656 1002017
rect 262220 1002040 262272 1002046
rect 260708 1002008 260710 1002017
rect 261850 1002008 261906 1002017
rect 260654 1001943 260710 1001952
rect 260932 1001972 260984 1001978
rect 259828 1001914 259880 1001920
rect 262220 1001982 262272 1001988
rect 261850 1001943 261906 1001952
rect 260932 1001914 260984 1001920
rect 260944 996130 260972 1001914
rect 261864 997762 261892 1001943
rect 261852 997756 261904 997762
rect 261852 997698 261904 997704
rect 260932 996124 260984 996130
rect 260932 996066 260984 996072
rect 262232 996062 262260 1001982
rect 262876 996130 262904 1002186
rect 264244 1002176 264296 1002182
rect 264244 1002118 264296 1002124
rect 263600 1002108 263652 1002114
rect 263600 1002050 263652 1002056
rect 263506 1002008 263562 1002017
rect 263506 1001943 263508 1001952
rect 263560 1001943 263562 1001952
rect 263508 1001914 263560 1001920
rect 263612 996198 263640 1002050
rect 264256 996198 264284 1002118
rect 267002 1002008 267058 1002017
rect 265624 1001972 265676 1001978
rect 267002 1001943 267058 1001952
rect 265624 1001914 265676 1001920
rect 263600 996192 263652 996198
rect 263600 996134 263652 996140
rect 264244 996192 264296 996198
rect 264244 996134 264296 996140
rect 262864 996124 262916 996130
rect 262864 996066 262916 996072
rect 262220 996056 262272 996062
rect 262220 995998 262272 996004
rect 245658 995007 245714 995016
rect 257344 995036 257396 995042
rect 232872 994978 232924 994984
rect 245672 992934 245700 995007
rect 257344 994978 257396 994984
rect 245660 992928 245712 992934
rect 245660 992870 245712 992876
rect 251456 992928 251508 992934
rect 251456 992870 251508 992876
rect 235632 991500 235684 991506
rect 235632 991442 235684 991448
rect 228364 984768 228416 984774
rect 228364 984710 228416 984716
rect 235644 983620 235672 991442
rect 251468 983634 251496 992870
rect 265636 986678 265664 1001914
rect 265624 986672 265676 986678
rect 265624 986614 265676 986620
rect 267016 985998 267044 1001943
rect 268396 996062 268424 1006810
rect 280804 1006324 280856 1006330
rect 280804 1006266 280856 1006272
rect 300216 1006324 300268 1006330
rect 300216 1006266 300268 1006272
rect 269764 1006120 269816 1006126
rect 269764 1006062 269816 1006068
rect 268476 1006052 268528 1006058
rect 268476 1005994 268528 1006000
rect 268488 997286 268516 1005994
rect 268476 997280 268528 997286
rect 268476 997222 268528 997228
rect 268384 996056 268436 996062
rect 268384 995998 268436 996004
rect 269776 990146 269804 1006062
rect 279332 997824 279384 997830
rect 279332 997766 279384 997772
rect 270316 997280 270368 997286
rect 270314 997248 270316 997257
rect 270368 997248 270370 997257
rect 270314 997183 270370 997192
rect 279344 995654 279372 997766
rect 279332 995648 279384 995654
rect 279332 995590 279384 995596
rect 269764 990140 269816 990146
rect 269764 990082 269816 990088
rect 268108 986672 268160 986678
rect 268108 986614 268160 986620
rect 267004 985992 267056 985998
rect 267004 985934 267056 985940
rect 251468 983606 251850 983634
rect 268120 983620 268148 986614
rect 280816 984842 280844 1006266
rect 300124 1006256 300176 1006262
rect 300124 1006198 300176 1006204
rect 298744 1006188 298796 1006194
rect 298744 1006130 298796 1006136
rect 298192 999184 298244 999190
rect 298192 999126 298244 999132
rect 298098 997792 298154 997801
rect 298020 997750 298098 997778
rect 284392 995852 284444 995858
rect 284392 995794 284444 995800
rect 294880 995852 294932 995858
rect 294880 995794 294932 995800
rect 284404 995738 284432 995794
rect 287978 995752 288034 995761
rect 284142 995710 284432 995738
rect 287822 995710 287978 995738
rect 291750 995752 291806 995761
rect 291502 995710 291750 995738
rect 287978 995687 288034 995696
rect 293590 995752 293646 995761
rect 293342 995710 293590 995738
rect 291750 995687 291806 995696
rect 294892 995738 294920 995794
rect 298020 995790 298048 997750
rect 298098 997727 298154 997736
rect 298204 995858 298232 999126
rect 298376 997756 298428 997762
rect 298376 997698 298428 997704
rect 298388 997257 298416 997698
rect 298374 997248 298430 997257
rect 298374 997183 298430 997192
rect 298284 996668 298336 996674
rect 298284 996610 298336 996616
rect 298192 995852 298244 995858
rect 298192 995794 298244 995800
rect 297272 995784 297324 995790
rect 294538 995710 294920 995738
rect 297022 995732 297272 995738
rect 297022 995726 297324 995732
rect 298008 995784 298060 995790
rect 298008 995726 298060 995732
rect 297022 995710 297312 995726
rect 293590 995687 293646 995696
rect 291106 995616 291162 995625
rect 290858 995574 291106 995602
rect 291106 995551 291162 995560
rect 292394 995480 292450 995489
rect 282840 995042 282868 995452
rect 283484 995217 283512 995452
rect 283470 995208 283526 995217
rect 283470 995143 283526 995152
rect 285968 995081 285996 995452
rect 286520 995110 286548 995452
rect 287164 995178 287192 995452
rect 290292 995353 290320 995452
rect 292146 995438 292394 995466
rect 295338 995480 295394 995489
rect 295182 995438 295338 995466
rect 292394 995415 292450 995424
rect 295338 995415 295394 995424
rect 290278 995344 290334 995353
rect 290278 995279 290334 995288
rect 298296 995217 298324 996610
rect 298756 996305 298784 1006130
rect 298928 1006120 298980 1006126
rect 298928 1006062 298980 1006068
rect 298742 996296 298798 996305
rect 298742 996231 298798 996240
rect 298940 995625 298968 1006062
rect 299020 996396 299072 996402
rect 299020 996338 299072 996344
rect 298926 995616 298982 995625
rect 298926 995551 298982 995560
rect 299032 995489 299060 996338
rect 300136 995897 300164 1006198
rect 300228 996674 300256 1006266
rect 300216 996668 300268 996674
rect 300216 996610 300268 996616
rect 300122 995888 300178 995897
rect 300122 995823 300178 995832
rect 299018 995480 299074 995489
rect 299018 995415 299074 995424
rect 300320 995353 300348 1006946
rect 426348 1006936 426400 1006942
rect 426346 1006904 426348 1006913
rect 429568 1006936 429620 1006942
rect 426400 1006904 426402 1006913
rect 426346 1006839 426402 1006848
rect 427174 1006904 427230 1006913
rect 429568 1006878 429620 1006884
rect 427174 1006839 427176 1006848
rect 427228 1006839 427230 1006848
rect 427176 1006810 427228 1006816
rect 425152 1006800 425204 1006806
rect 425150 1006768 425152 1006777
rect 425204 1006768 425206 1006777
rect 425150 1006703 425206 1006712
rect 427542 1006768 427598 1006777
rect 427542 1006703 427544 1006712
rect 427596 1006703 427598 1006712
rect 427544 1006674 427596 1006680
rect 428004 1006664 428056 1006670
rect 428002 1006632 428004 1006641
rect 428056 1006632 428058 1006641
rect 429580 1006602 429608 1006878
rect 440884 1006868 440936 1006874
rect 440884 1006810 440936 1006816
rect 428002 1006567 428058 1006576
rect 429568 1006596 429620 1006602
rect 429568 1006538 429620 1006544
rect 423496 1006528 423548 1006534
rect 423494 1006496 423496 1006505
rect 423548 1006496 423550 1006505
rect 423494 1006431 423550 1006440
rect 428370 1006496 428426 1006505
rect 428426 1006466 428504 1006482
rect 428426 1006460 428516 1006466
rect 428426 1006454 428464 1006460
rect 428370 1006431 428426 1006440
rect 428464 1006402 428516 1006408
rect 301504 1006392 301556 1006398
rect 310152 1006392 310204 1006398
rect 301504 1006334 301556 1006340
rect 308126 1006360 308182 1006369
rect 301516 996402 301544 1006334
rect 308126 1006295 308128 1006304
rect 308180 1006295 308182 1006304
rect 310150 1006360 310152 1006369
rect 425980 1006392 426032 1006398
rect 310204 1006360 310206 1006369
rect 310150 1006295 310206 1006304
rect 423862 1006360 423918 1006369
rect 423862 1006295 423864 1006304
rect 308128 1006266 308180 1006272
rect 423916 1006295 423918 1006304
rect 425978 1006360 425980 1006369
rect 426032 1006360 426034 1006369
rect 425978 1006295 426034 1006304
rect 423864 1006266 423916 1006272
rect 357348 1006256 357400 1006262
rect 306102 1006224 306158 1006233
rect 306102 1006159 306104 1006168
rect 306156 1006159 306158 1006168
rect 357346 1006224 357348 1006233
rect 374644 1006256 374696 1006262
rect 357400 1006224 357402 1006233
rect 357346 1006159 357402 1006168
rect 361394 1006224 361450 1006233
rect 430028 1006256 430080 1006262
rect 374644 1006198 374696 1006204
rect 424690 1006224 424746 1006233
rect 361394 1006159 361396 1006168
rect 306104 1006130 306156 1006136
rect 361448 1006159 361450 1006168
rect 369216 1006188 369268 1006194
rect 361396 1006130 361448 1006136
rect 369216 1006130 369268 1006136
rect 305644 1006120 305696 1006126
rect 304078 1006088 304134 1006097
rect 303528 1006052 303580 1006058
rect 304078 1006023 304080 1006032
rect 303528 1005994 303580 1006000
rect 304132 1006023 304134 1006032
rect 304906 1006088 304962 1006097
rect 304906 1006023 304908 1006032
rect 304080 1005994 304132 1006000
rect 304960 1006023 304962 1006032
rect 305642 1006088 305644 1006097
rect 358544 1006120 358596 1006126
rect 305696 1006088 305698 1006097
rect 305642 1006023 305698 1006032
rect 306470 1006088 306526 1006097
rect 310610 1006088 310666 1006097
rect 306470 1006023 306472 1006032
rect 304908 1005994 304960 1006000
rect 306524 1006023 306526 1006032
rect 307024 1006052 307076 1006058
rect 306472 1005994 306524 1006000
rect 310610 1006023 310612 1006032
rect 307024 1005994 307076 1006000
rect 310664 1006023 310666 1006032
rect 314658 1006088 314714 1006097
rect 354494 1006088 354550 1006097
rect 314658 1006023 314660 1006032
rect 310612 1005994 310664 1006000
rect 314712 1006023 314714 1006032
rect 330484 1006052 330536 1006058
rect 314660 1005994 314712 1006000
rect 330484 1005994 330536 1006000
rect 353116 1006052 353168 1006058
rect 355230 1006088 355286 1006097
rect 354550 1006046 355230 1006074
rect 354494 1006023 354496 1006032
rect 353116 1005994 353168 1006000
rect 354548 1006023 354550 1006032
rect 355230 1006023 355286 1006032
rect 356058 1006088 356114 1006097
rect 356058 1006023 356060 1006032
rect 354496 1005994 354548 1006000
rect 356112 1006023 356114 1006032
rect 358542 1006088 358544 1006097
rect 358596 1006088 358598 1006097
rect 358542 1006023 358598 1006032
rect 360844 1006052 360896 1006058
rect 356060 1005994 356112 1006000
rect 360844 1005994 360896 1006000
rect 302884 1001972 302936 1001978
rect 302884 1001914 302936 1001920
rect 302896 997121 302924 1001914
rect 303252 997824 303304 997830
rect 303250 997792 303252 997801
rect 303304 997792 303306 997801
rect 303250 997727 303306 997736
rect 302882 997112 302938 997121
rect 302882 997047 302938 997056
rect 301504 996396 301556 996402
rect 301504 996338 301556 996344
rect 300306 995344 300362 995353
rect 300306 995279 300362 995288
rect 298282 995208 298338 995217
rect 287152 995172 287204 995178
rect 298282 995143 298338 995152
rect 287152 995114 287204 995120
rect 286508 995104 286560 995110
rect 285954 995072 286010 995081
rect 282828 995036 282880 995042
rect 286508 995046 286560 995052
rect 285954 995007 286010 995016
rect 282828 994978 282880 994984
rect 303540 991506 303568 1005994
rect 304448 1004896 304500 1004902
rect 304448 1004838 304500 1004844
rect 306930 1004864 306986 1004873
rect 304264 1004828 304316 1004834
rect 304264 1004770 304316 1004776
rect 304276 995761 304304 1004770
rect 304262 995752 304318 995761
rect 304262 995687 304318 995696
rect 304460 995178 304488 1004838
rect 306930 1004799 306932 1004808
rect 306984 1004799 306986 1004808
rect 306932 1004770 306984 1004776
rect 305828 1004760 305880 1004766
rect 305828 1004702 305880 1004708
rect 305644 1004692 305696 1004698
rect 305644 1004634 305696 1004640
rect 305274 1002008 305330 1002017
rect 305274 1001943 305276 1001952
rect 305328 1001943 305330 1001952
rect 305276 1001914 305328 1001920
rect 304448 995172 304500 995178
rect 304448 995114 304500 995120
rect 305656 995110 305684 1004634
rect 305840 997830 305868 1004702
rect 305828 997824 305880 997830
rect 305828 997766 305880 997772
rect 307036 995994 307064 1005994
rect 307300 1004896 307352 1004902
rect 307298 1004864 307300 1004873
rect 307352 1004864 307354 1004873
rect 307298 1004799 307354 1004808
rect 308588 1004760 308640 1004766
rect 307758 1004728 307814 1004737
rect 307758 1004663 307760 1004672
rect 307812 1004663 307814 1004672
rect 308586 1004728 308588 1004737
rect 308640 1004728 308642 1004737
rect 308586 1004663 308642 1004672
rect 307760 1004634 307812 1004640
rect 311440 1002040 311492 1002046
rect 310150 1002008 310206 1002017
rect 310150 1001943 310152 1001952
rect 310204 1001943 310206 1001952
rect 311438 1002008 311440 1002017
rect 313372 1002040 313424 1002046
rect 311492 1002008 311494 1002017
rect 313372 1001982 313424 1001988
rect 311438 1001943 311494 1001952
rect 311900 1001972 311952 1001978
rect 310152 1001914 310204 1001920
rect 311900 1001914 311952 1001920
rect 307024 995988 307076 995994
rect 307024 995930 307076 995936
rect 305644 995104 305696 995110
rect 305644 995046 305696 995052
rect 311912 995042 311940 1001914
rect 312176 997960 312228 997966
rect 312174 997928 312176 997937
rect 312228 997928 312230 997937
rect 312174 997863 312230 997872
rect 313004 997824 313056 997830
rect 313002 997792 313004 997801
rect 313056 997792 313058 997801
rect 313002 997727 313058 997736
rect 313384 996130 313412 1001982
rect 327540 999184 327592 999190
rect 327540 999126 327592 999132
rect 314936 997960 314988 997966
rect 313830 997928 313886 997937
rect 314936 997902 314988 997908
rect 313830 997863 313832 997872
rect 313884 997863 313886 997872
rect 313832 997834 313884 997840
rect 314752 997824 314804 997830
rect 314752 997766 314804 997772
rect 314764 996198 314792 997766
rect 314752 996192 314804 996198
rect 314752 996134 314804 996140
rect 313372 996124 313424 996130
rect 313372 996066 313424 996072
rect 314948 996062 314976 997902
rect 316040 997892 316092 997898
rect 316040 997834 316092 997840
rect 315120 997824 315172 997830
rect 315118 997792 315120 997801
rect 315172 997792 315174 997801
rect 316052 997762 316080 997834
rect 319444 997824 319496 997830
rect 318062 997792 318118 997801
rect 315118 997727 315174 997736
rect 316040 997756 316092 997762
rect 319444 997766 319496 997772
rect 318062 997727 318118 997736
rect 316040 997698 316092 997704
rect 314936 996056 314988 996062
rect 314936 995998 314988 996004
rect 316408 995648 316460 995654
rect 316408 995590 316460 995596
rect 311900 995036 311952 995042
rect 311900 994978 311952 994984
rect 303528 991500 303580 991506
rect 303528 991442 303580 991448
rect 300492 990140 300544 990146
rect 300492 990082 300544 990088
rect 284300 985992 284352 985998
rect 284300 985934 284352 985940
rect 280804 984836 280856 984842
rect 280804 984778 280856 984784
rect 284312 983620 284340 985934
rect 300504 983620 300532 990082
rect 316420 983634 316448 995590
rect 318076 985998 318104 997727
rect 319456 997150 319484 997766
rect 319444 997144 319496 997150
rect 319444 997086 319496 997092
rect 327552 997082 327580 999126
rect 327540 997076 327592 997082
rect 327540 997018 327592 997024
rect 330496 987426 330524 1005994
rect 332600 997144 332652 997150
rect 332600 997086 332652 997092
rect 330484 987420 330536 987426
rect 330484 987362 330536 987368
rect 318064 985992 318116 985998
rect 318064 985934 318116 985940
rect 332612 983634 332640 997086
rect 353128 992934 353156 1005994
rect 354508 1005963 354536 1005994
rect 360566 1005408 360622 1005417
rect 360566 1005343 360568 1005352
rect 360620 1005343 360622 1005352
rect 360568 1005314 360620 1005320
rect 356520 1005304 356572 1005310
rect 356518 1005272 356520 1005281
rect 356572 1005272 356574 1005281
rect 356518 1005207 356574 1005216
rect 354588 1004692 354640 1004698
rect 354588 1004634 354640 1004640
rect 354600 998442 354628 1004634
rect 356520 1004624 356572 1004630
rect 356518 1004592 356520 1004601
rect 356572 1004592 356574 1004601
rect 356518 1004527 356574 1004536
rect 358084 1003944 358136 1003950
rect 358082 1003912 358084 1003921
rect 358136 1003912 358138 1003921
rect 358082 1003847 358138 1003856
rect 357072 1002040 357124 1002046
rect 358912 1002040 358964 1002046
rect 357072 1001982 357124 1001988
rect 357346 1002008 357402 1002017
rect 355784 1001972 355836 1001978
rect 355784 1001914 355836 1001920
rect 355796 998510 355824 1001914
rect 355784 998504 355836 998510
rect 355784 998446 355836 998452
rect 354588 998436 354640 998442
rect 354588 998378 354640 998384
rect 357084 995042 357112 1001982
rect 357346 1001943 357402 1001952
rect 358542 1002008 358598 1002017
rect 358910 1002008 358912 1002017
rect 358964 1002008 358966 1002017
rect 358542 1001943 358544 1001952
rect 357360 998782 357388 1001943
rect 358596 1001943 358598 1001952
rect 358728 1001972 358780 1001978
rect 358544 1001914 358596 1001920
rect 358910 1001943 358966 1001952
rect 359370 1002008 359426 1002017
rect 359370 1001943 359372 1001952
rect 358728 1001914 358780 1001920
rect 359424 1001943 359426 1001952
rect 360198 1002008 360254 1002017
rect 360198 1001943 360200 1001952
rect 359372 1001914 359424 1001920
rect 360252 1001943 360254 1001952
rect 360200 1001914 360252 1001920
rect 357348 998776 357400 998782
rect 357348 998718 357400 998724
rect 358740 998578 358768 1001914
rect 360200 998776 360252 998782
rect 360200 998718 360252 998724
rect 358728 998572 358780 998578
rect 358728 998514 358780 998520
rect 360212 995353 360240 998718
rect 360856 998646 360884 1005994
rect 363420 1004896 363472 1004902
rect 361762 1004864 361818 1004873
rect 361762 1004799 361764 1004808
rect 361816 1004799 361818 1004808
rect 363418 1004864 363420 1004873
rect 366364 1004896 366416 1004902
rect 363472 1004864 363474 1004873
rect 366364 1004838 366416 1004844
rect 363418 1004799 363474 1004808
rect 364984 1004828 365036 1004834
rect 361764 1004770 361816 1004776
rect 364984 1004770 365036 1004776
rect 364248 1004760 364300 1004766
rect 362590 1004728 362646 1004737
rect 362590 1004663 362592 1004672
rect 362644 1004663 362646 1004672
rect 364246 1004728 364248 1004737
rect 364300 1004728 364302 1004737
rect 364246 1004663 364302 1004672
rect 362592 1004634 362644 1004640
rect 361028 1002040 361080 1002046
rect 361026 1002008 361028 1002017
rect 363604 1002040 363656 1002046
rect 361080 1002008 361082 1002017
rect 363604 1001982 363656 1001988
rect 361026 1001943 361082 1001952
rect 362224 1001972 362276 1001978
rect 362224 1001914 362276 1001920
rect 360844 998640 360896 998646
rect 360844 998582 360896 998588
rect 360198 995344 360254 995353
rect 360198 995279 360254 995288
rect 362236 995217 362264 1001914
rect 363616 995489 363644 1001982
rect 364996 995994 365024 1004770
rect 365168 1004692 365220 1004698
rect 365168 1004634 365220 1004640
rect 365076 1002040 365128 1002046
rect 365074 1002008 365076 1002017
rect 365128 1002008 365130 1002017
rect 365074 1001943 365130 1001952
rect 365180 997014 365208 1004634
rect 365442 1002008 365498 1002017
rect 365442 1001943 365444 1001952
rect 365496 1001943 365498 1001952
rect 365444 1001914 365496 1001920
rect 365168 997008 365220 997014
rect 365168 996950 365220 996956
rect 366376 996130 366404 1004838
rect 366548 1004760 366600 1004766
rect 366548 1004702 366600 1004708
rect 366560 997393 366588 1004702
rect 369122 1002008 369178 1002017
rect 367744 1001972 367796 1001978
rect 369122 1001943 369178 1001952
rect 367744 1001914 367796 1001920
rect 367376 998640 367428 998646
rect 367376 998582 367428 998588
rect 366546 997384 366602 997393
rect 366546 997319 366602 997328
rect 366364 996124 366416 996130
rect 366364 996066 366416 996072
rect 367388 996062 367416 998582
rect 367376 996056 367428 996062
rect 367376 995998 367428 996004
rect 364984 995988 365036 995994
rect 364984 995930 365036 995936
rect 363602 995480 363658 995489
rect 363602 995415 363658 995424
rect 362222 995208 362278 995217
rect 362222 995143 362278 995152
rect 357072 995036 357124 995042
rect 357072 994978 357124 994984
rect 353116 992928 353168 992934
rect 353116 992870 353168 992876
rect 365444 987420 365496 987426
rect 365444 987362 365496 987368
rect 349160 985992 349212 985998
rect 349160 985934 349212 985940
rect 316420 983606 316802 983634
rect 332612 983606 332994 983634
rect 349172 983620 349200 985934
rect 365456 983620 365484 987362
rect 367756 986066 367784 1001914
rect 367836 997076 367888 997082
rect 367836 997018 367888 997024
rect 367848 991574 367876 997018
rect 367836 991568 367888 991574
rect 367836 991510 367888 991516
rect 367744 986060 367796 986066
rect 367744 986002 367796 986008
rect 369136 985998 369164 1001943
rect 369228 998374 369256 1006130
rect 371884 1006120 371936 1006126
rect 371884 1006062 371936 1006068
rect 370504 1002040 370556 1002046
rect 370504 1001982 370556 1001988
rect 369216 998368 369268 998374
rect 369216 998310 369268 998316
rect 369214 997384 369270 997393
rect 369214 997319 369216 997328
rect 369268 997319 369270 997328
rect 369216 997290 369268 997296
rect 369216 995512 369268 995518
rect 369214 995480 369216 995489
rect 369268 995480 369270 995489
rect 369214 995415 369270 995424
rect 370516 990146 370544 1001982
rect 371896 996282 371924 1006062
rect 372436 998572 372488 998578
rect 372436 998514 372488 998520
rect 372344 998368 372396 998374
rect 372342 998336 372344 998345
rect 372396 998336 372398 998345
rect 372342 998271 372398 998280
rect 372344 997348 372396 997354
rect 372344 997290 372396 997296
rect 372356 997257 372384 997290
rect 372342 997248 372398 997257
rect 372342 997183 372398 997192
rect 372344 997008 372396 997014
rect 372342 996976 372344 996985
rect 372396 996976 372398 996985
rect 372342 996911 372398 996920
rect 372342 996296 372398 996305
rect 371896 996254 372342 996282
rect 372342 996231 372398 996240
rect 372448 995625 372476 998514
rect 374656 995897 374684 1006198
rect 424690 1006159 424692 1006168
rect 424744 1006159 424746 1006168
rect 430026 1006224 430028 1006233
rect 430080 1006224 430082 1006233
rect 430026 1006159 430082 1006168
rect 424692 1006130 424744 1006136
rect 425520 1006120 425572 1006126
rect 422666 1006088 422722 1006097
rect 420736 1006052 420788 1006058
rect 422666 1006023 422668 1006032
rect 420736 1005994 420788 1006000
rect 422720 1006023 422722 1006032
rect 425518 1006088 425520 1006097
rect 425572 1006088 425574 1006097
rect 425518 1006023 425574 1006032
rect 422668 1005994 422720 1006000
rect 380164 1005372 380216 1005378
rect 380164 1005314 380216 1005320
rect 377404 1005304 377456 1005310
rect 377404 1005246 377456 1005252
rect 377416 996169 377444 1005246
rect 378324 1003944 378376 1003950
rect 378324 1003886 378376 1003892
rect 377402 996160 377458 996169
rect 377402 996095 377458 996104
rect 374642 995888 374698 995897
rect 374642 995823 374698 995832
rect 378336 995761 378364 1003886
rect 380176 998646 380204 1005314
rect 420748 1001978 420776 1005994
rect 428832 1005440 428884 1005446
rect 428830 1005408 428832 1005417
rect 428884 1005408 428886 1005417
rect 428830 1005343 428886 1005352
rect 432878 1005408 432934 1005417
rect 432878 1005343 432880 1005352
rect 432932 1005343 432934 1005352
rect 432880 1005314 432932 1005320
rect 432512 1005304 432564 1005310
rect 432510 1005272 432512 1005281
rect 432564 1005272 432566 1005281
rect 432510 1005207 432566 1005216
rect 421470 1002008 421526 1002017
rect 420736 1001972 420788 1001978
rect 421470 1001943 421472 1001952
rect 420736 1001914 420788 1001920
rect 421524 1001943 421526 1001952
rect 424322 1002008 424378 1002017
rect 426346 1002008 426402 1002017
rect 424322 1001943 424324 1001952
rect 421472 1001914 421524 1001920
rect 424376 1001943 424378 1001952
rect 425704 1001972 425756 1001978
rect 424324 1001914 424376 1001920
rect 426346 1001943 426402 1001952
rect 425704 1001914 425756 1001920
rect 380164 998640 380216 998646
rect 380164 998582 380216 998588
rect 383568 998640 383620 998646
rect 383620 998588 383700 998594
rect 383568 998582 383700 998588
rect 383580 998566 383700 998582
rect 383384 998504 383436 998510
rect 383384 998446 383436 998452
rect 381544 996056 381596 996062
rect 381544 995998 381596 996004
rect 381556 995926 381584 995998
rect 382108 995994 382320 996010
rect 382096 995988 382332 995994
rect 382148 995982 382280 995988
rect 382096 995930 382148 995936
rect 382280 995930 382332 995936
rect 381544 995920 381596 995926
rect 381544 995862 381596 995868
rect 383396 995858 383424 998446
rect 383568 998436 383620 998442
rect 383568 998378 383620 998384
rect 383474 998336 383530 998345
rect 383474 998271 383530 998280
rect 383384 995852 383436 995858
rect 383384 995794 383436 995800
rect 378322 995752 378378 995761
rect 383488 995722 383516 998271
rect 383580 997801 383608 998378
rect 383566 997792 383622 997801
rect 383566 997727 383622 997736
rect 383672 995790 383700 998566
rect 400128 997824 400180 997830
rect 400128 997766 400180 997772
rect 399944 997756 399996 997762
rect 399944 997698 399996 997704
rect 399956 997257 399984 997698
rect 400036 997688 400088 997694
rect 400036 997630 400088 997636
rect 399942 997248 399998 997257
rect 399942 997183 399998 997192
rect 400048 996985 400076 997630
rect 400034 996976 400090 996985
rect 400034 996911 400090 996920
rect 400140 995858 400168 997766
rect 385040 995852 385092 995858
rect 385040 995794 385092 995800
rect 393596 995852 393648 995858
rect 393596 995794 393648 995800
rect 396632 995852 396684 995858
rect 396632 995794 396684 995800
rect 400128 995852 400180 995858
rect 400128 995794 400180 995800
rect 383660 995784 383712 995790
rect 383660 995726 383712 995732
rect 384396 995784 384448 995790
rect 385052 995738 385080 995794
rect 388626 995752 388682 995761
rect 384448 995732 384698 995738
rect 384396 995726 384698 995732
rect 378322 995687 378378 995696
rect 383476 995716 383528 995722
rect 384408 995710 384698 995726
rect 385052 995710 385342 995738
rect 385696 995722 385986 995738
rect 385684 995716 385986 995722
rect 383476 995658 383528 995664
rect 385736 995710 385986 995716
rect 389362 995752 389418 995761
rect 388682 995710 389022 995738
rect 388626 995687 388682 995696
rect 392398 995752 392454 995761
rect 389418 995710 389666 995738
rect 389362 995687 389418 995696
rect 393410 995752 393466 995761
rect 392454 995710 392702 995738
rect 393346 995710 393410 995738
rect 392398 995687 392454 995696
rect 393608 995738 393636 995794
rect 396644 995738 396672 995794
rect 393608 995710 393990 995738
rect 396382 995710 396672 995738
rect 393410 995687 393466 995696
rect 385684 995658 385736 995664
rect 372434 995616 372490 995625
rect 372434 995551 372490 995560
rect 391938 995616 391994 995625
rect 391994 995574 392150 995602
rect 391938 995551 391994 995560
rect 372344 995512 372396 995518
rect 372342 995480 372344 995489
rect 372396 995480 372398 995489
rect 396722 995480 396778 995489
rect 372342 995415 372398 995424
rect 370780 995376 370832 995382
rect 370778 995344 370780 995353
rect 372344 995376 372396 995382
rect 370832 995344 370834 995353
rect 370778 995279 370834 995288
rect 372342 995344 372344 995353
rect 372396 995344 372398 995353
rect 372342 995279 372398 995288
rect 370780 995240 370832 995246
rect 370778 995208 370780 995217
rect 372344 995240 372396 995246
rect 370832 995208 370834 995217
rect 370778 995143 370834 995152
rect 372342 995208 372344 995217
rect 387812 995217 387840 995452
rect 388088 995438 388378 995466
rect 372396 995208 372398 995217
rect 372342 995143 372398 995152
rect 387798 995208 387854 995217
rect 387798 995143 387854 995152
rect 388088 995081 388116 995438
rect 395172 995353 395200 995452
rect 396778 995438 397026 995466
rect 396722 995415 396778 995424
rect 395158 995344 395214 995353
rect 395158 995279 395214 995288
rect 388074 995072 388130 995081
rect 398852 995042 398880 995452
rect 388074 995007 388130 995016
rect 398840 995036 398892 995042
rect 398840 994978 398892 994984
rect 420748 991574 420776 1001914
rect 425716 1001230 425744 1001914
rect 425704 1001224 425756 1001230
rect 425704 1001166 425756 1001172
rect 426360 999802 426388 1001943
rect 438768 1001224 438820 1001230
rect 438768 1001166 438820 1001172
rect 426348 999796 426400 999802
rect 426348 999738 426400 999744
rect 430854 998200 430910 998209
rect 430854 998135 430856 998144
rect 430908 998135 430910 998144
rect 436744 998164 436796 998170
rect 430856 998106 430908 998112
rect 436744 998106 436796 998112
rect 429660 998096 429712 998102
rect 429658 998064 429660 998073
rect 431960 998096 432012 998102
rect 429712 998064 429714 998073
rect 428464 998028 428516 998034
rect 429658 997999 429714 998008
rect 430854 998064 430910 998073
rect 430854 997999 430856 998008
rect 428464 997970 428516 997976
rect 430908 997999 430910 998008
rect 431682 998064 431738 998073
rect 431960 998038 432012 998044
rect 431682 997999 431684 998008
rect 430856 997970 430908 997976
rect 431736 997999 431738 998008
rect 431684 997970 431736 997976
rect 428476 996130 428504 997970
rect 430396 997960 430448 997966
rect 429198 997928 429254 997937
rect 429198 997863 429200 997872
rect 429252 997863 429254 997872
rect 430394 997928 430396 997937
rect 430448 997928 430450 997937
rect 430394 997863 430450 997872
rect 431224 997892 431276 997898
rect 429200 997834 429252 997840
rect 431224 997834 431276 997840
rect 431236 996198 431264 997834
rect 431224 996192 431276 996198
rect 431224 996134 431276 996140
rect 428464 996124 428516 996130
rect 428464 996066 428516 996072
rect 431972 995994 432000 998038
rect 433984 998028 434036 998034
rect 433984 997970 434036 997976
rect 432144 997960 432196 997966
rect 432050 997928 432106 997937
rect 432144 997902 432196 997908
rect 432050 997863 432052 997872
rect 432104 997863 432106 997872
rect 432052 997834 432104 997840
rect 432156 997754 432184 997902
rect 433432 997892 433484 997898
rect 433432 997834 433484 997840
rect 433444 997762 433472 997834
rect 432064 997726 432184 997754
rect 433432 997756 433484 997762
rect 432064 997694 432092 997726
rect 433432 997698 433484 997704
rect 432052 997688 432104 997694
rect 432052 997630 432104 997636
rect 433996 997393 434024 997970
rect 435362 997792 435418 997801
rect 435362 997727 435418 997736
rect 433982 997384 434038 997393
rect 433982 997319 434038 997328
rect 431960 995988 432012 995994
rect 431960 995930 432012 995936
rect 381636 991568 381688 991574
rect 381636 991510 381688 991516
rect 420736 991568 420788 991574
rect 420736 991510 420788 991516
rect 370504 990140 370556 990146
rect 370504 990082 370556 990088
rect 369124 985992 369176 985998
rect 369124 985934 369176 985940
rect 381648 983620 381676 991510
rect 435376 990146 435404 997727
rect 436558 997384 436614 997393
rect 436558 997319 436614 997328
rect 436572 997286 436600 997319
rect 436560 997280 436612 997286
rect 436560 997222 436612 997228
rect 436756 995994 436784 998106
rect 436744 995988 436796 995994
rect 436744 995930 436796 995936
rect 438780 995382 438808 1001166
rect 440240 997756 440292 997762
rect 440240 997698 440292 997704
rect 439688 997280 439740 997286
rect 439686 997248 439688 997257
rect 439740 997248 439742 997257
rect 439686 997183 439742 997192
rect 438768 995376 438820 995382
rect 439688 995376 439740 995382
rect 438768 995318 438820 995324
rect 439686 995344 439688 995353
rect 439740 995344 439742 995353
rect 439686 995279 439742 995288
rect 440252 994294 440280 997698
rect 440896 995217 440924 1006810
rect 469864 1006800 469916 1006806
rect 469864 1006742 469916 1006748
rect 443644 1006732 443696 1006738
rect 443644 1006674 443696 1006680
rect 441620 1006596 441672 1006602
rect 441620 1006538 441672 1006544
rect 441632 998442 441660 1006538
rect 441620 998436 441672 998442
rect 441620 998378 441672 998384
rect 443656 998345 443684 1006674
rect 448612 1006664 448664 1006670
rect 448612 1006606 448664 1006612
rect 446404 1006528 446456 1006534
rect 446404 1006470 446456 1006476
rect 446312 999796 446364 999802
rect 446312 999738 446364 999744
rect 443642 998336 443698 998345
rect 443642 998271 443698 998280
rect 440882 995208 440938 995217
rect 440882 995143 440938 995152
rect 446324 995081 446352 999738
rect 446416 999122 446444 1006470
rect 448520 1005440 448572 1005446
rect 448520 1005382 448572 1005388
rect 446404 999116 446456 999122
rect 446404 999058 446456 999064
rect 448532 998510 448560 1005382
rect 448624 1003950 448652 1006606
rect 457444 1006460 457496 1006466
rect 457444 1006402 457496 1006408
rect 451924 1006392 451976 1006398
rect 451924 1006334 451976 1006340
rect 448612 1003944 448664 1003950
rect 448612 1003886 448664 1003892
rect 448612 999116 448664 999122
rect 448612 999058 448664 999064
rect 448520 998504 448572 998510
rect 448520 998446 448572 998452
rect 448624 996305 448652 999058
rect 448610 996296 448666 996305
rect 448610 996231 448666 996240
rect 451936 995489 451964 1006334
rect 454684 1006324 454736 1006330
rect 454684 1006266 454736 1006272
rect 454696 996169 454724 1006266
rect 454682 996160 454738 996169
rect 454682 996095 454738 996104
rect 451922 995480 451978 995489
rect 451922 995415 451978 995424
rect 446310 995072 446366 995081
rect 457456 995042 457484 1006402
rect 468484 1006256 468536 1006262
rect 468484 1006198 468536 1006204
rect 460204 1006188 460256 1006194
rect 460204 1006130 460256 1006136
rect 460216 995110 460244 1006130
rect 464988 1006120 465040 1006126
rect 464988 1006062 465040 1006068
rect 462320 1005372 462372 1005378
rect 462320 1005314 462372 1005320
rect 460204 995104 460256 995110
rect 460204 995046 460256 995052
rect 446310 995007 446366 995016
rect 457444 995036 457496 995042
rect 457444 994978 457496 994984
rect 440240 994288 440292 994294
rect 440240 994230 440292 994236
rect 446128 994288 446180 994294
rect 446128 994230 446180 994236
rect 430304 990140 430356 990146
rect 430304 990082 430356 990088
rect 435364 990140 435416 990146
rect 435364 990082 435416 990088
rect 397828 986060 397880 986066
rect 397828 986002 397880 986008
rect 397840 983620 397868 986002
rect 414112 985992 414164 985998
rect 414112 985934 414164 985940
rect 414124 983620 414152 985934
rect 430316 983620 430344 990082
rect 446140 983634 446168 994230
rect 462332 983634 462360 1005314
rect 464804 1003944 464856 1003950
rect 464804 1003886 464856 1003892
rect 464816 998782 464844 1003886
rect 465000 1001978 465028 1006062
rect 467104 1005304 467156 1005310
rect 467104 1005246 467156 1005252
rect 464988 1001972 465040 1001978
rect 464988 1001914 465040 1001920
rect 464804 998776 464856 998782
rect 464804 998718 464856 998724
rect 467116 985998 467144 1005246
rect 468496 996062 468524 1006198
rect 468484 996056 468536 996062
rect 468484 995998 468536 996004
rect 469876 995625 469904 1006742
rect 508686 1006496 508742 1006505
rect 508686 1006431 508688 1006440
rect 508740 1006431 508742 1006440
rect 515404 1006460 515456 1006466
rect 508688 1006402 508740 1006408
rect 515404 1006402 515456 1006408
rect 501326 1006360 501382 1006369
rect 501326 1006295 501328 1006304
rect 501380 1006295 501382 1006304
rect 501328 1006266 501380 1006272
rect 505836 1006256 505888 1006262
rect 505834 1006224 505836 1006233
rect 514760 1006256 514812 1006262
rect 505888 1006224 505890 1006233
rect 514760 1006198 514812 1006204
rect 505834 1006159 505890 1006168
rect 498108 1006120 498160 1006126
rect 499672 1006120 499724 1006126
rect 498108 1006062 498160 1006068
rect 499670 1006088 499672 1006097
rect 504548 1006120 504600 1006126
rect 499724 1006088 499726 1006097
rect 498120 1001994 498148 1006062
rect 499670 1006023 499726 1006032
rect 504546 1006088 504548 1006097
rect 504600 1006088 504602 1006097
rect 504546 1006023 504602 1006032
rect 505374 1006088 505430 1006097
rect 505374 1006023 505376 1006032
rect 505428 1006023 505430 1006032
rect 505376 1005994 505428 1006000
rect 509882 1005408 509938 1005417
rect 509882 1005343 509884 1005352
rect 509936 1005343 509938 1005352
rect 509884 1005314 509936 1005320
rect 502892 1005304 502944 1005310
rect 502890 1005272 502892 1005281
rect 502944 1005272 502946 1005281
rect 502890 1005207 502946 1005216
rect 501694 1004864 501750 1004873
rect 499212 1004828 499264 1004834
rect 501694 1004799 501696 1004808
rect 499212 1004770 499264 1004776
rect 501748 1004799 501750 1004808
rect 501696 1004770 501748 1004776
rect 498474 1002008 498530 1002017
rect 472532 1001972 472584 1001978
rect 472532 1001914 472584 1001920
rect 498028 1001966 498474 1001994
rect 472440 998776 472492 998782
rect 472440 998718 472492 998724
rect 472348 998572 472400 998578
rect 472348 998514 472400 998520
rect 469862 995616 469918 995625
rect 472360 995586 472388 998514
rect 472452 995722 472480 998718
rect 472544 995858 472572 1001914
rect 472624 998368 472676 998374
rect 472624 998310 472676 998316
rect 472714 998336 472770 998345
rect 472532 995852 472584 995858
rect 472532 995794 472584 995800
rect 472636 995790 472664 998310
rect 472714 998271 472770 998280
rect 472624 995784 472676 995790
rect 472624 995726 472676 995732
rect 472440 995716 472492 995722
rect 472440 995658 472492 995664
rect 472728 995654 472756 998271
rect 488908 997756 488960 997762
rect 488908 997698 488960 997704
rect 488920 997257 488948 997698
rect 488906 997248 488962 997257
rect 488906 997183 488962 997192
rect 477684 995852 477736 995858
rect 477684 995794 477736 995800
rect 474004 995784 474056 995790
rect 473372 995722 473662 995738
rect 477696 995738 477724 995794
rect 481546 995752 481602 995761
rect 474056 995732 474306 995738
rect 474004 995726 474306 995732
rect 473360 995716 473662 995722
rect 473412 995710 473662 995716
rect 474016 995710 474306 995726
rect 477696 995710 477986 995738
rect 482650 995752 482706 995761
rect 481602 995710 481666 995738
rect 481546 995687 481602 995696
rect 485594 995752 485650 995761
rect 482706 995710 482954 995738
rect 485346 995710 485594 995738
rect 482650 995687 482706 995696
rect 485594 995687 485650 995696
rect 473360 995658 473412 995664
rect 472716 995648 472768 995654
rect 476396 995648 476448 995654
rect 472716 995590 472768 995596
rect 474752 995586 474950 995602
rect 483754 995616 483810 995625
rect 476448 995596 476790 995602
rect 476396 995590 476790 995596
rect 469862 995551 469918 995560
rect 472348 995580 472400 995586
rect 472348 995522 472400 995528
rect 474740 995580 474950 995586
rect 474792 995574 474950 995580
rect 476408 995574 476790 995590
rect 483810 995574 484150 995602
rect 483754 995551 483810 995560
rect 474740 995522 474792 995528
rect 476946 995480 477002 995489
rect 477002 995438 477342 995466
rect 476946 995415 477002 995424
rect 478616 995353 478644 995452
rect 478602 995344 478658 995353
rect 478602 995279 478658 995288
rect 481100 995217 481128 995452
rect 481086 995208 481142 995217
rect 481086 995143 481142 995152
rect 482296 995110 482324 995452
rect 482284 995104 482336 995110
rect 482284 995046 482336 995052
rect 485976 995042 486004 995452
rect 487816 995081 487844 995452
rect 487802 995072 487858 995081
rect 485964 995036 486016 995042
rect 487802 995007 487858 995016
rect 485964 994978 486016 994984
rect 498028 993002 498056 1001966
rect 498474 1001943 498530 1001952
rect 499224 995042 499252 1004770
rect 499488 1004760 499540 1004766
rect 500500 1004760 500552 1004766
rect 499488 1004702 499540 1004708
rect 500498 1004728 500500 1004737
rect 504364 1004760 504416 1004766
rect 500552 1004728 500554 1004737
rect 499396 1004556 499448 1004562
rect 499396 1004498 499448 1004504
rect 499408 999802 499436 1004498
rect 499500 1003542 499528 1004702
rect 504364 1004702 504416 1004708
rect 500498 1004663 500554 1004672
rect 500500 1004624 500552 1004630
rect 500498 1004592 500500 1004601
rect 500552 1004592 500554 1004601
rect 500498 1004527 500554 1004536
rect 501326 1004592 501382 1004601
rect 501326 1004527 501328 1004536
rect 501380 1004527 501382 1004536
rect 501328 1004498 501380 1004504
rect 499488 1003536 499540 1003542
rect 499488 1003478 499540 1003484
rect 500960 1003536 501012 1003542
rect 500960 1003478 501012 1003484
rect 500868 1002040 500920 1002046
rect 500868 1001982 500920 1001988
rect 499396 999796 499448 999802
rect 499396 999738 499448 999744
rect 500880 998510 500908 1001982
rect 500868 998504 500920 998510
rect 500868 998446 500920 998452
rect 500972 995217 501000 1003478
rect 502522 1002144 502578 1002153
rect 502522 1002079 502524 1002088
rect 502576 1002079 502578 1002088
rect 502524 1002050 502576 1002056
rect 503352 1002040 503404 1002046
rect 502890 1002008 502946 1002017
rect 502156 1001972 502208 1001978
rect 502890 1001943 502892 1001952
rect 502156 1001914 502208 1001920
rect 502944 1001943 502946 1001952
rect 503350 1002008 503352 1002017
rect 503404 1002008 503406 1002017
rect 503350 1001943 503406 1001952
rect 502892 1001914 502944 1001920
rect 502168 998442 502196 1001914
rect 504272 999796 504324 999802
rect 504272 999738 504324 999744
rect 502156 998436 502208 998442
rect 502156 998378 502208 998384
rect 500958 995208 501014 995217
rect 504284 995178 504312 999738
rect 500958 995143 501014 995152
rect 504272 995172 504324 995178
rect 504272 995114 504324 995120
rect 504376 995110 504404 1004702
rect 514772 1004154 514800 1006198
rect 514760 1004148 514812 1004154
rect 514760 1004090 514812 1004096
rect 505100 1002108 505152 1002114
rect 505100 1002050 505152 1002056
rect 505006 1002008 505062 1002017
rect 505006 1001943 505008 1001952
rect 505060 1001943 505062 1001952
rect 505008 1001914 505060 1001920
rect 505112 999802 505140 1002050
rect 506664 1001972 506716 1001978
rect 506664 1001914 506716 1001920
rect 505100 999796 505152 999802
rect 505100 999738 505152 999744
rect 506676 998306 506704 1001914
rect 513288 998504 513340 998510
rect 513288 998446 513340 998452
rect 506664 998300 506716 998306
rect 506664 998242 506716 998248
rect 507032 998096 507084 998102
rect 507030 998064 507032 998073
rect 510068 998096 510120 998102
rect 507084 998064 507086 998073
rect 507030 997999 507086 998008
rect 508226 998064 508282 998073
rect 510068 998038 510120 998044
rect 508226 997999 508228 998008
rect 508280 997999 508282 998008
rect 508228 997970 508280 997976
rect 507860 997960 507912 997966
rect 506202 997928 506258 997937
rect 506202 997863 506204 997872
rect 506256 997863 506258 997872
rect 507858 997928 507860 997937
rect 509884 997960 509936 997966
rect 507912 997928 507914 997937
rect 509054 997928 509110 997937
rect 507858 997863 507914 997872
rect 508504 997892 508556 997898
rect 506204 997834 506256 997840
rect 509884 997902 509936 997908
rect 509054 997863 509056 997872
rect 508504 997834 508556 997840
rect 509108 997863 509110 997872
rect 509056 997834 509108 997840
rect 507400 997824 507452 997830
rect 506570 997792 506626 997801
rect 506570 997727 506626 997736
rect 507398 997792 507400 997801
rect 507452 997792 507454 997801
rect 507398 997727 507454 997736
rect 506584 996198 506612 997727
rect 508516 996198 508544 997834
rect 509240 997824 509292 997830
rect 509516 997824 509568 997830
rect 509240 997766 509292 997772
rect 509514 997792 509516 997801
rect 509568 997792 509570 997801
rect 506572 996192 506624 996198
rect 506572 996134 506624 996140
rect 508504 996192 508556 996198
rect 508504 996134 508556 996140
rect 509252 996062 509280 997766
rect 509514 997727 509570 997736
rect 509896 996130 509924 997902
rect 509884 996124 509936 996130
rect 509884 996066 509936 996072
rect 510080 996062 510108 998038
rect 510896 998028 510948 998034
rect 510896 997970 510948 997976
rect 510712 997892 510764 997898
rect 510712 997834 510764 997840
rect 510724 997762 510752 997834
rect 510712 997756 510764 997762
rect 510712 997698 510764 997704
rect 509240 996056 509292 996062
rect 509240 995998 509292 996004
rect 510068 996056 510120 996062
rect 510068 995998 510120 996004
rect 510908 995994 510936 997970
rect 512642 997792 512698 997801
rect 512642 997727 512698 997736
rect 510896 995988 510948 995994
rect 510896 995930 510948 995936
rect 511078 995888 511134 995897
rect 511078 995823 511134 995832
rect 504364 995104 504416 995110
rect 504364 995046 504416 995052
rect 499212 995036 499264 995042
rect 499212 994978 499264 994984
rect 498016 992996 498068 993002
rect 498016 992938 498068 992944
rect 478972 990140 479024 990146
rect 478972 990082 479024 990088
rect 467104 985992 467156 985998
rect 467104 985934 467156 985940
rect 446140 983606 446522 983634
rect 462332 983606 462806 983634
rect 478984 983620 479012 990082
rect 495164 985992 495216 985998
rect 495164 985934 495216 985940
rect 495176 983620 495204 985934
rect 511092 983634 511120 995823
rect 512656 987426 512684 997727
rect 513300 995518 513328 998446
rect 514024 997824 514076 997830
rect 514024 997766 514076 997772
rect 513288 995512 513340 995518
rect 513288 995454 513340 995460
rect 514036 990146 514064 997766
rect 515416 997286 515444 1006402
rect 551928 1006392 551980 1006398
rect 551926 1006360 551928 1006369
rect 574744 1006392 574796 1006398
rect 551980 1006360 551982 1006369
rect 517520 1006324 517572 1006330
rect 551926 1006295 551982 1006304
rect 553950 1006360 554006 1006369
rect 574744 1006334 574796 1006340
rect 553950 1006295 553952 1006304
rect 517520 1006266 517572 1006272
rect 554004 1006295 554006 1006304
rect 563796 1006324 563848 1006330
rect 553952 1006266 554004 1006272
rect 563796 1006266 563848 1006272
rect 515956 999796 516008 999802
rect 515956 999738 516008 999744
rect 515404 997280 515456 997286
rect 515404 997222 515456 997228
rect 515968 995654 515996 999738
rect 517532 998442 517560 1006266
rect 555976 1006256 556028 1006262
rect 555974 1006224 555976 1006233
rect 556028 1006224 556030 1006233
rect 520832 1006188 520884 1006194
rect 555974 1006159 556030 1006168
rect 557170 1006224 557226 1006233
rect 557170 1006159 557172 1006168
rect 520832 1006130 520884 1006136
rect 557224 1006159 557226 1006168
rect 557172 1006130 557224 1006136
rect 517612 1005304 517664 1005310
rect 517612 1005246 517664 1005252
rect 517624 998510 517652 1005246
rect 517980 1004148 518032 1004154
rect 517980 1004090 518032 1004096
rect 517612 998504 517664 998510
rect 517992 998481 518020 1004090
rect 517612 998446 517664 998452
rect 517978 998472 518034 998481
rect 516048 998436 516100 998442
rect 516048 998378 516100 998384
rect 517520 998436 517572 998442
rect 517978 998407 518034 998416
rect 517520 998378 517572 998384
rect 516060 995790 516088 998378
rect 516690 998336 516746 998345
rect 516690 998271 516692 998280
rect 516744 998271 516746 998280
rect 516692 998242 516744 998248
rect 516692 997280 516744 997286
rect 516690 997248 516692 997257
rect 516744 997248 516746 997257
rect 516690 997183 516746 997192
rect 520844 995858 520872 1006130
rect 522304 1006120 522356 1006126
rect 522304 1006062 522356 1006068
rect 549168 1006120 549220 1006126
rect 550272 1006120 550324 1006126
rect 549168 1006062 549220 1006068
rect 550270 1006088 550272 1006097
rect 551100 1006120 551152 1006126
rect 550324 1006088 550326 1006097
rect 520924 1005372 520976 1005378
rect 520924 1005314 520976 1005320
rect 520832 995852 520884 995858
rect 520832 995794 520884 995800
rect 516048 995784 516100 995790
rect 516692 995784 516744 995790
rect 516048 995726 516100 995732
rect 516690 995752 516692 995761
rect 516744 995752 516746 995761
rect 516690 995687 516746 995696
rect 515956 995648 516008 995654
rect 516692 995648 516744 995654
rect 515956 995590 516008 995596
rect 516690 995616 516692 995625
rect 516744 995616 516746 995625
rect 516690 995551 516746 995560
rect 516692 995512 516744 995518
rect 516690 995480 516692 995489
rect 516744 995480 516746 995489
rect 516690 995415 516746 995424
rect 515220 995376 515272 995382
rect 515218 995344 515220 995353
rect 516692 995376 516744 995382
rect 515272 995344 515274 995353
rect 515218 995279 515274 995288
rect 516690 995344 516692 995353
rect 516744 995344 516746 995353
rect 516690 995279 516746 995288
rect 515218 995208 515274 995217
rect 515218 995143 515220 995152
rect 515272 995143 515274 995152
rect 516690 995208 516746 995217
rect 516690 995143 516692 995152
rect 515220 995114 515272 995120
rect 516744 995143 516746 995152
rect 516692 995114 516744 995120
rect 514024 990140 514076 990146
rect 514024 990082 514076 990088
rect 512644 987420 512696 987426
rect 512644 987362 512696 987368
rect 520936 985794 520964 1005314
rect 522316 995314 522344 1006062
rect 523868 998504 523920 998510
rect 523868 998446 523920 998452
rect 523958 998472 524014 998481
rect 523776 998436 523828 998442
rect 523776 998378 523828 998384
rect 523788 995722 523816 998378
rect 523880 995926 523908 998446
rect 523958 998407 524014 998416
rect 523972 996441 524000 998407
rect 524050 998336 524106 998345
rect 524050 998271 524106 998280
rect 523958 996432 524014 996441
rect 523958 996367 524014 996376
rect 523868 995920 523920 995926
rect 523868 995862 523920 995868
rect 524064 995790 524092 998271
rect 540336 997824 540388 997830
rect 540336 997766 540388 997772
rect 540348 995858 540376 997766
rect 540888 997688 540940 997694
rect 540888 997630 540940 997636
rect 540900 997257 540928 997630
rect 540886 997248 540942 997257
rect 540886 997183 540942 997192
rect 527916 995852 527968 995858
rect 527916 995794 527968 995800
rect 528560 995852 528612 995858
rect 528560 995794 528612 995800
rect 536840 995852 536892 995858
rect 536840 995794 536892 995800
rect 540336 995852 540388 995858
rect 540336 995794 540388 995800
rect 524052 995784 524104 995790
rect 524052 995726 524104 995732
rect 524788 995784 524840 995790
rect 525338 995752 525394 995761
rect 524840 995732 525090 995738
rect 524788 995726 525090 995732
rect 523776 995716 523828 995722
rect 524800 995710 525090 995726
rect 526166 995752 526222 995761
rect 525394 995710 525734 995738
rect 525338 995687 525394 995696
rect 527928 995738 527956 995794
rect 528572 995738 528600 995794
rect 536852 995738 536880 995794
rect 526222 995710 526378 995738
rect 527928 995710 528218 995738
rect 528572 995710 528770 995738
rect 529768 995722 530058 995738
rect 529756 995716 530058 995722
rect 526166 995687 526222 995696
rect 523776 995658 523828 995664
rect 529808 995710 530058 995716
rect 536774 995710 536880 995738
rect 529756 995658 529808 995664
rect 529018 995616 529074 995625
rect 529074 995574 529414 995602
rect 529018 995551 529074 995560
rect 538954 995480 539010 995489
rect 532160 995438 532542 995466
rect 532712 995438 533094 995466
rect 532160 995353 532188 995438
rect 532146 995344 532202 995353
rect 522304 995308 522356 995314
rect 532146 995279 532202 995288
rect 522304 995250 522356 995256
rect 532606 995208 532662 995217
rect 532712 995194 532740 995438
rect 532662 995166 532740 995194
rect 533724 995178 533752 995452
rect 533712 995172 533764 995178
rect 532606 995143 532662 995152
rect 533712 995114 533764 995120
rect 534368 995110 534396 995452
rect 534356 995104 534408 995110
rect 534356 995046 534408 995052
rect 535564 995042 535592 995452
rect 537404 995314 537432 995452
rect 539010 995438 539258 995466
rect 538954 995415 539010 995424
rect 537392 995308 537444 995314
rect 537392 995250 537444 995256
rect 535552 995036 535604 995042
rect 535552 994978 535604 994984
rect 549180 991642 549208 1006062
rect 550270 1006023 550326 1006032
rect 551098 1006088 551100 1006097
rect 556804 1006120 556856 1006126
rect 551152 1006088 551154 1006097
rect 551098 1006023 551154 1006032
rect 553122 1006088 553178 1006097
rect 556802 1006088 556804 1006097
rect 556856 1006088 556858 1006097
rect 553122 1006023 553124 1006032
rect 553176 1006023 553178 1006032
rect 556712 1006052 556764 1006058
rect 553124 1005994 553176 1006000
rect 556802 1006023 556858 1006032
rect 563704 1006052 563756 1006058
rect 556712 1005994 556764 1006000
rect 563704 1005994 563756 1006000
rect 556344 1004760 556396 1004766
rect 556342 1004728 556344 1004737
rect 556396 1004728 556398 1004737
rect 556342 1004663 556398 1004672
rect 552754 1002688 552810 1002697
rect 552754 1002623 552756 1002632
rect 552808 1002623 552810 1002632
rect 552756 1002594 552808 1002600
rect 552296 1002584 552348 1002590
rect 552294 1002552 552296 1002561
rect 552348 1002552 552350 1002561
rect 552294 1002487 552350 1002496
rect 554778 1002144 554834 1002153
rect 553216 1002108 553268 1002114
rect 554778 1002079 554780 1002088
rect 553216 1002050 553268 1002056
rect 554832 1002079 554834 1002088
rect 554780 1002050 554832 1002056
rect 551744 1002040 551796 1002046
rect 551744 1001982 551796 1001988
rect 553122 1002008 553178 1002017
rect 550548 1001972 550600 1001978
rect 550548 1001914 550600 1001920
rect 550560 998646 550588 1001914
rect 551756 999802 551784 1001982
rect 553122 1001943 553124 1001952
rect 553176 1001943 553178 1001952
rect 553124 1001914 553176 1001920
rect 551744 999796 551796 999802
rect 551744 999738 551796 999744
rect 550548 998640 550600 998646
rect 550548 998582 550600 998588
rect 553228 997490 553256 1002050
rect 553952 1002040 554004 1002046
rect 553950 1002008 553952 1002017
rect 554004 1002008 554006 1002017
rect 553950 1001943 554006 1001952
rect 554318 1002008 554374 1002017
rect 555146 1002008 555202 1002017
rect 554318 1001943 554374 1001952
rect 554700 1001966 555146 1001994
rect 554332 997626 554360 1001943
rect 554320 997620 554372 997626
rect 554320 997562 554372 997568
rect 554700 997558 554728 1001966
rect 555146 1001943 555202 1001952
rect 556160 998640 556212 998646
rect 556160 998582 556212 998588
rect 554688 997552 554740 997558
rect 554688 997494 554740 997500
rect 553216 997484 553268 997490
rect 553216 997426 553268 997432
rect 556172 995042 556200 998582
rect 556724 997150 556752 1005994
rect 559748 1004760 559800 1004766
rect 557630 1004728 557686 1004737
rect 559748 1004702 559800 1004708
rect 557630 1004663 557632 1004672
rect 557684 1004663 557686 1004672
rect 559564 1004692 559616 1004698
rect 557632 1004634 557684 1004640
rect 559564 1004634 559616 1004640
rect 559196 1002312 559248 1002318
rect 559194 1002280 559196 1002289
rect 559248 1002280 559250 1002289
rect 559194 1002215 559250 1002224
rect 558460 1002176 558512 1002182
rect 558458 1002144 558460 1002153
rect 558512 1002144 558514 1002153
rect 558458 1002079 558514 1002088
rect 558000 1002040 558052 1002046
rect 557998 1002008 558000 1002017
rect 558052 1002008 558054 1002017
rect 557998 1001943 558054 1001952
rect 558826 1002008 558882 1002017
rect 558826 1001943 558828 1001952
rect 558880 1001943 558882 1001952
rect 558828 1001914 558880 1001920
rect 556712 997144 556764 997150
rect 556712 997086 556764 997092
rect 559576 995654 559604 1004634
rect 559654 1002280 559710 1002289
rect 559654 1002215 559656 1002224
rect 559708 1002215 559710 1002224
rect 559656 1002186 559708 1002192
rect 559760 997762 559788 1004702
rect 562324 1002312 562376 1002318
rect 562324 1002254 562376 1002260
rect 561772 1002244 561824 1002250
rect 561772 1002186 561824 1002192
rect 560944 1002176 560996 1002182
rect 560022 1002144 560078 1002153
rect 561312 1002176 561364 1002182
rect 560944 1002118 560996 1002124
rect 561310 1002144 561312 1002153
rect 561364 1002144 561366 1002153
rect 560022 1002079 560024 1002088
rect 560076 1002079 560078 1002088
rect 560024 1002050 560076 1002056
rect 560392 1002040 560444 1002046
rect 560852 1002040 560904 1002046
rect 560392 1001982 560444 1001988
rect 560482 1002008 560538 1002017
rect 560300 1001972 560352 1001978
rect 560300 1001914 560352 1001920
rect 559748 997756 559800 997762
rect 559748 997698 559800 997704
rect 560312 996062 560340 1001914
rect 560404 996198 560432 1001982
rect 560482 1001943 560484 1001952
rect 560536 1001943 560538 1001952
rect 560850 1002008 560852 1002017
rect 560904 1002008 560906 1002017
rect 560850 1001943 560906 1001952
rect 560484 1001914 560536 1001920
rect 560392 996192 560444 996198
rect 560392 996134 560444 996140
rect 560300 996056 560352 996062
rect 560300 995998 560352 996004
rect 559564 995648 559616 995654
rect 559564 995590 559616 995596
rect 556160 995036 556212 995042
rect 556160 994978 556212 994984
rect 560956 991710 560984 1002118
rect 561310 1002079 561366 1002088
rect 561496 997552 561548 997558
rect 561496 997494 561548 997500
rect 561508 996962 561536 997494
rect 561588 997484 561640 997490
rect 561588 997426 561640 997432
rect 561600 997370 561628 997426
rect 561678 997384 561734 997393
rect 561600 997342 561678 997370
rect 561678 997319 561734 997328
rect 561678 996976 561734 996985
rect 561508 996934 561678 996962
rect 561678 996911 561734 996920
rect 561784 996130 561812 1002186
rect 562232 999796 562284 999802
rect 562232 999738 562284 999744
rect 562244 997558 562272 999738
rect 562232 997552 562284 997558
rect 562232 997494 562284 997500
rect 561772 996124 561824 996130
rect 561772 996066 561824 996072
rect 560944 991704 560996 991710
rect 560944 991646 560996 991652
rect 549168 991636 549220 991642
rect 549168 991578 549220 991584
rect 562336 990146 562364 1002254
rect 562508 1002108 562560 1002114
rect 562508 1002050 562560 1002056
rect 562520 993070 562548 1002050
rect 563060 1001972 563112 1001978
rect 563060 1001914 563112 1001920
rect 563072 997694 563100 1001914
rect 563716 999802 563744 1005994
rect 563808 1000142 563836 1006266
rect 570604 1006256 570656 1006262
rect 570604 1006198 570656 1006204
rect 564346 1006088 564402 1006097
rect 564346 1006023 564402 1006032
rect 564360 1005310 564388 1006023
rect 564348 1005304 564400 1005310
rect 564348 1005246 564400 1005252
rect 565912 1002652 565964 1002658
rect 565912 1002594 565964 1002600
rect 565084 1002040 565136 1002046
rect 565084 1001982 565136 1001988
rect 563796 1000136 563848 1000142
rect 563796 1000078 563848 1000084
rect 563704 999796 563756 999802
rect 563704 999738 563756 999744
rect 563060 997688 563112 997694
rect 563060 997630 563112 997636
rect 564990 997384 565046 997393
rect 564990 997319 565046 997328
rect 565004 997286 565032 997319
rect 564992 997280 565044 997286
rect 564992 997222 565044 997228
rect 564990 996976 565046 996985
rect 564990 996911 564992 996920
rect 565044 996911 565046 996920
rect 564992 996882 565044 996888
rect 562508 993064 562560 993070
rect 562508 993006 562560 993012
rect 560116 990140 560168 990146
rect 560116 990082 560168 990088
rect 562324 990140 562376 990146
rect 562324 990082 562376 990088
rect 543832 987420 543884 987426
rect 543832 987362 543884 987368
rect 520924 985788 520976 985794
rect 520924 985730 520976 985736
rect 527640 985788 527692 985794
rect 527640 985730 527692 985736
rect 511092 983606 511474 983634
rect 527652 983620 527680 985730
rect 543844 983620 543872 987362
rect 560128 983620 560156 990082
rect 565096 987426 565124 1001982
rect 565820 1000136 565872 1000142
rect 565820 1000078 565872 1000084
rect 565832 997694 565860 1000078
rect 565924 1000074 565952 1002594
rect 568672 1002584 568724 1002590
rect 568672 1002526 568724 1002532
rect 566464 1002176 566516 1002182
rect 566464 1002118 566516 1002124
rect 565912 1000068 565964 1000074
rect 565912 1000010 565964 1000016
rect 565820 997688 565872 997694
rect 565820 997630 565872 997636
rect 566476 988786 566504 1002118
rect 568120 997280 568172 997286
rect 568118 997248 568120 997257
rect 568172 997248 568174 997257
rect 568118 997183 568174 997192
rect 568120 996940 568172 996946
rect 568120 996882 568172 996888
rect 568132 996849 568160 996882
rect 568118 996840 568174 996849
rect 568118 996775 568174 996784
rect 568684 995110 568712 1002526
rect 568764 1000068 568816 1000074
rect 568764 1000010 568816 1000016
rect 568776 997490 568804 1000010
rect 568764 997484 568816 997490
rect 568764 997426 568816 997432
rect 570616 997082 570644 1006198
rect 573364 1006120 573416 1006126
rect 573364 1006062 573416 1006068
rect 571984 1005304 572036 1005310
rect 571984 1005246 572036 1005252
rect 570604 997076 570656 997082
rect 570604 997018 570656 997024
rect 568672 995104 568724 995110
rect 568672 995046 568724 995052
rect 566464 988780 566516 988786
rect 566464 988722 566516 988728
rect 565084 987420 565136 987426
rect 565084 987362 565136 987368
rect 571996 985998 572024 1005246
rect 572720 999796 572772 999802
rect 572720 999738 572772 999744
rect 572732 997286 572760 999738
rect 573376 997422 573404 1006062
rect 573364 997416 573416 997422
rect 573364 997358 573416 997364
rect 572720 997280 572772 997286
rect 572720 997222 572772 997228
rect 574756 995246 574784 1006334
rect 612740 1000544 612792 1000550
rect 612740 1000486 612792 1000492
rect 625528 1000544 625580 1000550
rect 625528 1000486 625580 1000492
rect 575572 997824 575624 997830
rect 575572 997766 575624 997772
rect 607128 997824 607180 997830
rect 607128 997766 607180 997772
rect 575584 997506 575612 997766
rect 607140 997626 607168 997766
rect 607128 997620 607180 997626
rect 607128 997562 607180 997568
rect 575584 997478 575704 997506
rect 575202 997248 575258 997257
rect 575202 997183 575204 997192
rect 575256 997183 575258 997192
rect 575204 997154 575256 997160
rect 575480 996872 575532 996878
rect 575478 996840 575480 996849
rect 575532 996840 575534 996849
rect 575478 996775 575534 996784
rect 574744 995240 574796 995246
rect 574744 995182 574796 995188
rect 575676 992234 575704 997478
rect 612752 997422 612780 1000486
rect 618168 999184 618220 999190
rect 618168 999126 618220 999132
rect 625436 999184 625488 999190
rect 625436 999126 625488 999132
rect 614120 998028 614172 998034
rect 614120 997970 614172 997976
rect 614132 997558 614160 997970
rect 614120 997552 614172 997558
rect 614120 997494 614172 997500
rect 618180 997490 618208 999126
rect 623688 997688 623740 997694
rect 623688 997630 623740 997636
rect 618168 997484 618220 997490
rect 618168 997426 618220 997432
rect 612740 997416 612792 997422
rect 612740 997358 612792 997364
rect 585140 997280 585192 997286
rect 580906 997248 580962 997257
rect 580906 997183 580908 997192
rect 580960 997183 580962 997192
rect 585138 997248 585140 997257
rect 590936 997280 590988 997286
rect 585192 997248 585194 997257
rect 585138 997183 585194 997192
rect 590934 997248 590936 997257
rect 590988 997248 590990 997257
rect 590934 997183 590990 997192
rect 620284 997212 620336 997218
rect 580908 997154 580960 997160
rect 620284 997154 620336 997160
rect 605932 997144 605984 997150
rect 605932 997086 605984 997092
rect 580724 996872 580776 996878
rect 580722 996840 580724 996849
rect 585508 996872 585560 996878
rect 580776 996840 580778 996849
rect 580722 996775 580778 996784
rect 585506 996840 585508 996849
rect 590568 996872 590620 996878
rect 585560 996840 585562 996849
rect 585506 996775 585562 996784
rect 590566 996840 590568 996849
rect 590620 996840 590622 996849
rect 590566 996775 590622 996784
rect 605944 996305 605972 997086
rect 605930 996296 605986 996305
rect 605930 996231 605986 996240
rect 620296 995178 620324 997154
rect 622400 997076 622452 997082
rect 622400 997018 622452 997024
rect 620284 995172 620336 995178
rect 620284 995114 620336 995120
rect 622412 995081 622440 997018
rect 623700 996713 623728 997630
rect 623686 996704 623742 996713
rect 623686 996639 623742 996648
rect 625448 995994 625476 999126
rect 625436 995988 625488 995994
rect 625436 995930 625488 995936
rect 625540 995586 625568 1000486
rect 625620 998028 625672 998034
rect 625620 997970 625672 997976
rect 625632 995722 625660 997970
rect 625712 997960 625764 997966
rect 625712 997902 625764 997908
rect 625724 995790 625752 997902
rect 625804 997824 625856 997830
rect 625804 997766 625856 997772
rect 625816 995858 625844 997766
rect 625894 996704 625950 996713
rect 625894 996639 625950 996648
rect 625908 995926 625936 996639
rect 625896 995920 625948 995926
rect 625896 995862 625948 995868
rect 625804 995852 625856 995858
rect 625804 995794 625856 995800
rect 626540 995852 626592 995858
rect 626540 995794 626592 995800
rect 630864 995852 630916 995858
rect 630864 995794 630916 995800
rect 631508 995852 631560 995858
rect 631508 995794 631560 995800
rect 625712 995784 625764 995790
rect 625712 995726 625764 995732
rect 626552 995738 626580 995794
rect 627184 995784 627236 995790
rect 625620 995716 625672 995722
rect 626552 995710 626888 995738
rect 630876 995738 630904 995794
rect 631520 995738 631548 995794
rect 633990 995752 634046 995761
rect 627236 995732 627532 995738
rect 627184 995726 627532 995732
rect 627196 995710 627532 995726
rect 630232 995722 630568 995738
rect 630220 995716 630568 995722
rect 625620 995658 625672 995664
rect 630272 995710 630568 995716
rect 630876 995710 631212 995738
rect 631520 995710 631856 995738
rect 640798 995752 640854 995761
rect 634046 995710 634340 995738
rect 633990 995687 634046 995696
rect 640854 995710 641056 995738
rect 640798 995687 640854 995696
rect 630220 995658 630272 995664
rect 661684 995648 661736 995654
rect 635186 995616 635242 995625
rect 627932 995586 628176 995602
rect 625528 995580 625580 995586
rect 625528 995522 625580 995528
rect 627920 995580 628176 995586
rect 627972 995574 628176 995580
rect 635242 995574 635536 995602
rect 661684 995590 661736 995596
rect 635186 995551 635242 995560
rect 627920 995522 627972 995528
rect 629680 995438 630016 995466
rect 634832 995438 634892 995466
rect 629680 995081 629708 995438
rect 634832 995110 634860 995438
rect 636166 995246 636194 995452
rect 637040 995438 637376 995466
rect 638572 995438 638908 995466
rect 636154 995240 636206 995246
rect 636154 995182 636206 995188
rect 634820 995104 634872 995110
rect 622398 995072 622454 995081
rect 622398 995007 622454 995016
rect 629666 995072 629722 995081
rect 634820 995046 634872 995052
rect 637040 995042 637068 995438
rect 638880 995058 638908 995438
rect 638972 995438 639216 995466
rect 638972 995178 639000 995438
rect 638960 995172 639012 995178
rect 638960 995114 639012 995120
rect 629666 995007 629722 995016
rect 637028 995036 637080 995042
rect 638880 995030 639000 995058
rect 637028 994978 637080 994984
rect 638972 994945 639000 995030
rect 638958 994936 639014 994945
rect 638958 994871 639014 994880
rect 640798 994936 640854 994945
rect 640798 994871 640854 994880
rect 575676 992206 575888 992234
rect 571984 985992 572036 985998
rect 571984 985934 572036 985940
rect 575860 983634 575888 992206
rect 592500 988780 592552 988786
rect 592500 988722 592552 988728
rect 575860 983606 576334 983634
rect 592512 983620 592540 988722
rect 624976 987420 625028 987426
rect 624976 987362 625028 987368
rect 608784 985992 608836 985998
rect 608784 985934 608836 985940
rect 608796 983620 608824 985934
rect 624988 983620 625016 987362
rect 640812 983634 640840 994871
rect 660304 993064 660356 993070
rect 660304 993006 660356 993012
rect 658924 991704 658976 991710
rect 658924 991646 658976 991652
rect 650000 984836 650052 984842
rect 650000 984778 650052 984784
rect 640812 983606 641194 983634
rect 62118 976032 62174 976041
rect 62118 975967 62174 975976
rect 62132 975730 62160 975967
rect 62120 975724 62172 975730
rect 62120 975666 62172 975672
rect 62118 962976 62174 962985
rect 62118 962911 62174 962920
rect 62132 961926 62160 962911
rect 62120 961920 62172 961926
rect 62120 961862 62172 961868
rect 62118 949920 62174 949929
rect 62118 949855 62174 949864
rect 62132 947374 62160 949855
rect 62120 947368 62172 947374
rect 62120 947310 62172 947316
rect 55862 939856 55918 939865
rect 55862 939791 55918 939800
rect 45744 937032 45796 937038
rect 62120 937032 62172 937038
rect 45744 936974 45796 936980
rect 62118 937000 62120 937009
rect 62172 937000 62174 937009
rect 62118 936935 62174 936944
rect 44178 934552 44234 934561
rect 44178 934487 44234 934496
rect 42890 934144 42946 934153
rect 42890 934079 42946 934088
rect 42798 933736 42854 933745
rect 42798 933671 42854 933680
rect 47584 932204 47636 932210
rect 47584 932146 47636 932152
rect 44824 870868 44876 870874
rect 44824 870810 44876 870816
rect 43628 858424 43680 858430
rect 43628 858366 43680 858372
rect 41892 823846 42012 823874
rect 41800 819182 41920 819210
rect 41708 816734 41828 816762
rect 41694 816640 41750 816649
rect 41524 816598 41694 816626
rect 41694 816575 41750 816584
rect 41800 814065 41828 816734
rect 41892 815697 41920 819182
rect 41878 815688 41934 815697
rect 41878 815623 41934 815632
rect 41984 814881 42012 823846
rect 43536 818372 43588 818378
rect 43536 818314 43588 818320
rect 41970 814872 42026 814881
rect 41970 814807 42026 814816
rect 41786 814056 41842 814065
rect 41786 813991 41842 814000
rect 40682 813240 40738 813249
rect 40682 813175 40738 813184
rect 33782 812424 33838 812433
rect 33782 812359 33838 812368
rect 33046 810384 33102 810393
rect 33046 810319 33102 810328
rect 32402 809160 32458 809169
rect 32402 809095 32458 809104
rect 32416 801106 32444 809095
rect 33060 802505 33088 810319
rect 33046 802496 33102 802505
rect 33046 802431 33102 802440
rect 32404 801100 32456 801106
rect 32404 801042 32456 801048
rect 33796 801009 33824 812359
rect 34426 810792 34482 810801
rect 34426 810727 34482 810736
rect 34440 802641 34468 810727
rect 35162 808752 35218 808761
rect 35162 808687 35218 808696
rect 34426 802632 34482 802641
rect 34426 802567 34482 802576
rect 35176 801174 35204 808687
rect 39854 807328 39910 807337
rect 39854 807263 39856 807272
rect 39908 807263 39910 807272
rect 39856 807230 39908 807236
rect 40696 801689 40724 813175
rect 42154 812832 42210 812841
rect 42154 812767 42210 812776
rect 41786 811608 41842 811617
rect 40776 811572 40828 811578
rect 41786 811543 41788 811552
rect 40776 811514 40828 811520
rect 41840 811543 41842 811552
rect 41788 811514 41840 811520
rect 40682 801680 40738 801689
rect 40682 801615 40738 801624
rect 35164 801168 35216 801174
rect 35164 801110 35216 801116
rect 33782 801000 33838 801009
rect 33782 800935 33838 800944
rect 40788 800562 40816 811514
rect 42062 809568 42118 809577
rect 42062 809503 42118 809512
rect 41788 807288 41840 807294
rect 41788 807230 41840 807236
rect 41800 806313 41828 807230
rect 41786 806304 41842 806313
rect 41786 806239 41842 806248
rect 42076 803826 42104 809503
rect 42168 803894 42196 812767
rect 42338 811200 42394 811209
rect 42338 811135 42394 811144
rect 42156 803888 42208 803894
rect 42156 803830 42208 803836
rect 42064 803820 42116 803826
rect 42064 803762 42116 803768
rect 40776 800556 40828 800562
rect 40776 800498 40828 800504
rect 42352 800018 42380 811135
rect 42798 809976 42854 809985
rect 42798 809911 42854 809920
rect 42616 803888 42668 803894
rect 42616 803830 42668 803836
rect 42156 800012 42208 800018
rect 42156 799954 42208 799960
rect 42340 800012 42392 800018
rect 42340 799954 42392 799960
rect 42168 799445 42196 799954
rect 42628 798182 42656 803830
rect 42708 803820 42760 803826
rect 42708 803762 42760 803768
rect 42156 798176 42208 798182
rect 42156 798118 42208 798124
rect 42616 798176 42668 798182
rect 42616 798118 42668 798124
rect 42168 797605 42196 798118
rect 42156 797292 42208 797298
rect 42156 797234 42208 797240
rect 42168 796960 42196 797234
rect 42430 796784 42486 796793
rect 42430 796719 42486 796728
rect 42156 796340 42208 796346
rect 42156 796282 42208 796288
rect 42168 795765 42196 796282
rect 42444 795054 42472 796719
rect 42720 796346 42748 803762
rect 42708 796340 42760 796346
rect 42708 796282 42760 796288
rect 42708 796204 42760 796210
rect 42708 796146 42760 796152
rect 42156 795048 42208 795054
rect 42156 794990 42208 794996
rect 42432 795048 42484 795054
rect 42432 794990 42484 794996
rect 42168 794580 42196 794990
rect 42432 794912 42484 794918
rect 42432 794854 42484 794860
rect 42156 794300 42208 794306
rect 42156 794242 42208 794248
rect 42168 793900 42196 794242
rect 42156 793824 42208 793830
rect 42156 793766 42208 793772
rect 42168 793288 42196 793766
rect 42444 793218 42472 794854
rect 42720 794306 42748 796146
rect 42708 794300 42760 794306
rect 42708 794242 42760 794248
rect 42708 794164 42760 794170
rect 42708 794106 42760 794112
rect 42156 793212 42208 793218
rect 42156 793154 42208 793160
rect 42432 793212 42484 793218
rect 42432 793154 42484 793160
rect 42168 792744 42196 793154
rect 42432 793076 42484 793082
rect 42432 793018 42484 793024
rect 42338 792024 42394 792033
rect 42338 791959 42394 791968
rect 42156 790696 42208 790702
rect 42156 790638 42208 790644
rect 42168 790228 42196 790638
rect 42156 790152 42208 790158
rect 42156 790094 42208 790100
rect 42168 789616 42196 790094
rect 42352 789478 42380 791959
rect 42444 790158 42472 793018
rect 42720 792010 42748 794106
rect 42812 793082 42840 809911
rect 43442 806304 43498 806313
rect 43442 806239 43498 806248
rect 43076 801168 43128 801174
rect 43076 801110 43128 801116
rect 42892 801100 42944 801106
rect 42892 801042 42944 801048
rect 42904 796210 42932 801042
rect 42984 800556 43036 800562
rect 42984 800498 43036 800504
rect 42892 796204 42944 796210
rect 42892 796146 42944 796152
rect 42892 794980 42944 794986
rect 42892 794922 42944 794928
rect 42904 793830 42932 794922
rect 42996 794918 43024 800498
rect 42984 794912 43036 794918
rect 42984 794854 43036 794860
rect 43088 794170 43116 801110
rect 43168 799060 43220 799066
rect 43168 799002 43220 799008
rect 43180 797298 43208 799002
rect 43168 797292 43220 797298
rect 43168 797234 43220 797240
rect 43076 794164 43128 794170
rect 43076 794106 43128 794112
rect 42892 793824 42944 793830
rect 42892 793766 42944 793772
rect 42800 793076 42852 793082
rect 42800 793018 42852 793024
rect 42720 791982 42840 792010
rect 42706 791888 42762 791897
rect 42706 791823 42762 791832
rect 42432 790152 42484 790158
rect 42432 790094 42484 790100
rect 42156 789472 42208 789478
rect 42156 789414 42208 789420
rect 42340 789472 42392 789478
rect 42340 789414 42392 789420
rect 42168 788936 42196 789414
rect 42720 788866 42748 791823
rect 42812 790702 42840 791982
rect 42800 790696 42852 790702
rect 42800 790638 42852 790644
rect 42156 788860 42208 788866
rect 42156 788802 42208 788808
rect 42708 788860 42760 788866
rect 42708 788802 42760 788808
rect 42168 788392 42196 788802
rect 42706 788216 42762 788225
rect 42706 788151 42762 788160
rect 42430 788080 42486 788089
rect 42430 788015 42486 788024
rect 42444 787030 42472 788015
rect 42156 787024 42208 787030
rect 42156 786966 42208 786972
rect 42432 787024 42484 787030
rect 42432 786966 42484 786972
rect 42168 786556 42196 786966
rect 41786 786176 41842 786185
rect 41786 786111 41842 786120
rect 41800 785944 41828 786111
rect 42720 785670 42748 788151
rect 42156 785664 42208 785670
rect 42156 785606 42208 785612
rect 42708 785664 42760 785670
rect 42708 785606 42760 785612
rect 42168 785264 42196 785606
rect 8588 775132 8616 775268
rect 9048 775132 9076 775268
rect 9508 775132 9536 775268
rect 9968 775132 9996 775268
rect 10428 775132 10456 775268
rect 10888 775132 10916 775268
rect 11348 775132 11376 775268
rect 11808 775132 11836 775268
rect 12268 775132 12296 775268
rect 12728 775132 12756 775268
rect 13188 775132 13216 775268
rect 13648 775132 13676 775268
rect 14108 775132 14136 775268
rect 35806 774344 35862 774353
rect 35806 774279 35862 774288
rect 35820 774246 35848 774279
rect 35808 774240 35860 774246
rect 35808 774182 35860 774188
rect 42798 772032 42854 772041
rect 42798 771967 42854 771976
rect 33782 769448 33838 769457
rect 33782 769383 33838 769392
rect 32402 768632 32458 768641
rect 32402 768567 32458 768576
rect 31022 767816 31078 767825
rect 31022 767751 31078 767760
rect 30378 764144 30434 764153
rect 30378 764079 30434 764088
rect 30392 763337 30420 764079
rect 30378 763328 30434 763337
rect 30378 763263 30434 763272
rect 31036 759694 31064 767751
rect 31024 759688 31076 759694
rect 31024 759630 31076 759636
rect 32416 758334 32444 768567
rect 32494 766592 32550 766601
rect 32494 766527 32550 766536
rect 32508 758402 32536 766527
rect 33796 758538 33824 769383
rect 40682 769040 40738 769049
rect 40682 768975 40738 768984
rect 35162 767408 35218 767417
rect 35162 767343 35218 767352
rect 33784 758532 33836 758538
rect 33784 758474 33836 758480
rect 32496 758396 32548 758402
rect 32496 758338 32548 758344
rect 32404 758328 32456 758334
rect 35176 758305 35204 767343
rect 32404 758270 32456 758276
rect 35162 758296 35218 758305
rect 35162 758231 35218 758240
rect 40696 757761 40724 768975
rect 41510 762920 41566 762929
rect 41510 762855 41566 762864
rect 41524 761802 41552 762855
rect 41512 761796 41564 761802
rect 41512 761738 41564 761744
rect 41880 759688 41932 759694
rect 41880 759630 41932 759636
rect 40682 757752 40738 757761
rect 40682 757687 40738 757696
rect 41892 757042 41920 759630
rect 42432 758532 42484 758538
rect 42432 758474 42484 758480
rect 41880 757036 41932 757042
rect 41880 756978 41932 756984
rect 41880 756764 41932 756770
rect 41880 756706 41932 756712
rect 41892 756226 41920 756706
rect 42444 755546 42472 758474
rect 42708 758396 42760 758402
rect 42708 758338 42760 758344
rect 42720 756537 42748 758338
rect 42706 756528 42762 756537
rect 42706 756463 42762 756472
rect 42432 755540 42484 755546
rect 42432 755482 42484 755488
rect 42156 755472 42208 755478
rect 42156 755414 42208 755420
rect 42168 755206 42196 755414
rect 42616 755268 42668 755274
rect 42616 755210 42668 755216
rect 42156 755200 42208 755206
rect 42156 755142 42208 755148
rect 42156 754928 42208 754934
rect 42156 754870 42208 754876
rect 42168 754392 42196 754870
rect 42064 754112 42116 754118
rect 42064 754054 42116 754060
rect 42076 753780 42104 754054
rect 41786 753128 41842 753137
rect 41786 753063 41842 753072
rect 41800 752556 41828 753063
rect 41786 751768 41842 751777
rect 41786 751703 41842 751712
rect 41800 751369 41828 751703
rect 42156 751120 42208 751126
rect 42156 751062 42208 751068
rect 42168 750720 42196 751062
rect 41786 750408 41842 750417
rect 41786 750343 41842 750352
rect 41800 750108 41828 750343
rect 42156 749828 42208 749834
rect 42156 749770 42208 749776
rect 42168 749529 42196 749770
rect 42076 746978 42104 747048
rect 42064 746972 42116 746978
rect 42064 746914 42116 746920
rect 42156 746972 42208 746978
rect 42156 746914 42208 746920
rect 42168 746401 42196 746914
rect 42628 746706 42656 755210
rect 42706 749320 42762 749329
rect 42706 749255 42762 749264
rect 42720 746978 42748 749255
rect 42708 746972 42760 746978
rect 42708 746914 42760 746920
rect 42708 746836 42760 746842
rect 42708 746778 42760 746784
rect 42616 746700 42668 746706
rect 42616 746642 42668 746648
rect 42614 746600 42670 746609
rect 42614 746535 42670 746544
rect 42156 746088 42208 746094
rect 42156 746030 42208 746036
rect 42168 745756 42196 746030
rect 42156 745476 42208 745482
rect 42156 745418 42208 745424
rect 42168 745212 42196 745418
rect 42156 743776 42208 743782
rect 42156 743718 42208 743724
rect 42168 743376 42196 743718
rect 42628 743306 42656 746535
rect 42720 746094 42748 746778
rect 42708 746088 42760 746094
rect 42708 746030 42760 746036
rect 42708 745952 42760 745958
rect 42708 745894 42760 745900
rect 42720 743782 42748 745894
rect 42708 743776 42760 743782
rect 42708 743718 42760 743724
rect 42156 743300 42208 743306
rect 42156 743242 42208 743248
rect 42616 743300 42668 743306
rect 42616 743242 42668 743248
rect 42168 742696 42196 743242
rect 41786 742384 41842 742393
rect 41786 742319 41842 742328
rect 41800 742084 41828 742319
rect 8588 731884 8616 732020
rect 9048 731884 9076 732020
rect 9508 731884 9536 732020
rect 9968 731884 9996 732020
rect 10428 731884 10456 732020
rect 10888 731884 10916 732020
rect 11348 731884 11376 732020
rect 11808 731884 11836 732020
rect 12268 731884 12296 732020
rect 12728 731884 12756 732020
rect 13188 731884 13216 732020
rect 13648 731884 13676 732020
rect 14108 731884 14136 732020
rect 31392 731400 31444 731406
rect 31392 731342 31444 731348
rect 31404 730289 31432 731342
rect 31576 731332 31628 731338
rect 31576 731274 31628 731280
rect 31482 731096 31538 731105
rect 31482 731031 31484 731040
rect 31536 731031 31538 731040
rect 31484 731002 31536 731008
rect 31588 730697 31616 731274
rect 31668 731196 31720 731202
rect 31668 731138 31720 731144
rect 31680 731105 31708 731138
rect 31666 731096 31722 731105
rect 31666 731031 31722 731040
rect 31574 730688 31630 730697
rect 31574 730623 31630 730632
rect 31390 730280 31446 730289
rect 31390 730215 31446 730224
rect 42812 729337 42840 771967
rect 42890 767136 42946 767145
rect 42890 767071 42946 767080
rect 42904 746842 42932 767071
rect 42982 765912 43038 765921
rect 42982 765847 43038 765856
rect 42996 751126 43024 765847
rect 43168 758328 43220 758334
rect 43168 758270 43220 758276
rect 43180 755274 43208 758270
rect 43260 756288 43312 756294
rect 43260 756230 43312 756236
rect 43168 755268 43220 755274
rect 43168 755210 43220 755216
rect 43272 754118 43300 756230
rect 43260 754112 43312 754118
rect 43260 754054 43312 754060
rect 43076 752140 43128 752146
rect 43076 752082 43128 752088
rect 42984 751120 43036 751126
rect 42984 751062 43036 751068
rect 43088 749834 43116 752082
rect 43076 749828 43128 749834
rect 43076 749770 43128 749776
rect 42984 749420 43036 749426
rect 42984 749362 43036 749368
rect 42996 747046 43024 749362
rect 42984 747040 43036 747046
rect 42984 746982 43036 746988
rect 42892 746836 42944 746842
rect 42892 746778 42944 746784
rect 43076 746700 43128 746706
rect 43076 746642 43128 746648
rect 43088 745482 43116 746642
rect 43076 745476 43128 745482
rect 43076 745418 43128 745424
rect 42798 729328 42854 729337
rect 42798 729263 42854 729272
rect 42798 727288 42854 727297
rect 42798 727223 42854 727232
rect 31022 726608 31078 726617
rect 31022 726543 31078 726552
rect 31036 715465 31064 726543
rect 40682 726200 40738 726209
rect 40682 726135 40738 726144
rect 33782 725384 33838 725393
rect 33782 725319 33838 725328
rect 33796 715601 33824 725319
rect 34426 723344 34482 723353
rect 34426 723279 34482 723288
rect 33782 715592 33838 715601
rect 34440 715562 34468 723279
rect 33782 715527 33838 715536
rect 34428 715556 34480 715562
rect 34428 715498 34480 715504
rect 31022 715456 31078 715465
rect 31022 715391 31078 715400
rect 40696 714814 40724 726135
rect 42154 725248 42210 725257
rect 42154 725183 42210 725192
rect 40866 724568 40922 724577
rect 40866 724503 40922 724512
rect 40774 723344 40830 723353
rect 40774 723279 40830 723288
rect 40684 714808 40736 714814
rect 40684 714750 40736 714756
rect 40788 714105 40816 723279
rect 40880 716242 40908 724503
rect 42062 724024 42118 724033
rect 42062 723959 42118 723968
rect 41510 720896 41566 720905
rect 41510 720831 41566 720840
rect 41524 719710 41552 720831
rect 41512 719704 41564 719710
rect 41510 719672 41512 719681
rect 41564 719672 41566 719681
rect 41510 719607 41566 719616
rect 40868 716236 40920 716242
rect 40868 716178 40920 716184
rect 41880 716236 41932 716242
rect 41880 716178 41932 716184
rect 40774 714096 40830 714105
rect 40774 714031 40830 714040
rect 41892 713862 41920 716178
rect 41880 713856 41932 713862
rect 42076 713833 42104 723959
rect 42168 716922 42196 725183
rect 42156 716916 42208 716922
rect 42156 716858 42208 716864
rect 42524 716916 42576 716922
rect 42524 716858 42576 716864
rect 42156 715556 42208 715562
rect 42156 715498 42208 715504
rect 42168 713862 42196 715498
rect 42432 714808 42484 714814
rect 42432 714750 42484 714756
rect 42156 713856 42208 713862
rect 41880 713798 41932 713804
rect 42062 713824 42118 713833
rect 42156 713798 42208 713804
rect 42062 713759 42118 713768
rect 41880 713584 41932 713590
rect 41880 713526 41932 713532
rect 41892 713048 41920 713526
rect 42444 713289 42472 714750
rect 42430 713280 42486 713289
rect 42430 713215 42486 713224
rect 42536 712337 42564 716858
rect 42522 712328 42578 712337
rect 42522 712263 42578 712272
rect 42524 712156 42576 712162
rect 42524 712098 42576 712104
rect 42154 711784 42210 711793
rect 42154 711719 42210 711728
rect 42168 711212 42196 711719
rect 42536 711006 42564 712098
rect 42524 711000 42576 711006
rect 42524 710942 42576 710948
rect 42156 710932 42208 710938
rect 42156 710874 42208 710880
rect 42168 710561 42196 710874
rect 42522 710832 42578 710841
rect 42522 710767 42578 710776
rect 41786 709880 41842 709889
rect 41786 709815 41842 709824
rect 41800 709376 41828 709815
rect 42536 708626 42564 710767
rect 42156 708620 42208 708626
rect 42156 708562 42208 708568
rect 42524 708620 42576 708626
rect 42524 708562 42576 708568
rect 42168 708152 42196 708562
rect 42522 708520 42578 708529
rect 42522 708455 42578 708464
rect 42156 708076 42208 708082
rect 42156 708018 42208 708024
rect 42168 707540 42196 708018
rect 42156 707260 42208 707266
rect 42156 707202 42208 707208
rect 42168 706860 42196 707202
rect 42536 706790 42564 708455
rect 42156 706784 42208 706790
rect 42156 706726 42208 706732
rect 42524 706784 42576 706790
rect 42524 706726 42576 706732
rect 42168 706316 42196 706726
rect 42522 706616 42578 706625
rect 42522 706551 42578 706560
rect 42536 706058 42564 706551
rect 42444 706030 42564 706058
rect 42246 704984 42302 704993
rect 42246 704919 42302 704928
rect 42064 704268 42116 704274
rect 42064 704210 42116 704216
rect 42076 703868 42104 704210
rect 42156 703588 42208 703594
rect 42156 703530 42208 703536
rect 42168 703188 42196 703530
rect 42064 702908 42116 702914
rect 42064 702850 42116 702856
rect 42076 702576 42104 702850
rect 42260 702574 42288 704919
rect 42444 703050 42472 706030
rect 42432 703044 42484 703050
rect 42432 702986 42484 702992
rect 42430 702944 42486 702953
rect 42430 702879 42486 702888
rect 42248 702568 42300 702574
rect 42248 702510 42300 702516
rect 42064 702296 42116 702302
rect 42064 702238 42116 702244
rect 42076 702032 42104 702238
rect 42444 700466 42472 702879
rect 42156 700460 42208 700466
rect 42156 700402 42208 700408
rect 42432 700460 42484 700466
rect 42432 700402 42484 700408
rect 42168 700165 42196 700402
rect 42156 699916 42208 699922
rect 42156 699858 42208 699864
rect 42168 699516 42196 699858
rect 41786 699408 41842 699417
rect 41786 699343 41842 699352
rect 41800 698904 41828 699343
rect 35716 692096 35768 692102
rect 35716 692038 35768 692044
rect 8588 688772 8616 688908
rect 9048 688772 9076 688908
rect 9508 688772 9536 688908
rect 9968 688772 9996 688908
rect 10428 688772 10456 688908
rect 10888 688772 10916 688908
rect 11348 688772 11376 688908
rect 11808 688772 11836 688908
rect 12268 688772 12296 688908
rect 12728 688772 12756 688908
rect 13188 688772 13216 688908
rect 13648 688772 13676 688908
rect 14108 688772 14136 688908
rect 35622 688392 35678 688401
rect 35622 688327 35678 688336
rect 35636 687818 35664 688327
rect 35624 687812 35676 687818
rect 35624 687754 35676 687760
rect 35728 687313 35756 692038
rect 35808 687948 35860 687954
rect 35808 687890 35860 687896
rect 35820 687721 35848 687890
rect 35806 687712 35862 687721
rect 35806 687647 35862 687656
rect 35714 687304 35770 687313
rect 35714 687239 35770 687248
rect 42812 684457 42840 727223
rect 42890 724432 42946 724441
rect 42890 724367 42946 724376
rect 42904 699922 42932 724367
rect 42982 722392 43038 722401
rect 42982 722327 43038 722336
rect 42996 712094 43024 722327
rect 42996 712066 43116 712094
rect 42984 711000 43036 711006
rect 42984 710942 43036 710948
rect 42996 703594 43024 710942
rect 43088 704274 43116 712066
rect 43168 709368 43220 709374
rect 43168 709310 43220 709316
rect 43180 708082 43208 709310
rect 43168 708076 43220 708082
rect 43168 708018 43220 708024
rect 43076 704268 43128 704274
rect 43076 704210 43128 704216
rect 42984 703588 43036 703594
rect 42984 703530 43036 703536
rect 42892 699916 42944 699922
rect 42892 699858 42944 699864
rect 42798 684448 42854 684457
rect 42798 684383 42854 684392
rect 42798 684040 42854 684049
rect 42798 683975 42854 683984
rect 39302 683632 39358 683641
rect 39302 683567 39358 683576
rect 32402 682816 32458 682825
rect 32402 682751 32458 682760
rect 31022 681592 31078 681601
rect 31022 681527 31078 681536
rect 30470 676866 30526 676875
rect 30470 676801 30526 676810
rect 31036 672790 31064 681527
rect 31024 672784 31076 672790
rect 31024 672726 31076 672732
rect 32416 671401 32444 682751
rect 35162 680368 35218 680377
rect 35162 680303 35218 680312
rect 35176 672858 35204 680303
rect 35164 672852 35216 672858
rect 35164 672794 35216 672800
rect 32402 671392 32458 671401
rect 32402 671327 32458 671336
rect 39316 670993 39344 683567
rect 41694 683088 41750 683097
rect 40684 683052 40736 683058
rect 41694 683023 41696 683032
rect 40684 682994 40736 683000
rect 41748 683023 41750 683032
rect 41696 682994 41748 683000
rect 39302 670984 39358 670993
rect 40696 670954 40724 682994
rect 41694 681864 41750 681873
rect 40776 681828 40828 681834
rect 41694 681799 41696 681808
rect 40776 681770 40828 681776
rect 41748 681799 41750 681808
rect 41696 681770 41748 681776
rect 40788 671022 40816 681770
rect 41970 680776 42026 680785
rect 41970 680711 42026 680720
rect 41880 672784 41932 672790
rect 41880 672726 41932 672732
rect 40776 671016 40828 671022
rect 40776 670958 40828 670964
rect 39302 670919 39358 670928
rect 40684 670948 40736 670954
rect 40684 670890 40736 670896
rect 41892 670614 41920 672726
rect 41984 670614 42012 680711
rect 42432 672852 42484 672858
rect 42432 672794 42484 672800
rect 42064 671016 42116 671022
rect 42064 670958 42116 670964
rect 42076 670721 42104 670958
rect 42062 670712 42118 670721
rect 42062 670647 42118 670656
rect 41880 670608 41932 670614
rect 41880 670550 41932 670556
rect 41972 670608 42024 670614
rect 41972 670550 42024 670556
rect 41880 670404 41932 670410
rect 41880 670346 41932 670352
rect 41892 669868 41920 670346
rect 42444 670177 42472 672794
rect 42708 670948 42760 670954
rect 42708 670890 42760 670896
rect 42430 670168 42486 670177
rect 42430 670103 42486 670112
rect 42720 669497 42748 670890
rect 42706 669488 42762 669497
rect 42706 669423 42762 669432
rect 42708 669384 42760 669390
rect 42708 669326 42760 669332
rect 42062 668536 42118 668545
rect 42062 668471 42118 668480
rect 42076 668032 42104 668471
rect 42720 667894 42748 669326
rect 42156 667888 42208 667894
rect 42156 667830 42208 667836
rect 42708 667888 42760 667894
rect 42708 667830 42760 667836
rect 42168 667352 42196 667830
rect 42708 667752 42760 667758
rect 42708 667694 42760 667700
rect 42720 666738 42748 667694
rect 42156 666732 42208 666738
rect 42156 666674 42208 666680
rect 42708 666732 42760 666738
rect 42708 666674 42760 666680
rect 42168 666165 42196 666674
rect 42708 666528 42760 666534
rect 42708 666470 42760 666476
rect 41786 665408 41842 665417
rect 41786 665343 41842 665352
rect 41800 664972 41828 665343
rect 41786 664592 41842 664601
rect 41786 664527 41842 664536
rect 41800 664325 41828 664527
rect 42720 664222 42748 666470
rect 42156 664216 42208 664222
rect 42156 664158 42208 664164
rect 42708 664216 42760 664222
rect 42708 664158 42760 664164
rect 42168 663680 42196 664158
rect 42062 663368 42118 663377
rect 42062 663303 42118 663312
rect 42076 663136 42104 663303
rect 42706 661328 42762 661337
rect 42706 661263 42762 661272
rect 42156 661088 42208 661094
rect 42156 661030 42208 661036
rect 42168 660620 42196 661030
rect 42154 660512 42210 660521
rect 42154 660447 42210 660456
rect 42168 660008 42196 660447
rect 42522 660376 42578 660385
rect 42522 660311 42578 660320
rect 42156 659728 42208 659734
rect 42156 659670 42208 659676
rect 42168 659357 42196 659670
rect 42156 659048 42208 659054
rect 42156 658990 42208 658996
rect 42168 658784 42196 658990
rect 42338 658336 42394 658345
rect 42338 658271 42394 658280
rect 42156 657280 42208 657286
rect 42156 657222 42208 657228
rect 42168 656948 42196 657222
rect 42156 656872 42208 656878
rect 42156 656814 42208 656820
rect 42168 656336 42196 656814
rect 42352 656198 42380 658271
rect 42536 657286 42564 660311
rect 42720 659054 42748 661263
rect 42708 659048 42760 659054
rect 42708 658990 42760 658996
rect 42524 657280 42576 657286
rect 42524 657222 42576 657228
rect 42156 656192 42208 656198
rect 42156 656134 42208 656140
rect 42340 656192 42392 656198
rect 42340 656134 42392 656140
rect 42168 655656 42196 656134
rect 8588 645524 8616 645660
rect 9048 645524 9076 645660
rect 9508 645524 9536 645660
rect 9968 645524 9996 645660
rect 10428 645524 10456 645660
rect 10888 645524 10916 645660
rect 11348 645524 11376 645660
rect 11808 645524 11836 645660
rect 12268 645524 12296 645660
rect 12728 645524 12756 645660
rect 13188 645524 13216 645660
rect 13648 645524 13676 645660
rect 14108 645524 14136 645660
rect 35622 644736 35678 644745
rect 35622 644671 35678 644680
rect 35806 644736 35862 644745
rect 35806 644671 35862 644680
rect 35636 644570 35664 644671
rect 35820 644638 35848 644671
rect 35808 644632 35860 644638
rect 35808 644574 35860 644580
rect 35624 644564 35676 644570
rect 35624 644506 35676 644512
rect 42812 641481 42840 683975
rect 42890 679144 42946 679153
rect 42890 679079 42946 679088
rect 42904 668658 42932 679079
rect 42982 678736 43038 678745
rect 42982 678671 43038 678680
rect 42996 673454 43024 678671
rect 42996 673426 43116 673454
rect 42984 670608 43036 670614
rect 42984 670550 43036 670556
rect 42996 668778 43024 670550
rect 42984 668772 43036 668778
rect 42984 668714 43036 668720
rect 42904 668630 43024 668658
rect 42892 668568 42944 668574
rect 42892 668510 42944 668516
rect 42904 659734 42932 668510
rect 42996 663794 43024 668630
rect 43088 666534 43116 673426
rect 43076 666528 43128 666534
rect 43076 666470 43128 666476
rect 42996 663766 43116 663794
rect 43088 661094 43116 663766
rect 43076 661088 43128 661094
rect 43076 661030 43128 661036
rect 42892 659728 42944 659734
rect 42892 659670 42944 659676
rect 42892 658300 42944 658306
rect 42892 658242 42944 658248
rect 42904 656878 42932 658242
rect 42892 656872 42944 656878
rect 42892 656814 42944 656820
rect 42798 641472 42854 641481
rect 42798 641407 42854 641416
rect 33782 639840 33838 639849
rect 33782 639775 33838 639784
rect 32402 638208 32458 638217
rect 32402 638143 32458 638152
rect 32416 629950 32444 638143
rect 32404 629944 32456 629950
rect 32404 629886 32456 629892
rect 33796 628590 33824 639775
rect 40682 639432 40738 639441
rect 40682 639367 40738 639376
rect 35162 637800 35218 637809
rect 35162 637735 35218 637744
rect 35176 629921 35204 637735
rect 35162 629912 35218 629921
rect 35162 629847 35218 629856
rect 40696 629105 40724 639367
rect 40866 639024 40922 639033
rect 40866 638959 40922 638968
rect 40682 629096 40738 629105
rect 40682 629031 40738 629040
rect 40880 628969 40908 638959
rect 42798 638616 42854 638625
rect 42798 638551 42854 638560
rect 41050 637392 41106 637401
rect 41050 637327 41106 637336
rect 41064 629241 41092 637327
rect 41788 629944 41840 629950
rect 41788 629886 41840 629892
rect 41050 629232 41106 629241
rect 41050 629167 41106 629176
rect 40866 628960 40922 628969
rect 40866 628895 40922 628904
rect 33784 628584 33836 628590
rect 33784 628526 33836 628532
rect 41800 627434 41828 629886
rect 42524 628584 42576 628590
rect 42524 628526 42576 628532
rect 41788 627428 41840 627434
rect 41788 627370 41840 627376
rect 41788 627088 41840 627094
rect 41788 627030 41840 627036
rect 41800 626620 41828 627030
rect 42536 625326 42564 628526
rect 42156 625320 42208 625326
rect 42156 625262 42208 625268
rect 42524 625320 42576 625326
rect 42524 625262 42576 625268
rect 42168 624784 42196 625262
rect 42522 625152 42578 625161
rect 42522 625087 42578 625096
rect 42156 624708 42208 624714
rect 42156 624650 42208 624656
rect 42168 624172 42196 624650
rect 42536 623898 42564 625087
rect 42524 623892 42576 623898
rect 42524 623834 42576 623840
rect 42522 623792 42578 623801
rect 42522 623727 42578 623736
rect 42156 623484 42208 623490
rect 42156 623426 42208 623432
rect 42168 622948 42196 623426
rect 42536 622198 42564 623727
rect 42064 622192 42116 622198
rect 42064 622134 42116 622140
rect 42524 622192 42576 622198
rect 42524 622134 42576 622140
rect 42076 621792 42104 622134
rect 42812 622062 42840 638551
rect 42890 635760 42946 635769
rect 42890 635695 42946 635704
rect 42524 622056 42576 622062
rect 42524 621998 42576 622004
rect 42800 622056 42852 622062
rect 42800 621998 42852 622004
rect 41786 621480 41842 621489
rect 41786 621415 41842 621424
rect 41800 621112 41828 621415
rect 42064 620832 42116 620838
rect 42064 620774 42116 620780
rect 42076 620500 42104 620774
rect 42536 620362 42564 621998
rect 42064 620356 42116 620362
rect 42064 620298 42116 620304
rect 42524 620356 42576 620362
rect 42524 620298 42576 620304
rect 42076 619956 42104 620298
rect 42904 620226 42932 635695
rect 43074 635352 43130 635361
rect 43074 635287 43130 635296
rect 42984 626612 43036 626618
rect 42984 626554 43036 626560
rect 42996 624714 43024 626554
rect 42984 624708 43036 624714
rect 42984 624650 43036 624656
rect 43088 620838 43116 635287
rect 43076 620832 43128 620838
rect 43076 620774 43128 620780
rect 42524 620220 42576 620226
rect 42524 620162 42576 620168
rect 42892 620220 42944 620226
rect 42892 620162 42944 620168
rect 42246 619032 42302 619041
rect 42246 618967 42302 618976
rect 42156 617908 42208 617914
rect 42156 617850 42208 617856
rect 42168 617440 42196 617850
rect 42064 617160 42116 617166
rect 42064 617102 42116 617108
rect 42076 616828 42104 617102
rect 42260 616162 42288 618967
rect 42536 617914 42564 620162
rect 42524 617908 42576 617914
rect 42524 617850 42576 617856
rect 42524 617772 42576 617778
rect 42524 617714 42576 617720
rect 42536 617166 42564 617714
rect 42524 617160 42576 617166
rect 42524 617102 42576 617108
rect 42522 616856 42578 616865
rect 42522 616791 42578 616800
rect 42182 616134 42288 616162
rect 42246 616040 42302 616049
rect 42246 615975 42302 615984
rect 42260 615618 42288 615975
rect 42182 615590 42288 615618
rect 41878 614136 41934 614145
rect 41878 614071 41934 614080
rect 41892 613768 41920 614071
rect 42536 613494 42564 616791
rect 42156 613488 42208 613494
rect 42156 613430 42208 613436
rect 42524 613488 42576 613494
rect 42524 613430 42576 613436
rect 42168 613121 42196 613430
rect 41786 612776 41842 612785
rect 41786 612711 41842 612720
rect 41800 612476 41828 612711
rect 8588 602276 8616 602412
rect 9048 602276 9076 602412
rect 9508 602276 9536 602412
rect 9968 602276 9996 602412
rect 10428 602276 10456 602412
rect 10888 602276 10916 602412
rect 11348 602276 11376 602412
rect 11808 602276 11836 602412
rect 12268 602276 12296 602412
rect 12728 602276 12756 602412
rect 13188 602276 13216 602412
rect 13648 602276 13676 602412
rect 14108 602276 14136 602412
rect 35806 601896 35862 601905
rect 35806 601831 35862 601840
rect 35820 601730 35848 601831
rect 35808 601724 35860 601730
rect 35808 601666 35860 601672
rect 35808 601588 35860 601594
rect 35808 601530 35860 601536
rect 35716 601520 35768 601526
rect 35820 601497 35848 601530
rect 35716 601462 35768 601468
rect 35806 601488 35862 601497
rect 35728 600681 35756 601462
rect 35806 601423 35862 601432
rect 35808 601384 35860 601390
rect 35808 601326 35860 601332
rect 35820 601089 35848 601326
rect 35806 601080 35862 601089
rect 35806 601015 35862 601024
rect 35714 600672 35770 600681
rect 35714 600607 35770 600616
rect 42798 597680 42854 597689
rect 42798 597615 42854 597624
rect 39302 597000 39358 597009
rect 39302 596935 39358 596944
rect 33782 594960 33838 594969
rect 33782 594895 33838 594904
rect 32402 593328 32458 593337
rect 32402 593263 32458 593272
rect 32416 585818 32444 593263
rect 33796 585886 33824 594895
rect 33784 585880 33836 585886
rect 33784 585822 33836 585828
rect 32404 585812 32456 585818
rect 32404 585754 32456 585760
rect 39316 585177 39344 596935
rect 40682 596592 40738 596601
rect 40682 596527 40738 596536
rect 39302 585168 39358 585177
rect 39302 585103 39358 585112
rect 40696 584594 40724 596527
rect 40774 595776 40830 595785
rect 40774 595711 40830 595720
rect 40788 584662 40816 595711
rect 42062 594008 42118 594017
rect 42062 593943 42118 593952
rect 41510 591288 41566 591297
rect 41510 591223 41566 591232
rect 41524 590073 41552 591223
rect 41510 590064 41566 590073
rect 41510 589999 41566 590008
rect 41524 589966 41552 589999
rect 41512 589960 41564 589966
rect 41512 589902 41564 589908
rect 41880 585880 41932 585886
rect 41880 585822 41932 585828
rect 41788 585812 41840 585818
rect 41788 585754 41840 585760
rect 40776 584656 40828 584662
rect 40776 584598 40828 584604
rect 40684 584588 40736 584594
rect 40684 584530 40736 584536
rect 41800 584225 41828 585754
rect 41892 584254 41920 585822
rect 41972 584588 42024 584594
rect 41972 584530 42024 584536
rect 41880 584248 41932 584254
rect 41786 584216 41842 584225
rect 41984 584225 42012 584530
rect 42076 584254 42104 593943
rect 42432 584656 42484 584662
rect 42432 584598 42484 584604
rect 42064 584248 42116 584254
rect 41880 584190 41932 584196
rect 41970 584216 42026 584225
rect 41786 584151 41842 584160
rect 42064 584190 42116 584196
rect 41970 584151 42026 584160
rect 41880 583976 41932 583982
rect 41880 583918 41932 583924
rect 41892 583440 41920 583918
rect 42444 583681 42472 584598
rect 42708 584248 42760 584254
rect 42708 584190 42760 584196
rect 42430 583672 42486 583681
rect 42430 583607 42486 583616
rect 41970 582176 42026 582185
rect 41970 582111 42026 582120
rect 41984 581604 42012 582111
rect 42156 581324 42208 581330
rect 42156 581266 42208 581272
rect 42168 580961 42196 581266
rect 41786 580272 41842 580281
rect 41786 580207 41842 580216
rect 41800 579768 41828 580207
rect 41786 579048 41842 579057
rect 41786 578983 41842 578992
rect 41800 578544 41828 578983
rect 42156 578468 42208 578474
rect 42156 578410 42208 578416
rect 42168 578218 42196 578410
rect 42076 578190 42196 578218
rect 42076 577932 42104 578190
rect 41786 577552 41842 577561
rect 41786 577487 41842 577496
rect 41800 577281 41828 577487
rect 42156 576972 42208 576978
rect 42156 576914 42208 576920
rect 42168 576708 42196 576914
rect 42720 576881 42748 584190
rect 42706 576872 42762 576881
rect 42706 576807 42762 576816
rect 42432 576360 42484 576366
rect 42432 576302 42484 576308
rect 42338 575920 42394 575929
rect 42338 575855 42394 575864
rect 42156 574592 42208 574598
rect 42156 574534 42208 574540
rect 42168 574260 42196 574534
rect 42352 574122 42380 575855
rect 42444 574598 42472 576302
rect 42432 574592 42484 574598
rect 42432 574534 42484 574540
rect 42156 574116 42208 574122
rect 42156 574058 42208 574064
rect 42340 574116 42392 574122
rect 42340 574058 42392 574064
rect 42168 573580 42196 574058
rect 42338 573744 42394 573753
rect 42338 573679 42394 573688
rect 42156 573504 42208 573510
rect 42156 573446 42208 573452
rect 42168 572968 42196 573446
rect 41970 572792 42026 572801
rect 41970 572727 42026 572736
rect 41984 572424 42012 572727
rect 42352 571538 42380 573679
rect 42706 571568 42762 571577
rect 42340 571532 42392 571538
rect 42706 571503 42762 571512
rect 42340 571474 42392 571480
rect 42064 570920 42116 570926
rect 42064 570862 42116 570868
rect 42076 570588 42104 570862
rect 42154 570480 42210 570489
rect 42154 570415 42210 570424
rect 42168 569908 42196 570415
rect 42720 569634 42748 571503
rect 42064 569628 42116 569634
rect 42064 569570 42116 569576
rect 42708 569628 42760 569634
rect 42708 569570 42760 569576
rect 42076 569296 42104 569570
rect 35624 562352 35676 562358
rect 35624 562294 35676 562300
rect 8588 559164 8616 559300
rect 9048 559164 9076 559300
rect 9508 559164 9536 559300
rect 9968 559164 9996 559300
rect 10428 559164 10456 559300
rect 10888 559164 10916 559300
rect 11348 559164 11376 559300
rect 11808 559164 11836 559300
rect 12268 559164 12296 559300
rect 12728 559164 12756 559300
rect 13188 559164 13216 559300
rect 13648 559164 13676 559300
rect 14108 559164 14136 559300
rect 35636 558385 35664 562294
rect 35622 558376 35678 558385
rect 35806 558376 35862 558385
rect 35622 558311 35678 558320
rect 35716 558340 35768 558346
rect 35806 558311 35862 558320
rect 35716 558282 35768 558288
rect 35728 557977 35756 558282
rect 35820 558210 35848 558311
rect 35808 558204 35860 558210
rect 35808 558146 35860 558152
rect 35714 557968 35770 557977
rect 35714 557903 35770 557912
rect 42812 554849 42840 597615
rect 42890 594416 42946 594425
rect 42890 594351 42946 594360
rect 42904 581670 42932 594351
rect 42982 592784 43038 592793
rect 42982 592719 43038 592728
rect 42892 581664 42944 581670
rect 42892 581606 42944 581612
rect 42892 579692 42944 579698
rect 42892 579634 42944 579640
rect 42904 578474 42932 579634
rect 42892 578468 42944 578474
rect 42892 578410 42944 578416
rect 42996 576366 43024 592719
rect 43076 581664 43128 581670
rect 43076 581606 43128 581612
rect 42984 576360 43036 576366
rect 42984 576302 43036 576308
rect 43088 573510 43116 581606
rect 43168 578264 43220 578270
rect 43168 578206 43220 578212
rect 43180 576978 43208 578206
rect 43168 576972 43220 576978
rect 43168 576914 43220 576920
rect 43076 573504 43128 573510
rect 43076 573446 43128 573452
rect 42982 556880 43038 556889
rect 42982 556815 43038 556824
rect 42890 556064 42946 556073
rect 42890 555999 42946 556008
rect 42798 554840 42854 554849
rect 42798 554775 42854 554784
rect 42904 554690 42932 555999
rect 42812 554662 42932 554690
rect 40866 553888 40922 553897
rect 40866 553823 40922 553832
rect 40682 553480 40738 553489
rect 40682 553415 40738 553424
rect 32402 552664 32458 552673
rect 32402 552599 32458 552608
rect 31022 551848 31078 551857
rect 31022 551783 31078 551792
rect 31036 543046 31064 551783
rect 31666 548176 31722 548185
rect 31666 548111 31722 548120
rect 31680 547194 31708 548111
rect 31668 547188 31720 547194
rect 31668 547130 31720 547136
rect 31024 543040 31076 543046
rect 31024 542982 31076 542988
rect 32416 542881 32444 552599
rect 35808 547188 35860 547194
rect 35808 547130 35860 547136
rect 35820 546961 35848 547130
rect 35806 546952 35862 546961
rect 35806 546887 35862 546896
rect 32402 542872 32458 542881
rect 32402 542807 32458 542816
rect 40696 542366 40724 553415
rect 40774 552256 40830 552265
rect 40774 552191 40830 552200
rect 40684 542360 40736 542366
rect 40788 542337 40816 552191
rect 40880 545193 40908 553823
rect 40958 553072 41014 553081
rect 40958 553007 41014 553016
rect 40866 545184 40922 545193
rect 40866 545119 40922 545128
rect 40972 543017 41000 553007
rect 41788 543040 41840 543046
rect 40958 543008 41014 543017
rect 41788 542982 41840 542988
rect 40958 542943 41014 542952
rect 40684 542302 40736 542308
rect 40774 542328 40830 542337
rect 40774 542263 40830 542272
rect 41800 541074 41828 542982
rect 42708 542360 42760 542366
rect 42708 542302 42760 542308
rect 41788 541068 41840 541074
rect 41788 541010 41840 541016
rect 41788 540796 41840 540802
rect 41788 540738 41840 540744
rect 41800 540260 41828 540738
rect 42720 538966 42748 542302
rect 42064 538960 42116 538966
rect 42064 538902 42116 538908
rect 42708 538960 42760 538966
rect 42708 538902 42760 538908
rect 42076 538424 42104 538902
rect 42156 538212 42208 538218
rect 42156 538154 42208 538160
rect 42168 537744 42196 538154
rect 42064 537124 42116 537130
rect 42064 537066 42116 537072
rect 42076 536588 42104 537066
rect 42616 536852 42668 536858
rect 42616 536794 42668 536800
rect 42628 536042 42656 536794
rect 42616 536036 42668 536042
rect 42616 535978 42668 535984
rect 42614 535936 42670 535945
rect 42614 535871 42670 535880
rect 42156 535832 42208 535838
rect 42156 535774 42208 535780
rect 42168 535364 42196 535774
rect 42064 535288 42116 535294
rect 42064 535230 42116 535236
rect 42076 534752 42104 535230
rect 41786 534576 41842 534585
rect 41786 534511 41842 534520
rect 41800 534072 41828 534511
rect 42628 534002 42656 535871
rect 42156 533996 42208 534002
rect 42156 533938 42208 533944
rect 42616 533996 42668 534002
rect 42616 533938 42668 533944
rect 42168 533528 42196 533938
rect 42614 533896 42670 533905
rect 42614 533831 42670 533840
rect 42338 532672 42394 532681
rect 42338 532607 42394 532616
rect 42156 531480 42208 531486
rect 42156 531422 42208 531428
rect 42168 531045 42196 531422
rect 41786 530768 41842 530777
rect 41786 530703 41842 530712
rect 41800 530400 41828 530703
rect 42156 530120 42208 530126
rect 42156 530062 42208 530068
rect 42168 529757 42196 530062
rect 42352 529650 42380 532607
rect 42628 531486 42656 533831
rect 42616 531480 42668 531486
rect 42616 531422 42668 531428
rect 42616 531344 42668 531350
rect 42616 531286 42668 531292
rect 42628 530126 42656 531286
rect 42616 530120 42668 530126
rect 42616 530062 42668 530068
rect 42340 529644 42392 529650
rect 42340 529586 42392 529592
rect 42338 529544 42394 529553
rect 42156 529508 42208 529514
rect 42338 529479 42394 529488
rect 42156 529450 42208 529456
rect 42168 529205 42196 529450
rect 42076 527270 42104 527340
rect 42352 527270 42380 529479
rect 42614 529408 42670 529417
rect 42614 529343 42670 529352
rect 42064 527264 42116 527270
rect 42064 527206 42116 527212
rect 42340 527264 42392 527270
rect 42340 527206 42392 527212
rect 42156 527196 42208 527202
rect 42156 527138 42208 527144
rect 42168 526728 42196 527138
rect 42628 526658 42656 529343
rect 42156 526652 42208 526658
rect 42156 526594 42208 526600
rect 42616 526652 42668 526658
rect 42616 526594 42668 526600
rect 42168 526077 42196 526594
rect 40684 518968 40736 518974
rect 40684 518910 40736 518916
rect 40696 432614 40724 518910
rect 40868 497480 40920 497486
rect 40868 497422 40920 497428
rect 40684 432608 40736 432614
rect 40684 432550 40736 432556
rect 8588 431596 8616 431664
rect 9048 431596 9076 431664
rect 9508 431596 9536 431664
rect 9968 431596 9996 431664
rect 10428 431596 10456 431664
rect 10888 431596 10916 431664
rect 11348 431596 11376 431664
rect 11808 431596 11836 431664
rect 12268 431596 12296 431664
rect 12728 431596 12756 431664
rect 13188 431596 13216 431664
rect 13648 431596 13676 431664
rect 14108 431596 14136 431664
rect 40880 430166 40908 497422
rect 41788 432608 41840 432614
rect 41788 432550 41840 432556
rect 41800 430545 41828 432550
rect 41786 430536 41842 430545
rect 41786 430471 41842 430480
rect 40868 430160 40920 430166
rect 41788 430160 41840 430166
rect 40868 430102 40920 430108
rect 41786 430128 41788 430137
rect 41840 430128 41842 430137
rect 41786 430063 41842 430072
rect 42812 428913 42840 554662
rect 42996 554554 43024 556815
rect 42904 554526 43024 554554
rect 42904 429729 42932 554526
rect 42982 551168 43038 551177
rect 42982 551103 43038 551112
rect 42996 531350 43024 551103
rect 43074 549944 43130 549953
rect 43074 549879 43130 549888
rect 43088 535294 43116 549879
rect 43168 539640 43220 539646
rect 43168 539582 43220 539588
rect 43180 538218 43208 539582
rect 43168 538212 43220 538218
rect 43168 538154 43220 538160
rect 43076 535288 43128 535294
rect 43076 535230 43128 535236
rect 42984 531344 43036 531350
rect 42984 531286 43036 531292
rect 42984 528624 43036 528630
rect 42984 528566 43036 528572
rect 42996 527202 43024 528566
rect 42984 527196 43036 527202
rect 42984 527138 43036 527144
rect 43350 430944 43406 430953
rect 43350 430879 43406 430888
rect 43364 430642 43392 430879
rect 43352 430636 43404 430642
rect 43352 430578 43404 430584
rect 42890 429720 42946 429729
rect 42890 429655 42946 429664
rect 42798 428904 42854 428913
rect 42798 428839 42854 428848
rect 43166 427680 43222 427689
rect 43166 427615 43222 427624
rect 42890 426864 42946 426873
rect 42890 426799 42946 426808
rect 41786 426456 41842 426465
rect 41786 426391 41842 426400
rect 41800 425746 41828 426391
rect 40776 425740 40828 425746
rect 40776 425682 40828 425688
rect 41788 425740 41840 425746
rect 41788 425682 41840 425688
rect 35162 425232 35218 425241
rect 35162 425167 35218 425176
rect 32402 424416 32458 424425
rect 32402 424351 32458 424360
rect 31022 422376 31078 422385
rect 31022 422311 31078 422320
rect 31036 414730 31064 422311
rect 32416 414866 32444 424351
rect 32404 414860 32456 414866
rect 32404 414802 32456 414808
rect 31024 414724 31076 414730
rect 31024 414666 31076 414672
rect 35176 414633 35204 425167
rect 40788 425077 40816 425682
rect 40774 425068 40830 425077
rect 40774 425003 40830 425012
rect 41326 425068 41382 425077
rect 41326 425003 41382 425012
rect 41340 418033 41368 425003
rect 42798 421968 42854 421977
rect 42798 421903 42854 421912
rect 41786 419520 41842 419529
rect 41786 419455 41788 419464
rect 41840 419455 41842 419464
rect 41788 419426 41840 419432
rect 41326 418024 41382 418033
rect 41326 417959 41382 417968
rect 41880 414860 41932 414866
rect 41880 414802 41932 414808
rect 35162 414624 35218 414633
rect 35162 414559 35218 414568
rect 41892 413438 41920 414802
rect 42524 414724 42576 414730
rect 42524 414666 42576 414672
rect 41880 413432 41932 413438
rect 41880 413374 41932 413380
rect 41880 413160 41932 413166
rect 41880 413102 41932 413108
rect 41892 412624 41920 413102
rect 42154 411224 42210 411233
rect 42154 411159 42210 411168
rect 42168 410788 42196 411159
rect 42156 410712 42208 410718
rect 42156 410654 42208 410660
rect 42168 410176 42196 410654
rect 41786 409456 41842 409465
rect 41786 409391 41842 409400
rect 41800 408952 41828 409391
rect 42064 408196 42116 408202
rect 42064 408138 42116 408144
rect 42076 407796 42104 408138
rect 42536 407658 42564 414666
rect 42156 407652 42208 407658
rect 42156 407594 42208 407600
rect 42524 407652 42576 407658
rect 42524 407594 42576 407600
rect 42168 407116 42196 407594
rect 42064 406836 42116 406842
rect 42064 406778 42116 406784
rect 42076 406504 42104 406778
rect 41786 406328 41842 406337
rect 41786 406263 41842 406272
rect 41800 405929 41828 406263
rect 42812 403918 42840 421903
rect 42156 403912 42208 403918
rect 42156 403854 42208 403860
rect 42800 403912 42852 403918
rect 42800 403854 42852 403860
rect 42168 403444 42196 403854
rect 42156 402960 42208 402966
rect 42156 402902 42208 402908
rect 42168 402801 42196 402902
rect 41786 402520 41842 402529
rect 41786 402455 41842 402464
rect 41800 402152 41828 402455
rect 41970 401840 42026 401849
rect 41970 401775 42026 401784
rect 41984 401608 42012 401775
rect 41786 400072 41842 400081
rect 41786 400007 41842 400016
rect 41800 399772 41828 400007
rect 41786 399664 41842 399673
rect 41786 399599 41842 399608
rect 41800 399121 41828 399599
rect 41786 398848 41842 398857
rect 41786 398783 41842 398792
rect 41800 398480 41828 398783
rect 8588 388348 8616 388484
rect 9048 388348 9076 388484
rect 9508 388348 9536 388484
rect 9968 388348 9996 388484
rect 10428 388348 10456 388484
rect 10888 388348 10916 388484
rect 11348 388348 11376 388484
rect 11808 388348 11836 388484
rect 12268 388348 12296 388484
rect 12728 388348 12756 388484
rect 13188 388348 13216 388484
rect 13648 388348 13676 388484
rect 14108 388348 14136 388484
rect 35716 387796 35768 387802
rect 35716 387738 35768 387744
rect 35624 387524 35676 387530
rect 35624 387466 35676 387472
rect 35636 387161 35664 387466
rect 35622 387152 35678 387161
rect 35622 387087 35678 387096
rect 35728 386753 35756 387738
rect 35808 387660 35860 387666
rect 35808 387602 35860 387608
rect 35820 387569 35848 387602
rect 35806 387560 35862 387569
rect 35806 387495 35862 387504
rect 35808 387388 35860 387394
rect 35808 387330 35860 387336
rect 35820 387161 35848 387330
rect 35806 387152 35862 387161
rect 35806 387087 35862 387096
rect 35714 386744 35770 386753
rect 35714 386679 35770 386688
rect 42904 384033 42932 426799
rect 43074 421152 43130 421161
rect 43074 421087 43130 421096
rect 43088 408202 43116 421087
rect 43076 408196 43128 408202
rect 43076 408138 43128 408144
rect 43180 384849 43208 427615
rect 43166 384840 43222 384849
rect 43166 384775 43222 384784
rect 42890 384024 42946 384033
rect 42890 383959 42946 383968
rect 42798 383616 42854 383625
rect 42798 383551 42854 383560
rect 40866 382664 40922 382673
rect 40866 382599 40922 382608
rect 37922 381440 37978 381449
rect 37922 381375 37978 381384
rect 31022 381032 31078 381041
rect 31022 380967 31078 380976
rect 31036 371890 31064 380967
rect 33782 378176 33838 378185
rect 33782 378111 33838 378120
rect 33796 371929 33824 378111
rect 35806 377360 35862 377369
rect 35806 377295 35862 377304
rect 35820 376038 35848 377295
rect 35808 376032 35860 376038
rect 35808 375974 35860 375980
rect 33782 371920 33838 371929
rect 31024 371884 31076 371890
rect 33782 371855 33838 371864
rect 31024 371826 31076 371832
rect 37936 371385 37964 381375
rect 40682 379400 40738 379409
rect 40682 379335 40738 379344
rect 37922 371376 37978 371385
rect 37922 371311 37978 371320
rect 40696 370598 40724 379335
rect 40880 371278 40908 382599
rect 41510 376136 41566 376145
rect 41510 376071 41566 376080
rect 41524 376038 41552 376071
rect 41512 376032 41564 376038
rect 41512 375974 41564 375980
rect 42340 371884 42392 371890
rect 42340 371826 42392 371832
rect 40868 371272 40920 371278
rect 40868 371214 40920 371220
rect 40684 370592 40736 370598
rect 40684 370534 40736 370540
rect 41788 370592 41840 370598
rect 41788 370534 41840 370540
rect 41800 370297 41828 370534
rect 41786 370288 41842 370297
rect 41786 370223 41842 370232
rect 42352 369714 42380 371826
rect 42708 371272 42760 371278
rect 42708 371214 42760 371220
rect 42156 369708 42208 369714
rect 42156 369650 42208 369656
rect 42340 369708 42392 369714
rect 42340 369650 42392 369656
rect 42168 369444 42196 369650
rect 42720 368150 42748 371214
rect 42156 368144 42208 368150
rect 42156 368086 42208 368092
rect 42708 368144 42760 368150
rect 42708 368086 42760 368092
rect 42168 367608 42196 368086
rect 42168 366858 42196 366961
rect 42156 366852 42208 366858
rect 42156 366794 42208 366800
rect 42708 366852 42760 366858
rect 42708 366794 42760 366800
rect 41878 366344 41934 366353
rect 41878 366279 41934 366288
rect 41892 365772 41920 366279
rect 42156 365016 42208 365022
rect 42156 364958 42208 364964
rect 42168 364548 42196 364958
rect 42156 364336 42208 364342
rect 42156 364278 42208 364284
rect 42168 363936 42196 364278
rect 42720 364274 42748 366794
rect 42708 364268 42760 364274
rect 42708 364210 42760 364216
rect 41970 363760 42026 363769
rect 41970 363695 42026 363704
rect 41984 363256 42012 363695
rect 41786 362944 41842 362953
rect 41786 362879 41842 362888
rect 41800 362712 41828 362879
rect 42064 360732 42116 360738
rect 42064 360674 42116 360680
rect 42076 360264 42104 360674
rect 41786 360088 41842 360097
rect 41786 360023 41842 360032
rect 41800 359584 41828 360023
rect 42156 359508 42208 359514
rect 42156 359450 42208 359456
rect 42168 358972 42196 359450
rect 41786 358728 41842 358737
rect 41786 358663 41842 358672
rect 41800 358428 41828 358663
rect 41786 356960 41842 356969
rect 41786 356895 41842 356904
rect 41800 356592 41828 356895
rect 42156 356040 42208 356046
rect 42156 355982 42208 355988
rect 42168 355912 42196 355982
rect 41786 355736 41842 355745
rect 41786 355671 41842 355680
rect 41800 355300 41828 355671
rect 8588 345100 8616 345236
rect 9048 345100 9076 345236
rect 9508 345100 9536 345236
rect 9968 345100 9996 345236
rect 10428 345100 10456 345236
rect 10888 345100 10916 345236
rect 11348 345100 11376 345236
rect 11808 345100 11836 345236
rect 12268 345100 12296 345236
rect 12728 345100 12756 345236
rect 13188 345100 13216 345236
rect 13648 345100 13676 345236
rect 14108 345100 14136 345236
rect 35716 344480 35768 344486
rect 35716 344422 35768 344428
rect 35622 344312 35678 344321
rect 35622 344247 35678 344256
rect 35636 344214 35664 344247
rect 35624 344208 35676 344214
rect 35624 344150 35676 344156
rect 35728 343913 35756 344422
rect 35808 344344 35860 344350
rect 35806 344312 35808 344321
rect 35860 344312 35862 344321
rect 35806 344247 35862 344256
rect 35714 343904 35770 343913
rect 35714 343839 35770 343848
rect 42812 340921 42840 383551
rect 42890 380352 42946 380361
rect 42890 380287 42946 380296
rect 42904 359514 42932 380287
rect 42982 378720 43038 378729
rect 42982 378655 43038 378664
rect 42996 360738 43024 378655
rect 43074 377904 43130 377913
rect 43074 377839 43130 377848
rect 43088 365022 43116 377839
rect 43076 365016 43128 365022
rect 43076 364958 43128 364964
rect 42984 360732 43036 360738
rect 42984 360674 43036 360680
rect 42892 359508 42944 359514
rect 42892 359450 42944 359456
rect 42798 340912 42854 340921
rect 42798 340847 42854 340856
rect 42798 340504 42854 340513
rect 42798 340439 42854 340448
rect 40866 339416 40922 339425
rect 40866 339351 40922 339360
rect 40682 338192 40738 338201
rect 40682 338127 40738 338136
rect 30378 334112 30434 334121
rect 30378 334047 30434 334056
rect 30392 333305 30420 334047
rect 30378 333296 30434 333305
rect 30378 333231 30380 333240
rect 30432 333231 30434 333240
rect 30380 333202 30432 333208
rect 30392 333171 30420 333202
rect 40696 328409 40724 338127
rect 40880 334121 40908 339351
rect 40866 334112 40922 334121
rect 40866 334047 40922 334056
rect 40682 328400 40738 328409
rect 40682 328335 40738 328344
rect 42064 326800 42116 326806
rect 42064 326742 42116 326748
rect 42076 326264 42104 326742
rect 41786 324864 41842 324873
rect 41786 324799 41842 324808
rect 41800 324428 41828 324799
rect 42168 323338 42196 323748
rect 42156 323332 42208 323338
rect 42156 323274 42208 323280
rect 42616 323332 42668 323338
rect 42616 323274 42668 323280
rect 42064 322924 42116 322930
rect 42064 322866 42116 322872
rect 42076 322592 42104 322866
rect 42628 321570 42656 323274
rect 42616 321564 42668 321570
rect 42616 321506 42668 321512
rect 42156 321496 42208 321502
rect 42156 321438 42208 321444
rect 42168 321368 42196 321438
rect 41786 321192 41842 321201
rect 41786 321127 41842 321136
rect 41800 320725 41828 321127
rect 42168 320006 42196 320076
rect 42156 320000 42208 320006
rect 41970 319968 42026 319977
rect 42156 319942 42208 319948
rect 41970 319903 42026 319912
rect 41984 319532 42012 319903
rect 41786 317384 41842 317393
rect 41786 317319 41842 317328
rect 41800 317045 41828 317319
rect 42156 316736 42208 316742
rect 42156 316678 42208 316684
rect 42168 316404 42196 316678
rect 41786 315888 41842 315897
rect 41786 315823 41842 315832
rect 41800 315757 41828 315823
rect 41786 315480 41842 315489
rect 41786 315415 41842 315424
rect 41800 315180 41828 315415
rect 41878 313848 41934 313857
rect 41878 313783 41934 313792
rect 41892 313344 41920 313783
rect 41786 313168 41842 313177
rect 41786 313103 41842 313112
rect 41800 312732 41828 313103
rect 41786 312352 41842 312361
rect 41786 312287 41842 312296
rect 41800 312052 41828 312287
rect 41972 307080 42024 307086
rect 41972 307022 42024 307028
rect 8588 301988 8616 302124
rect 9048 301988 9076 302124
rect 9508 301988 9536 302124
rect 9968 301988 9996 302124
rect 10428 301988 10456 302124
rect 10888 301988 10916 302124
rect 11348 301988 11376 302124
rect 11808 301988 11836 302124
rect 12268 301988 12296 302124
rect 12728 301988 12756 302124
rect 13188 301988 13216 302124
rect 13648 301988 13676 302124
rect 14108 301988 14136 302124
rect 41984 300937 42012 307022
rect 42062 301336 42118 301345
rect 42062 301271 42118 301280
rect 42076 300966 42104 301271
rect 42064 300960 42116 300966
rect 41970 300928 42026 300937
rect 42064 300902 42116 300908
rect 41970 300863 42026 300872
rect 42812 297673 42840 340439
rect 43074 338056 43130 338065
rect 43074 337991 43130 338000
rect 42982 336424 43038 336433
rect 42982 336359 43038 336368
rect 42890 334792 42946 334801
rect 42890 334727 42946 334736
rect 42904 321502 42932 334727
rect 42996 322930 43024 336359
rect 43088 326806 43116 337991
rect 43076 326800 43128 326806
rect 43076 326742 43128 326748
rect 42984 322924 43036 322930
rect 42984 322866 43036 322872
rect 42892 321496 42944 321502
rect 42892 321438 42944 321444
rect 43074 298888 43130 298897
rect 43074 298823 43130 298832
rect 42798 297664 42854 297673
rect 42798 297599 42854 297608
rect 33782 296440 33838 296449
rect 33782 296375 33838 296384
rect 33796 284889 33824 296375
rect 42430 294808 42486 294817
rect 42430 294743 42486 294752
rect 33782 284880 33838 284889
rect 33782 284815 33838 284824
rect 42444 283626 42472 294743
rect 42982 293176 43038 293185
rect 42982 293111 43038 293120
rect 42890 291952 42946 291961
rect 42890 291887 42946 291896
rect 42156 283620 42208 283626
rect 42156 283562 42208 283568
rect 42432 283620 42484 283626
rect 42432 283562 42484 283568
rect 42168 283045 42196 283562
rect 41786 281480 41842 281489
rect 41786 281415 41842 281424
rect 41800 281180 41828 281415
rect 42156 281104 42208 281110
rect 42156 281046 42208 281052
rect 42168 280568 42196 281046
rect 42156 279880 42208 279886
rect 42156 279822 42208 279828
rect 42168 279344 42196 279822
rect 42706 278760 42762 278769
rect 42706 278695 42762 278704
rect 42064 278656 42116 278662
rect 42064 278598 42116 278604
rect 42076 278188 42104 278598
rect 41800 277409 41828 277508
rect 41786 277400 41842 277409
rect 41786 277335 41842 277344
rect 42156 277160 42208 277166
rect 42156 277102 42208 277108
rect 42168 276896 42196 277102
rect 41786 276720 41842 276729
rect 41786 276655 41842 276664
rect 41800 276352 41828 276655
rect 42156 274304 42208 274310
rect 42156 274246 42208 274252
rect 42168 273836 42196 274246
rect 42064 273352 42116 273358
rect 42064 273294 42116 273300
rect 42076 273224 42104 273294
rect 42720 273086 42748 278695
rect 42904 277166 42932 291887
rect 42996 279886 43024 293111
rect 42984 279880 43036 279886
rect 42984 279822 43036 279828
rect 42892 277160 42944 277166
rect 42892 277102 42944 277108
rect 42156 273080 42208 273086
rect 42156 273022 42208 273028
rect 42708 273080 42760 273086
rect 42708 273022 42760 273028
rect 42168 272544 42196 273022
rect 41786 272368 41842 272377
rect 41786 272303 41842 272312
rect 41800 272000 41828 272303
rect 41970 270464 42026 270473
rect 41970 270399 42026 270408
rect 41984 270164 42012 270399
rect 41786 269784 41842 269793
rect 41786 269719 41842 269728
rect 41800 269521 41828 269719
rect 41786 269104 41842 269113
rect 41786 269039 41842 269048
rect 41800 268872 41828 269039
rect 8588 258740 8616 258876
rect 9048 258740 9076 258876
rect 9508 258740 9536 258876
rect 9968 258740 9996 258876
rect 10428 258740 10456 258876
rect 10888 258740 10916 258876
rect 11348 258740 11376 258876
rect 11808 258740 11836 258876
rect 12268 258740 12296 258876
rect 12728 258740 12756 258876
rect 13188 258740 13216 258876
rect 13648 258740 13676 258876
rect 14108 258740 14136 258876
rect 35806 258360 35862 258369
rect 35806 258295 35862 258304
rect 35820 258126 35848 258295
rect 35808 258120 35860 258126
rect 35808 258062 35860 258068
rect 31668 258052 31720 258058
rect 31668 257994 31720 258000
rect 31680 257961 31708 257994
rect 31666 257952 31722 257961
rect 31576 257916 31628 257922
rect 31666 257887 31722 257896
rect 31576 257858 31628 257864
rect 31588 257145 31616 257858
rect 31668 257780 31720 257786
rect 31668 257722 31720 257728
rect 31680 257553 31708 257722
rect 31666 257544 31722 257553
rect 31666 257479 31722 257488
rect 31574 257136 31630 257145
rect 31574 257071 31630 257080
rect 42890 256456 42946 256465
rect 42890 256391 42946 256400
rect 31022 251832 31078 251841
rect 31022 251767 31078 251776
rect 31036 243545 31064 251767
rect 42706 251560 42762 251569
rect 42706 251495 42762 251504
rect 39946 250608 40002 250617
rect 39946 250543 40002 250552
rect 35806 246528 35862 246537
rect 35806 246463 35862 246472
rect 35820 245682 35848 246463
rect 35808 245676 35860 245682
rect 35808 245618 35860 245624
rect 31022 243536 31078 243545
rect 31022 243471 31078 243480
rect 39960 241641 39988 250543
rect 42720 245818 42748 251495
rect 42798 245848 42854 245857
rect 42432 245812 42484 245818
rect 42432 245754 42484 245760
rect 42708 245812 42760 245818
rect 42798 245783 42854 245792
rect 42708 245754 42760 245760
rect 40038 244624 40094 244633
rect 40038 244559 40094 244568
rect 40052 244225 40080 244559
rect 40038 244216 40094 244225
rect 40038 244151 40094 244160
rect 40498 243536 40554 243545
rect 40498 243471 40554 243480
rect 39946 241632 40002 241641
rect 39946 241567 40002 241576
rect 40512 240961 40540 243471
rect 40498 240952 40554 240961
rect 40498 240887 40554 240896
rect 42444 240378 42472 245754
rect 42706 245712 42762 245721
rect 42706 245647 42762 245656
rect 42156 240372 42208 240378
rect 42156 240314 42208 240320
rect 42432 240372 42484 240378
rect 42432 240314 42484 240320
rect 42168 239836 42196 240314
rect 42720 238921 42748 245647
rect 42706 238912 42762 238921
rect 42706 238847 42762 238856
rect 42708 238808 42760 238814
rect 42708 238750 42760 238756
rect 41878 238504 41934 238513
rect 41878 238439 41934 238448
rect 41892 238000 41920 238439
rect 42720 237969 42748 238750
rect 42812 238105 42840 245783
rect 42798 238096 42854 238105
rect 42798 238031 42854 238040
rect 42706 237960 42762 237969
rect 42706 237895 42762 237904
rect 41786 236736 41842 236745
rect 41786 236671 41842 236680
rect 41800 236164 41828 236671
rect 42156 235408 42208 235414
rect 42156 235350 42208 235356
rect 42168 234969 42196 235350
rect 41786 234832 41842 234841
rect 41786 234767 41842 234776
rect 41800 234328 41828 234767
rect 42156 234048 42208 234054
rect 42156 233990 42208 233996
rect 42168 233681 42196 233990
rect 41786 233336 41842 233345
rect 41786 233271 41842 233280
rect 41800 233104 41828 233271
rect 41800 230489 41828 230656
rect 41786 230480 41842 230489
rect 41786 230415 41842 230424
rect 42064 230376 42116 230382
rect 42064 230318 42116 230324
rect 42076 229976 42104 230318
rect 42154 229936 42210 229945
rect 42154 229871 42210 229880
rect 42168 229364 42196 229871
rect 41786 228984 41842 228993
rect 41786 228919 41842 228928
rect 41800 228820 41828 228919
rect 42062 227352 42118 227361
rect 42062 227287 42118 227296
rect 42076 226984 42104 227287
rect 42156 226704 42208 226710
rect 42156 226646 42208 226652
rect 42168 226304 42196 226646
rect 41786 226128 41842 226137
rect 41786 226063 41842 226072
rect 41800 225692 41828 226063
rect 35716 218952 35768 218958
rect 35716 218894 35768 218900
rect 35624 217320 35676 217326
rect 35624 217262 35676 217268
rect 8588 215492 8616 215628
rect 9048 215492 9076 215628
rect 9508 215492 9536 215628
rect 9968 215492 9996 215628
rect 10428 215492 10456 215628
rect 10888 215492 10916 215628
rect 11348 215492 11376 215628
rect 11808 215492 11836 215628
rect 12268 215492 12296 215628
rect 12728 215492 12756 215628
rect 13188 215492 13216 215628
rect 13648 215492 13676 215628
rect 14108 215492 14136 215628
rect 35636 214713 35664 217262
rect 35622 214704 35678 214713
rect 35622 214639 35678 214648
rect 35728 214305 35756 218894
rect 35806 214704 35862 214713
rect 35806 214639 35862 214648
rect 35820 214606 35848 214639
rect 35808 214600 35860 214606
rect 35808 214542 35860 214548
rect 35714 214296 35770 214305
rect 35714 214231 35770 214240
rect 40868 214260 40920 214266
rect 40868 214202 40920 214208
rect 40684 214124 40736 214130
rect 40684 214066 40736 214072
rect 31206 210216 31262 210225
rect 31206 210151 31262 210160
rect 31022 209808 31078 209817
rect 31022 209743 31078 209752
rect 31036 199481 31064 209743
rect 31022 199472 31078 199481
rect 31022 199407 31078 199416
rect 31220 199345 31248 210151
rect 39302 208584 39358 208593
rect 39302 208519 39358 208528
rect 35806 203280 35862 203289
rect 35806 203215 35862 203224
rect 35820 202910 35848 203215
rect 35808 202904 35860 202910
rect 35808 202846 35860 202852
rect 31206 199336 31262 199345
rect 31206 199271 31262 199280
rect 39316 197713 39344 208519
rect 40696 204513 40724 214066
rect 40880 204921 40908 214202
rect 42800 214192 42852 214198
rect 42800 214134 42852 214140
rect 41788 214056 41840 214062
rect 41788 213998 41840 214004
rect 41328 213988 41380 213994
rect 41328 213930 41380 213936
rect 41340 211041 41368 213930
rect 41800 211721 41828 213998
rect 42812 212537 42840 214134
rect 42904 213761 42932 256391
rect 43088 256057 43116 298823
rect 43456 278186 43484 806239
rect 43548 710938 43576 818314
rect 43640 773673 43668 858366
rect 44270 815280 44326 815289
rect 44270 815215 44326 815224
rect 44178 813648 44234 813657
rect 44178 813583 44234 813592
rect 43626 773664 43682 773673
rect 43626 773599 43682 773608
rect 44192 770817 44220 813583
rect 44284 772449 44312 815215
rect 44362 808344 44418 808353
rect 44362 808279 44418 808288
rect 44376 794986 44404 808279
rect 44364 794980 44416 794986
rect 44364 794922 44416 794928
rect 44730 772848 44786 772857
rect 44730 772783 44786 772792
rect 44270 772440 44326 772449
rect 44270 772375 44326 772384
rect 44178 770808 44234 770817
rect 44178 770743 44234 770752
rect 44638 770400 44694 770409
rect 44638 770335 44694 770344
rect 44362 769992 44418 770001
rect 44362 769927 44418 769936
rect 44376 745958 44404 769927
rect 44454 768360 44510 768369
rect 44454 768295 44510 768304
rect 44468 752146 44496 768295
rect 44546 765504 44602 765513
rect 44546 765439 44602 765448
rect 44456 752140 44508 752146
rect 44456 752082 44508 752088
rect 44560 749426 44588 765439
rect 44548 749420 44600 749426
rect 44548 749362 44600 749368
rect 44364 745952 44416 745958
rect 44364 745894 44416 745900
rect 44178 728920 44234 728929
rect 44178 728855 44234 728864
rect 43536 710932 43588 710938
rect 43536 710874 43588 710880
rect 44192 686089 44220 728855
rect 44652 727705 44680 770335
rect 44744 731406 44772 772783
rect 44836 756294 44864 870810
rect 46204 767372 46256 767378
rect 46204 767314 46256 767320
rect 44824 756288 44876 756294
rect 44824 756230 44876 756236
rect 44916 753568 44968 753574
rect 44916 753510 44968 753516
rect 44732 731400 44784 731406
rect 44732 731342 44784 731348
rect 44638 727696 44694 727705
rect 44638 727631 44694 727640
rect 44546 722800 44602 722809
rect 44546 722735 44602 722744
rect 44362 721984 44418 721993
rect 44362 721919 44418 721928
rect 44376 707266 44404 721919
rect 44560 709374 44588 722735
rect 44824 714876 44876 714882
rect 44824 714818 44876 714824
rect 44548 709368 44600 709374
rect 44548 709310 44600 709316
rect 44364 707260 44416 707266
rect 44364 707202 44416 707208
rect 44270 686488 44326 686497
rect 44270 686423 44326 686432
rect 44178 686080 44234 686089
rect 44178 686015 44234 686024
rect 44178 685672 44234 685681
rect 44178 685607 44234 685616
rect 43536 662448 43588 662454
rect 43536 662390 43588 662396
rect 43548 581330 43576 662390
rect 44192 643113 44220 685607
rect 44284 643793 44312 686423
rect 44362 681184 44418 681193
rect 44362 681119 44418 681128
rect 44376 658306 44404 681119
rect 44454 679960 44510 679969
rect 44454 679895 44510 679904
rect 44468 667962 44496 679895
rect 44456 667956 44508 667962
rect 44456 667898 44508 667904
rect 44364 658300 44416 658306
rect 44364 658242 44416 658248
rect 44270 643784 44326 643793
rect 44270 643719 44326 643728
rect 44362 643240 44418 643249
rect 44362 643175 44418 643184
rect 44178 643104 44234 643113
rect 44178 643039 44234 643048
rect 44178 642288 44234 642297
rect 44178 642223 44234 642232
rect 43628 623824 43680 623830
rect 43628 623766 43680 623772
rect 43640 601662 43668 623766
rect 43628 601656 43680 601662
rect 43628 601598 43680 601604
rect 44086 599856 44142 599865
rect 44086 599791 44142 599800
rect 44100 599570 44128 599791
rect 44192 599729 44220 642223
rect 44270 640792 44326 640801
rect 44270 640727 44326 640736
rect 44178 599720 44234 599729
rect 44178 599655 44234 599664
rect 44100 599542 44220 599570
rect 43536 581324 43588 581330
rect 43536 581266 43588 581272
rect 43536 571396 43588 571402
rect 43536 571338 43588 571344
rect 43548 562358 43576 571338
rect 43536 562352 43588 562358
rect 43536 562294 43588 562300
rect 44192 557297 44220 599542
rect 44284 598097 44312 640727
rect 44376 601526 44404 643175
rect 44454 636984 44510 636993
rect 44454 636919 44510 636928
rect 44468 618322 44496 636919
rect 44836 626618 44864 714818
rect 44928 692102 44956 753510
rect 44916 692096 44968 692102
rect 44916 692038 44968 692044
rect 46216 669390 46244 767314
rect 46204 669384 46256 669390
rect 46204 669326 46256 669332
rect 44824 626612 44876 626618
rect 44824 626554 44876 626560
rect 44456 618316 44508 618322
rect 44456 618258 44508 618264
rect 44824 610020 44876 610026
rect 44824 609962 44876 609968
rect 44364 601520 44416 601526
rect 44364 601462 44416 601468
rect 44546 599312 44602 599321
rect 44546 599247 44602 599256
rect 44270 598088 44326 598097
rect 44270 598023 44326 598032
rect 44362 595640 44418 595649
rect 44362 595575 44418 595584
rect 44376 578270 44404 595575
rect 44454 593192 44510 593201
rect 44454 593127 44510 593136
rect 44468 579698 44496 593127
rect 44456 579692 44508 579698
rect 44456 579634 44508 579640
rect 44364 578264 44416 578270
rect 44364 578206 44416 578212
rect 44178 557288 44234 557297
rect 44178 557223 44234 557232
rect 44560 556481 44588 599247
rect 44546 556472 44602 556481
rect 44546 556407 44602 556416
rect 44178 555248 44234 555257
rect 44178 555183 44234 555192
rect 44192 428097 44220 555183
rect 44638 554432 44694 554441
rect 44638 554367 44694 554376
rect 44362 551576 44418 551585
rect 44362 551511 44418 551520
rect 44376 528630 44404 551511
rect 44546 550352 44602 550361
rect 44546 550287 44602 550296
rect 44454 548720 44510 548729
rect 44454 548655 44510 548664
rect 44468 536858 44496 548655
rect 44560 538286 44588 550287
rect 44548 538280 44600 538286
rect 44548 538222 44600 538228
rect 44456 536852 44508 536858
rect 44456 536794 44508 536800
rect 44364 528624 44416 528630
rect 44364 528566 44416 528572
rect 44362 429312 44418 429321
rect 44362 429247 44418 429256
rect 44270 428496 44326 428505
rect 44270 428431 44326 428440
rect 44178 428088 44234 428097
rect 44178 428023 44234 428032
rect 44284 427938 44312 428431
rect 44192 427910 44312 427938
rect 43536 401668 43588 401674
rect 43536 401610 43588 401616
rect 43548 281110 43576 401610
rect 43628 389224 43680 389230
rect 43628 389166 43680 389172
rect 43640 300529 43668 389166
rect 44192 385665 44220 427910
rect 44376 427814 44404 429247
rect 44284 427786 44404 427814
rect 44284 387802 44312 427786
rect 44652 427281 44680 554367
rect 44836 539646 44864 609962
rect 46204 597576 46256 597582
rect 46204 597518 46256 597524
rect 46216 558346 46244 597518
rect 46204 558340 46256 558346
rect 46204 558282 46256 558288
rect 44824 539640 44876 539646
rect 44824 539582 44876 539588
rect 44916 440292 44968 440298
rect 44916 440234 44968 440240
rect 44638 427272 44694 427281
rect 44638 427207 44694 427216
rect 44362 423192 44418 423201
rect 44362 423127 44418 423136
rect 44376 402966 44404 423127
rect 44454 421560 44510 421569
rect 44454 421495 44510 421504
rect 44468 406842 44496 421495
rect 44824 419484 44876 419490
rect 44824 419426 44876 419432
rect 44456 406836 44508 406842
rect 44456 406778 44508 406784
rect 44364 402960 44416 402966
rect 44364 402902 44416 402908
rect 44272 387796 44324 387802
rect 44272 387738 44324 387744
rect 44270 386064 44326 386073
rect 44270 385999 44326 386008
rect 44178 385656 44234 385665
rect 44178 385591 44234 385600
rect 44178 384432 44234 384441
rect 44178 384367 44234 384376
rect 44192 341737 44220 384367
rect 44284 343369 44312 385999
rect 44638 385248 44694 385257
rect 44638 385183 44694 385192
rect 44454 380760 44510 380769
rect 44454 380695 44510 380704
rect 44468 356046 44496 380695
rect 44546 379128 44602 379137
rect 44546 379063 44602 379072
rect 44560 364342 44588 379063
rect 44548 364336 44600 364342
rect 44548 364278 44600 364284
rect 44456 356040 44508 356046
rect 44456 355982 44508 355988
rect 44270 343360 44326 343369
rect 44270 343295 44326 343304
rect 44362 342952 44418 342961
rect 44362 342887 44418 342896
rect 44270 342136 44326 342145
rect 44270 342071 44326 342080
rect 44178 341728 44234 341737
rect 44178 341663 44234 341672
rect 44284 341578 44312 342071
rect 44192 341550 44312 341578
rect 43720 322992 43772 322998
rect 43720 322934 43772 322940
rect 43626 300520 43682 300529
rect 43626 300455 43682 300464
rect 43628 298172 43680 298178
rect 43628 298114 43680 298120
rect 43536 281104 43588 281110
rect 43536 281046 43588 281052
rect 43444 278180 43496 278186
rect 43444 278122 43496 278128
rect 43074 256048 43130 256057
rect 43074 255983 43130 255992
rect 43074 255640 43130 255649
rect 43074 255575 43130 255584
rect 42982 250336 43038 250345
rect 42982 250271 43038 250280
rect 42996 230382 43024 250271
rect 42984 230376 43036 230382
rect 42984 230318 43036 230324
rect 42890 213752 42946 213761
rect 42890 213687 42946 213696
rect 43088 212945 43116 255575
rect 43166 241632 43222 241641
rect 43166 241567 43222 241576
rect 43180 238814 43208 241567
rect 43168 238808 43220 238814
rect 43168 238750 43220 238756
rect 43640 214606 43668 298114
rect 43732 258058 43760 322934
rect 44192 299305 44220 341550
rect 44376 341442 44404 342887
rect 44652 342553 44680 385183
rect 44638 342544 44694 342553
rect 44638 342479 44694 342488
rect 44284 341414 44404 341442
rect 44284 300121 44312 341414
rect 44362 341320 44418 341329
rect 44362 341255 44418 341264
rect 44270 300112 44326 300121
rect 44270 300047 44326 300056
rect 44178 299296 44234 299305
rect 44178 299231 44234 299240
rect 44376 298489 44404 341255
rect 44454 336832 44510 336841
rect 44454 336767 44510 336776
rect 44468 316742 44496 336767
rect 44546 335200 44602 335209
rect 44546 335135 44602 335144
rect 44560 320006 44588 335135
rect 44548 320000 44600 320006
rect 44548 319942 44600 319948
rect 44456 316736 44508 316742
rect 44456 316678 44508 316684
rect 44730 299704 44786 299713
rect 44730 299639 44786 299648
rect 44362 298480 44418 298489
rect 44362 298415 44418 298424
rect 44270 298072 44326 298081
rect 44270 298007 44326 298016
rect 44178 291544 44234 291553
rect 44178 291479 44234 291488
rect 43994 291136 44050 291145
rect 43994 291071 44050 291080
rect 43810 290728 43866 290737
rect 43810 290663 43866 290672
rect 43720 258052 43772 258058
rect 43720 257994 43772 258000
rect 43824 231130 43852 290663
rect 44008 264246 44036 291071
rect 44192 278662 44220 291479
rect 44180 278656 44232 278662
rect 44180 278598 44232 278604
rect 43996 264240 44048 264246
rect 43996 264182 44048 264188
rect 44284 255241 44312 298007
rect 44638 297256 44694 297265
rect 44638 297191 44694 297200
rect 44454 293584 44510 293593
rect 44454 293519 44510 293528
rect 44468 273358 44496 293519
rect 44546 292360 44602 292369
rect 44546 292295 44602 292304
rect 44560 274310 44588 292295
rect 44548 274304 44600 274310
rect 44548 274246 44600 274252
rect 44456 273352 44508 273358
rect 44456 273294 44508 273300
rect 44270 255232 44326 255241
rect 44270 255167 44326 255176
rect 44546 254824 44602 254833
rect 44546 254759 44602 254768
rect 44270 254008 44326 254017
rect 44270 253943 44326 253952
rect 43812 231124 43864 231130
rect 43812 231066 43864 231072
rect 43628 214600 43680 214606
rect 43628 214542 43680 214548
rect 43074 212936 43130 212945
rect 43074 212871 43130 212880
rect 42798 212528 42854 212537
rect 42798 212463 42854 212472
rect 41786 211712 41842 211721
rect 41786 211647 41842 211656
rect 44284 211313 44312 253943
rect 44362 251152 44418 251161
rect 44362 251087 44418 251096
rect 44376 226710 44404 251087
rect 44454 248704 44510 248713
rect 44454 248639 44510 248648
rect 44468 234054 44496 248639
rect 44560 248414 44588 254759
rect 44652 254425 44680 297191
rect 44744 257922 44772 299639
rect 44836 278050 44864 419426
rect 44928 344486 44956 440234
rect 46204 349172 46256 349178
rect 46204 349114 46256 349120
rect 44916 344480 44968 344486
rect 44916 344422 44968 344428
rect 44916 336796 44968 336802
rect 44916 336738 44968 336744
rect 44824 278044 44876 278050
rect 44824 277986 44876 277992
rect 44928 258126 44956 336738
rect 45006 289912 45062 289921
rect 45006 289847 45062 289856
rect 44916 258120 44968 258126
rect 44916 258062 44968 258068
rect 44732 257916 44784 257922
rect 44732 257858 44784 257864
rect 44638 254416 44694 254425
rect 44638 254351 44694 254360
rect 44560 248386 44680 248414
rect 44546 248296 44602 248305
rect 44546 248231 44602 248240
rect 44560 235414 44588 248231
rect 44548 235408 44600 235414
rect 44548 235350 44600 235356
rect 44456 234048 44508 234054
rect 44456 233990 44508 233996
rect 44364 226704 44416 226710
rect 44364 226646 44416 226652
rect 44652 212129 44680 248386
rect 45020 218754 45048 289847
rect 46216 257786 46244 349114
rect 46296 284368 46348 284374
rect 46296 284310 46348 284316
rect 46204 257780 46256 257786
rect 46204 257722 46256 257728
rect 45008 218748 45060 218754
rect 45008 218690 45060 218696
rect 46308 217326 46336 284310
rect 47596 218890 47624 932146
rect 62118 923808 62174 923817
rect 62118 923743 62174 923752
rect 62132 923302 62160 923743
rect 47676 923296 47728 923302
rect 47676 923238 47728 923244
rect 62120 923296 62172 923302
rect 62120 923238 62172 923244
rect 47688 799066 47716 923238
rect 62118 910752 62174 910761
rect 62118 910687 62174 910696
rect 62132 909498 62160 910687
rect 54484 909492 54536 909498
rect 54484 909434 54536 909440
rect 62120 909492 62172 909498
rect 62120 909434 62172 909440
rect 51724 897048 51776 897054
rect 51724 896990 51776 896996
rect 48964 884672 49016 884678
rect 48964 884614 49016 884620
rect 48976 817562 49004 884614
rect 50344 832176 50396 832182
rect 50344 832118 50396 832124
rect 48964 817556 49016 817562
rect 48964 817498 49016 817504
rect 49056 805996 49108 806002
rect 49056 805938 49108 805944
rect 47676 799060 47728 799066
rect 47676 799002 47728 799008
rect 48964 761796 49016 761802
rect 48964 761738 49016 761744
rect 47676 727320 47728 727326
rect 47676 727262 47728 727268
rect 47688 687954 47716 727262
rect 47676 687948 47728 687954
rect 47676 687890 47728 687896
rect 47676 674892 47728 674898
rect 47676 674834 47728 674840
rect 47688 644638 47716 674834
rect 47676 644632 47728 644638
rect 47676 644574 47728 644580
rect 47676 636268 47728 636274
rect 47676 636210 47728 636216
rect 47688 601730 47716 636210
rect 47676 601724 47728 601730
rect 47676 601666 47728 601672
rect 47768 583772 47820 583778
rect 47768 583714 47820 583720
rect 47780 558210 47808 583714
rect 47768 558204 47820 558210
rect 47768 558146 47820 558152
rect 47676 557592 47728 557598
rect 47676 557534 47728 557540
rect 47688 410718 47716 557534
rect 47676 410712 47728 410718
rect 47676 410654 47728 410660
rect 47676 375420 47728 375426
rect 47676 375362 47728 375368
rect 47688 300966 47716 375362
rect 47676 300960 47728 300966
rect 47676 300902 47728 300908
rect 48976 231402 49004 761738
rect 49068 731270 49096 805938
rect 50356 773945 50384 832118
rect 51736 817426 51764 896990
rect 53104 844620 53156 844626
rect 53104 844562 53156 844568
rect 51724 817420 51776 817426
rect 51724 817362 51776 817368
rect 51724 779748 51776 779754
rect 51724 779690 51776 779696
rect 50342 773936 50398 773945
rect 50342 773871 50398 773880
rect 50436 741124 50488 741130
rect 50436 741066 50488 741072
rect 49056 731264 49108 731270
rect 49056 731206 49108 731212
rect 50344 719704 50396 719710
rect 50344 719646 50396 719652
rect 49056 688696 49108 688702
rect 49056 688638 49108 688644
rect 49068 644570 49096 688638
rect 49056 644564 49108 644570
rect 49056 644506 49108 644512
rect 49056 506524 49108 506530
rect 49056 506466 49108 506472
rect 49068 364274 49096 506466
rect 49056 364268 49108 364274
rect 49056 364210 49108 364216
rect 49056 333260 49108 333266
rect 49056 333202 49108 333208
rect 48964 231396 49016 231402
rect 48964 231338 49016 231344
rect 49068 231198 49096 333202
rect 50356 231470 50384 719646
rect 50448 687818 50476 741066
rect 51736 731134 51764 779690
rect 53116 774246 53144 844562
rect 54496 816921 54524 909434
rect 62118 897832 62174 897841
rect 62118 897767 62174 897776
rect 62132 897054 62160 897767
rect 62120 897048 62172 897054
rect 62120 896990 62172 896996
rect 62118 884776 62174 884785
rect 62118 884711 62174 884720
rect 62132 884678 62160 884711
rect 62120 884672 62172 884678
rect 62120 884614 62172 884620
rect 62118 871720 62174 871729
rect 62118 871655 62174 871664
rect 62132 870874 62160 871655
rect 62120 870868 62172 870874
rect 62120 870810 62172 870816
rect 62118 858664 62174 858673
rect 62118 858599 62174 858608
rect 62132 858430 62160 858599
rect 62120 858424 62172 858430
rect 62120 858366 62172 858372
rect 62118 845608 62174 845617
rect 62118 845543 62174 845552
rect 62132 844626 62160 845543
rect 62120 844620 62172 844626
rect 62120 844562 62172 844568
rect 62118 832552 62174 832561
rect 62118 832487 62174 832496
rect 62132 832182 62160 832487
rect 62120 832176 62172 832182
rect 62120 832118 62172 832124
rect 62118 819496 62174 819505
rect 62118 819431 62174 819440
rect 62132 818378 62160 819431
rect 62120 818372 62172 818378
rect 62120 818314 62172 818320
rect 54482 816912 54538 816921
rect 54482 816847 54538 816856
rect 62118 806576 62174 806585
rect 62118 806511 62174 806520
rect 62132 806002 62160 806511
rect 62120 805996 62172 806002
rect 62120 805938 62172 805944
rect 62118 793656 62174 793665
rect 62118 793591 62174 793600
rect 62132 793558 62160 793591
rect 54484 793552 54536 793558
rect 54484 793494 54536 793500
rect 62120 793552 62172 793558
rect 62120 793494 62172 793500
rect 53104 774240 53156 774246
rect 53104 774182 53156 774188
rect 51724 731128 51776 731134
rect 51724 731070 51776 731076
rect 54496 730998 54524 793494
rect 62118 780464 62174 780473
rect 62118 780399 62174 780408
rect 62132 779754 62160 780399
rect 62120 779748 62172 779754
rect 62120 779690 62172 779696
rect 62118 767408 62174 767417
rect 62118 767343 62120 767352
rect 62172 767343 62174 767352
rect 62120 767314 62172 767320
rect 62118 754352 62174 754361
rect 62118 754287 62174 754296
rect 62132 753574 62160 754287
rect 62120 753568 62172 753574
rect 62120 753510 62172 753516
rect 62118 741296 62174 741305
rect 62118 741231 62174 741240
rect 62132 741130 62160 741231
rect 62120 741124 62172 741130
rect 62120 741066 62172 741072
rect 54484 730992 54536 730998
rect 54484 730934 54536 730940
rect 62118 728240 62174 728249
rect 62118 728175 62174 728184
rect 62132 727326 62160 728175
rect 62120 727320 62172 727326
rect 62120 727262 62172 727268
rect 62118 715320 62174 715329
rect 62118 715255 62174 715264
rect 62132 714882 62160 715255
rect 62120 714876 62172 714882
rect 62120 714818 62172 714824
rect 62762 702264 62818 702273
rect 62762 702199 62818 702208
rect 62118 689208 62174 689217
rect 62118 689143 62174 689152
rect 62132 688702 62160 689143
rect 62120 688696 62172 688702
rect 62120 688638 62172 688644
rect 50436 687812 50488 687818
rect 50436 687754 50488 687760
rect 51724 676864 51776 676870
rect 51724 676806 51776 676812
rect 50528 480276 50580 480282
rect 50528 480218 50580 480224
rect 50436 454096 50488 454102
rect 50436 454038 50488 454044
rect 50448 321570 50476 454038
rect 50540 387666 50568 480218
rect 50528 387660 50580 387666
rect 50528 387602 50580 387608
rect 50436 321564 50488 321570
rect 50436 321506 50488 321512
rect 50344 231464 50396 231470
rect 50344 231406 50396 231412
rect 51736 231266 51764 676806
rect 62118 676152 62174 676161
rect 62118 676087 62174 676096
rect 62132 674898 62160 676087
rect 62120 674892 62172 674898
rect 62120 674834 62172 674840
rect 62118 663096 62174 663105
rect 62118 663031 62174 663040
rect 62132 662454 62160 663031
rect 62120 662448 62172 662454
rect 62120 662390 62172 662396
rect 54484 650072 54536 650078
rect 62120 650072 62172 650078
rect 54484 650014 54536 650020
rect 62118 650040 62120 650049
rect 62172 650040 62174 650049
rect 53102 633448 53158 633457
rect 53102 633383 53158 633392
rect 51816 532772 51868 532778
rect 51816 532714 51868 532720
rect 51828 430642 51856 532714
rect 51816 430636 51868 430642
rect 51816 430578 51868 430584
rect 51816 415472 51868 415478
rect 51816 415414 51868 415420
rect 51828 344350 51856 415414
rect 51908 362976 51960 362982
rect 51908 362918 51960 362924
rect 51816 344344 51868 344350
rect 51816 344286 51868 344292
rect 51920 307086 51948 362918
rect 51908 307080 51960 307086
rect 51908 307022 51960 307028
rect 51724 231260 51776 231266
rect 51724 231202 51776 231208
rect 49056 231192 49108 231198
rect 49056 231134 49108 231140
rect 52736 225616 52788 225622
rect 52736 225558 52788 225564
rect 52460 220788 52512 220794
rect 52460 220730 52512 220736
rect 52472 219434 52500 220730
rect 52288 219406 52500 219434
rect 47584 218884 47636 218890
rect 47584 218826 47636 218832
rect 46296 217320 46348 217326
rect 46296 217262 46348 217268
rect 52184 217320 52236 217326
rect 52184 217262 52236 217268
rect 48964 214396 49016 214402
rect 48964 214338 49016 214344
rect 46572 214328 46624 214334
rect 46572 214270 46624 214276
rect 46584 213353 46612 214270
rect 46570 213344 46626 213353
rect 46570 213279 46626 213288
rect 44638 212120 44694 212129
rect 44638 212055 44694 212064
rect 44270 211304 44326 211313
rect 44270 211239 44326 211248
rect 41326 211032 41382 211041
rect 41326 210967 41382 210976
rect 42798 209264 42854 209273
rect 42798 209199 42854 209208
rect 40866 204912 40922 204921
rect 40866 204847 40922 204856
rect 40682 204504 40738 204513
rect 40682 204439 40738 204448
rect 39302 197704 39358 197713
rect 39302 197639 39358 197648
rect 41878 197160 41934 197169
rect 41878 197095 41934 197104
rect 41892 196656 41920 197095
rect 41786 195256 41842 195265
rect 41786 195191 41842 195200
rect 41800 194820 41828 195191
rect 42064 193180 42116 193186
rect 42064 193122 42116 193128
rect 42076 192984 42104 193122
rect 42064 191684 42116 191690
rect 42064 191626 42116 191632
rect 42076 191148 42104 191626
rect 42168 191622 42196 191760
rect 42156 191616 42208 191622
rect 42156 191558 42208 191564
rect 42156 190868 42208 190874
rect 42156 190810 42208 190816
rect 42168 190468 42196 190810
rect 41786 190224 41842 190233
rect 41786 190159 41842 190168
rect 41800 189924 41828 190159
rect 42156 187672 42208 187678
rect 42156 187614 42208 187620
rect 42168 187445 42196 187614
rect 41786 187368 41842 187377
rect 41786 187303 41842 187312
rect 41800 186796 41828 187303
rect 42064 186312 42116 186318
rect 42064 186254 42116 186260
rect 42076 186184 42104 186254
rect 42812 185910 42840 209199
rect 44178 208040 44234 208049
rect 44178 207975 44234 207984
rect 42890 207632 42946 207641
rect 42890 207567 42946 207576
rect 42904 186318 42932 207567
rect 42982 206408 43038 206417
rect 42982 206343 43038 206352
rect 42996 191690 43024 206343
rect 43074 205592 43130 205601
rect 43074 205527 43130 205536
rect 42984 191684 43036 191690
rect 42984 191626 43036 191632
rect 43088 190874 43116 205527
rect 43076 190868 43128 190874
rect 43076 190810 43128 190816
rect 42892 186312 42944 186318
rect 42892 186254 42944 186260
rect 42156 185904 42208 185910
rect 42156 185846 42208 185852
rect 42800 185904 42852 185910
rect 42800 185846 42852 185852
rect 42168 185605 42196 185846
rect 41786 184104 41842 184113
rect 41786 184039 41842 184048
rect 41800 183765 41828 184039
rect 44192 183462 44220 207975
rect 44454 206816 44510 206825
rect 44454 206751 44510 206760
rect 44270 206000 44326 206009
rect 44270 205935 44326 205944
rect 44284 187678 44312 205935
rect 44362 205184 44418 205193
rect 44362 205119 44418 205128
rect 44376 191622 44404 205119
rect 44468 193186 44496 206751
rect 48976 202910 49004 214338
rect 48964 202904 49016 202910
rect 48964 202846 49016 202852
rect 44456 193180 44508 193186
rect 44456 193122 44508 193128
rect 44364 191616 44416 191622
rect 44364 191558 44416 191564
rect 44272 187672 44324 187678
rect 44272 187614 44324 187620
rect 42156 183456 42208 183462
rect 42156 183398 42208 183404
rect 44180 183456 44232 183462
rect 44180 183398 44232 183404
rect 42168 183124 42196 183398
rect 41786 183016 41842 183025
rect 41786 182951 41842 182960
rect 41800 182477 41828 182951
rect 52196 51746 52224 217262
rect 52288 53174 52316 219406
rect 52748 217410 52776 225558
rect 53116 218385 53144 633383
rect 54496 601390 54524 650014
rect 62118 649975 62174 649984
rect 62776 643521 62804 702199
rect 62762 643512 62818 643521
rect 62762 643447 62818 643456
rect 62118 637120 62174 637129
rect 62118 637055 62174 637064
rect 62132 636274 62160 637055
rect 62120 636268 62172 636274
rect 62120 636210 62172 636216
rect 62118 624064 62174 624073
rect 62118 623999 62174 624008
rect 62132 623830 62160 623999
rect 62120 623824 62172 623830
rect 62120 623766 62172 623772
rect 62118 611008 62174 611017
rect 62118 610943 62174 610952
rect 62132 610026 62160 610943
rect 62120 610020 62172 610026
rect 62120 609962 62172 609968
rect 54484 601384 54536 601390
rect 54484 601326 54536 601332
rect 62118 597952 62174 597961
rect 62118 597887 62174 597896
rect 62132 597582 62160 597887
rect 62120 597576 62172 597582
rect 62120 597518 62172 597524
rect 54484 589960 54536 589966
rect 54484 589902 54536 589908
rect 53196 492720 53248 492726
rect 53196 492662 53248 492668
rect 53208 387530 53236 492662
rect 53196 387524 53248 387530
rect 53196 387466 53248 387472
rect 53196 376032 53248 376038
rect 53196 375974 53248 375980
rect 53208 278118 53236 375974
rect 53196 278112 53248 278118
rect 53196 278054 53248 278060
rect 54496 231334 54524 589902
rect 62118 584896 62174 584905
rect 62118 584831 62174 584840
rect 62132 583778 62160 584831
rect 62120 583772 62172 583778
rect 62120 583714 62172 583720
rect 62118 571840 62174 571849
rect 62118 571775 62174 571784
rect 62132 571402 62160 571775
rect 62120 571396 62172 571402
rect 62120 571338 62172 571344
rect 62118 558784 62174 558793
rect 62118 558719 62174 558728
rect 62132 557598 62160 558719
rect 62120 557592 62172 557598
rect 62120 557534 62172 557540
rect 55864 547188 55916 547194
rect 55864 547130 55916 547136
rect 54576 427848 54628 427854
rect 54576 427790 54628 427796
rect 54588 344214 54616 427790
rect 54576 344208 54628 344214
rect 54576 344150 54628 344156
rect 54484 231328 54536 231334
rect 54484 231270 54536 231276
rect 54392 228472 54444 228478
rect 54392 228414 54444 228420
rect 53656 228404 53708 228410
rect 53656 228346 53708 228352
rect 53102 218376 53158 218385
rect 53102 218311 53158 218320
rect 53668 217410 53696 228346
rect 54404 217410 54432 228414
rect 55034 222864 55090 222873
rect 55034 222799 55090 222808
rect 55048 217410 55076 222799
rect 55876 218822 55904 547130
rect 62762 545864 62818 545873
rect 62762 545799 62818 545808
rect 62118 532808 62174 532817
rect 62118 532743 62120 532752
rect 62172 532743 62174 532752
rect 62120 532714 62172 532720
rect 62118 519752 62174 519761
rect 62118 519687 62174 519696
rect 62132 518974 62160 519687
rect 62120 518968 62172 518974
rect 62120 518910 62172 518916
rect 62118 506696 62174 506705
rect 62118 506631 62174 506640
rect 62132 506530 62160 506631
rect 62120 506524 62172 506530
rect 62120 506466 62172 506472
rect 62776 497486 62804 545799
rect 62764 497480 62816 497486
rect 62764 497422 62816 497428
rect 62118 493640 62174 493649
rect 62118 493575 62174 493584
rect 62132 492726 62160 493575
rect 62120 492720 62172 492726
rect 62120 492662 62172 492668
rect 62118 480584 62174 480593
rect 62118 480519 62174 480528
rect 62132 480282 62160 480519
rect 62120 480276 62172 480282
rect 62120 480218 62172 480224
rect 62118 467528 62174 467537
rect 62118 467463 62174 467472
rect 62132 466478 62160 467463
rect 55956 466472 56008 466478
rect 55956 466414 56008 466420
rect 62120 466472 62172 466478
rect 62120 466414 62172 466420
rect 55968 387394 55996 466414
rect 62118 454608 62174 454617
rect 62118 454543 62174 454552
rect 62132 454102 62160 454543
rect 62120 454096 62172 454102
rect 62120 454038 62172 454044
rect 62118 441552 62174 441561
rect 62118 441487 62174 441496
rect 62132 440298 62160 441487
rect 62120 440292 62172 440298
rect 62120 440234 62172 440240
rect 62118 428496 62174 428505
rect 62118 428431 62174 428440
rect 62132 427854 62160 428431
rect 62120 427848 62172 427854
rect 62120 427790 62172 427796
rect 62120 415472 62172 415478
rect 62118 415440 62120 415449
rect 62172 415440 62174 415449
rect 62118 415375 62174 415384
rect 62118 402384 62174 402393
rect 62118 402319 62174 402328
rect 62132 401674 62160 402319
rect 62120 401668 62172 401674
rect 62120 401610 62172 401616
rect 62118 389328 62174 389337
rect 62118 389263 62174 389272
rect 62132 389230 62160 389263
rect 62120 389224 62172 389230
rect 62120 389166 62172 389172
rect 55956 387388 56008 387394
rect 55956 387330 56008 387336
rect 62118 376272 62174 376281
rect 62118 376207 62174 376216
rect 62132 375426 62160 376207
rect 62120 375420 62172 375426
rect 62120 375362 62172 375368
rect 62118 363352 62174 363361
rect 62118 363287 62174 363296
rect 62132 362982 62160 363287
rect 62120 362976 62172 362982
rect 62120 362918 62172 362924
rect 62118 350296 62174 350305
rect 62118 350231 62174 350240
rect 62132 349178 62160 350231
rect 62120 349172 62172 349178
rect 62120 349114 62172 349120
rect 62118 337240 62174 337249
rect 62118 337175 62174 337184
rect 62132 336802 62160 337175
rect 62120 336796 62172 336802
rect 62120 336738 62172 336744
rect 62118 324184 62174 324193
rect 62118 324119 62174 324128
rect 62132 322998 62160 324119
rect 62120 322992 62172 322998
rect 62120 322934 62172 322940
rect 62118 311128 62174 311137
rect 62118 311063 62174 311072
rect 62132 310554 62160 311063
rect 55956 310548 56008 310554
rect 55956 310490 56008 310496
rect 62120 310548 62172 310554
rect 62120 310490 62172 310496
rect 55968 218958 55996 310490
rect 62118 298208 62174 298217
rect 62118 298143 62120 298152
rect 62172 298143 62174 298152
rect 62120 298114 62172 298120
rect 62118 285152 62174 285161
rect 62118 285087 62174 285096
rect 62132 284374 62160 285087
rect 62120 284368 62172 284374
rect 62120 284310 62172 284316
rect 647252 278310 647542 278338
rect 65918 277766 66208 277794
rect 66180 268394 66208 277766
rect 67008 275398 67036 277780
rect 66996 275392 67048 275398
rect 66996 275334 67048 275340
rect 68204 271182 68232 277780
rect 68192 271176 68244 271182
rect 68192 271118 68244 271124
rect 69400 268462 69428 277780
rect 70596 274718 70624 277780
rect 71792 275330 71820 277780
rect 71780 275324 71832 275330
rect 71780 275266 71832 275272
rect 70584 274712 70636 274718
rect 70584 274654 70636 274660
rect 72988 272542 73016 277780
rect 74092 274922 74120 277780
rect 75302 277766 75868 277794
rect 76498 277766 77156 277794
rect 74080 274916 74132 274922
rect 74080 274858 74132 274864
rect 73804 274712 73856 274718
rect 73804 274654 73856 274660
rect 72976 272536 73028 272542
rect 72976 272478 73028 272484
rect 69388 268456 69440 268462
rect 69388 268398 69440 268404
rect 66168 268388 66220 268394
rect 66168 268330 66220 268336
rect 73816 267034 73844 274654
rect 75840 268530 75868 277766
rect 77128 270026 77156 277766
rect 77208 274916 77260 274922
rect 77208 274858 77260 274864
rect 77220 272610 77248 274858
rect 77208 272604 77260 272610
rect 77208 272546 77260 272552
rect 77116 270020 77168 270026
rect 77116 269962 77168 269968
rect 77680 268598 77708 277780
rect 78876 272746 78904 277780
rect 78864 272740 78916 272746
rect 78864 272682 78916 272688
rect 80072 268666 80100 277780
rect 81268 275466 81296 277780
rect 82386 277766 82768 277794
rect 81256 275460 81308 275466
rect 81256 275402 81308 275408
rect 82740 268734 82768 277766
rect 83568 271590 83596 277780
rect 84764 272678 84792 277780
rect 84752 272672 84804 272678
rect 84752 272614 84804 272620
rect 83556 271584 83608 271590
rect 83556 271526 83608 271532
rect 85960 269890 85988 277780
rect 85948 269884 86000 269890
rect 85948 269826 86000 269832
rect 87156 268802 87184 277780
rect 88352 274990 88380 277780
rect 88340 274984 88392 274990
rect 88340 274926 88392 274932
rect 89548 273970 89576 277780
rect 90652 275534 90680 277780
rect 91862 277766 92428 277794
rect 90640 275528 90692 275534
rect 90640 275470 90692 275476
rect 90364 274984 90416 274990
rect 90364 274926 90416 274932
rect 89536 273964 89588 273970
rect 89536 273906 89588 273912
rect 87144 268796 87196 268802
rect 87144 268738 87196 268744
rect 82728 268728 82780 268734
rect 82728 268670 82780 268676
rect 80060 268660 80112 268666
rect 80060 268602 80112 268608
rect 77668 268592 77720 268598
rect 77668 268534 77720 268540
rect 75828 268524 75880 268530
rect 75828 268466 75880 268472
rect 90376 267102 90404 274926
rect 92400 268870 92428 277766
rect 93044 275602 93072 277780
rect 93032 275596 93084 275602
rect 93032 275538 93084 275544
rect 94240 272814 94268 277780
rect 94228 272808 94280 272814
rect 94228 272750 94280 272756
rect 95436 268938 95464 277780
rect 96632 274854 96660 277780
rect 96620 274848 96672 274854
rect 96620 274790 96672 274796
rect 97736 274038 97764 277780
rect 98946 277766 99328 277794
rect 97724 274032 97776 274038
rect 97724 273974 97776 273980
rect 99300 269006 99328 277766
rect 100128 275670 100156 277780
rect 100116 275664 100168 275670
rect 100116 275606 100168 275612
rect 100024 274848 100076 274854
rect 100024 274790 100076 274796
rect 99288 269000 99340 269006
rect 99288 268942 99340 268948
rect 95424 268932 95476 268938
rect 95424 268874 95476 268880
rect 92388 268864 92440 268870
rect 92388 268806 92440 268812
rect 100036 267170 100064 274790
rect 101324 272882 101352 277780
rect 101312 272876 101364 272882
rect 101312 272818 101364 272824
rect 102520 269074 102548 277780
rect 103716 274718 103744 277780
rect 103704 274712 103756 274718
rect 103704 274654 103756 274660
rect 104912 271250 104940 277780
rect 106030 277766 106228 277794
rect 104900 271244 104952 271250
rect 104900 271186 104952 271192
rect 102508 269068 102560 269074
rect 102508 269010 102560 269016
rect 106200 268326 106228 277766
rect 107212 275738 107240 277780
rect 108422 277766 108988 277794
rect 109618 277766 110368 277794
rect 107200 275732 107252 275738
rect 107200 275674 107252 275680
rect 106924 274712 106976 274718
rect 106924 274654 106976 274660
rect 106188 268320 106240 268326
rect 106188 268262 106240 268268
rect 106936 267238 106964 274654
rect 108960 269822 108988 277766
rect 108948 269816 109000 269822
rect 108948 269758 109000 269764
rect 110340 268258 110368 277766
rect 110800 270366 110828 277780
rect 111996 274106 112024 277780
rect 113192 274174 113220 277780
rect 113180 274168 113232 274174
rect 113180 274110 113232 274116
rect 111984 274100 112036 274106
rect 111984 274042 112036 274048
rect 114296 271454 114324 277780
rect 115506 277766 115888 277794
rect 114284 271448 114336 271454
rect 114284 271390 114336 271396
rect 110788 270360 110840 270366
rect 110788 270302 110840 270308
rect 110328 268252 110380 268258
rect 110328 268194 110380 268200
rect 115860 268190 115888 277766
rect 116688 271318 116716 277780
rect 117884 272950 117912 277780
rect 117872 272944 117924 272950
rect 117872 272886 117924 272892
rect 116676 271312 116728 271318
rect 116676 271254 116728 271260
rect 119080 269890 119108 277780
rect 120276 273018 120304 277780
rect 121380 274378 121408 277780
rect 122590 277766 122788 277794
rect 121368 274372 121420 274378
rect 121368 274314 121420 274320
rect 120264 273012 120316 273018
rect 120264 272954 120316 272960
rect 122760 269958 122788 277766
rect 123772 274242 123800 277780
rect 124982 277766 125548 277794
rect 126178 277766 126928 277794
rect 123760 274236 123812 274242
rect 123760 274178 123812 274184
rect 125520 270026 125548 277766
rect 126900 270094 126928 277766
rect 127360 271386 127388 277780
rect 128556 274582 128584 277780
rect 129660 277394 129688 277780
rect 130870 277766 131068 277794
rect 132066 277766 132448 277794
rect 133262 277766 133828 277794
rect 134458 277766 135208 277794
rect 129568 277366 129688 277394
rect 128544 274576 128596 274582
rect 128544 274518 128596 274524
rect 127348 271380 127400 271386
rect 127348 271322 127400 271328
rect 129568 270162 129596 277366
rect 129556 270156 129608 270162
rect 129556 270098 129608 270104
rect 126888 270088 126940 270094
rect 126888 270030 126940 270036
rect 124220 270020 124272 270026
rect 124220 269962 124272 269968
rect 125508 270020 125560 270026
rect 125508 269962 125560 269968
rect 122748 269952 122800 269958
rect 122748 269894 122800 269900
rect 116492 269884 116544 269890
rect 116492 269826 116544 269832
rect 119068 269884 119120 269890
rect 119068 269826 119120 269832
rect 115848 268184 115900 268190
rect 115848 268126 115900 268132
rect 116504 267374 116532 269826
rect 124232 267578 124260 269962
rect 131040 268122 131068 277766
rect 131028 268116 131080 268122
rect 131028 268058 131080 268064
rect 124220 267572 124272 267578
rect 124220 267514 124272 267520
rect 116492 267368 116544 267374
rect 116492 267310 116544 267316
rect 132420 267306 132448 277766
rect 133800 270230 133828 277766
rect 133788 270224 133840 270230
rect 133788 270166 133840 270172
rect 135180 268054 135208 277766
rect 135640 271522 135668 277780
rect 136836 271658 136864 277780
rect 137940 274310 137968 277780
rect 139150 277766 139348 277794
rect 140346 277766 140728 277794
rect 137928 274304 137980 274310
rect 137928 274246 137980 274252
rect 136824 271652 136876 271658
rect 136824 271594 136876 271600
rect 135628 271516 135680 271522
rect 135628 271458 135680 271464
rect 135168 268048 135220 268054
rect 135168 267990 135220 267996
rect 139320 267442 139348 277766
rect 140700 270298 140728 277766
rect 141528 273086 141556 277780
rect 142724 276010 142752 277780
rect 142712 276004 142764 276010
rect 142712 275946 142764 275952
rect 141516 273080 141568 273086
rect 141516 273022 141568 273028
rect 143920 270366 143948 277780
rect 145024 271726 145052 277780
rect 145012 271720 145064 271726
rect 145012 271662 145064 271668
rect 140780 270360 140832 270366
rect 140780 270302 140832 270308
rect 143908 270360 143960 270366
rect 143908 270302 143960 270308
rect 140688 270292 140740 270298
rect 140688 270234 140740 270240
rect 140792 267714 140820 270302
rect 146220 269686 146248 277780
rect 147430 277766 147628 277794
rect 147600 270434 147628 277766
rect 148612 274446 148640 277780
rect 149822 277766 150388 277794
rect 148600 274440 148652 274446
rect 148600 274382 148652 274388
rect 147588 270428 147640 270434
rect 147588 270370 147640 270376
rect 146208 269680 146260 269686
rect 146208 269622 146260 269628
rect 140780 267708 140832 267714
rect 140780 267650 140832 267656
rect 150360 267510 150388 277766
rect 151004 274514 151032 277780
rect 150992 274508 151044 274514
rect 150992 274450 151044 274456
rect 152200 273154 152228 277780
rect 153304 275942 153332 277780
rect 153292 275936 153344 275942
rect 153292 275878 153344 275884
rect 152188 273148 152240 273154
rect 152188 273090 152240 273096
rect 154500 270502 154528 277780
rect 155696 271794 155724 277780
rect 156906 277766 157288 277794
rect 155684 271788 155736 271794
rect 155684 271730 155736 271736
rect 154488 270496 154540 270502
rect 154488 270438 154540 270444
rect 157260 267646 157288 277766
rect 158088 273222 158116 277780
rect 159284 274650 159312 277780
rect 160480 275806 160508 277780
rect 160468 275800 160520 275806
rect 160468 275742 160520 275748
rect 159272 274644 159324 274650
rect 159272 274586 159324 274592
rect 158076 273216 158128 273222
rect 158076 273158 158128 273164
rect 161584 271862 161612 277780
rect 162780 272474 162808 277780
rect 163990 277766 164188 277794
rect 162768 272468 162820 272474
rect 162768 272410 162820 272416
rect 161572 271856 161624 271862
rect 161572 271798 161624 271804
rect 157248 267640 157300 267646
rect 157248 267582 157300 267588
rect 150348 267504 150400 267510
rect 150348 267446 150400 267452
rect 139308 267436 139360 267442
rect 139308 267378 139360 267384
rect 132408 267300 132460 267306
rect 132408 267242 132460 267248
rect 106924 267232 106976 267238
rect 106924 267174 106976 267180
rect 100024 267164 100076 267170
rect 100024 267106 100076 267112
rect 90364 267096 90416 267102
rect 90364 267038 90416 267044
rect 73804 267028 73856 267034
rect 73804 266970 73856 266976
rect 164160 266966 164188 277766
rect 165172 271590 165200 277780
rect 164884 271584 164936 271590
rect 164884 271526 164936 271532
rect 165160 271584 165212 271590
rect 165160 271526 165212 271532
rect 164148 266960 164200 266966
rect 164148 266902 164200 266908
rect 164896 266762 164924 271526
rect 166368 271114 166396 277780
rect 167564 275874 167592 277780
rect 167552 275868 167604 275874
rect 167552 275810 167604 275816
rect 166356 271108 166408 271114
rect 166356 271050 166408 271056
rect 168668 271046 168696 277780
rect 169864 273834 169892 277780
rect 171060 277394 171088 277780
rect 170968 277366 171088 277394
rect 169852 273828 169904 273834
rect 169852 273770 169904 273776
rect 168656 271040 168708 271046
rect 168656 270982 168708 270988
rect 170968 266898 170996 277366
rect 172256 273902 172284 277780
rect 173466 277766 173848 277794
rect 172244 273896 172296 273902
rect 172244 273838 172296 273844
rect 173820 269618 173848 277766
rect 174648 275262 174676 277780
rect 174636 275256 174688 275262
rect 174636 275198 174688 275204
rect 175844 270978 175872 277780
rect 175832 270972 175884 270978
rect 175832 270914 175884 270920
rect 173808 269612 173860 269618
rect 173808 269554 173860 269560
rect 176948 269550 176976 277780
rect 178144 275126 178172 277780
rect 178132 275120 178184 275126
rect 178132 275062 178184 275068
rect 177580 269680 177632 269686
rect 177580 269622 177632 269628
rect 176936 269544 176988 269550
rect 176936 269486 176988 269492
rect 170956 266892 171008 266898
rect 170956 266834 171008 266840
rect 177592 266830 177620 269622
rect 179340 269618 179368 277780
rect 180550 277766 180748 277794
rect 179328 269612 179380 269618
rect 179328 269554 179380 269560
rect 180720 269550 180748 277766
rect 181168 276004 181220 276010
rect 181168 275946 181220 275952
rect 180708 269544 180760 269550
rect 180708 269486 180760 269492
rect 181180 267918 181208 275946
rect 181732 275194 181760 277780
rect 181720 275188 181772 275194
rect 181720 275130 181772 275136
rect 182928 272270 182956 277780
rect 184138 277766 184888 277794
rect 182916 272264 182968 272270
rect 182916 272206 182968 272212
rect 184860 269482 184888 277766
rect 185228 276010 185256 277780
rect 185216 276004 185268 276010
rect 185216 275946 185268 275952
rect 185584 275392 185636 275398
rect 185584 275334 185636 275340
rect 185596 273562 185624 275334
rect 185584 273556 185636 273562
rect 185584 273498 185636 273504
rect 186424 270842 186452 277780
rect 187620 272406 187648 277780
rect 188816 275398 188844 277780
rect 190026 277766 190408 277794
rect 188804 275392 188856 275398
rect 188804 275334 188856 275340
rect 187608 272400 187660 272406
rect 187608 272342 187660 272348
rect 186412 270836 186464 270842
rect 186412 270778 186464 270784
rect 184848 269476 184900 269482
rect 184848 269418 184900 269424
rect 190380 267986 190408 277766
rect 191208 272746 191236 277780
rect 191104 272740 191156 272746
rect 191104 272682 191156 272688
rect 191196 272740 191248 272746
rect 191196 272682 191248 272688
rect 190368 267980 190420 267986
rect 190368 267922 190420 267928
rect 181168 267912 181220 267918
rect 181168 267854 181220 267860
rect 177580 266824 177632 266830
rect 177580 266766 177632 266772
rect 164884 266756 164936 266762
rect 164884 266698 164936 266704
rect 191116 266490 191144 272682
rect 192312 270910 192340 277780
rect 192484 273556 192536 273562
rect 192484 273498 192536 273504
rect 192300 270904 192352 270910
rect 192300 270846 192352 270852
rect 192392 268388 192444 268394
rect 192392 268330 192444 268336
rect 191104 266484 191156 266490
rect 191104 266426 191156 266432
rect 192404 264316 192432 268330
rect 192496 264330 192524 273498
rect 193508 272338 193536 277780
rect 193864 275324 193916 275330
rect 193864 275266 193916 275272
rect 193496 272332 193548 272338
rect 193496 272274 193548 272280
rect 193220 271176 193272 271182
rect 193220 271118 193272 271124
rect 192496 264302 192786 264330
rect 193232 264316 193260 271118
rect 193680 268456 193732 268462
rect 193680 268398 193732 268404
rect 193692 264316 193720 268398
rect 193876 266422 193904 275266
rect 194704 273766 194732 277780
rect 194692 273760 194744 273766
rect 194692 273702 194744 273708
rect 194692 272604 194744 272610
rect 194692 272546 194744 272552
rect 194140 267028 194192 267034
rect 194140 266970 194192 266976
rect 193864 266416 193916 266422
rect 193864 266358 193916 266364
rect 194152 264316 194180 266970
rect 194600 266416 194652 266422
rect 194600 266358 194652 266364
rect 194612 264316 194640 266358
rect 194704 265606 194732 272546
rect 195900 272542 195928 277780
rect 195980 275120 196032 275126
rect 195980 275062 196032 275068
rect 194784 272536 194836 272542
rect 194784 272478 194836 272484
rect 195888 272536 195940 272542
rect 195888 272478 195940 272484
rect 194692 265600 194744 265606
rect 194692 265542 194744 265548
rect 194796 264330 194824 272478
rect 195428 268524 195480 268530
rect 195428 268466 195480 268472
rect 194796 264302 195086 264330
rect 195440 264316 195468 268466
rect 195992 268394 196020 275062
rect 196716 274576 196768 274582
rect 196716 274518 196768 274524
rect 196624 274372 196676 274378
rect 196624 274314 196676 274320
rect 196532 268592 196584 268598
rect 196532 268534 196584 268540
rect 195980 268388 196032 268394
rect 195980 268330 196032 268336
rect 196348 267572 196400 267578
rect 196348 267514 196400 267520
rect 195612 265600 195664 265606
rect 195612 265542 195664 265548
rect 195624 264330 195652 265542
rect 195624 264302 195914 264330
rect 196360 264316 196388 267514
rect 196544 264330 196572 268534
rect 196636 266626 196664 274314
rect 196728 267578 196756 274518
rect 197096 273698 197124 277780
rect 197820 275460 197872 275466
rect 197820 275402 197872 275408
rect 197084 273692 197136 273698
rect 197084 273634 197136 273640
rect 197268 268660 197320 268666
rect 197268 268602 197320 268608
rect 196716 267572 196768 267578
rect 196716 267514 196768 267520
rect 196624 266620 196676 266626
rect 196624 266562 196676 266568
rect 196544 264302 196834 264330
rect 197280 264316 197308 268602
rect 197728 266484 197780 266490
rect 197728 266426 197780 266432
rect 197740 264316 197768 266426
rect 197832 264330 197860 275402
rect 198292 274378 198320 277780
rect 199488 274582 199516 277780
rect 199476 274576 199528 274582
rect 199476 274518 199528 274524
rect 198280 274372 198332 274378
rect 198280 274314 198332 274320
rect 200488 273964 200540 273970
rect 200488 273906 200540 273912
rect 198924 272672 198976 272678
rect 198924 272614 198976 272620
rect 198556 268728 198608 268734
rect 198556 268670 198608 268676
rect 197832 264302 198122 264330
rect 198568 264316 198596 268670
rect 198936 264330 198964 272614
rect 200396 268796 200448 268802
rect 200396 268738 200448 268744
rect 199936 267368 199988 267374
rect 199936 267310 199988 267316
rect 199476 266756 199528 266762
rect 199476 266698 199528 266704
rect 198936 264302 199042 264330
rect 199488 264316 199516 266698
rect 199948 264316 199976 267310
rect 200408 264316 200436 268738
rect 200500 264330 200528 273906
rect 200592 271182 200620 277780
rect 201408 275596 201460 275602
rect 201408 275538 201460 275544
rect 200856 271448 200908 271454
rect 200856 271390 200908 271396
rect 200580 271176 200632 271182
rect 200580 271118 200632 271124
rect 200868 267238 200896 271390
rect 201420 268802 201448 275538
rect 201684 275528 201736 275534
rect 201684 275470 201736 275476
rect 201592 272808 201644 272814
rect 201592 272750 201644 272756
rect 201408 268796 201460 268802
rect 201408 268738 201460 268744
rect 200764 267232 200816 267238
rect 200764 267174 200816 267180
rect 200856 267232 200908 267238
rect 200856 267174 200908 267180
rect 200776 266762 200804 267174
rect 201224 267096 201276 267102
rect 201224 267038 201276 267044
rect 200764 266756 200816 266762
rect 200764 266698 200816 266704
rect 200500 264302 200790 264330
rect 201236 264316 201264 267038
rect 201604 265606 201632 272750
rect 201592 265600 201644 265606
rect 201592 265542 201644 265548
rect 201696 264316 201724 275470
rect 201788 272610 201816 277780
rect 201776 272604 201828 272610
rect 201776 272546 201828 272552
rect 202984 271454 203012 277780
rect 203616 274032 203668 274038
rect 203616 273974 203668 273980
rect 202972 271448 203024 271454
rect 202972 271390 203024 271396
rect 203524 268932 203576 268938
rect 203524 268874 203576 268880
rect 202144 268864 202196 268870
rect 202144 268806 202196 268812
rect 202156 264316 202184 268806
rect 203064 268796 203116 268802
rect 203064 268738 203116 268744
rect 202420 267028 202472 267034
rect 202420 266970 202472 266976
rect 202432 266626 202460 266970
rect 202420 266620 202472 266626
rect 202420 266562 202472 266568
rect 202236 265600 202288 265606
rect 202236 265542 202288 265548
rect 202248 264330 202276 265542
rect 202248 264302 202630 264330
rect 203076 264316 203104 268738
rect 203536 264316 203564 268874
rect 203628 264330 203656 273974
rect 204180 272814 204208 277780
rect 204904 275936 204956 275942
rect 204904 275878 204956 275884
rect 204812 272876 204864 272882
rect 204812 272818 204864 272824
rect 204168 272808 204220 272814
rect 204168 272750 204220 272756
rect 204444 269000 204496 269006
rect 204444 268942 204496 268948
rect 204352 267164 204404 267170
rect 204352 267106 204404 267112
rect 203628 264302 203918 264330
rect 204364 264316 204392 267106
rect 204456 264330 204484 268942
rect 204824 267734 204852 272818
rect 204916 268802 204944 275878
rect 205376 273970 205404 277780
rect 205824 275664 205876 275670
rect 205824 275606 205876 275612
rect 205364 273964 205416 273970
rect 205364 273906 205416 273912
rect 204904 268796 204956 268802
rect 204904 268738 204956 268744
rect 204824 267706 204944 267734
rect 204916 264330 204944 267706
rect 205836 264330 205864 275606
rect 206572 272678 206600 277780
rect 207020 275256 207072 275262
rect 207020 275198 207072 275204
rect 206560 272672 206612 272678
rect 206560 272614 206612 272620
rect 206284 271244 206336 271250
rect 206284 271186 206336 271192
rect 206192 269068 206244 269074
rect 206192 269010 206244 269016
rect 204456 264302 204838 264330
rect 204916 264302 205298 264330
rect 205758 264302 205864 264330
rect 206204 264316 206232 269010
rect 206296 264330 206324 271186
rect 207032 268734 207060 275198
rect 207768 274718 207796 277780
rect 208400 275732 208452 275738
rect 208400 275674 208452 275680
rect 207756 274712 207808 274718
rect 207756 274654 207808 274660
rect 207940 269816 207992 269822
rect 207940 269758 207992 269764
rect 207020 268728 207072 268734
rect 207020 268670 207072 268676
rect 207480 268320 207532 268326
rect 207480 268262 207532 268268
rect 207020 266756 207072 266762
rect 207020 266698 207072 266704
rect 206296 264302 206586 264330
rect 207032 264316 207060 266698
rect 207492 264316 207520 268262
rect 207952 264316 207980 269758
rect 208412 264316 208440 275674
rect 208872 275330 208900 277780
rect 210068 275602 210096 277780
rect 211278 277766 211384 277794
rect 210056 275596 210108 275602
rect 210056 275538 210108 275544
rect 208860 275324 208912 275330
rect 208860 275266 208912 275272
rect 210608 274712 210660 274718
rect 210608 274654 210660 274660
rect 209964 274168 210016 274174
rect 209964 274110 210016 274116
rect 208952 274100 209004 274106
rect 208952 274042 209004 274048
rect 208860 268252 208912 268258
rect 208860 268194 208912 268200
rect 208872 264316 208900 268194
rect 208964 264330 208992 274042
rect 209688 267708 209740 267714
rect 209688 267650 209740 267656
rect 208964 264302 209254 264330
rect 209700 264316 209728 267650
rect 209976 264330 210004 274110
rect 210620 268462 210648 274654
rect 211252 271312 211304 271318
rect 211252 271254 211304 271260
rect 210608 268456 210660 268462
rect 210608 268398 210660 268404
rect 210608 268184 210660 268190
rect 210608 268126 210660 268132
rect 209976 264302 210174 264330
rect 210620 264316 210648 268126
rect 211068 267096 211120 267102
rect 211068 267038 211120 267044
rect 211080 264316 211108 267038
rect 211264 264330 211292 271254
rect 211356 268530 211384 277766
rect 212460 275670 212488 277780
rect 213656 275738 213684 277780
rect 214866 277766 215248 277794
rect 213644 275732 213696 275738
rect 213644 275674 213696 275680
rect 212448 275664 212500 275670
rect 212448 275606 212500 275612
rect 213184 275188 213236 275194
rect 213184 275130 213236 275136
rect 212724 273012 212776 273018
rect 212724 272954 212776 272960
rect 211988 272944 212040 272950
rect 211988 272886 212040 272892
rect 211896 269884 211948 269890
rect 211896 269826 211948 269832
rect 211344 268524 211396 268530
rect 211344 268466 211396 268472
rect 211264 264302 211554 264330
rect 211908 264316 211936 269826
rect 212000 264330 212028 272886
rect 212736 264330 212764 272954
rect 213196 267102 213224 275130
rect 214104 274236 214156 274242
rect 214104 274178 214156 274184
rect 213276 269952 213328 269958
rect 213276 269894 213328 269900
rect 213184 267096 213236 267102
rect 213184 267038 213236 267044
rect 212000 264302 212382 264330
rect 212736 264302 212842 264330
rect 213288 264316 213316 269894
rect 213736 267028 213788 267034
rect 213736 266970 213788 266976
rect 213748 264316 213776 266970
rect 214116 264330 214144 274178
rect 214656 270088 214708 270094
rect 214656 270030 214708 270036
rect 214116 264302 214222 264330
rect 214668 264316 214696 270030
rect 215024 270020 215076 270026
rect 215024 269962 215076 269968
rect 215036 264316 215064 269962
rect 215220 268666 215248 277766
rect 215956 275466 215984 277780
rect 215944 275460 215996 275466
rect 215944 275402 215996 275408
rect 215852 275392 215904 275398
rect 215852 275334 215904 275340
rect 215484 271380 215536 271386
rect 215484 271322 215536 271328
rect 215208 268660 215260 268666
rect 215208 268602 215260 268608
rect 215496 264316 215524 271322
rect 215668 270156 215720 270162
rect 215668 270098 215720 270104
rect 215680 264330 215708 270098
rect 215864 267102 215892 275334
rect 216956 270224 217008 270230
rect 216956 270166 217008 270172
rect 216864 268116 216916 268122
rect 216864 268058 216916 268064
rect 216404 267572 216456 267578
rect 216404 267514 216456 267520
rect 215852 267096 215904 267102
rect 215852 267038 215904 267044
rect 215680 264302 215970 264330
rect 216416 264316 216444 267514
rect 216876 264316 216904 268058
rect 216968 264330 216996 270166
rect 217152 268598 217180 277780
rect 217324 276004 217376 276010
rect 217324 275946 217376 275952
rect 217140 268592 217192 268598
rect 217140 268534 217192 268540
rect 217336 267238 217364 275946
rect 218244 271652 218296 271658
rect 218244 271594 218296 271600
rect 218152 268048 218204 268054
rect 218152 267990 218204 267996
rect 217692 267300 217744 267306
rect 217692 267242 217744 267248
rect 217324 267232 217376 267238
rect 217324 267174 217376 267180
rect 216968 264302 217350 264330
rect 217704 264316 217732 267242
rect 218164 264316 218192 267990
rect 218256 264330 218284 271594
rect 218348 268870 218376 277780
rect 219544 273018 219572 277780
rect 220636 275800 220688 275806
rect 220636 275742 220688 275748
rect 219624 274304 219676 274310
rect 219624 274246 219676 274252
rect 219532 273012 219584 273018
rect 219532 272954 219584 272960
rect 218704 271516 218756 271522
rect 218704 271458 218756 271464
rect 218336 268864 218388 268870
rect 218336 268806 218388 268812
rect 218716 264330 218744 271458
rect 219636 264330 219664 274246
rect 220648 270298 220676 275742
rect 220740 275398 220768 277780
rect 221950 277766 222148 277794
rect 220728 275392 220780 275398
rect 220728 275334 220780 275340
rect 220820 273080 220872 273086
rect 220820 273022 220872 273028
rect 219992 270292 220044 270298
rect 219992 270234 220044 270240
rect 220636 270292 220688 270298
rect 220636 270234 220688 270240
rect 218256 264302 218638 264330
rect 218716 264302 219098 264330
rect 219558 264302 219664 264330
rect 220004 264316 220032 270234
rect 220360 267436 220412 267442
rect 220360 267378 220412 267384
rect 220372 264316 220400 267378
rect 220832 264316 220860 273022
rect 221280 270360 221332 270366
rect 221280 270302 221332 270308
rect 221292 264316 221320 270302
rect 222120 269006 222148 277766
rect 223028 275732 223080 275738
rect 223028 275674 223080 275680
rect 222752 274440 222804 274446
rect 222752 274382 222804 274388
rect 222292 271720 222344 271726
rect 222292 271662 222344 271668
rect 222108 269000 222160 269006
rect 222108 268942 222160 268948
rect 221740 267912 221792 267918
rect 221740 267854 221792 267860
rect 221752 264316 221780 267854
rect 222304 264330 222332 271662
rect 222660 270428 222712 270434
rect 222660 270370 222712 270376
rect 222226 264302 222332 264330
rect 222672 264316 222700 270370
rect 222764 267734 222792 274382
rect 223040 274038 223068 275674
rect 223132 275534 223160 277780
rect 223212 275868 223264 275874
rect 223212 275810 223264 275816
rect 223120 275528 223172 275534
rect 223120 275470 223172 275476
rect 223028 274032 223080 274038
rect 223028 273974 223080 273980
rect 223224 269142 223252 275810
rect 223764 274508 223816 274514
rect 223764 274450 223816 274456
rect 223672 273148 223724 273154
rect 223672 273090 223724 273096
rect 223212 269136 223264 269142
rect 223212 269078 223264 269084
rect 222764 267706 223160 267734
rect 223028 266824 223080 266830
rect 223028 266766 223080 266772
rect 223040 264316 223068 266766
rect 223132 264330 223160 267706
rect 223684 265606 223712 273090
rect 223672 265600 223724 265606
rect 223672 265542 223724 265548
rect 223776 264330 223804 274450
rect 224236 271250 224264 277780
rect 224960 275664 225012 275670
rect 224960 275606 225012 275612
rect 224972 271522 225000 275606
rect 224960 271516 225012 271522
rect 224960 271458 225012 271464
rect 224224 271244 224276 271250
rect 224224 271186 224276 271192
rect 225328 270496 225380 270502
rect 225328 270438 225380 270444
rect 224408 267504 224460 267510
rect 224408 267446 224460 267452
rect 223132 264302 223514 264330
rect 223776 264302 223974 264330
rect 224420 264316 224448 267446
rect 224500 265600 224552 265606
rect 224500 265542 224552 265548
rect 224512 264330 224540 265542
rect 224512 264302 224894 264330
rect 225340 264316 225368 270438
rect 225432 268938 225460 277780
rect 226340 273216 226392 273222
rect 226340 273158 226392 273164
rect 225604 272264 225656 272270
rect 225604 272206 225656 272212
rect 225420 268932 225472 268938
rect 225420 268874 225472 268880
rect 225616 267306 225644 272206
rect 226156 271788 226208 271794
rect 226156 271730 226208 271736
rect 225788 268796 225840 268802
rect 225788 268738 225840 268744
rect 225604 267300 225656 267306
rect 225604 267242 225656 267248
rect 225800 264316 225828 268738
rect 226168 264316 226196 271730
rect 226352 264330 226380 273158
rect 226628 271318 226656 277780
rect 227824 274718 227852 277780
rect 227812 274712 227864 274718
rect 227812 274654 227864 274660
rect 226892 274644 226944 274650
rect 226892 274586 226944 274592
rect 226904 273254 226932 274586
rect 226904 273226 227208 273254
rect 226616 271312 226668 271318
rect 226616 271254 226668 271260
rect 227076 267640 227128 267646
rect 227076 267582 227128 267588
rect 226352 264302 226642 264330
rect 227088 264316 227116 267582
rect 227180 264330 227208 273226
rect 228824 272468 228876 272474
rect 228824 272410 228876 272416
rect 227996 271856 228048 271862
rect 227996 271798 228048 271804
rect 227628 270836 227680 270842
rect 227628 270778 227680 270784
rect 227640 267374 227668 270778
rect 227628 267368 227680 267374
rect 227628 267310 227680 267316
rect 227180 264302 227562 264330
rect 228008 264316 228036 271798
rect 228456 270292 228508 270298
rect 228456 270234 228508 270240
rect 228468 264316 228496 270234
rect 228836 264316 228864 272410
rect 229020 268802 229048 277780
rect 229928 274712 229980 274718
rect 229928 274654 229980 274660
rect 229284 271584 229336 271590
rect 229284 271526 229336 271532
rect 229008 268796 229060 268802
rect 229008 268738 229060 268744
rect 229296 264316 229324 271526
rect 229940 269822 229968 274654
rect 230216 271386 230244 277780
rect 231412 274106 231440 277780
rect 232530 277766 233188 277794
rect 231768 275596 231820 275602
rect 231768 275538 231820 275544
rect 231400 274100 231452 274106
rect 231400 274042 231452 274048
rect 231032 273828 231084 273834
rect 231032 273770 231084 273776
rect 231044 273254 231072 273770
rect 231044 273226 231256 273254
rect 230204 271380 230256 271386
rect 230204 271322 230256 271328
rect 230204 271108 230256 271114
rect 230204 271050 230256 271056
rect 229928 269816 229980 269822
rect 229928 269758 229980 269764
rect 229744 266824 229796 266830
rect 229744 266766 229796 266772
rect 229756 264316 229784 266766
rect 230216 264316 230244 271050
rect 230664 271040 230716 271046
rect 230664 270982 230716 270988
rect 230480 267980 230532 267986
rect 230480 267922 230532 267928
rect 230492 266490 230520 267922
rect 230480 266484 230532 266490
rect 230480 266426 230532 266432
rect 230676 264316 230704 270982
rect 231124 269136 231176 269142
rect 231124 269078 231176 269084
rect 231136 264316 231164 269078
rect 231228 264330 231256 273226
rect 231780 270162 231808 275538
rect 232044 273896 232096 273902
rect 232044 273838 232096 273844
rect 231768 270156 231820 270162
rect 231768 270098 231820 270104
rect 232056 264330 232084 273838
rect 232872 269748 232924 269754
rect 232872 269690 232924 269696
rect 232412 266756 232464 266762
rect 232412 266698 232464 266704
rect 231228 264302 231518 264330
rect 231978 264302 232084 264330
rect 232424 264316 232452 266698
rect 232884 264316 232912 269690
rect 233160 267170 233188 277766
rect 233332 270972 233384 270978
rect 233332 270914 233384 270920
rect 233148 267164 233200 267170
rect 233148 267106 233200 267112
rect 233344 264316 233372 270914
rect 233712 269890 233740 277780
rect 234908 275602 234936 277780
rect 234896 275596 234948 275602
rect 234896 275538 234948 275544
rect 234620 275324 234672 275330
rect 234620 275266 234672 275272
rect 234632 270230 234660 275266
rect 235264 272400 235316 272406
rect 235264 272342 235316 272348
rect 234620 270224 234672 270230
rect 234620 270166 234672 270172
rect 233700 269884 233752 269890
rect 233700 269826 233752 269832
rect 234160 269680 234212 269686
rect 234160 269622 234212 269628
rect 233792 268728 233844 268734
rect 233792 268670 233844 268676
rect 233804 264316 233832 268670
rect 234172 264316 234200 269622
rect 234620 269612 234672 269618
rect 234620 269554 234672 269560
rect 234632 264316 234660 269554
rect 235080 268388 235132 268394
rect 235080 268330 235132 268336
rect 235092 264316 235120 268330
rect 235276 266422 235304 272342
rect 236104 270026 236132 277780
rect 237300 277394 237328 277780
rect 238510 277766 238708 277794
rect 237208 277366 237328 277394
rect 236736 272944 236788 272950
rect 236736 272886 236788 272892
rect 236092 270020 236144 270026
rect 236092 269962 236144 269968
rect 235540 269544 235592 269550
rect 235540 269486 235592 269492
rect 235264 266416 235316 266422
rect 235264 266358 235316 266364
rect 235552 264316 235580 269486
rect 236644 269000 236696 269006
rect 236644 268942 236696 268948
rect 236656 267306 236684 268942
rect 236748 267510 236776 272886
rect 237208 269958 237236 277366
rect 238024 273692 238076 273698
rect 238024 273634 238076 273640
rect 237196 269952 237248 269958
rect 237196 269894 237248 269900
rect 236920 269476 236972 269482
rect 236920 269418 236972 269424
rect 236736 267504 236788 267510
rect 236736 267446 236788 267452
rect 236000 267300 236052 267306
rect 236000 267242 236052 267248
rect 236644 267300 236696 267306
rect 236644 267242 236696 267248
rect 236012 264316 236040 267242
rect 236460 267028 236512 267034
rect 236460 266970 236512 266976
rect 236472 264316 236500 266970
rect 236932 264316 236960 269418
rect 237288 267368 237340 267374
rect 237288 267310 237340 267316
rect 237300 264316 237328 267310
rect 238036 267238 238064 273634
rect 237748 267232 237800 267238
rect 237748 267174 237800 267180
rect 238024 267232 238076 267238
rect 238024 267174 238076 267180
rect 237760 264316 237788 267174
rect 238680 267034 238708 277766
rect 239600 275330 239628 277780
rect 240810 277766 241468 277794
rect 242006 277766 242296 277794
rect 240048 275460 240100 275466
rect 240048 275402 240100 275408
rect 239588 275324 239640 275330
rect 239588 275266 239640 275272
rect 239220 272808 239272 272814
rect 239220 272750 239272 272756
rect 238852 270904 238904 270910
rect 238852 270846 238904 270852
rect 238668 267028 238720 267034
rect 238668 266970 238720 266976
rect 238668 266484 238720 266490
rect 238668 266426 238720 266432
rect 238208 266416 238260 266422
rect 238208 266358 238260 266364
rect 238220 264316 238248 266358
rect 238680 264316 238708 266426
rect 238864 265606 238892 270846
rect 239128 267096 239180 267102
rect 239128 267038 239180 267044
rect 238852 265600 238904 265606
rect 238852 265542 238904 265548
rect 239140 264316 239168 267038
rect 239232 264330 239260 272750
rect 240060 272746 240088 275402
rect 240140 273760 240192 273766
rect 240140 273702 240192 273708
rect 240048 272740 240100 272746
rect 240048 272682 240100 272688
rect 239312 268864 239364 268870
rect 239312 268806 239364 268812
rect 239324 267102 239352 268806
rect 239312 267096 239364 267102
rect 239312 267038 239364 267044
rect 240152 265606 240180 273702
rect 240968 272536 241020 272542
rect 240968 272478 241020 272484
rect 240232 272332 240284 272338
rect 240232 272274 240284 272280
rect 240244 267734 240272 272274
rect 240244 267706 240364 267734
rect 239680 265600 239732 265606
rect 239680 265542 239732 265548
rect 240140 265600 240192 265606
rect 240140 265542 240192 265548
rect 239692 264330 239720 265542
rect 240336 264330 240364 267706
rect 240508 265600 240560 265606
rect 240508 265542 240560 265548
rect 240520 264330 240548 265542
rect 240980 264330 241008 272478
rect 241440 270094 241468 277766
rect 242072 274576 242124 274582
rect 242072 274518 242124 274524
rect 241612 274372 241664 274378
rect 241612 274314 241664 274320
rect 241428 270088 241480 270094
rect 241428 270030 241480 270036
rect 241624 267734 241652 274314
rect 241624 267706 241928 267734
rect 241796 267232 241848 267238
rect 241796 267174 241848 267180
rect 239232 264302 239614 264330
rect 239692 264302 239982 264330
rect 240336 264302 240442 264330
rect 240520 264302 240902 264330
rect 240980 264302 241362 264330
rect 241808 264316 241836 267174
rect 241900 264330 241928 267706
rect 242084 264602 242112 274518
rect 242268 271182 242296 277766
rect 243188 274174 243216 277780
rect 244280 275528 244332 275534
rect 244280 275470 244332 275476
rect 243360 275392 243412 275398
rect 243360 275334 243412 275340
rect 243176 274168 243228 274174
rect 243176 274110 243228 274116
rect 243176 272604 243228 272610
rect 243176 272546 243228 272552
rect 242992 271448 243044 271454
rect 242992 271390 243044 271396
rect 242164 271176 242216 271182
rect 242164 271118 242216 271124
rect 242256 271176 242308 271182
rect 242256 271118 242308 271124
rect 242176 266422 242204 271118
rect 242164 266416 242216 266422
rect 242164 266358 242216 266364
rect 243004 265606 243032 271390
rect 243084 266416 243136 266422
rect 243084 266358 243136 266364
rect 242992 265600 243044 265606
rect 242992 265542 243044 265548
rect 242084 264574 242388 264602
rect 242360 264330 242388 264574
rect 241900 264302 242282 264330
rect 242360 264302 242650 264330
rect 243096 264316 243124 266358
rect 243188 264330 243216 272546
rect 243372 267782 243400 275334
rect 244292 273902 244320 275470
rect 244384 275398 244412 277780
rect 244372 275392 244424 275398
rect 244372 275334 244424 275340
rect 244556 273964 244608 273970
rect 244556 273906 244608 273912
rect 244280 273896 244332 273902
rect 244280 273838 244332 273844
rect 244372 272672 244424 272678
rect 244372 272614 244424 272620
rect 244188 268660 244240 268666
rect 244188 268602 244240 268608
rect 243360 267776 243412 267782
rect 243360 267718 243412 267724
rect 244200 266422 244228 268602
rect 244188 266416 244240 266422
rect 244188 266358 244240 266364
rect 244384 265606 244412 272614
rect 244464 267504 244516 267510
rect 244464 267446 244516 267452
rect 243636 265600 243688 265606
rect 243636 265542 243688 265548
rect 244372 265600 244424 265606
rect 244372 265542 244424 265548
rect 243648 264330 243676 265542
rect 243188 264302 243570 264330
rect 243648 264302 244030 264330
rect 244476 264316 244504 267446
rect 244568 264330 244596 273906
rect 245580 272542 245608 277780
rect 245660 275596 245712 275602
rect 245660 275538 245712 275544
rect 245568 272536 245620 272542
rect 245568 272478 245620 272484
rect 245292 268932 245344 268938
rect 245292 268874 245344 268880
rect 245304 267238 245332 268874
rect 245672 268666 245700 275538
rect 246776 272610 246804 277780
rect 247894 277766 248368 277794
rect 249090 277766 249748 277794
rect 247224 274032 247276 274038
rect 247224 273974 247276 273980
rect 246764 272604 246816 272610
rect 246764 272546 246816 272552
rect 246212 270224 246264 270230
rect 246212 270166 246264 270172
rect 245660 268660 245712 268666
rect 245660 268602 245712 268608
rect 245752 268456 245804 268462
rect 245752 268398 245804 268404
rect 245292 267232 245344 267238
rect 245292 267174 245344 267180
rect 245016 265600 245068 265606
rect 245016 265542 245068 265548
rect 245028 264330 245056 265542
rect 244568 264302 244950 264330
rect 245028 264302 245318 264330
rect 245764 264316 245792 268398
rect 246224 264316 246252 270166
rect 246672 270156 246724 270162
rect 246672 270098 246724 270104
rect 246684 264316 246712 270098
rect 247132 268524 247184 268530
rect 247132 268466 247184 268472
rect 247144 264316 247172 268466
rect 247236 265606 247264 273974
rect 247316 271516 247368 271522
rect 247316 271458 247368 271464
rect 247224 265600 247276 265606
rect 247224 265542 247276 265548
rect 247328 264330 247356 271458
rect 248340 268394 248368 277766
rect 248604 272740 248656 272746
rect 248604 272682 248656 272688
rect 248328 268388 248380 268394
rect 248328 268330 248380 268336
rect 248420 266416 248472 266422
rect 248420 266358 248472 266364
rect 247684 265600 247736 265606
rect 247684 265542 247736 265548
rect 247696 264330 247724 265542
rect 247328 264302 247618 264330
rect 247696 264302 248078 264330
rect 248432 264316 248460 266358
rect 248616 264330 248644 272682
rect 249340 268592 249392 268598
rect 249340 268534 249392 268540
rect 248616 264302 248906 264330
rect 249352 264316 249380 268534
rect 249720 268462 249748 277766
rect 250272 275806 250300 277780
rect 250260 275800 250312 275806
rect 250260 275742 250312 275748
rect 251180 275800 251232 275806
rect 251180 275742 251232 275748
rect 251192 273970 251220 275742
rect 251468 275738 251496 277780
rect 251456 275732 251508 275738
rect 251456 275674 251508 275680
rect 252376 275732 252428 275738
rect 252376 275674 252428 275680
rect 251180 273964 251232 273970
rect 251180 273906 251232 273912
rect 251364 273896 251416 273902
rect 251364 273838 251416 273844
rect 249984 272876 250036 272882
rect 249984 272818 250036 272824
rect 249708 268456 249760 268462
rect 249708 268398 249760 268404
rect 249800 267096 249852 267102
rect 249800 267038 249852 267044
rect 249812 264316 249840 267038
rect 249996 264330 250024 272818
rect 251272 271244 251324 271250
rect 251272 271186 251324 271192
rect 250720 267776 250772 267782
rect 250720 267718 250772 267724
rect 249996 264302 250286 264330
rect 250732 264316 250760 267718
rect 251088 267300 251140 267306
rect 251088 267242 251140 267248
rect 251100 264316 251128 267242
rect 251284 265606 251312 271186
rect 251272 265600 251324 265606
rect 251272 265542 251324 265548
rect 251376 264330 251404 273838
rect 252388 267102 252416 275674
rect 252664 274922 252692 277780
rect 252928 275324 252980 275330
rect 252928 275266 252980 275272
rect 252652 274916 252704 274922
rect 252652 274858 252704 274864
rect 252940 271658 252968 275266
rect 252928 271652 252980 271658
rect 252928 271594 252980 271600
rect 252744 271312 252796 271318
rect 252744 271254 252796 271260
rect 252468 267232 252520 267238
rect 252468 267174 252520 267180
rect 252376 267096 252428 267102
rect 252376 267038 252428 267044
rect 251732 265600 251784 265606
rect 251732 265542 251784 265548
rect 251744 264330 251772 265542
rect 251376 264302 251574 264330
rect 251744 264302 252034 264330
rect 252480 264316 252508 267174
rect 252756 264330 252784 271254
rect 253860 271250 253888 277780
rect 255070 277766 255268 277794
rect 256174 277766 256648 277794
rect 257370 277766 258028 277794
rect 254308 274100 254360 274106
rect 254308 274042 254360 274048
rect 254032 271380 254084 271386
rect 254032 271322 254084 271328
rect 253848 271244 253900 271250
rect 253848 271186 253900 271192
rect 253388 269816 253440 269822
rect 253388 269758 253440 269764
rect 252756 264302 252954 264330
rect 253400 264316 253428 269758
rect 253756 268796 253808 268802
rect 253756 268738 253808 268744
rect 253768 264316 253796 268738
rect 254044 264330 254072 271322
rect 254320 264330 254348 274042
rect 255240 267170 255268 277766
rect 256424 270020 256476 270026
rect 256424 269962 256476 269968
rect 255596 269884 255648 269890
rect 255596 269826 255648 269832
rect 255136 267164 255188 267170
rect 255136 267106 255188 267112
rect 255228 267164 255280 267170
rect 255228 267106 255280 267112
rect 254044 264302 254242 264330
rect 254320 264302 254702 264330
rect 255148 264316 255176 267106
rect 255608 264316 255636 269826
rect 256056 268660 256108 268666
rect 256056 268602 256108 268608
rect 256068 264316 256096 268602
rect 256436 264316 256464 269962
rect 256620 267238 256648 277766
rect 257436 271652 257488 271658
rect 257436 271594 257488 271600
rect 256884 269952 256936 269958
rect 256884 269894 256936 269900
rect 256608 267232 256660 267238
rect 256608 267174 256660 267180
rect 256896 264316 256924 269894
rect 257344 267028 257396 267034
rect 257344 266970 257396 266976
rect 257356 264316 257384 266970
rect 257448 264330 257476 271594
rect 258000 267034 258028 277766
rect 258552 275806 258580 277780
rect 258540 275800 258592 275806
rect 258540 275742 258592 275748
rect 259368 275392 259420 275398
rect 259368 275334 259420 275340
rect 258632 274168 258684 274174
rect 258632 274110 258684 274116
rect 258264 271176 258316 271182
rect 258264 271118 258316 271124
rect 258080 270088 258132 270094
rect 258080 270030 258132 270036
rect 257988 267028 258040 267034
rect 257988 266970 258040 266976
rect 258092 264330 258120 270030
rect 258276 267734 258304 271118
rect 258644 267734 258672 274110
rect 259380 267734 259408 275334
rect 259748 275330 259776 277780
rect 259736 275324 259788 275330
rect 259736 275266 259788 275272
rect 260944 274922 260972 277780
rect 262140 274990 262168 277780
rect 262128 274984 262180 274990
rect 262128 274926 262180 274932
rect 260932 274916 260984 274922
rect 260932 274858 260984 274864
rect 263244 274718 263272 277780
rect 264440 274786 264468 277780
rect 265650 277766 266308 277794
rect 264612 275800 264664 275806
rect 264612 275742 264664 275748
rect 264428 274780 264480 274786
rect 264428 274722 264480 274728
rect 263232 274712 263284 274718
rect 263232 274654 263284 274660
rect 262404 274644 262456 274650
rect 262404 274586 262456 274592
rect 261484 273964 261536 273970
rect 261484 273906 261536 273912
rect 259644 272604 259696 272610
rect 259644 272546 259696 272552
rect 258276 267706 258396 267734
rect 258644 267706 258856 267734
rect 259380 267706 259500 267734
rect 258368 264330 258396 267706
rect 258828 264330 258856 267706
rect 259472 264330 259500 267706
rect 259656 265606 259684 272546
rect 259736 272536 259788 272542
rect 259736 272478 259788 272484
rect 259644 265600 259696 265606
rect 259644 265542 259696 265548
rect 259748 264330 259776 272478
rect 261392 268456 261444 268462
rect 261392 268398 261444 268404
rect 260932 268388 260984 268394
rect 260932 268330 260984 268336
rect 260196 265600 260248 265606
rect 260196 265542 260248 265548
rect 260208 264330 260236 265542
rect 257448 264302 257830 264330
rect 258092 264302 258290 264330
rect 258368 264302 258750 264330
rect 258828 264302 259210 264330
rect 259472 264302 259578 264330
rect 259748 264302 260038 264330
rect 260208 264302 260498 264330
rect 260944 264316 260972 268330
rect 261404 264316 261432 268398
rect 261496 264330 261524 273906
rect 262312 271244 262364 271250
rect 262312 271186 262364 271192
rect 262220 267096 262272 267102
rect 262220 267038 262272 267044
rect 261496 264302 261878 264330
rect 262232 264316 262260 267038
rect 262324 265606 262352 271186
rect 262312 265600 262364 265606
rect 262312 265542 262364 265548
rect 262416 264330 262444 274586
rect 264060 267232 264112 267238
rect 264060 267174 264112 267180
rect 263600 267164 263652 267170
rect 263600 267106 263652 267112
rect 262772 265600 262824 265606
rect 262772 265542 262824 265548
rect 262784 264330 262812 265542
rect 262416 264302 262706 264330
rect 262784 264302 263166 264330
rect 263612 264316 263640 267106
rect 264072 264316 264100 267174
rect 264520 267028 264572 267034
rect 264520 266970 264572 266976
rect 264532 264316 264560 266970
rect 264624 264330 264652 275742
rect 265072 275324 265124 275330
rect 265072 275266 265124 275272
rect 264980 274984 265032 274990
rect 264980 274926 265032 274932
rect 264992 265606 265020 274926
rect 264980 265600 265032 265606
rect 264980 265542 265032 265548
rect 265084 264330 265112 275266
rect 265440 274916 265492 274922
rect 265440 274858 265492 274864
rect 265452 264330 265480 274858
rect 266280 274666 266308 277766
rect 266728 274780 266780 274786
rect 266728 274722 266780 274728
rect 266452 274712 266504 274718
rect 266280 274638 266400 274666
rect 266452 274654 266504 274660
rect 266372 265606 266400 274638
rect 265900 265600 265952 265606
rect 265900 265542 265952 265548
rect 266360 265600 266412 265606
rect 266360 265542 266412 265548
rect 265912 264330 265940 265542
rect 266464 264330 266492 274654
rect 266740 267734 266768 274722
rect 266832 274718 266860 277780
rect 268042 277766 268148 277794
rect 266820 274712 266872 274718
rect 266820 274654 266872 274660
rect 267740 274712 267792 274718
rect 267740 274654 267792 274660
rect 266740 267706 266860 267734
rect 266832 264330 266860 267706
rect 267280 265600 267332 265606
rect 267280 265542 267332 265548
rect 267292 264330 267320 265542
rect 267752 264330 267780 274654
rect 268120 264330 268148 277766
rect 269224 267734 269252 277780
rect 269040 267706 269252 267734
rect 269408 277766 270434 277794
rect 270512 277766 271538 277794
rect 272168 277766 272734 277794
rect 273272 277766 273930 277794
rect 274652 277766 275126 277794
rect 269040 264330 269068 267706
rect 264624 264302 264914 264330
rect 265084 264302 265374 264330
rect 265452 264302 265834 264330
rect 265912 264302 266294 264330
rect 266464 264302 266754 264330
rect 266832 264302 267214 264330
rect 267292 264302 267582 264330
rect 267752 264302 268042 264330
rect 268120 264302 268502 264330
rect 268962 264302 269068 264330
rect 269408 264316 269436 277766
rect 270512 267734 270540 277766
rect 270236 267706 270540 267734
rect 270236 264330 270264 267706
rect 272064 267504 272116 267510
rect 272064 267446 272116 267452
rect 271604 266620 271656 266626
rect 271604 266562 271656 266568
rect 271144 266552 271196 266558
rect 271144 266494 271196 266500
rect 270684 266484 270736 266490
rect 270684 266426 270736 266432
rect 270316 266416 270368 266422
rect 270316 266358 270368 266364
rect 269882 264302 270264 264330
rect 270328 264316 270356 266358
rect 270696 264316 270724 266426
rect 271156 264316 271184 266494
rect 271616 264316 271644 266562
rect 272076 264316 272104 267446
rect 272168 266422 272196 277766
rect 273168 274168 273220 274174
rect 273168 274110 273220 274116
rect 272524 266892 272576 266898
rect 272524 266834 272576 266840
rect 272156 266416 272208 266422
rect 272156 266358 272208 266364
rect 272536 264316 272564 266834
rect 273180 264330 273208 274110
rect 273272 266490 273300 277766
rect 274180 272536 274232 272542
rect 274180 272478 274232 272484
rect 273352 270088 273404 270094
rect 273352 270030 273404 270036
rect 273260 266484 273312 266490
rect 273260 266426 273312 266432
rect 273010 264302 273208 264330
rect 273364 264316 273392 270030
rect 274192 264330 274220 272478
rect 274272 268456 274324 268462
rect 274272 268398 274324 268404
rect 273838 264302 274220 264330
rect 274284 264316 274312 268398
rect 274652 266558 274680 277766
rect 274732 270020 274784 270026
rect 274732 269962 274784 269968
rect 274640 266552 274692 266558
rect 274640 266494 274692 266500
rect 274744 264316 274772 269962
rect 276020 269952 276072 269958
rect 276020 269894 276072 269900
rect 275652 268388 275704 268394
rect 275652 268330 275704 268336
rect 275192 266552 275244 266558
rect 275192 266494 275244 266500
rect 275204 264316 275232 266494
rect 275664 264316 275692 268330
rect 276032 264316 276060 269894
rect 276308 266626 276336 277780
rect 277504 277394 277532 277780
rect 277412 277366 277532 277394
rect 277780 277766 278714 277794
rect 277308 274032 277360 274038
rect 277308 273974 277360 273980
rect 276940 267300 276992 267306
rect 276940 267242 276992 267248
rect 276296 266620 276348 266626
rect 276296 266562 276348 266568
rect 276480 266416 276532 266422
rect 276480 266358 276532 266364
rect 276492 264316 276520 266358
rect 276952 264316 276980 267242
rect 277320 266422 277348 273974
rect 277412 267510 277440 277366
rect 277400 267504 277452 267510
rect 277400 267446 277452 267452
rect 277780 266898 277808 277766
rect 279804 274174 279832 277780
rect 280172 277766 281014 277794
rect 279792 274168 279844 274174
rect 279792 274110 279844 274116
rect 279424 273284 279476 273290
rect 279424 273226 279476 273232
rect 277860 269884 277912 269890
rect 277860 269826 277912 269832
rect 277768 266892 277820 266898
rect 277768 266834 277820 266840
rect 277400 266620 277452 266626
rect 277400 266562 277452 266568
rect 277308 266416 277360 266422
rect 277308 266358 277360 266364
rect 277412 264316 277440 266562
rect 277872 264316 277900 269826
rect 279148 269816 279200 269822
rect 279148 269758 279200 269764
rect 278688 268796 278740 268802
rect 278688 268738 278740 268744
rect 278320 267028 278372 267034
rect 278320 266970 278372 266976
rect 278332 264316 278360 266970
rect 278700 264316 278728 268738
rect 279160 264316 279188 269758
rect 279436 266558 279464 273226
rect 279976 271312 280028 271318
rect 279976 271254 280028 271260
rect 279424 266552 279476 266558
rect 279424 266494 279476 266500
rect 279988 264330 280016 271254
rect 280172 270094 280200 277766
rect 282196 272542 282224 277780
rect 282932 277766 283406 277794
rect 284312 277766 284602 277794
rect 282828 272740 282880 272746
rect 282828 272682 282880 272688
rect 282184 272536 282236 272542
rect 282184 272478 282236 272484
rect 281356 271244 281408 271250
rect 281356 271186 281408 271192
rect 280160 270088 280212 270094
rect 280160 270030 280212 270036
rect 280528 268660 280580 268666
rect 280528 268602 280580 268608
rect 280540 266626 280568 268602
rect 280528 266620 280580 266626
rect 280528 266562 280580 266568
rect 280988 266620 281040 266626
rect 280988 266562 281040 266568
rect 280068 266484 280120 266490
rect 280068 266426 280120 266432
rect 279634 264302 280016 264330
rect 280080 264316 280108 266426
rect 280528 266416 280580 266422
rect 280528 266358 280580 266364
rect 280540 264316 280568 266358
rect 281000 264316 281028 266562
rect 281368 266422 281396 271186
rect 282736 270088 282788 270094
rect 282736 270030 282788 270036
rect 281448 268524 281500 268530
rect 281448 268466 281500 268472
rect 281356 266416 281408 266422
rect 281356 266358 281408 266364
rect 281460 264316 281488 268466
rect 282748 267306 282776 270030
rect 282736 267300 282788 267306
rect 282736 267242 282788 267248
rect 282276 266688 282328 266694
rect 282276 266630 282328 266636
rect 281816 266416 281868 266422
rect 281816 266358 281868 266364
rect 281828 264316 281856 266358
rect 282288 264316 282316 266630
rect 282840 264330 282868 272682
rect 282932 268462 282960 277766
rect 284024 271176 284076 271182
rect 284024 271118 284076 271124
rect 283012 268592 283064 268598
rect 283012 268534 283064 268540
rect 282920 268456 282972 268462
rect 282920 268398 282972 268404
rect 283024 266422 283052 268534
rect 283196 267640 283248 267646
rect 283196 267582 283248 267588
rect 283012 266416 283064 266422
rect 283012 266358 283064 266364
rect 282762 264302 282868 264330
rect 283208 264316 283236 267582
rect 284036 264330 284064 271118
rect 284312 270026 284340 277766
rect 285784 273290 285812 277780
rect 285876 277766 286902 277794
rect 287072 277766 288098 277794
rect 285772 273284 285824 273290
rect 285772 273226 285824 273232
rect 285588 272672 285640 272678
rect 285588 272614 285640 272620
rect 284300 270020 284352 270026
rect 284300 269962 284352 269968
rect 284852 268864 284904 268870
rect 284852 268806 284904 268812
rect 284484 267572 284536 267578
rect 284484 267514 284536 267520
rect 284116 266416 284168 266422
rect 284116 266358 284168 266364
rect 283682 264302 284064 264330
rect 284128 264316 284156 266358
rect 284496 264316 284524 267514
rect 284864 266490 284892 268806
rect 284944 267708 284996 267714
rect 284944 267650 284996 267656
rect 284852 266484 284904 266490
rect 284852 266426 284904 266432
rect 284956 264316 284984 267650
rect 285600 264330 285628 272614
rect 285876 268394 285904 277766
rect 286876 272536 286928 272542
rect 286876 272478 286928 272484
rect 286784 268456 286836 268462
rect 286784 268398 286836 268404
rect 285864 268388 285916 268394
rect 285864 268330 285916 268336
rect 286232 268388 286284 268394
rect 286232 268330 286284 268336
rect 286244 264330 286272 268330
rect 286324 267164 286376 267170
rect 286324 267106 286376 267112
rect 285430 264302 285628 264330
rect 285890 264302 286272 264330
rect 286336 264316 286364 267106
rect 286796 266422 286824 268398
rect 286784 266416 286836 266422
rect 286784 266358 286836 266364
rect 286888 264330 286916 272478
rect 287072 269958 287100 277766
rect 289084 274304 289136 274310
rect 289084 274246 289136 274252
rect 287704 273964 287756 273970
rect 287704 273906 287756 273912
rect 287060 269952 287112 269958
rect 287060 269894 287112 269900
rect 287716 266694 287744 273906
rect 288348 272604 288400 272610
rect 288348 272546 288400 272552
rect 287796 271788 287848 271794
rect 287796 271730 287848 271736
rect 287808 267034 287836 271730
rect 288072 267436 288124 267442
rect 288072 267378 288124 267384
rect 287796 267028 287848 267034
rect 287796 266970 287848 266976
rect 287704 266688 287756 266694
rect 287704 266630 287756 266636
rect 287612 266484 287664 266490
rect 287612 266426 287664 266432
rect 287152 266416 287204 266422
rect 287152 266358 287204 266364
rect 286810 264302 286916 264330
rect 287164 264316 287192 266358
rect 287624 264316 287652 266426
rect 288084 264316 288112 267378
rect 288360 266422 288388 272546
rect 288532 267504 288584 267510
rect 288532 267446 288584 267452
rect 288348 266416 288400 266422
rect 288348 266358 288400 266364
rect 288544 264316 288572 267446
rect 288992 267232 289044 267238
rect 288992 267174 289044 267180
rect 289004 264316 289032 267174
rect 289096 266490 289124 274246
rect 289280 274038 289308 277780
rect 289832 277766 290490 277794
rect 291212 277766 291686 277794
rect 292592 277766 292882 277794
rect 289268 274032 289320 274038
rect 289268 273974 289320 273980
rect 289176 272876 289228 272882
rect 289176 272818 289228 272824
rect 289188 266626 289216 272818
rect 289832 270094 289860 277766
rect 291016 274372 291068 274378
rect 291016 274314 291068 274320
rect 289820 270088 289872 270094
rect 289820 270030 289872 270036
rect 290924 268728 290976 268734
rect 290924 268670 290976 268676
rect 290936 267646 290964 268670
rect 290924 267640 290976 267646
rect 290924 267582 290976 267588
rect 289452 267368 289504 267374
rect 289452 267310 289504 267316
rect 289176 266620 289228 266626
rect 289176 266562 289228 266568
rect 289084 266484 289136 266490
rect 289084 266426 289136 266432
rect 289464 264316 289492 267310
rect 290740 267300 290792 267306
rect 290740 267242 290792 267248
rect 289820 266484 289872 266490
rect 289820 266426 289872 266432
rect 289832 264316 289860 266426
rect 290280 266416 290332 266422
rect 290280 266358 290332 266364
rect 290292 264316 290320 266358
rect 290752 264316 290780 267242
rect 291028 266490 291056 274314
rect 291108 274236 291160 274242
rect 291108 274178 291160 274184
rect 291016 266484 291068 266490
rect 291016 266426 291068 266432
rect 291120 266422 291148 274178
rect 291212 268666 291240 277766
rect 292488 274168 292540 274174
rect 292488 274110 292540 274116
rect 291844 272808 291896 272814
rect 291844 272750 291896 272756
rect 291200 268660 291252 268666
rect 291200 268602 291252 268608
rect 291476 268660 291528 268666
rect 291476 268602 291528 268608
rect 291488 267578 291516 268602
rect 291856 267714 291884 272750
rect 292120 269612 292172 269618
rect 292120 269554 292172 269560
rect 291844 267708 291896 267714
rect 291844 267650 291896 267656
rect 291476 267572 291528 267578
rect 291476 267514 291528 267520
rect 291660 266484 291712 266490
rect 291660 266426 291712 266432
rect 291108 266416 291160 266422
rect 291108 266358 291160 266364
rect 291200 266416 291252 266422
rect 291200 266358 291252 266364
rect 291212 264316 291240 266358
rect 291672 264316 291700 266426
rect 292132 264316 292160 269554
rect 292500 266422 292528 274110
rect 292592 269890 292620 277766
rect 294064 271794 294092 277780
rect 294156 277766 295182 277794
rect 295352 277766 296378 277794
rect 294052 271788 294104 271794
rect 294052 271730 294104 271736
rect 293868 270496 293920 270502
rect 293868 270438 293920 270444
rect 292580 269884 292632 269890
rect 292580 269826 292632 269832
rect 293408 269680 293460 269686
rect 293408 269622 293460 269628
rect 292580 267096 292632 267102
rect 292580 267038 292632 267044
rect 292488 266416 292540 266422
rect 292488 266358 292540 266364
rect 292592 264316 292620 267038
rect 292948 266756 293000 266762
rect 292948 266698 293000 266704
rect 292960 264316 292988 266698
rect 293420 264316 293448 269622
rect 293880 264316 293908 270438
rect 294156 268802 294184 277766
rect 295352 269822 295380 277766
rect 295984 274440 296036 274446
rect 295984 274382 296036 274388
rect 295340 269816 295392 269822
rect 295340 269758 295392 269764
rect 294788 269748 294840 269754
rect 294788 269690 294840 269696
rect 294144 268796 294196 268802
rect 294144 268738 294196 268744
rect 294328 266892 294380 266898
rect 294328 266834 294380 266840
rect 294340 264316 294368 266834
rect 294800 264316 294828 269690
rect 295248 267028 295300 267034
rect 295248 266970 295300 266976
rect 295260 264316 295288 266970
rect 295996 266490 296024 274382
rect 296444 274100 296496 274106
rect 296444 274042 296496 274048
rect 296076 270428 296128 270434
rect 296076 270370 296128 270376
rect 295984 266484 296036 266490
rect 295984 266426 296036 266432
rect 295616 266416 295668 266422
rect 295616 266358 295668 266364
rect 295628 264316 295656 266358
rect 296088 264316 296116 270370
rect 296456 264330 296484 274042
rect 296536 271856 296588 271862
rect 296536 271798 296588 271804
rect 296548 266422 296576 271798
rect 297560 271318 297588 277780
rect 298112 277766 298770 277794
rect 297824 271788 297876 271794
rect 297824 271730 297876 271736
rect 297548 271312 297600 271318
rect 297548 271254 297600 271260
rect 297456 270156 297508 270162
rect 297456 270098 297508 270104
rect 296536 266416 296588 266422
rect 296536 266358 296588 266364
rect 296996 266416 297048 266422
rect 296996 266358 297048 266364
rect 296456 264302 296562 264330
rect 297008 264316 297036 266358
rect 297468 264316 297496 270098
rect 297836 266422 297864 271730
rect 297916 270360 297968 270366
rect 297916 270302 297968 270308
rect 297824 266416 297876 266422
rect 297824 266358 297876 266364
rect 297928 264316 297956 270302
rect 298112 268870 298140 277766
rect 299952 271250 299980 277780
rect 300768 274032 300820 274038
rect 300768 273974 300820 273980
rect 300124 273216 300176 273222
rect 300124 273158 300176 273164
rect 299940 271244 299992 271250
rect 299940 271186 299992 271192
rect 298744 270292 298796 270298
rect 298744 270234 298796 270240
rect 298100 268864 298152 268870
rect 298100 268806 298152 268812
rect 298284 267640 298336 267646
rect 298284 267582 298336 267588
rect 298296 264316 298324 267582
rect 298756 264316 298784 270234
rect 299204 267708 299256 267714
rect 299204 267650 299256 267656
rect 299216 264316 299244 267650
rect 299664 267572 299716 267578
rect 299664 267514 299716 267520
rect 299676 264316 299704 267514
rect 300136 267442 300164 273158
rect 300400 270224 300452 270230
rect 300400 270166 300452 270172
rect 300124 267436 300176 267442
rect 300124 267378 300176 267384
rect 300412 264330 300440 270166
rect 300780 264330 300808 273974
rect 301148 272882 301176 277780
rect 302344 277394 302372 277780
rect 302252 277366 302372 277394
rect 302436 277766 303462 277794
rect 301504 273148 301556 273154
rect 301504 273090 301556 273096
rect 301136 272876 301188 272882
rect 301136 272818 301188 272824
rect 301412 270088 301464 270094
rect 301412 270030 301464 270036
rect 300952 266416 301004 266422
rect 300952 266358 301004 266364
rect 300150 264302 300440 264330
rect 300610 264302 300808 264330
rect 300964 264316 300992 266358
rect 301424 264316 301452 270030
rect 301516 267510 301544 273090
rect 302148 271720 302200 271726
rect 302148 271662 302200 271668
rect 301504 267504 301556 267510
rect 301504 267446 301556 267452
rect 301872 266756 301924 266762
rect 301872 266698 301924 266704
rect 301884 264316 301912 266698
rect 302160 266422 302188 271662
rect 302252 268530 302280 277366
rect 302436 268598 302464 277766
rect 304644 273970 304672 277780
rect 304632 273964 304684 273970
rect 304632 273906 304684 273912
rect 304724 273964 304776 273970
rect 304724 273906 304776 273912
rect 304264 273896 304316 273902
rect 304264 273838 304316 273844
rect 303252 269952 303304 269958
rect 303252 269894 303304 269900
rect 302424 268592 302476 268598
rect 302424 268534 302476 268540
rect 302240 268524 302292 268530
rect 302240 268466 302292 268472
rect 302332 268184 302384 268190
rect 302332 268126 302384 268132
rect 302148 266416 302200 266422
rect 302148 266358 302200 266364
rect 302344 264316 302372 268126
rect 302792 266484 302844 266490
rect 302792 266426 302844 266432
rect 302804 264316 302832 266426
rect 303264 264316 303292 269894
rect 303712 268252 303764 268258
rect 303712 268194 303764 268200
rect 303724 264316 303752 268194
rect 304276 267374 304304 273838
rect 304264 267368 304316 267374
rect 304264 267310 304316 267316
rect 304080 266416 304132 266422
rect 304080 266358 304132 266364
rect 304092 264316 304120 266358
rect 304736 264330 304764 273906
rect 305840 272746 305868 277780
rect 306392 277766 307050 277794
rect 305828 272740 305880 272746
rect 305828 272682 305880 272688
rect 304816 271652 304868 271658
rect 304816 271594 304868 271600
rect 304828 266422 304856 271594
rect 306288 271584 306340 271590
rect 306288 271526 306340 271532
rect 306012 270020 306064 270026
rect 306012 269962 306064 269968
rect 305920 269884 305972 269890
rect 305920 269826 305972 269832
rect 305000 267436 305052 267442
rect 305000 267378 305052 267384
rect 304816 266416 304868 266422
rect 304816 266358 304868 266364
rect 304566 264302 304764 264330
rect 305012 264316 305040 267378
rect 305460 266416 305512 266422
rect 305460 266358 305512 266364
rect 305472 264316 305500 266358
rect 305932 264316 305960 269826
rect 306024 266490 306052 269962
rect 306012 266484 306064 266490
rect 306012 266426 306064 266432
rect 306300 266422 306328 271526
rect 306392 268734 306420 277766
rect 307024 273284 307076 273290
rect 307024 273226 307076 273232
rect 306380 268728 306432 268734
rect 306380 268670 306432 268676
rect 306380 267504 306432 267510
rect 306380 267446 306432 267452
rect 306288 266416 306340 266422
rect 306288 266358 306340 266364
rect 306392 264316 306420 267446
rect 307036 267170 307064 273226
rect 307576 271516 307628 271522
rect 307576 271458 307628 271464
rect 307484 271448 307536 271454
rect 307484 271390 307536 271396
rect 307024 267164 307076 267170
rect 307024 267106 307076 267112
rect 306748 266416 306800 266422
rect 306748 266358 306800 266364
rect 306760 264316 306788 266358
rect 307496 264330 307524 271390
rect 307588 266422 307616 271458
rect 308232 271182 308260 277780
rect 309152 277766 309442 277794
rect 308956 271380 309008 271386
rect 308956 271322 309008 271328
rect 308220 271176 308272 271182
rect 308220 271118 308272 271124
rect 307760 269544 307812 269550
rect 307760 269486 307812 269492
rect 307668 268320 307720 268326
rect 307668 268262 307720 268268
rect 307576 266416 307628 266422
rect 307576 266358 307628 266364
rect 307234 264302 307524 264330
rect 307680 264316 307708 268262
rect 307772 267306 307800 269486
rect 308588 267368 308640 267374
rect 308588 267310 308640 267316
rect 307760 267300 307812 267306
rect 307760 267242 307812 267248
rect 308128 266416 308180 266422
rect 308128 266358 308180 266364
rect 308140 264316 308168 266358
rect 308600 264316 308628 267310
rect 308968 266422 308996 271322
rect 309048 269000 309100 269006
rect 309048 268942 309100 268948
rect 308956 266416 309008 266422
rect 308956 266358 309008 266364
rect 309060 264316 309088 268942
rect 309152 268462 309180 277766
rect 309784 273692 309836 273698
rect 309784 273634 309836 273640
rect 309140 268456 309192 268462
rect 309140 268398 309192 268404
rect 309796 267238 309824 273634
rect 310336 271312 310388 271318
rect 310336 271254 310388 271260
rect 309784 267232 309836 267238
rect 309784 267174 309836 267180
rect 309876 266688 309928 266694
rect 309876 266630 309928 266636
rect 309416 266416 309468 266422
rect 309416 266358 309468 266364
rect 309428 264316 309456 266358
rect 309888 264316 309916 266630
rect 310348 266422 310376 271254
rect 310428 268932 310480 268938
rect 310428 268874 310480 268880
rect 310336 266416 310388 266422
rect 310336 266358 310388 266364
rect 310440 264330 310468 268874
rect 310532 268666 310560 277780
rect 311164 274644 311216 274650
rect 311164 274586 311216 274592
rect 310520 268660 310572 268666
rect 310520 268602 310572 268608
rect 311176 266898 311204 274586
rect 311728 272814 311756 277780
rect 312452 274576 312504 274582
rect 312452 274518 312504 274524
rect 311716 272808 311768 272814
rect 311716 272750 311768 272756
rect 311716 271244 311768 271250
rect 311716 271186 311768 271192
rect 311256 267300 311308 267306
rect 311256 267242 311308 267248
rect 311164 266892 311216 266898
rect 311164 266834 311216 266840
rect 310796 266416 310848 266422
rect 310796 266358 310848 266364
rect 310362 264302 310468 264330
rect 310808 264316 310836 266358
rect 311268 264316 311296 267242
rect 311728 266422 311756 271186
rect 311808 268864 311860 268870
rect 311808 268806 311860 268812
rect 311716 266416 311768 266422
rect 311716 266358 311768 266364
rect 311820 264330 311848 268806
rect 312464 266966 312492 274518
rect 312924 272678 312952 277780
rect 313292 277766 314134 277794
rect 312912 272672 312964 272678
rect 312912 272614 312964 272620
rect 313004 268796 313056 268802
rect 313004 268738 313056 268744
rect 312544 267232 312596 267238
rect 312544 267174 312596 267180
rect 312452 266960 312504 266966
rect 312452 266902 312504 266908
rect 312084 266484 312136 266490
rect 312084 266426 312136 266432
rect 311742 264302 311848 264330
rect 312096 264316 312124 266426
rect 312556 264316 312584 267174
rect 313016 264316 313044 268738
rect 313292 268394 313320 277766
rect 315316 273290 315344 277780
rect 315304 273284 315356 273290
rect 315304 273226 315356 273232
rect 314476 273080 314528 273086
rect 314476 273022 314528 273028
rect 314292 273012 314344 273018
rect 314292 272954 314344 272960
rect 313280 268388 313332 268394
rect 313280 268330 313332 268336
rect 313464 266416 313516 266422
rect 313464 266358 313516 266364
rect 313476 264316 313504 266358
rect 314304 264330 314332 272954
rect 314384 268728 314436 268734
rect 314384 268670 314436 268676
rect 313950 264302 314332 264330
rect 314396 264316 314424 268670
rect 314488 266422 314516 273022
rect 315856 272944 315908 272950
rect 315856 272886 315908 272892
rect 315304 271176 315356 271182
rect 315304 271118 315356 271124
rect 315212 267164 315264 267170
rect 315212 267106 315264 267112
rect 314476 266416 314528 266422
rect 314476 266358 314528 266364
rect 314844 266416 314896 266422
rect 314844 266358 314896 266364
rect 314856 264316 314884 266358
rect 315224 264316 315252 267106
rect 315316 266490 315344 271118
rect 315672 268660 315724 268666
rect 315672 268602 315724 268608
rect 315304 266484 315356 266490
rect 315304 266426 315356 266432
rect 315684 264316 315712 268602
rect 315868 266422 315896 272886
rect 316512 272542 316540 277780
rect 316684 273760 316736 273766
rect 316684 273702 316736 273708
rect 316500 272536 316552 272542
rect 316500 272478 316552 272484
rect 316696 267102 316724 273702
rect 317236 272876 317288 272882
rect 317236 272818 317288 272824
rect 317052 268592 317104 268598
rect 317052 268534 317104 268540
rect 316684 267096 316736 267102
rect 316684 267038 316736 267044
rect 316592 266484 316644 266490
rect 316592 266426 316644 266432
rect 315856 266416 315908 266422
rect 315856 266358 315908 266364
rect 316132 266416 316184 266422
rect 316132 266358 316184 266364
rect 316144 264316 316172 266358
rect 316604 264316 316632 266426
rect 317064 264316 317092 268534
rect 317248 266422 317276 272818
rect 317708 272610 317736 277780
rect 318812 274310 318840 277780
rect 318800 274304 318852 274310
rect 318800 274246 318852 274252
rect 319444 273828 319496 273834
rect 319444 273770 319496 273776
rect 318616 272740 318668 272746
rect 318616 272682 318668 272688
rect 317696 272604 317748 272610
rect 317696 272546 317748 272552
rect 318340 268524 318392 268530
rect 318340 268466 318392 268472
rect 317880 267096 317932 267102
rect 317880 267038 317932 267044
rect 317236 266416 317288 266422
rect 317236 266358 317288 266364
rect 317512 266416 317564 266422
rect 317512 266358 317564 266364
rect 317524 264316 317552 266358
rect 317892 264316 317920 267038
rect 318352 264316 318380 268466
rect 318628 266422 318656 272682
rect 319456 267034 319484 273770
rect 320008 273222 320036 277780
rect 320824 274508 320876 274514
rect 320824 274450 320876 274456
rect 319996 273216 320048 273222
rect 319996 273158 320048 273164
rect 319996 272672 320048 272678
rect 319996 272614 320048 272620
rect 319720 268456 319772 268462
rect 319720 268398 319772 268404
rect 319444 267028 319496 267034
rect 319444 266970 319496 266976
rect 319260 266552 319312 266558
rect 319260 266494 319312 266500
rect 318616 266416 318668 266422
rect 318616 266358 318668 266364
rect 318800 266416 318852 266422
rect 318800 266358 318852 266364
rect 318812 264316 318840 266358
rect 319272 264316 319300 266494
rect 319732 264316 319760 268398
rect 320008 266422 320036 272614
rect 320836 267714 320864 274450
rect 321204 273154 321232 277780
rect 322204 274304 322256 274310
rect 322204 274246 322256 274252
rect 321192 273148 321244 273154
rect 321192 273090 321244 273096
rect 321376 272604 321428 272610
rect 321376 272546 321428 272552
rect 320824 267708 320876 267714
rect 320824 267650 320876 267656
rect 320548 267028 320600 267034
rect 320548 266970 320600 266976
rect 319996 266416 320048 266422
rect 319996 266358 320048 266364
rect 320180 266416 320232 266422
rect 320180 266358 320232 266364
rect 320192 264316 320220 266358
rect 320560 264316 320588 266970
rect 321008 266960 321060 266966
rect 321008 266902 321060 266908
rect 321020 264316 321048 266902
rect 321388 266422 321416 272546
rect 321468 272536 321520 272542
rect 321468 272478 321520 272484
rect 321376 266416 321428 266422
rect 321376 266358 321428 266364
rect 321480 264316 321508 272478
rect 321928 269816 321980 269822
rect 321928 269758 321980 269764
rect 321940 264316 321968 269758
rect 322216 266830 322244 274246
rect 322400 273698 322428 277780
rect 323596 273902 323624 277780
rect 324792 274378 324820 277780
rect 324780 274372 324832 274378
rect 324780 274314 324832 274320
rect 325988 274242 326016 277780
rect 326988 276344 327040 276350
rect 326988 276286 327040 276292
rect 325976 274236 326028 274242
rect 325976 274178 326028 274184
rect 323584 273896 323636 273902
rect 323584 273838 323636 273844
rect 322388 273692 322440 273698
rect 322388 273634 322440 273640
rect 324964 273488 325016 273494
rect 324964 273430 325016 273436
rect 322664 272808 322716 272814
rect 322664 272750 322716 272756
rect 322296 270972 322348 270978
rect 322296 270914 322348 270920
rect 322308 267646 322336 270914
rect 322388 268388 322440 268394
rect 322388 268330 322440 268336
rect 322296 267640 322348 267646
rect 322296 267582 322348 267588
rect 322204 266824 322256 266830
rect 322204 266766 322256 266772
rect 322400 264316 322428 268330
rect 322676 264330 322704 272750
rect 324136 272128 324188 272134
rect 324136 272070 324188 272076
rect 323584 269272 323636 269278
rect 323584 269214 323636 269220
rect 323216 269068 323268 269074
rect 323216 269010 323268 269016
rect 322676 264302 322874 264330
rect 323228 264316 323256 269010
rect 323596 266694 323624 269214
rect 323676 267640 323728 267646
rect 323676 267582 323728 267588
rect 323584 266688 323636 266694
rect 323584 266630 323636 266636
rect 323688 264316 323716 267582
rect 324148 264316 324176 272070
rect 324976 266558 325004 273430
rect 325608 272196 325660 272202
rect 325608 272138 325660 272144
rect 324964 266552 325016 266558
rect 324964 266494 325016 266500
rect 324596 266416 324648 266422
rect 324596 266358 324648 266364
rect 324608 264316 324636 266358
rect 325056 265192 325108 265198
rect 325056 265134 325108 265140
rect 325068 264316 325096 265134
rect 325620 264330 325648 272138
rect 326344 271040 326396 271046
rect 326344 270982 326396 270988
rect 326356 267578 326384 270982
rect 326896 270700 326948 270706
rect 326896 270642 326948 270648
rect 326344 267572 326396 267578
rect 326344 267514 326396 267520
rect 325976 266824 326028 266830
rect 325976 266766 326028 266772
rect 325542 264302 325648 264330
rect 325988 264316 326016 266766
rect 326344 266552 326396 266558
rect 326344 266494 326396 266500
rect 326356 264316 326384 266494
rect 326908 264330 326936 270642
rect 327000 266558 327028 276286
rect 327092 269550 327120 277780
rect 328288 274174 328316 277780
rect 329484 274446 329512 277780
rect 329852 277766 330694 277794
rect 329748 276412 329800 276418
rect 329748 276354 329800 276360
rect 329472 274440 329524 274446
rect 329472 274382 329524 274388
rect 328276 274168 328328 274174
rect 328276 274110 328328 274116
rect 329104 272264 329156 272270
rect 329104 272206 329156 272212
rect 328368 272060 328420 272066
rect 328368 272002 328420 272008
rect 327080 269544 327132 269550
rect 327080 269486 327132 269492
rect 328184 266620 328236 266626
rect 328184 266562 328236 266568
rect 326988 266552 327040 266558
rect 326988 266494 327040 266500
rect 327264 266552 327316 266558
rect 327264 266494 327316 266500
rect 326830 264302 326936 264330
rect 327276 264316 327304 266494
rect 327724 265260 327776 265266
rect 327724 265202 327776 265208
rect 327736 264316 327764 265202
rect 328196 264316 328224 266562
rect 328380 266558 328408 272002
rect 328644 266756 328696 266762
rect 328644 266698 328696 266704
rect 328368 266552 328420 266558
rect 328368 266494 328420 266500
rect 328656 264316 328684 266698
rect 329116 266626 329144 272206
rect 329656 270768 329708 270774
rect 329656 270710 329708 270716
rect 329104 266620 329156 266626
rect 329104 266562 329156 266568
rect 329012 266552 329064 266558
rect 329012 266494 329064 266500
rect 329024 264316 329052 266494
rect 329668 264330 329696 270710
rect 329760 266558 329788 276354
rect 329852 269618 329880 277766
rect 330760 276480 330812 276486
rect 330760 276422 330812 276428
rect 330668 274984 330720 274990
rect 330668 274926 330720 274932
rect 329840 269612 329892 269618
rect 329840 269554 329892 269560
rect 330680 266558 330708 274926
rect 329748 266552 329800 266558
rect 329748 266494 329800 266500
rect 329932 266552 329984 266558
rect 329932 266494 329984 266500
rect 330668 266552 330720 266558
rect 330668 266494 330720 266500
rect 329498 264302 329696 264330
rect 329944 264316 329972 266494
rect 330772 264330 330800 276422
rect 331876 273766 331904 277780
rect 333072 274650 333100 277780
rect 333992 277766 334190 277794
rect 333888 276548 333940 276554
rect 333888 276490 333940 276496
rect 333796 275460 333848 275466
rect 333796 275402 333848 275408
rect 333060 274644 333112 274650
rect 333060 274586 333112 274592
rect 331864 273760 331916 273766
rect 331864 273702 331916 273708
rect 332508 272332 332560 272338
rect 332508 272274 332560 272280
rect 331128 268048 331180 268054
rect 331128 267990 331180 267996
rect 331140 267646 331168 267990
rect 331128 267640 331180 267646
rect 331128 267582 331180 267588
rect 330852 267572 330904 267578
rect 330852 267514 330904 267520
rect 330418 264302 330800 264330
rect 330864 264316 330892 267514
rect 331312 266892 331364 266898
rect 331312 266834 331364 266840
rect 331324 264316 331352 266834
rect 331680 265328 331732 265334
rect 331680 265270 331732 265276
rect 331692 264316 331720 265270
rect 332520 264330 332548 272274
rect 333808 266626 333836 275402
rect 332600 266620 332652 266626
rect 332600 266562 332652 266568
rect 333796 266620 333848 266626
rect 333796 266562 333848 266568
rect 332166 264302 332548 264330
rect 332612 264316 332640 266562
rect 333900 266558 333928 276490
rect 333992 269686 334020 277766
rect 335268 276616 335320 276622
rect 335268 276558 335320 276564
rect 335176 275052 335228 275058
rect 335176 274994 335228 275000
rect 333980 269680 334032 269686
rect 333980 269622 334032 269628
rect 334072 266824 334124 266830
rect 334072 266766 334124 266772
rect 334808 266824 334860 266830
rect 334808 266766 334860 266772
rect 334084 266558 334112 266766
rect 334256 266756 334308 266762
rect 334256 266698 334308 266704
rect 333060 266552 333112 266558
rect 333060 266494 333112 266500
rect 333888 266552 333940 266558
rect 333888 266494 333940 266500
rect 334072 266552 334124 266558
rect 334072 266494 334124 266500
rect 333072 264316 333100 266494
rect 333520 265396 333572 265402
rect 333520 265338 333572 265344
rect 333532 264316 333560 265338
rect 334268 264330 334296 266698
rect 334348 265464 334400 265470
rect 334348 265406 334400 265412
rect 334006 264302 334296 264330
rect 334360 264316 334388 265406
rect 334820 264316 334848 266766
rect 335188 264330 335216 274994
rect 335280 266830 335308 276558
rect 335372 270502 335400 277780
rect 336568 274582 336596 277780
rect 336752 277766 337778 277794
rect 336556 274576 336608 274582
rect 336556 274518 336608 274524
rect 336004 271108 336056 271114
rect 336004 271050 336056 271056
rect 335360 270496 335412 270502
rect 335360 270438 335412 270444
rect 335728 269340 335780 269346
rect 335728 269282 335780 269288
rect 335360 268116 335412 268122
rect 335360 268058 335412 268064
rect 335372 267510 335400 268058
rect 335360 267504 335412 267510
rect 335360 267446 335412 267452
rect 335268 266824 335320 266830
rect 335268 266766 335320 266772
rect 335188 264302 335294 264330
rect 335740 264316 335768 269282
rect 336016 267442 336044 271050
rect 336752 269754 336780 277766
rect 337844 275188 337896 275194
rect 337844 275130 337896 275136
rect 336740 269748 336792 269754
rect 336740 269690 336792 269696
rect 337108 269408 337160 269414
rect 337108 269350 337160 269356
rect 336004 267436 336056 267442
rect 336004 267378 336056 267384
rect 336648 266892 336700 266898
rect 336648 266834 336700 266840
rect 336188 265532 336240 265538
rect 336188 265474 336240 265480
rect 336200 264316 336228 265474
rect 336660 264316 336688 266834
rect 337120 264316 337148 269350
rect 337476 266824 337528 266830
rect 337476 266766 337528 266772
rect 337488 264316 337516 266766
rect 337856 264330 337884 275130
rect 338960 273834 338988 277780
rect 339408 277636 339460 277642
rect 339408 277578 339460 277584
rect 338948 273828 339000 273834
rect 338948 273770 339000 273776
rect 337936 270836 337988 270842
rect 337936 270778 337988 270784
rect 337948 266830 337976 270778
rect 338396 269476 338448 269482
rect 338396 269418 338448 269424
rect 337936 266824 337988 266830
rect 337936 266766 337988 266772
rect 337856 264302 337962 264330
rect 338408 264316 338436 269418
rect 339420 267734 339448 277578
rect 340156 271862 340184 277780
rect 340892 277766 341366 277794
rect 340604 275256 340656 275262
rect 340604 275198 340656 275204
rect 340144 271856 340196 271862
rect 340144 271798 340196 271804
rect 339776 269544 339828 269550
rect 339776 269486 339828 269492
rect 339236 267706 339448 267734
rect 339236 264330 339264 267706
rect 339316 267436 339368 267442
rect 339316 267378 339368 267384
rect 338882 264302 339264 264330
rect 339328 264316 339356 267378
rect 339788 264316 339816 269486
rect 340144 266824 340196 266830
rect 340144 266766 340196 266772
rect 340156 264316 340184 266766
rect 340616 264316 340644 275198
rect 340696 273556 340748 273562
rect 340696 273498 340748 273504
rect 340708 266830 340736 273498
rect 340892 270434 340920 277766
rect 342456 274106 342484 277780
rect 343364 275868 343416 275874
rect 343364 275810 343416 275816
rect 342444 274100 342496 274106
rect 342444 274042 342496 274048
rect 341892 273624 341944 273630
rect 341892 273566 341944 273572
rect 340880 270428 340932 270434
rect 340880 270370 340932 270376
rect 341064 269612 341116 269618
rect 341064 269554 341116 269560
rect 340696 266824 340748 266830
rect 340696 266766 340748 266772
rect 341076 264316 341104 269554
rect 341904 264330 341932 273566
rect 342444 269680 342496 269686
rect 342444 269622 342496 269628
rect 342168 267912 342220 267918
rect 342168 267854 342220 267860
rect 341984 267708 342036 267714
rect 341984 267650 342036 267656
rect 341550 264302 341932 264330
rect 341996 264316 342024 267650
rect 342180 266966 342208 267854
rect 342168 266960 342220 266966
rect 342168 266902 342220 266908
rect 342456 264316 342484 269622
rect 342812 266824 342864 266830
rect 342812 266766 342864 266772
rect 342824 264316 342852 266766
rect 343376 264330 343404 275810
rect 343456 273692 343508 273698
rect 343456 273634 343508 273640
rect 343468 266830 343496 273634
rect 343652 271794 343680 277780
rect 343836 277766 344862 277794
rect 345032 277766 346058 277794
rect 343640 271788 343692 271794
rect 343640 271730 343692 271736
rect 343836 270162 343864 277766
rect 344560 273760 344612 273766
rect 344560 273702 344612 273708
rect 344284 270632 344336 270638
rect 344284 270574 344336 270580
rect 343824 270156 343876 270162
rect 343824 270098 343876 270104
rect 344008 270156 344060 270162
rect 344008 270098 344060 270104
rect 343456 266824 343508 266830
rect 343456 266766 343508 266772
rect 344020 264330 344048 270098
rect 344296 267374 344324 270574
rect 344284 267368 344336 267374
rect 344284 267310 344336 267316
rect 344572 264330 344600 273702
rect 345032 270366 345060 277766
rect 346124 276004 346176 276010
rect 346124 275946 346176 275952
rect 345020 270360 345072 270366
rect 345020 270302 345072 270308
rect 345112 269748 345164 269754
rect 345112 269690 345164 269696
rect 344652 266892 344704 266898
rect 344652 266834 344704 266840
rect 343298 264302 343404 264330
rect 343758 264302 344048 264330
rect 344218 264302 344600 264330
rect 344664 264316 344692 266834
rect 345124 264316 345152 269690
rect 345480 266960 345532 266966
rect 345480 266902 345532 266908
rect 345492 264316 345520 266902
rect 346136 264330 346164 275946
rect 346216 273828 346268 273834
rect 346216 273770 346268 273776
rect 346228 266966 346256 273770
rect 347240 270978 347268 277780
rect 347792 277766 348450 277794
rect 347688 273896 347740 273902
rect 347688 273838 347740 273844
rect 347228 270972 347280 270978
rect 347228 270914 347280 270920
rect 346768 270496 346820 270502
rect 346768 270438 346820 270444
rect 346400 267368 346452 267374
rect 346400 267310 346452 267316
rect 346216 266960 346268 266966
rect 346216 266902 346268 266908
rect 346412 266898 346440 267310
rect 346400 266892 346452 266898
rect 346400 266834 346452 266840
rect 346780 264330 346808 270438
rect 347320 267640 347372 267646
rect 347320 267582 347372 267588
rect 346860 267368 346912 267374
rect 346860 267310 346912 267316
rect 345966 264302 346164 264330
rect 346426 264302 346808 264330
rect 346872 264316 346900 267310
rect 347332 264316 347360 267582
rect 347700 267374 347728 273838
rect 347792 270298 347820 277766
rect 348792 275936 348844 275942
rect 348792 275878 348844 275884
rect 348056 270428 348108 270434
rect 348056 270370 348108 270376
rect 347780 270292 347832 270298
rect 347780 270234 347832 270240
rect 347688 267368 347740 267374
rect 347688 267310 347740 267316
rect 348068 264330 348096 270370
rect 348240 267368 348292 267374
rect 348240 267310 348292 267316
rect 347806 264302 348096 264330
rect 348252 264316 348280 267310
rect 348804 264330 348832 275878
rect 349632 274514 349660 277780
rect 350448 274644 350500 274650
rect 350448 274586 350500 274592
rect 349620 274508 349672 274514
rect 349620 274450 349672 274456
rect 348976 274168 349028 274174
rect 348976 274110 349028 274116
rect 348988 267374 349016 274110
rect 349068 270360 349120 270366
rect 349068 270302 349120 270308
rect 348976 267368 349028 267374
rect 348976 267310 349028 267316
rect 348634 264302 348832 264330
rect 349080 264316 349108 270302
rect 350262 270192 350318 270201
rect 350262 270127 350318 270136
rect 349988 267504 350040 267510
rect 349988 267446 350040 267452
rect 349528 267368 349580 267374
rect 349528 267310 349580 267316
rect 349540 264316 349568 267310
rect 350000 264316 350028 267446
rect 350276 264330 350304 270127
rect 350354 268968 350410 268977
rect 350354 268903 350410 268912
rect 350368 267578 350396 268903
rect 350356 267572 350408 267578
rect 350356 267514 350408 267520
rect 350460 267374 350488 274586
rect 350736 271046 350764 277780
rect 351828 277364 351880 277370
rect 351828 277306 351880 277312
rect 351736 274576 351788 274582
rect 351736 274518 351788 274524
rect 350724 271040 350776 271046
rect 350724 270982 350776 270988
rect 351644 270564 351696 270570
rect 351644 270506 351696 270512
rect 350448 267368 350500 267374
rect 350448 267310 350500 267316
rect 350908 267368 350960 267374
rect 350908 267310 350960 267316
rect 350276 264302 350474 264330
rect 350920 264316 350948 267310
rect 351656 264330 351684 270506
rect 351748 267374 351776 274518
rect 351736 267368 351788 267374
rect 351736 267310 351788 267316
rect 351840 264330 351868 277306
rect 351932 270230 351960 277780
rect 353128 274038 353156 277780
rect 353208 274508 353260 274514
rect 353208 274450 353260 274456
rect 353116 274032 353168 274038
rect 353116 273974 353168 273980
rect 351920 270224 351972 270230
rect 351920 270166 351972 270172
rect 352656 267504 352708 267510
rect 352656 267446 352708 267452
rect 352196 267368 352248 267374
rect 352196 267310 352248 267316
rect 351302 264302 351684 264330
rect 351762 264302 351868 264330
rect 352208 264316 352236 267310
rect 352668 264316 352696 267446
rect 353220 267374 353248 274450
rect 354324 271726 354352 277780
rect 354692 277766 355534 277794
rect 354588 277296 354640 277302
rect 354588 277238 354640 277244
rect 354496 275800 354548 275806
rect 354496 275742 354548 275748
rect 354404 274440 354456 274446
rect 354404 274382 354456 274388
rect 354312 271720 354364 271726
rect 354312 271662 354364 271668
rect 354416 267374 354444 274382
rect 353208 267368 353260 267374
rect 353208 267310 353260 267316
rect 353576 267368 353628 267374
rect 353576 267310 353628 267316
rect 354404 267368 354456 267374
rect 354404 267310 354456 267316
rect 353116 265600 353168 265606
rect 353116 265542 353168 265548
rect 353128 264316 353156 265542
rect 353588 264316 353616 267310
rect 354508 264602 354536 275742
rect 354324 264574 354536 264602
rect 354324 264330 354352 264574
rect 354600 264330 354628 277238
rect 354692 270094 354720 277766
rect 355968 274372 356020 274378
rect 355968 274314 356020 274320
rect 354680 270088 354732 270094
rect 354680 270030 354732 270036
rect 354680 267844 354732 267850
rect 354680 267786 354732 267792
rect 354692 266422 354720 267786
rect 355324 267436 355376 267442
rect 355324 267378 355376 267384
rect 354680 266416 354732 266422
rect 354680 266358 354732 266364
rect 354864 266416 354916 266422
rect 354864 266358 354916 266364
rect 353970 264302 354352 264330
rect 354430 264302 354628 264330
rect 354876 264316 354904 266358
rect 355336 264316 355364 267378
rect 355980 266422 356008 274314
rect 356716 274310 356744 277780
rect 357452 277766 357926 277794
rect 358832 277766 359030 277794
rect 360226 277766 360332 277794
rect 357348 277228 357400 277234
rect 357348 277170 357400 277176
rect 357256 275732 357308 275738
rect 357256 275674 357308 275680
rect 356704 274304 356756 274310
rect 356704 274246 356756 274252
rect 357164 274304 357216 274310
rect 357164 274246 357216 274252
rect 357176 266422 357204 274246
rect 355968 266416 356020 266422
rect 355968 266358 356020 266364
rect 356244 266416 356296 266422
rect 356244 266358 356296 266364
rect 357164 266416 357216 266422
rect 357164 266358 357216 266364
rect 355784 266348 355836 266354
rect 355784 266290 355836 266296
rect 355796 264316 355824 266290
rect 356256 264316 356284 266358
rect 357268 264602 357296 275674
rect 356992 264574 357296 264602
rect 356992 264330 357020 264574
rect 357360 264330 357388 277170
rect 357452 268190 357480 277766
rect 357532 270292 357584 270298
rect 357532 270234 357584 270240
rect 357440 268184 357492 268190
rect 357440 268126 357492 268132
rect 356638 264302 357020 264330
rect 357098 264302 357388 264330
rect 357544 264316 357572 270234
rect 358832 270026 358860 277766
rect 360108 277160 360160 277166
rect 360108 277102 360160 277108
rect 360016 275664 360068 275670
rect 360016 275606 360068 275612
rect 359924 272400 359976 272406
rect 359924 272342 359976 272348
rect 358820 270020 358872 270026
rect 358820 269962 358872 269968
rect 357990 267472 358046 267481
rect 357990 267407 358046 267416
rect 358004 264316 358032 267407
rect 359936 266422 359964 272342
rect 358912 266416 358964 266422
rect 358912 266358 358964 266364
rect 359924 266416 359976 266422
rect 359924 266358 359976 266364
rect 358452 266280 358504 266286
rect 358452 266222 358504 266228
rect 358464 264316 358492 266222
rect 358924 264316 358952 266358
rect 360028 264602 360056 275606
rect 359660 264574 360056 264602
rect 359660 264330 359688 264574
rect 360120 264330 360148 277102
rect 360200 270224 360252 270230
rect 360200 270166 360252 270172
rect 359398 264302 359688 264330
rect 359766 264302 360148 264330
rect 360212 264316 360240 270166
rect 360304 269958 360332 277766
rect 360396 277766 361422 277794
rect 360292 269952 360344 269958
rect 360292 269894 360344 269900
rect 360396 268258 360424 277766
rect 362316 275596 362368 275602
rect 362316 275538 362368 275544
rect 360384 268252 360436 268258
rect 360384 268194 360436 268200
rect 361488 268184 361540 268190
rect 361488 268126 361540 268132
rect 360660 267368 360712 267374
rect 360660 267310 360712 267316
rect 360672 264316 360700 267310
rect 361500 267306 361528 268126
rect 361488 267300 361540 267306
rect 361488 267242 361540 267248
rect 361856 267232 361908 267238
rect 361856 267174 361908 267180
rect 361120 266212 361172 266218
rect 361120 266154 361172 266160
rect 361132 264316 361160 266154
rect 361868 264330 361896 267174
rect 362328 264330 362356 275538
rect 362604 271658 362632 277780
rect 362776 274236 362828 274242
rect 362776 274178 362828 274184
rect 362684 272468 362736 272474
rect 362684 272410 362736 272416
rect 362592 271652 362644 271658
rect 362592 271594 362644 271600
rect 362696 267238 362724 272410
rect 362684 267232 362736 267238
rect 362684 267174 362736 267180
rect 362408 266416 362460 266422
rect 362408 266358 362460 266364
rect 361606 264302 361896 264330
rect 362066 264302 362356 264330
rect 362420 264316 362448 266358
rect 362788 264330 362816 274178
rect 363800 273970 363828 277780
rect 363788 273964 363840 273970
rect 363788 273906 363840 273912
rect 364248 273216 364300 273222
rect 364248 273158 364300 273164
rect 364156 270972 364208 270978
rect 364156 270914 364208 270920
rect 362868 270904 362920 270910
rect 362868 270846 362920 270852
rect 362880 266422 362908 270846
rect 362960 268252 363012 268258
rect 362960 268194 363012 268200
rect 362972 267306 363000 268194
rect 362960 267300 363012 267306
rect 362960 267242 363012 267248
rect 363328 267300 363380 267306
rect 363328 267242 363380 267248
rect 362868 266416 362920 266422
rect 362868 266358 362920 266364
rect 362788 264302 362894 264330
rect 363340 264316 363368 267242
rect 364168 264330 364196 270914
rect 363814 264302 364196 264330
rect 364260 264316 364288 273158
rect 364996 271114 365024 277780
rect 365444 275528 365496 275534
rect 365444 275470 365496 275476
rect 364984 271108 365036 271114
rect 364984 271050 365036 271056
rect 365456 266422 365484 275470
rect 366100 271590 366128 277780
rect 367112 277766 367310 277794
rect 366088 271584 366140 271590
rect 366088 271526 366140 271532
rect 366824 271108 366876 271114
rect 366824 271050 366876 271056
rect 365536 271040 365588 271046
rect 365536 270982 365588 270988
rect 364708 266416 364760 266422
rect 364708 266358 364760 266364
rect 365444 266416 365496 266422
rect 365444 266358 365496 266364
rect 364720 264316 364748 266358
rect 365548 264738 365576 270982
rect 365628 270088 365680 270094
rect 365628 270030 365680 270036
rect 365456 264710 365576 264738
rect 365456 264330 365484 264710
rect 365640 264330 365668 270030
rect 365994 267336 366050 267345
rect 365994 267271 366050 267280
rect 365102 264302 365484 264330
rect 365562 264302 365668 264330
rect 366008 264316 366036 267271
rect 366836 264330 366864 271050
rect 367112 269890 367140 277766
rect 368386 275496 368442 275505
rect 368386 275431 368442 275440
rect 368112 271856 368164 271862
rect 368112 271798 368164 271804
rect 367100 269884 367152 269890
rect 367100 269826 367152 269832
rect 368020 267232 368072 267238
rect 368020 267174 368072 267180
rect 368032 266490 368060 267174
rect 368020 266484 368072 266490
rect 368020 266426 368072 266432
rect 367376 266416 367428 266422
rect 367376 266358 367428 266364
rect 367008 264512 367060 264518
rect 367008 264454 367060 264460
rect 367020 264330 367048 264454
rect 366482 264302 366864 264330
rect 366942 264302 367048 264330
rect 367388 264316 367416 266358
rect 368124 264330 368152 271798
rect 368202 268832 368258 268841
rect 368202 268767 368258 268776
rect 367770 264302 368152 264330
rect 368216 264316 368244 268767
rect 368400 266422 368428 275431
rect 368492 268122 368520 277780
rect 369320 277766 369702 277794
rect 369320 271522 369348 277766
rect 369768 273148 369820 273154
rect 369768 273090 369820 273096
rect 369492 271788 369544 271794
rect 369492 271730 369544 271736
rect 369308 271516 369360 271522
rect 369308 271458 369360 271464
rect 368480 268116 368532 268122
rect 368480 268058 368532 268064
rect 368664 266484 368716 266490
rect 368664 266426 368716 266432
rect 368388 266416 368440 266422
rect 368388 266358 368440 266364
rect 368676 264316 368704 266426
rect 369504 264330 369532 271730
rect 369676 267776 369728 267782
rect 369676 267718 369728 267724
rect 369688 267170 369716 267718
rect 369676 267164 369728 267170
rect 369676 267106 369728 267112
rect 369780 264330 369808 273090
rect 370780 271720 370832 271726
rect 370780 271662 370832 271668
rect 370044 266416 370096 266422
rect 370044 266358 370096 266364
rect 369150 264302 369532 264330
rect 369610 264302 369808 264330
rect 370056 264316 370084 266358
rect 370792 264330 370820 271662
rect 370884 271454 370912 277780
rect 371252 277766 372094 277794
rect 371146 275360 371202 275369
rect 371146 275295 371202 275304
rect 371056 274100 371108 274106
rect 371056 274042 371108 274048
rect 370872 271448 370924 271454
rect 370872 271390 370924 271396
rect 371068 264330 371096 274042
rect 371160 266422 371188 275295
rect 371252 268326 371280 277766
rect 372160 271652 372212 271658
rect 372160 271594 372212 271600
rect 371240 268320 371292 268326
rect 371240 268262 371292 268268
rect 371884 268320 371936 268326
rect 371884 268262 371936 268268
rect 371332 267232 371384 267238
rect 371332 267174 371384 267180
rect 371148 266416 371200 266422
rect 371148 266358 371200 266364
rect 370530 264302 370820 264330
rect 370898 264302 371096 264330
rect 371344 264316 371372 267174
rect 371896 267170 371924 268262
rect 371884 267164 371936 267170
rect 371884 267106 371936 267112
rect 372172 264330 372200 271594
rect 373276 271386 373304 277780
rect 373906 275224 373962 275233
rect 373906 275159 373962 275168
rect 373816 271584 373868 271590
rect 373816 271526 373868 271532
rect 373264 271380 373316 271386
rect 373264 271322 373316 271328
rect 372252 270020 372304 270026
rect 372252 269962 372304 269968
rect 371818 264302 372200 264330
rect 372264 264316 372292 269962
rect 372712 266416 372764 266422
rect 372712 266358 372764 266364
rect 372724 264316 372752 266358
rect 373172 266144 373224 266150
rect 373172 266086 373224 266092
rect 373184 264316 373212 266086
rect 373828 264330 373856 271526
rect 373920 266422 373948 275159
rect 374380 270638 374408 277780
rect 375392 277766 375590 277794
rect 375288 271516 375340 271522
rect 375288 271458 375340 271464
rect 374368 270632 374420 270638
rect 374368 270574 374420 270580
rect 374368 269952 374420 269958
rect 374368 269894 374420 269900
rect 373908 266416 373960 266422
rect 373908 266358 373960 266364
rect 374380 264330 374408 269894
rect 374460 266076 374512 266082
rect 374460 266018 374512 266024
rect 373566 264302 373856 264330
rect 374026 264302 374408 264330
rect 374472 264316 374500 266018
rect 375300 264330 375328 271458
rect 375392 269006 375420 277766
rect 375932 275120 375984 275126
rect 375932 275062 375984 275068
rect 375656 274032 375708 274038
rect 375656 273974 375708 273980
rect 375380 269000 375432 269006
rect 375380 268942 375432 268948
rect 375668 264330 375696 273974
rect 375944 270570 375972 275062
rect 376576 271448 376628 271454
rect 376576 271390 376628 271396
rect 376484 271380 376536 271386
rect 376484 271322 376536 271328
rect 375932 270564 375984 270570
rect 375932 270506 375984 270512
rect 376208 266416 376260 266422
rect 376208 266358 376260 266364
rect 375840 266008 375892 266014
rect 375840 265950 375892 265956
rect 374946 264302 375328 264330
rect 375406 264302 375696 264330
rect 375852 264316 375880 265950
rect 376220 264316 376248 266358
rect 376496 264330 376524 271322
rect 376588 266422 376616 271390
rect 376772 271318 376800 277780
rect 376956 277766 377982 277794
rect 378152 277766 379178 277794
rect 376760 271312 376812 271318
rect 376760 271254 376812 271260
rect 376956 269278 376984 277766
rect 377956 271312 378008 271318
rect 377956 271254 378008 271260
rect 376944 269272 376996 269278
rect 376944 269214 376996 269220
rect 376576 266416 376628 266422
rect 376576 266358 376628 266364
rect 377128 265940 377180 265946
rect 377128 265882 377180 265888
rect 376496 264302 376694 264330
rect 377140 264316 377168 265882
rect 377968 264330 377996 271254
rect 378048 269884 378100 269890
rect 378048 269826 378100 269832
rect 377614 264302 377996 264330
rect 378060 264316 378088 269826
rect 378152 268938 378180 277766
rect 379428 273964 379480 273970
rect 379428 273906 379480 273912
rect 379242 271416 379298 271425
rect 379242 271351 379298 271360
rect 378140 268932 378192 268938
rect 378140 268874 378192 268880
rect 378784 267232 378836 267238
rect 378784 267174 378836 267180
rect 378796 266490 378824 267174
rect 378784 266484 378836 266490
rect 378784 266426 378836 266432
rect 378508 265872 378560 265878
rect 378508 265814 378560 265820
rect 378520 264316 378548 265814
rect 379256 264330 379284 271351
rect 379440 264330 379468 273906
rect 380360 271250 380388 277780
rect 380912 277766 381570 277794
rect 382292 277766 382674 277794
rect 380348 271244 380400 271250
rect 380348 271186 380400 271192
rect 380624 271244 380676 271250
rect 380624 271186 380676 271192
rect 379796 265804 379848 265810
rect 379796 265746 379848 265752
rect 378902 264302 379284 264330
rect 379362 264302 379468 264330
rect 379808 264316 379836 265746
rect 380636 264330 380664 271186
rect 380912 268190 380940 277766
rect 382004 277024 382056 277030
rect 382004 276966 382056 276972
rect 380900 268184 380952 268190
rect 380900 268126 380952 268132
rect 380714 267064 380770 267073
rect 380714 266999 380770 267008
rect 380282 264302 380664 264330
rect 380728 264316 380756 266999
rect 382016 266422 382044 276966
rect 382094 271280 382150 271289
rect 382094 271215 382150 271224
rect 381176 266416 381228 266422
rect 381176 266358 381228 266364
rect 382004 266416 382056 266422
rect 382004 266358 382056 266364
rect 381188 264316 381216 266358
rect 382108 264602 382136 271215
rect 382188 268932 382240 268938
rect 382188 268874 382240 268880
rect 381924 264574 382136 264602
rect 381924 264330 381952 264574
rect 382200 264330 382228 268874
rect 382292 268870 382320 277766
rect 383856 271182 383884 277780
rect 385066 277766 385172 277794
rect 384948 277092 385000 277098
rect 384948 277034 385000 277040
rect 384580 276956 384632 276962
rect 384580 276898 384632 276904
rect 383844 271176 383896 271182
rect 383290 271144 383346 271153
rect 383844 271118 383896 271124
rect 383290 271079 383346 271088
rect 382280 268864 382332 268870
rect 382280 268806 382332 268812
rect 382464 265736 382516 265742
rect 382464 265678 382516 265684
rect 381662 264302 381952 264330
rect 382030 264302 382228 264330
rect 382476 264316 382504 265678
rect 383304 264330 383332 271079
rect 383382 270056 383438 270065
rect 383382 269991 383438 270000
rect 382950 264302 383332 264330
rect 383396 264316 383424 269991
rect 383844 266416 383896 266422
rect 383844 266358 383896 266364
rect 383856 264316 383884 266358
rect 384592 264330 384620 276898
rect 384960 266422 384988 277034
rect 385144 268258 385172 277766
rect 385236 277766 386262 277794
rect 385236 268802 385264 277766
rect 387248 276888 387300 276894
rect 387248 276830 387300 276836
rect 386234 273864 386290 273873
rect 386234 273799 386290 273808
rect 385224 268796 385276 268802
rect 385224 268738 385276 268744
rect 385132 268252 385184 268258
rect 385132 268194 385184 268200
rect 385132 267980 385184 267986
rect 385132 267922 385184 267928
rect 384948 266416 385000 266422
rect 384948 266358 385000 266364
rect 384948 264444 385000 264450
rect 384948 264386 385000 264392
rect 384960 264330 384988 264386
rect 384330 264302 384620 264330
rect 384698 264302 384988 264330
rect 385144 264316 385172 267922
rect 385592 265668 385644 265674
rect 385592 265610 385644 265616
rect 385604 264316 385632 265610
rect 386248 264330 386276 273799
rect 387064 271924 387116 271930
rect 387064 271866 387116 271872
rect 386512 268116 386564 268122
rect 386512 268058 386564 268064
rect 386078 264302 386276 264330
rect 386524 264316 386552 268058
rect 387076 267102 387104 271866
rect 387064 267096 387116 267102
rect 387064 267038 387116 267044
rect 387260 264330 387288 276830
rect 387444 273086 387472 277780
rect 387432 273080 387484 273086
rect 387432 273022 387484 273028
rect 388444 273080 388496 273086
rect 388444 273022 388496 273028
rect 388258 269920 388314 269929
rect 388258 269855 388314 269864
rect 387800 266484 387852 266490
rect 387800 266426 387852 266432
rect 387616 264376 387668 264382
rect 386998 264302 387288 264330
rect 387366 264324 387616 264330
rect 387366 264318 387668 264324
rect 387366 264302 387656 264318
rect 387812 264316 387840 266426
rect 388272 264316 388300 269855
rect 388456 267073 388484 273022
rect 388640 273018 388668 277780
rect 389192 277766 389758 277794
rect 389088 277568 389140 277574
rect 389088 277510 389140 277516
rect 388628 273012 388680 273018
rect 388628 272954 388680 272960
rect 388442 267064 388498 267073
rect 388442 266999 388498 267008
rect 389100 264330 389128 277510
rect 389192 268734 389220 277766
rect 389272 275324 389324 275330
rect 389272 275266 389324 275272
rect 389284 269822 389312 275266
rect 390940 272950 390968 277780
rect 391952 277766 392150 277794
rect 391756 276820 391808 276826
rect 391756 276762 391808 276768
rect 390928 272944 390980 272950
rect 390928 272886 390980 272892
rect 389272 269816 389324 269822
rect 389272 269758 389324 269764
rect 390008 269816 390060 269822
rect 390008 269758 390060 269764
rect 389180 268728 389232 268734
rect 389180 268670 389232 268676
rect 389180 268184 389232 268190
rect 389180 268126 389232 268132
rect 388746 264302 389128 264330
rect 389192 264316 389220 268126
rect 389638 265976 389694 265985
rect 389638 265911 389694 265920
rect 389652 264316 389680 265911
rect 390020 264316 390048 269758
rect 390468 268252 390520 268258
rect 390468 268194 390520 268200
rect 390480 264316 390508 268194
rect 391768 266422 391796 276762
rect 391952 267782 391980 277766
rect 392584 271176 392636 271182
rect 392584 271118 392636 271124
rect 391940 267776 391992 267782
rect 391940 267718 391992 267724
rect 392032 267776 392084 267782
rect 392032 267718 392084 267724
rect 392044 267594 392072 267718
rect 391860 267566 392072 267594
rect 390928 266416 390980 266422
rect 391756 266416 391808 266422
rect 390928 266358 390980 266364
rect 391386 266384 391442 266393
rect 390940 264316 390968 266358
rect 391756 266358 391808 266364
rect 391386 266319 391442 266328
rect 391400 264316 391428 266319
rect 391860 264316 391888 267566
rect 392596 266393 392624 271118
rect 393136 269000 393188 269006
rect 393136 268942 393188 268948
rect 392582 266384 392638 266393
rect 392582 266319 392638 266328
rect 392306 265840 392362 265849
rect 392306 265775 392362 265784
rect 392320 264316 392348 265775
rect 392794 264314 393084 264330
rect 393148 264316 393176 268942
rect 393332 268666 393360 277780
rect 394424 277500 394476 277506
rect 394424 277442 394476 277448
rect 393320 268660 393372 268666
rect 393320 268602 393372 268608
rect 393596 266484 393648 266490
rect 393596 266426 393648 266432
rect 393608 264316 393636 266426
rect 394436 264330 394464 277442
rect 394528 272882 394556 277780
rect 394712 277766 395738 277794
rect 396092 277766 396934 277794
rect 394608 276752 394660 276758
rect 394608 276694 394660 276700
rect 394516 272876 394568 272882
rect 394516 272818 394568 272824
rect 394620 272218 394648 276694
rect 394528 272190 394648 272218
rect 394528 266490 394556 272190
rect 394608 268864 394660 268870
rect 394608 268806 394660 268812
rect 394516 266484 394568 266490
rect 394516 266426 394568 266432
rect 394620 264330 394648 268806
rect 394712 268326 394740 277766
rect 395804 271992 395856 271998
rect 395804 271934 395856 271940
rect 395436 268796 395488 268802
rect 395436 268738 395488 268744
rect 394700 268320 394752 268326
rect 394700 268262 394752 268268
rect 394976 266484 395028 266490
rect 394976 266426 395028 266432
rect 392794 264308 393096 264314
rect 392794 264302 393044 264308
rect 394082 264302 394464 264330
rect 394542 264302 394648 264330
rect 394988 264316 395016 266426
rect 395448 264316 395476 268738
rect 395816 266490 395844 271934
rect 395896 268728 395948 268734
rect 395896 268670 395948 268676
rect 395804 266484 395856 266490
rect 395804 266426 395856 266432
rect 395908 264330 395936 268670
rect 396092 268598 396120 277766
rect 397276 273012 397328 273018
rect 397276 272954 397328 272960
rect 397184 268660 397236 268666
rect 397184 268602 397236 268608
rect 396080 268592 396132 268598
rect 396080 268534 396132 268540
rect 396264 266484 396316 266490
rect 396264 266426 396316 266432
rect 395830 264302 395936 264330
rect 396276 264316 396304 266426
rect 397196 264316 397224 268602
rect 397288 266490 397316 272954
rect 398024 272746 398052 277780
rect 398380 277432 398432 277438
rect 398380 277374 398432 277380
rect 398012 272740 398064 272746
rect 398012 272682 398064 272688
rect 397642 267744 397698 267753
rect 397642 267679 397698 267688
rect 397276 266484 397328 266490
rect 397276 266426 397328 266432
rect 397656 264316 397684 267679
rect 398392 264330 398420 277374
rect 398840 275392 398892 275398
rect 398840 275334 398892 275340
rect 398852 269074 398880 275334
rect 398932 272944 398984 272950
rect 398932 272886 398984 272892
rect 398840 269068 398892 269074
rect 398840 269010 398892 269016
rect 398470 268696 398526 268705
rect 398470 268631 398526 268640
rect 398130 264302 398420 264330
rect 398484 264316 398512 268631
rect 398944 264316 398972 272886
rect 399220 271930 399248 277780
rect 400232 277766 400430 277794
rect 399208 271924 399260 271930
rect 399208 271866 399260 271872
rect 399852 268592 399904 268598
rect 399852 268534 399904 268540
rect 399864 264316 399892 268534
rect 400232 268530 400260 277766
rect 400312 272876 400364 272882
rect 400312 272818 400364 272824
rect 400220 268524 400272 268530
rect 400220 268466 400272 268472
rect 400324 264316 400352 272818
rect 401612 272678 401640 277780
rect 402808 273494 402836 277780
rect 402992 277766 404018 277794
rect 402796 273488 402848 273494
rect 402796 273430 402848 273436
rect 402888 273488 402940 273494
rect 402888 273430 402940 273436
rect 401968 272740 402020 272746
rect 401968 272682 402020 272688
rect 401600 272672 401652 272678
rect 401600 272614 401652 272620
rect 401598 269784 401654 269793
rect 401598 269719 401654 269728
rect 401140 268524 401192 268530
rect 401140 268466 401192 268472
rect 400772 267028 400824 267034
rect 400772 266970 400824 266976
rect 400784 264316 400812 266970
rect 401152 264316 401180 268466
rect 401612 267050 401640 269719
rect 401520 267034 401640 267050
rect 401508 267028 401640 267034
rect 401560 267022 401640 267028
rect 401508 266970 401560 266976
rect 401980 264330 402008 272682
rect 402518 268560 402574 268569
rect 402518 268495 402574 268504
rect 402060 267096 402112 267102
rect 402060 267038 402112 267044
rect 401626 264302 402008 264330
rect 402072 264316 402100 267038
rect 402532 264316 402560 268495
rect 402900 267102 402928 273430
rect 402992 268462 403020 277766
rect 403440 274916 403492 274922
rect 403440 274858 403492 274864
rect 403256 272672 403308 272678
rect 403256 272614 403308 272620
rect 402980 268456 403032 268462
rect 402980 268398 403032 268404
rect 402888 267096 402940 267102
rect 402888 267038 402940 267044
rect 403268 264330 403296 272614
rect 403452 272066 403480 274858
rect 404266 272776 404322 272785
rect 404266 272711 404322 272720
rect 403440 272060 403492 272066
rect 403440 272002 403492 272008
rect 403900 268456 403952 268462
rect 403900 268398 403952 268404
rect 403438 267608 403494 267617
rect 403438 267543 403494 267552
rect 403006 264302 403296 264330
rect 403452 264316 403480 267543
rect 403912 264316 403940 268398
rect 404280 264316 404308 272711
rect 405200 272610 405228 277780
rect 405936 277766 406318 277794
rect 407132 277766 407514 277794
rect 405648 276072 405700 276078
rect 405648 276014 405700 276020
rect 405188 272604 405240 272610
rect 405188 272546 405240 272552
rect 405556 272604 405608 272610
rect 405556 272546 405608 272552
rect 405186 268424 405242 268433
rect 405186 268359 405242 268368
rect 404728 267096 404780 267102
rect 404728 267038 404780 267044
rect 404740 264316 404768 267038
rect 405200 264316 405228 268359
rect 405568 264330 405596 272546
rect 405660 267102 405688 276014
rect 405648 267096 405700 267102
rect 405648 267038 405700 267044
rect 405936 267034 405964 277766
rect 406934 272640 406990 272649
rect 406934 272575 406990 272584
rect 405924 267028 405976 267034
rect 405924 266970 405976 266976
rect 406108 267028 406160 267034
rect 406108 266970 406160 266976
rect 405568 264302 405674 264330
rect 406120 264316 406148 266970
rect 406566 265704 406622 265713
rect 406566 265639 406622 265648
rect 406580 264316 406608 265639
rect 406948 264316 406976 272575
rect 407132 267918 407160 277766
rect 408408 276684 408460 276690
rect 408408 276626 408460 276632
rect 408420 273254 408448 276626
rect 408236 273226 408448 273254
rect 407120 267912 407172 267918
rect 407120 267854 407172 267860
rect 407394 266384 407450 266393
rect 407394 266319 407450 266328
rect 407408 264316 407436 266319
rect 408236 264330 408264 273226
rect 408696 272542 408724 277780
rect 409892 275330 409920 277780
rect 409984 277766 411102 277794
rect 411824 277766 412298 277794
rect 409880 275324 409932 275330
rect 409880 275266 409932 275272
rect 409144 274848 409196 274854
rect 409144 274790 409196 274796
rect 408684 272536 408736 272542
rect 408314 272504 408370 272513
rect 408684 272478 408736 272484
rect 408314 272439 408370 272448
rect 407882 264302 408264 264330
rect 408328 264316 408356 272439
rect 408684 269068 408736 269074
rect 408684 269010 408736 269016
rect 408696 266490 408724 269010
rect 409156 266558 409184 274790
rect 409788 272536 409840 272542
rect 409788 272478 409840 272484
rect 409144 266552 409196 266558
rect 409144 266494 409196 266500
rect 408684 266484 408736 266490
rect 408684 266426 408736 266432
rect 408776 266484 408828 266490
rect 408776 266426 408828 266432
rect 408788 264316 408816 266426
rect 409234 265568 409290 265577
rect 409234 265503 409290 265512
rect 409248 264316 409276 265503
rect 409800 264330 409828 272478
rect 409984 268394 410012 277766
rect 411168 275324 411220 275330
rect 411168 275266 411220 275272
rect 411074 274000 411130 274009
rect 411074 273935 411130 273944
rect 409972 268388 410024 268394
rect 409972 268330 410024 268336
rect 410432 268388 410484 268394
rect 410432 268330 410484 268336
rect 410064 266416 410116 266422
rect 410444 266393 410472 268330
rect 410524 267096 410576 267102
rect 410524 267038 410576 267044
rect 410064 266358 410116 266364
rect 410430 266384 410486 266393
rect 409630 264302 409828 264330
rect 410076 264316 410104 266358
rect 410430 266319 410486 266328
rect 410536 264316 410564 267038
rect 411088 266422 411116 273935
rect 411076 266416 411128 266422
rect 411076 266358 411128 266364
rect 411180 264330 411208 275266
rect 411824 272814 411852 277766
rect 413388 275398 413416 277780
rect 414032 277766 414598 277794
rect 413376 275392 413428 275398
rect 413376 275334 413428 275340
rect 411812 272808 411864 272814
rect 411812 272750 411864 272756
rect 411904 272808 411956 272814
rect 411904 272750 411956 272756
rect 411916 267753 411944 272750
rect 414032 268138 414060 277766
rect 415780 272134 415808 277780
rect 416792 277766 416990 277794
rect 415768 272128 415820 272134
rect 415768 272070 415820 272076
rect 413940 268110 414060 268138
rect 413940 268054 413968 268110
rect 413928 268048 413980 268054
rect 413928 267990 413980 267996
rect 414020 268048 414072 268054
rect 414020 267990 414072 267996
rect 411902 267744 411958 267753
rect 411902 267679 411958 267688
rect 411442 267200 411498 267209
rect 411442 267135 411498 267144
rect 411010 264302 411208 264330
rect 411456 264316 411484 267135
rect 411902 267064 411958 267073
rect 411902 266999 411958 267008
rect 411916 264316 411944 266999
rect 414032 266626 414060 267990
rect 416792 267850 416820 277766
rect 416780 267844 416832 267850
rect 416780 267786 416832 267792
rect 414756 267096 414808 267102
rect 414808 267044 414980 267050
rect 414756 267038 414980 267044
rect 414768 267034 414980 267038
rect 414768 267028 414992 267034
rect 414768 267022 414940 267028
rect 414940 266970 414992 266976
rect 414020 266620 414072 266626
rect 414020 266562 414072 266568
rect 418172 265198 418200 277780
rect 419368 272202 419396 277780
rect 419540 275392 419592 275398
rect 419540 275334 419592 275340
rect 419552 274009 419580 275334
rect 420564 274854 420592 277780
rect 421668 276350 421696 277780
rect 421656 276344 421708 276350
rect 421656 276286 421708 276292
rect 420552 274848 420604 274854
rect 420552 274790 420604 274796
rect 419538 274000 419594 274009
rect 419538 273935 419594 273944
rect 419356 272196 419408 272202
rect 419356 272138 419408 272144
rect 420184 272196 420236 272202
rect 420184 272138 420236 272144
rect 420196 266694 420224 272138
rect 422864 270706 422892 277780
rect 424060 274922 424088 277780
rect 425072 277766 425270 277794
rect 424048 274916 424100 274922
rect 424048 274858 424100 274864
rect 422852 270700 422904 270706
rect 422852 270642 422904 270648
rect 420184 266688 420236 266694
rect 420184 266630 420236 266636
rect 425072 265266 425100 277766
rect 426452 272270 426480 277780
rect 426636 277766 427662 277794
rect 426440 272264 426492 272270
rect 426440 272206 426492 272212
rect 426636 268054 426664 277766
rect 428844 276418 428872 277780
rect 428832 276412 428884 276418
rect 428832 276354 428884 276360
rect 429948 270774 429976 277780
rect 431144 274990 431172 277780
rect 432340 276486 432368 277780
rect 433352 277766 433550 277794
rect 432328 276480 432380 276486
rect 432328 276422 432380 276428
rect 431132 274984 431184 274990
rect 431132 274926 431184 274932
rect 429936 270768 429988 270774
rect 429936 270710 429988 270716
rect 433352 268977 433380 277766
rect 434732 272202 434760 277780
rect 434916 277766 435942 277794
rect 434720 272196 434772 272202
rect 434720 272138 434772 272144
rect 433338 268968 433394 268977
rect 433338 268903 433394 268912
rect 426624 268048 426676 268054
rect 426624 267990 426676 267996
rect 434916 265334 434944 277766
rect 435364 272332 435416 272338
rect 435364 272274 435416 272280
rect 435376 266762 435404 272274
rect 437032 272270 437060 277780
rect 438228 275466 438256 277780
rect 439424 276554 439452 277780
rect 440252 277766 440634 277794
rect 439412 276548 439464 276554
rect 439412 276490 439464 276496
rect 438216 275460 438268 275466
rect 438216 275402 438268 275408
rect 438860 275460 438912 275466
rect 438860 275402 438912 275408
rect 438872 273494 438900 275402
rect 438860 273488 438912 273494
rect 438860 273430 438912 273436
rect 437020 272264 437072 272270
rect 437020 272206 437072 272212
rect 435364 266756 435416 266762
rect 435364 266698 435416 266704
rect 440252 265402 440280 277766
rect 441816 272338 441844 277780
rect 441804 272332 441856 272338
rect 441804 272274 441856 272280
rect 443012 265470 443040 277780
rect 444208 276622 444236 277780
rect 444196 276616 444248 276622
rect 444196 276558 444248 276564
rect 445312 275058 445340 277780
rect 445772 277766 446522 277794
rect 447152 277766 447718 277794
rect 448532 277766 448914 277794
rect 449912 277766 450110 277794
rect 445300 275052 445352 275058
rect 445300 274994 445352 275000
rect 445772 269346 445800 277766
rect 445760 269340 445812 269346
rect 445760 269282 445812 269288
rect 447152 265538 447180 277766
rect 448532 266830 448560 277766
rect 449912 269414 449940 277766
rect 451292 270842 451320 277780
rect 452488 275194 452516 277780
rect 452672 277766 453606 277794
rect 452476 275188 452528 275194
rect 452476 275130 452528 275136
rect 451280 270836 451332 270842
rect 451280 270778 451332 270784
rect 452672 269482 452700 277766
rect 454788 277642 454816 277780
rect 455432 277766 455998 277794
rect 456812 277766 457194 277794
rect 454776 277636 454828 277642
rect 454776 277578 454828 277584
rect 452660 269476 452712 269482
rect 452660 269418 452712 269424
rect 449900 269408 449952 269414
rect 449900 269350 449952 269356
rect 455432 266898 455460 277766
rect 456812 269550 456840 277766
rect 458376 273562 458404 277780
rect 459572 275262 459600 277780
rect 459664 277766 460690 277794
rect 459560 275256 459612 275262
rect 459560 275198 459612 275204
rect 458364 273556 458416 273562
rect 458364 273498 458416 273504
rect 459664 269618 459692 277766
rect 459744 275256 459796 275262
rect 459744 275198 459796 275204
rect 459652 269612 459704 269618
rect 459652 269554 459704 269560
rect 456800 269544 456852 269550
rect 456800 269486 456852 269492
rect 459756 267986 459784 275198
rect 461872 273630 461900 277780
rect 462332 277766 463082 277794
rect 463712 277766 464278 277794
rect 461860 273624 461912 273630
rect 461860 273566 461912 273572
rect 459744 267980 459796 267986
rect 459744 267922 459796 267928
rect 462332 267714 462360 277766
rect 463712 269686 463740 277766
rect 465460 273698 465488 277780
rect 466656 275874 466684 277780
rect 466644 275868 466696 275874
rect 466644 275810 466696 275816
rect 466736 275868 466788 275874
rect 466736 275810 466788 275816
rect 465448 273692 465500 273698
rect 465448 273634 465500 273640
rect 466748 271998 466776 275810
rect 466736 271992 466788 271998
rect 466736 271934 466788 271940
rect 467852 270162 467880 277780
rect 468956 273766 468984 277780
rect 469232 277766 470166 277794
rect 470612 277766 471362 277794
rect 468944 273760 468996 273766
rect 468944 273702 468996 273708
rect 467840 270156 467892 270162
rect 467840 270098 467892 270104
rect 463700 269680 463752 269686
rect 463700 269622 463752 269628
rect 469232 269618 469260 277766
rect 469312 270156 469364 270162
rect 469312 270098 469364 270104
rect 464712 269612 464764 269618
rect 464712 269554 464764 269560
rect 469220 269612 469272 269618
rect 469220 269554 469272 269560
rect 462320 267708 462372 267714
rect 462320 267650 462372 267656
rect 464724 266966 464752 269554
rect 469324 267617 469352 270098
rect 470612 269754 470640 277766
rect 472544 273834 472572 277780
rect 473740 276010 473768 277780
rect 474752 277766 474950 277794
rect 473728 276004 473780 276010
rect 473728 275946 473780 275952
rect 472532 273828 472584 273834
rect 472532 273770 472584 273776
rect 474752 270502 474780 277766
rect 476132 273902 476160 277780
rect 476316 277766 477250 277794
rect 477512 277766 478446 277794
rect 479352 277766 479642 277794
rect 476120 273896 476172 273902
rect 476120 273838 476172 273844
rect 474740 270496 474792 270502
rect 474740 270438 474792 270444
rect 470600 269748 470652 269754
rect 470600 269690 470652 269696
rect 476316 267646 476344 277766
rect 477512 270434 477540 277766
rect 479352 274174 479380 277766
rect 480824 275942 480852 277780
rect 481652 277766 482034 277794
rect 480812 275936 480864 275942
rect 480812 275878 480864 275884
rect 481180 275936 481232 275942
rect 481180 275878 481232 275884
rect 479340 274168 479392 274174
rect 479340 274110 479392 274116
rect 479524 274168 479576 274174
rect 479524 274110 479576 274116
rect 477500 270428 477552 270434
rect 477500 270370 477552 270376
rect 476304 267640 476356 267646
rect 469310 267608 469366 267617
rect 476304 267582 476356 267588
rect 469310 267543 469366 267552
rect 464712 266960 464764 266966
rect 464712 266902 464764 266908
rect 455420 266892 455472 266898
rect 455420 266834 455472 266840
rect 448520 266824 448572 266830
rect 448520 266766 448572 266772
rect 479536 266490 479564 274110
rect 481192 268122 481220 275878
rect 481652 270366 481680 277766
rect 483216 274650 483244 277780
rect 483400 277766 484334 277794
rect 484412 277766 485530 277794
rect 483204 274644 483256 274650
rect 483204 274586 483256 274592
rect 481640 270360 481692 270366
rect 481640 270302 481692 270308
rect 481180 268116 481232 268122
rect 481180 268058 481232 268064
rect 483400 267578 483428 277766
rect 484412 270201 484440 277766
rect 486712 274582 486740 277780
rect 487908 275126 487936 277780
rect 489104 277370 489132 277780
rect 489092 277364 489144 277370
rect 489092 277306 489144 277312
rect 487896 275120 487948 275126
rect 487896 275062 487948 275068
rect 486700 274576 486752 274582
rect 486700 274518 486752 274524
rect 490300 274514 490328 277780
rect 491496 277394 491524 277780
rect 491404 277366 491524 277394
rect 492232 277766 492614 277794
rect 490288 274508 490340 274514
rect 490288 274450 490340 274456
rect 491300 272332 491352 272338
rect 491300 272274 491352 272280
rect 484398 270192 484454 270201
rect 484398 270127 484454 270136
rect 483388 267572 483440 267578
rect 483388 267514 483440 267520
rect 479524 266484 479576 266490
rect 479524 266426 479576 266432
rect 491312 265606 491340 272274
rect 491404 267510 491432 277366
rect 492232 272338 492260 277766
rect 493324 274508 493376 274514
rect 493324 274450 493376 274456
rect 492220 272332 492272 272338
rect 492220 272274 492272 272280
rect 491392 267504 491444 267510
rect 493336 267481 493364 274450
rect 493796 274446 493824 277780
rect 494992 275806 495020 277780
rect 496188 277302 496216 277780
rect 496176 277296 496228 277302
rect 496176 277238 496228 277244
rect 494980 275800 495032 275806
rect 494980 275742 495032 275748
rect 495072 275800 495124 275806
rect 495072 275742 495124 275748
rect 493784 274440 493836 274446
rect 493784 274382 493836 274388
rect 495084 268190 495112 275742
rect 497384 274378 497412 277780
rect 498212 277766 498594 277794
rect 499592 277766 499790 277794
rect 497372 274372 497424 274378
rect 497372 274314 497424 274320
rect 495072 268184 495124 268190
rect 495072 268126 495124 268132
rect 491392 267446 491444 267452
rect 493322 267472 493378 267481
rect 498212 267442 498240 277766
rect 493322 267407 493378 267416
rect 498200 267436 498252 267442
rect 498200 267378 498252 267384
rect 499592 266354 499620 277766
rect 500880 274310 500908 277780
rect 502076 275738 502104 277780
rect 503272 277234 503300 277780
rect 503732 277766 504482 277794
rect 503260 277228 503312 277234
rect 503260 277170 503312 277176
rect 502064 275732 502116 275738
rect 502064 275674 502116 275680
rect 500868 274304 500920 274310
rect 500868 274246 500920 274252
rect 503732 270298 503760 277766
rect 505664 274514 505692 277780
rect 506492 277766 506874 277794
rect 505652 274508 505704 274514
rect 505652 274450 505704 274456
rect 503720 270292 503772 270298
rect 503720 270234 503772 270240
rect 499580 266348 499632 266354
rect 499580 266290 499632 266296
rect 506492 266286 506520 277766
rect 507860 275732 507912 275738
rect 507860 275674 507912 275680
rect 507872 268258 507900 275674
rect 507964 272406 507992 277780
rect 509160 275670 509188 277780
rect 510356 277166 510384 277780
rect 510632 277766 511566 277794
rect 512012 277766 512762 277794
rect 513392 277766 513958 277794
rect 510344 277160 510396 277166
rect 510344 277102 510396 277108
rect 509148 275664 509200 275670
rect 509148 275606 509200 275612
rect 507952 272400 508004 272406
rect 507952 272342 508004 272348
rect 510632 270230 510660 277766
rect 510620 270224 510672 270230
rect 510620 270166 510672 270172
rect 507860 268252 507912 268258
rect 507860 268194 507912 268200
rect 512012 267374 512040 277766
rect 512000 267368 512052 267374
rect 512000 267310 512052 267316
rect 506480 266280 506532 266286
rect 506480 266222 506532 266228
rect 513392 266218 513420 277766
rect 515140 272474 515168 277780
rect 516244 275602 516272 277780
rect 516232 275596 516284 275602
rect 516232 275538 516284 275544
rect 515128 272468 515180 272474
rect 515128 272410 515180 272416
rect 517440 270910 517468 277780
rect 518636 274242 518664 277780
rect 518912 277766 519846 277794
rect 518624 274236 518676 274242
rect 518624 274178 518676 274184
rect 517428 270904 517480 270910
rect 517428 270846 517480 270852
rect 518912 269142 518940 277766
rect 521028 270978 521056 277780
rect 522224 273222 522252 277780
rect 523420 275534 523448 277780
rect 523408 275528 523460 275534
rect 523408 275470 523460 275476
rect 523592 275528 523644 275534
rect 523592 275470 523644 275476
rect 522212 273216 522264 273222
rect 522212 273158 522264 273164
rect 521016 270972 521068 270978
rect 521016 270914 521068 270920
rect 518992 269340 519044 269346
rect 518992 269282 519044 269288
rect 516140 269136 516192 269142
rect 516140 269078 516192 269084
rect 518900 269136 518952 269142
rect 518900 269078 518952 269084
rect 516152 267306 516180 269078
rect 519004 267345 519032 269282
rect 523604 267782 523632 275470
rect 523684 274236 523736 274242
rect 523684 274178 523736 274184
rect 523592 267776 523644 267782
rect 523592 267718 523644 267724
rect 518990 267336 519046 267345
rect 516140 267300 516192 267306
rect 518990 267271 519046 267280
rect 516140 267242 516192 267248
rect 523696 267238 523724 274178
rect 524524 271046 524552 277780
rect 524616 277766 525734 277794
rect 525812 277766 526930 277794
rect 524512 271040 524564 271046
rect 524512 270982 524564 270988
rect 524616 270094 524644 277766
rect 524604 270088 524656 270094
rect 524604 270030 524656 270036
rect 525812 269346 525840 277766
rect 528112 271114 528140 277780
rect 528572 277766 529322 277794
rect 528100 271108 528152 271114
rect 528100 271050 528152 271056
rect 525800 269340 525852 269346
rect 525800 269282 525852 269288
rect 523684 267232 523736 267238
rect 523684 267174 523736 267180
rect 513380 266212 513432 266218
rect 513380 266154 513432 266160
rect 491300 265600 491352 265606
rect 491300 265542 491352 265548
rect 447140 265532 447192 265538
rect 447140 265474 447192 265480
rect 443000 265464 443052 265470
rect 443000 265406 443052 265412
rect 440240 265396 440292 265402
rect 440240 265338 440292 265344
rect 434904 265328 434956 265334
rect 434904 265270 434956 265276
rect 425060 265260 425112 265266
rect 425060 265202 425112 265208
rect 418160 265192 418212 265198
rect 418160 265134 418212 265140
rect 528572 264518 528600 277766
rect 530504 275505 530532 277780
rect 530490 275496 530546 275505
rect 530490 275431 530546 275440
rect 531608 271862 531636 277780
rect 532804 277394 532832 277780
rect 532712 277366 532832 277394
rect 531596 271856 531648 271862
rect 531596 271798 531648 271804
rect 532712 268841 532740 277366
rect 534000 274242 534028 277780
rect 533988 274236 534040 274242
rect 533988 274178 534040 274184
rect 535196 271794 535224 277780
rect 536392 273154 536420 277780
rect 537588 275369 537616 277780
rect 537574 275360 537630 275369
rect 537574 275295 537630 275304
rect 536380 273148 536432 273154
rect 536380 273090 536432 273096
rect 535184 271788 535236 271794
rect 535184 271730 535236 271736
rect 538784 271726 538812 277780
rect 539888 274106 539916 277780
rect 541084 277394 541112 277780
rect 540992 277366 541112 277394
rect 539876 274100 539928 274106
rect 539876 274042 539928 274048
rect 538772 271720 538824 271726
rect 538772 271662 538824 271668
rect 532698 268832 532754 268841
rect 532698 268767 532754 268776
rect 540992 267170 541020 277366
rect 542280 271658 542308 277780
rect 542372 277766 543490 277794
rect 542268 271652 542320 271658
rect 542268 271594 542320 271600
rect 542372 270026 542400 277766
rect 544672 275233 544700 277780
rect 545132 277766 545882 277794
rect 544658 275224 544714 275233
rect 544658 275159 544714 275168
rect 542360 270020 542412 270026
rect 542360 269962 542412 269968
rect 540980 267164 541032 267170
rect 540980 267106 541032 267112
rect 545132 266150 545160 277766
rect 547064 271590 547092 277780
rect 547892 277766 548182 277794
rect 547052 271584 547104 271590
rect 547052 271526 547104 271532
rect 547892 269958 547920 277766
rect 549364 277394 549392 277780
rect 549272 277366 549392 277394
rect 547880 269952 547932 269958
rect 547880 269894 547932 269900
rect 545120 266144 545172 266150
rect 545120 266086 545172 266092
rect 549272 266082 549300 277366
rect 550560 271522 550588 277780
rect 551756 274038 551784 277780
rect 552032 277766 552966 277794
rect 551744 274032 551796 274038
rect 551744 273974 551796 273980
rect 550548 271516 550600 271522
rect 550548 271458 550600 271464
rect 549260 266076 549312 266082
rect 549260 266018 549312 266024
rect 552032 266014 552060 277766
rect 554148 271454 554176 277780
rect 554136 271448 554188 271454
rect 554136 271390 554188 271396
rect 555252 271386 555280 277780
rect 556172 277766 556462 277794
rect 555240 271380 555292 271386
rect 555240 271322 555292 271328
rect 552020 266008 552072 266014
rect 552020 265950 552072 265956
rect 556172 265946 556200 277766
rect 557644 271318 557672 277780
rect 557736 277766 558854 277794
rect 558932 277766 560050 277794
rect 557632 271312 557684 271318
rect 557632 271254 557684 271260
rect 557736 269890 557764 277766
rect 557724 269884 557776 269890
rect 557724 269826 557776 269832
rect 556160 265940 556212 265946
rect 556160 265882 556212 265888
rect 558932 265878 558960 277766
rect 561232 271425 561260 277780
rect 562428 273970 562456 277780
rect 563072 277766 563546 277794
rect 562416 273964 562468 273970
rect 562416 273906 562468 273912
rect 561218 271416 561274 271425
rect 561218 271351 561274 271360
rect 558920 265872 558972 265878
rect 558920 265814 558972 265820
rect 563072 265810 563100 277766
rect 564728 271250 564756 277780
rect 565924 273086 565952 277780
rect 567120 277030 567148 277780
rect 567108 277024 567160 277030
rect 567108 276966 567160 276972
rect 565912 273080 565964 273086
rect 565912 273022 565964 273028
rect 568316 271289 568344 277780
rect 568592 277766 569526 277794
rect 569972 277766 570722 277794
rect 568302 271280 568358 271289
rect 564716 271244 564768 271250
rect 568302 271215 568358 271224
rect 564716 271186 564768 271192
rect 568592 268938 568620 277766
rect 568580 268932 568632 268938
rect 568580 268874 568632 268880
rect 563060 265804 563112 265810
rect 563060 265746 563112 265752
rect 569972 265742 570000 277766
rect 571812 271153 571840 277780
rect 572732 277766 573022 277794
rect 571798 271144 571854 271153
rect 571798 271079 571854 271088
rect 572732 270065 572760 277766
rect 574204 277098 574232 277780
rect 574192 277092 574244 277098
rect 574192 277034 574244 277040
rect 575400 276962 575428 277780
rect 575492 277766 576610 277794
rect 575388 276956 575440 276962
rect 575388 276898 575440 276904
rect 572718 270056 572774 270065
rect 572718 269991 572774 270000
rect 569960 265736 570012 265742
rect 569960 265678 570012 265684
rect 528560 264512 528612 264518
rect 528560 264454 528612 264460
rect 575492 264450 575520 277766
rect 577688 275732 577740 275738
rect 577688 275674 577740 275680
rect 577700 269006 577728 275674
rect 577792 275262 577820 277780
rect 578252 277766 578910 277794
rect 577780 275256 577832 275262
rect 577780 275198 577832 275204
rect 577688 269000 577740 269006
rect 577688 268942 577740 268948
rect 578252 265674 578280 277766
rect 580092 273873 580120 277780
rect 581288 275942 581316 277780
rect 582484 276894 582512 277780
rect 582576 277766 583694 277794
rect 583772 277766 584890 277794
rect 585152 277766 586086 277794
rect 582472 276888 582524 276894
rect 582472 276830 582524 276836
rect 581276 275936 581328 275942
rect 581276 275878 581328 275884
rect 581644 275596 581696 275602
rect 581644 275538 581696 275544
rect 580078 273864 580134 273873
rect 580078 273799 580134 273808
rect 581656 273018 581684 275538
rect 581644 273012 581696 273018
rect 581644 272954 581696 272960
rect 578240 265668 578292 265674
rect 578240 265610 578292 265616
rect 575480 264444 575532 264450
rect 575480 264386 575532 264392
rect 582576 264382 582604 277766
rect 583772 269074 583800 277766
rect 585152 269929 585180 277766
rect 587176 277574 587204 277780
rect 587164 277568 587216 277574
rect 587164 277510 587216 277516
rect 588372 275806 588400 277780
rect 589292 277766 589582 277794
rect 588360 275800 588412 275806
rect 588360 275742 588412 275748
rect 585138 269920 585194 269929
rect 585138 269855 585194 269864
rect 583760 269068 583812 269074
rect 583760 269010 583812 269016
rect 589292 265985 589320 277766
rect 590764 277394 590792 277780
rect 590672 277366 590792 277394
rect 590672 269822 590700 277366
rect 591960 275670 591988 277780
rect 593156 276826 593184 277780
rect 593144 276820 593196 276826
rect 593144 276762 593196 276768
rect 591948 275664 592000 275670
rect 591948 275606 592000 275612
rect 592040 275664 592092 275670
rect 592040 275606 592092 275612
rect 592052 275482 592080 275606
rect 591960 275454 592080 275482
rect 591960 272950 591988 275454
rect 591948 272944 592000 272950
rect 591948 272886 592000 272892
rect 594352 271182 594380 277780
rect 594812 277766 595470 277794
rect 596192 277766 596666 277794
rect 597572 277766 597862 277794
rect 594812 275618 594840 277766
rect 594720 275590 594840 275618
rect 594720 275534 594748 275590
rect 594708 275528 594760 275534
rect 594708 275470 594760 275476
rect 594800 275528 594852 275534
rect 594800 275470 594852 275476
rect 594812 272882 594840 275470
rect 594800 272876 594852 272882
rect 594800 272818 594852 272824
rect 594340 271176 594392 271182
rect 594340 271118 594392 271124
rect 590660 269816 590712 269822
rect 590660 269758 590712 269764
rect 589278 265976 589334 265985
rect 589278 265911 589334 265920
rect 596192 265849 596220 277766
rect 596178 265840 596234 265849
rect 596178 265775 596234 265784
rect 582564 264376 582616 264382
rect 582564 264318 582616 264324
rect 597572 264314 597600 277766
rect 599044 275738 599072 277780
rect 600240 276758 600268 277780
rect 601436 277506 601464 277780
rect 601712 277766 602554 277794
rect 601424 277500 601476 277506
rect 601424 277442 601476 277448
rect 600228 276752 600280 276758
rect 600228 276694 600280 276700
rect 599032 275732 599084 275738
rect 599032 275674 599084 275680
rect 601712 268870 601740 277766
rect 603736 275874 603764 277780
rect 604472 277766 604946 277794
rect 605852 277766 606142 277794
rect 603724 275868 603776 275874
rect 603724 275810 603776 275816
rect 601700 268864 601752 268870
rect 601700 268806 601752 268812
rect 604472 268802 604500 277766
rect 604460 268796 604512 268802
rect 604460 268738 604512 268744
rect 605852 268734 605880 277766
rect 607324 275602 607352 277780
rect 607416 277766 608534 277794
rect 608612 277766 609730 277794
rect 607312 275596 607364 275602
rect 607312 275538 607364 275544
rect 605840 268728 605892 268734
rect 605840 268670 605892 268676
rect 597560 264308 597612 264314
rect 393044 264250 393096 264256
rect 597560 264250 597612 264256
rect 396998 264208 397054 264217
rect 396750 264166 396998 264194
rect 401230 264208 401286 264217
rect 399418 264178 399800 264194
rect 399418 264172 399812 264178
rect 399418 264166 399760 264172
rect 396998 264143 397054 264152
rect 607416 264178 607444 277766
rect 608612 268666 608640 277766
rect 610820 272814 610848 277780
rect 612016 277438 612044 277780
rect 612752 277766 613226 277794
rect 612004 277432 612056 277438
rect 612004 277374 612056 277380
rect 610808 272808 610860 272814
rect 610808 272750 610860 272756
rect 612752 268705 612780 277766
rect 614408 275670 614436 277780
rect 615604 277394 615632 277780
rect 615512 277366 615632 277394
rect 615696 277766 616814 277794
rect 614396 275664 614448 275670
rect 614396 275606 614448 275612
rect 612738 268696 612794 268705
rect 608600 268660 608652 268666
rect 612738 268631 612794 268640
rect 608600 268602 608652 268608
rect 401230 264143 401232 264152
rect 399760 264114 399812 264120
rect 401284 264143 401286 264152
rect 607404 264172 607456 264178
rect 401232 264114 401284 264120
rect 607404 264114 607456 264120
rect 615512 264110 615540 277366
rect 615696 268598 615724 277766
rect 617996 275534 618024 277780
rect 618272 277766 619114 277794
rect 619652 277766 620310 277794
rect 617984 275528 618036 275534
rect 617984 275470 618036 275476
rect 618272 269793 618300 277766
rect 618258 269784 618314 269793
rect 618258 269719 618314 269728
rect 615684 268592 615736 268598
rect 615684 268534 615736 268540
rect 619652 268530 619680 277766
rect 621492 272746 621520 277780
rect 622688 275466 622716 277780
rect 623884 277394 623912 277780
rect 623792 277366 623912 277394
rect 622676 275460 622728 275466
rect 622676 275402 622728 275408
rect 621480 272740 621532 272746
rect 621480 272682 621532 272688
rect 623792 268569 623820 277366
rect 625080 272678 625108 277780
rect 625172 277766 626198 277794
rect 626552 277766 627394 277794
rect 625068 272672 625120 272678
rect 625068 272614 625120 272620
rect 625172 270162 625200 277766
rect 625160 270156 625212 270162
rect 625160 270098 625212 270104
rect 623778 268560 623834 268569
rect 619640 268524 619692 268530
rect 623778 268495 623834 268504
rect 619640 268466 619692 268472
rect 626552 268462 626580 277766
rect 628576 272785 628604 277780
rect 629772 276010 629800 277780
rect 630692 277766 630982 277794
rect 629760 276004 629812 276010
rect 629760 275946 629812 275952
rect 628562 272776 628618 272785
rect 628562 272711 628618 272720
rect 626540 268456 626592 268462
rect 630692 268433 630720 277766
rect 632164 272610 632192 277780
rect 632256 277766 633374 277794
rect 633452 277766 634478 277794
rect 632152 272604 632204 272610
rect 632152 272546 632204 272552
rect 626540 268398 626592 268404
rect 630678 268424 630734 268433
rect 630678 268359 630734 268368
rect 632256 267102 632284 277766
rect 632244 267096 632296 267102
rect 632244 267038 632296 267044
rect 633452 265713 633480 277766
rect 635660 272649 635688 277780
rect 636212 277766 636870 277794
rect 635646 272640 635702 272649
rect 635646 272575 635702 272584
rect 636212 268394 636240 277766
rect 638052 276690 638080 277780
rect 638040 276684 638092 276690
rect 638040 276626 638092 276632
rect 639248 272513 639276 277780
rect 640444 274174 640472 277780
rect 640536 277766 641654 277794
rect 640432 274168 640484 274174
rect 640432 274110 640484 274116
rect 639234 272504 639290 272513
rect 639234 272439 639290 272448
rect 636200 268388 636252 268394
rect 636200 268330 636252 268336
rect 633438 265704 633494 265713
rect 633438 265639 633494 265648
rect 640536 265577 640564 277766
rect 642744 272542 642772 277780
rect 643940 275398 643968 277780
rect 644492 277766 645150 277794
rect 643928 275392 643980 275398
rect 643928 275334 643980 275340
rect 642732 272536 642784 272542
rect 642732 272478 642784 272484
rect 644492 267034 644520 277766
rect 646332 275330 646360 277780
rect 646320 275324 646372 275330
rect 646320 275266 646372 275272
rect 647252 267209 647280 278310
rect 647332 278180 647384 278186
rect 647332 278122 647384 278128
rect 647238 267200 647294 267209
rect 647238 267135 647294 267144
rect 644480 267028 644532 267034
rect 644480 266970 644532 266976
rect 640522 265568 640578 265577
rect 640522 265503 640578 265512
rect 615500 264104 615552 264110
rect 615500 264046 615552 264052
rect 415306 262304 415362 262313
rect 415306 262239 415308 262248
rect 415360 262239 415362 262248
rect 572720 262268 572772 262274
rect 415308 262210 415360 262216
rect 572720 262210 572772 262216
rect 414202 259176 414258 259185
rect 414202 259111 414258 259120
rect 189078 258632 189134 258641
rect 189078 258567 189134 258576
rect 189092 258126 189120 258567
rect 414216 258126 414244 259111
rect 179420 258120 179472 258126
rect 179420 258062 179472 258068
rect 189080 258120 189132 258126
rect 189080 258062 189132 258068
rect 414204 258120 414256 258126
rect 414204 258062 414256 258068
rect 571524 258120 571576 258126
rect 571524 258062 571576 258068
rect 179432 251394 179460 258062
rect 415306 255912 415362 255921
rect 415306 255847 415362 255856
rect 415320 255338 415348 255847
rect 415308 255332 415360 255338
rect 415308 255274 415360 255280
rect 571432 255332 571484 255338
rect 571432 255274 571484 255280
rect 414386 252784 414442 252793
rect 414386 252719 414442 252728
rect 414400 252618 414428 252719
rect 414388 252612 414440 252618
rect 414388 252554 414440 252560
rect 173900 251388 173952 251394
rect 173900 251330 173952 251336
rect 179420 251388 179472 251394
rect 179420 251330 179472 251336
rect 173912 249354 173940 251330
rect 414202 249520 414258 249529
rect 414202 249455 414258 249464
rect 171784 249348 171836 249354
rect 171784 249290 171836 249296
rect 173900 249348 173952 249354
rect 173900 249290 173952 249296
rect 85026 247344 85082 247353
rect 85026 247279 85082 247288
rect 84842 247208 84898 247217
rect 84842 247143 84898 247152
rect 67548 231668 67600 231674
rect 67548 231610 67600 231616
rect 66902 229936 66958 229945
rect 66902 229871 66958 229880
rect 58622 229800 58678 229809
rect 58622 229735 58678 229744
rect 57612 226364 57664 226370
rect 57612 226306 57664 226312
rect 56048 225684 56100 225690
rect 56048 225626 56100 225632
rect 55956 218952 56008 218958
rect 55956 218894 56008 218900
rect 55864 218816 55916 218822
rect 55864 218758 55916 218764
rect 56060 217410 56088 225626
rect 56874 221504 56930 221513
rect 56874 221439 56930 221448
rect 56888 217410 56916 221439
rect 57624 220862 57652 226306
rect 57612 220856 57664 220862
rect 57612 220798 57664 220804
rect 58636 220658 58664 229735
rect 62120 229084 62172 229090
rect 62120 229026 62172 229032
rect 59266 226944 59322 226953
rect 59266 226879 59322 226888
rect 58714 223000 58770 223009
rect 58714 222935 58770 222944
rect 57612 220652 57664 220658
rect 57612 220594 57664 220600
rect 58624 220652 58676 220658
rect 58624 220594 58676 220600
rect 57624 217410 57652 220594
rect 58728 219434 58756 222935
rect 58636 219406 58756 219434
rect 58636 217410 58664 219406
rect 59280 217410 59308 226879
rect 62132 226370 62160 229026
rect 62762 227080 62818 227089
rect 62762 227015 62818 227024
rect 62120 226364 62172 226370
rect 62120 226306 62172 226312
rect 62026 224224 62082 224233
rect 62026 224159 62082 224168
rect 60280 221468 60332 221474
rect 60280 221410 60332 221416
rect 60292 217410 60320 221410
rect 61108 219564 61160 219570
rect 61108 219506 61160 219512
rect 61120 217410 61148 219506
rect 62040 217410 62068 224159
rect 62776 217410 62804 227015
rect 65340 222964 65392 222970
rect 65340 222906 65392 222912
rect 63408 221536 63460 221542
rect 63408 221478 63460 221484
rect 63420 217410 63448 221478
rect 64512 220108 64564 220114
rect 64512 220050 64564 220056
rect 64524 217410 64552 220050
rect 65352 217410 65380 222906
rect 66076 222896 66128 222902
rect 66076 222838 66128 222844
rect 66088 217410 66116 222838
rect 66916 219570 66944 229871
rect 67560 229158 67588 231610
rect 84856 231538 84884 247143
rect 85040 231606 85068 247279
rect 171796 241602 171824 249290
rect 414216 248470 414244 249455
rect 414204 248464 414256 248470
rect 414204 248406 414256 248412
rect 190366 248024 190422 248033
rect 190366 247959 190422 247968
rect 171784 241596 171836 241602
rect 171784 241538 171836 241544
rect 164884 241460 164936 241466
rect 164884 241402 164936 241408
rect 85028 231600 85080 231606
rect 85028 231542 85080 231548
rect 84844 231532 84896 231538
rect 84844 231474 84896 231480
rect 136364 230240 136416 230246
rect 136364 230182 136416 230188
rect 132408 229968 132460 229974
rect 132408 229910 132460 229916
rect 91744 229900 91796 229906
rect 91744 229842 91796 229848
rect 85396 229832 85448 229838
rect 85396 229774 85448 229780
rect 71688 229764 71740 229770
rect 71688 229706 71740 229712
rect 67548 229152 67600 229158
rect 67548 229094 67600 229100
rect 69478 224360 69534 224369
rect 69478 224295 69534 224304
rect 68744 223032 68796 223038
rect 68744 222974 68796 222980
rect 66994 221640 67050 221649
rect 66994 221575 67050 221584
rect 66904 219564 66956 219570
rect 66904 219506 66956 219512
rect 67008 217410 67036 221575
rect 67546 220144 67602 220153
rect 67546 220079 67602 220088
rect 67560 217410 67588 220079
rect 68756 217410 68784 222974
rect 69492 217410 69520 224295
rect 70214 221776 70270 221785
rect 70214 221711 70270 221720
rect 70228 217410 70256 221711
rect 71700 220794 71728 229706
rect 77944 228540 77996 228546
rect 77944 228482 77996 228488
rect 72974 227216 73030 227225
rect 72974 227151 73030 227160
rect 72054 224496 72110 224505
rect 72054 224431 72110 224440
rect 71228 220788 71280 220794
rect 71228 220730 71280 220736
rect 71688 220788 71740 220794
rect 71688 220730 71740 220736
rect 71240 217410 71268 220730
rect 72068 217410 72096 224431
rect 72988 217410 73016 227151
rect 76288 225752 76340 225758
rect 76288 225694 76340 225700
rect 75368 223100 75420 223106
rect 75368 223042 75420 223048
rect 73710 221912 73766 221921
rect 73710 221847 73766 221856
rect 73724 217410 73752 221847
rect 74446 220280 74502 220289
rect 74446 220215 74502 220224
rect 74460 217410 74488 220215
rect 75380 217410 75408 223042
rect 76300 217410 76328 225694
rect 77024 221604 77076 221610
rect 77024 221546 77076 221552
rect 77036 217410 77064 221546
rect 77956 217410 77984 228482
rect 82728 227180 82780 227186
rect 82728 227122 82780 227128
rect 78494 224632 78550 224641
rect 78494 224567 78550 224576
rect 78508 217410 78536 224567
rect 82176 223168 82228 223174
rect 82176 223110 82228 223116
rect 80428 221672 80480 221678
rect 80428 221614 80480 221620
rect 79600 220312 79652 220318
rect 79600 220254 79652 220260
rect 79612 217410 79640 220254
rect 80440 217410 80468 221614
rect 81256 220176 81308 220182
rect 81256 220118 81308 220124
rect 81268 217410 81296 220118
rect 82188 217410 82216 223110
rect 82740 217410 82768 227122
rect 83832 221740 83884 221746
rect 83832 221682 83884 221688
rect 83844 217410 83872 221682
rect 85408 220794 85436 229774
rect 91756 228546 91784 229842
rect 120816 229084 120868 229090
rect 120816 229026 120868 229032
rect 117228 229016 117280 229022
rect 117228 228958 117280 228964
rect 114192 228948 114244 228954
rect 114192 228890 114244 228896
rect 110696 228880 110748 228886
rect 110696 228822 110748 228828
rect 107476 228812 107528 228818
rect 107476 228754 107528 228760
rect 103980 228744 104032 228750
rect 103980 228686 104032 228692
rect 100668 228676 100720 228682
rect 100668 228618 100720 228624
rect 97264 228608 97316 228614
rect 97264 228550 97316 228556
rect 91744 228540 91796 228546
rect 91744 228482 91796 228488
rect 93768 228540 93820 228546
rect 93768 228482 93820 228488
rect 90546 228440 90602 228449
rect 90546 228375 90602 228384
rect 86866 228304 86922 228313
rect 86866 228239 86922 228248
rect 86316 225820 86368 225826
rect 86316 225762 86368 225768
rect 85488 221808 85540 221814
rect 85488 221750 85540 221756
rect 84660 220788 84712 220794
rect 84660 220730 84712 220736
rect 85396 220788 85448 220794
rect 85396 220730 85448 220736
rect 84672 217410 84700 220730
rect 85500 217410 85528 221750
rect 86328 217410 86356 225762
rect 86880 217410 86908 228239
rect 89534 225584 89590 225593
rect 89534 225519 89590 225528
rect 88156 224256 88208 224262
rect 88156 224198 88208 224204
rect 88168 217410 88196 224198
rect 88892 221876 88944 221882
rect 88892 221818 88944 221824
rect 88904 217410 88932 221818
rect 89548 217410 89576 225519
rect 90560 217410 90588 228375
rect 91376 227384 91428 227390
rect 91376 227326 91428 227332
rect 91388 217410 91416 227326
rect 93030 225720 93086 225729
rect 93030 225655 93086 225664
rect 92294 223136 92350 223145
rect 92294 223071 92350 223080
rect 92308 217410 92336 223071
rect 93044 217410 93072 225655
rect 93780 217410 93808 228482
rect 96528 225888 96580 225894
rect 96528 225830 96580 225836
rect 95608 223236 95660 223242
rect 95608 223178 95660 223184
rect 94780 220244 94832 220250
rect 94780 220186 94832 220192
rect 94792 217410 94820 220186
rect 95620 217410 95648 223178
rect 96540 217410 96568 225830
rect 97276 217410 97304 228550
rect 99840 225956 99892 225962
rect 99840 225898 99892 225904
rect 99010 223272 99066 223281
rect 99010 223207 99066 223216
rect 97816 219564 97868 219570
rect 97816 219506 97868 219512
rect 97828 217410 97856 219506
rect 99024 217410 99052 223207
rect 99852 217410 99880 225898
rect 100680 217410 100708 228618
rect 103244 226024 103296 226030
rect 103244 225966 103296 225972
rect 101496 224324 101548 224330
rect 101496 224266 101548 224272
rect 100760 222012 100812 222018
rect 100760 221954 100812 221960
rect 100772 220318 100800 221954
rect 100760 220312 100812 220318
rect 100760 220254 100812 220260
rect 101508 217410 101536 224266
rect 101956 223304 102008 223310
rect 101956 223246 102008 223252
rect 52440 217382 52776 217410
rect 53268 217382 53696 217410
rect 54096 217382 54432 217410
rect 54924 217382 55076 217410
rect 55752 217382 56088 217410
rect 56580 217382 56916 217410
rect 57408 217382 57652 217410
rect 58328 217382 58664 217410
rect 59156 217382 59308 217410
rect 59984 217382 60320 217410
rect 60812 217382 61148 217410
rect 61640 217382 62068 217410
rect 62468 217382 62804 217410
rect 63296 217382 63448 217410
rect 64216 217382 64552 217410
rect 65044 217382 65380 217410
rect 65872 217382 66116 217410
rect 66700 217382 67036 217410
rect 67528 217382 67588 217410
rect 68356 217382 68784 217410
rect 69184 217382 69520 217410
rect 70104 217382 70256 217410
rect 70932 217382 71268 217410
rect 71760 217382 72096 217410
rect 72588 217382 73016 217410
rect 73416 217382 73752 217410
rect 74244 217382 74488 217410
rect 75072 217382 75408 217410
rect 75992 217382 76328 217410
rect 76820 217382 77064 217410
rect 77648 217382 77984 217410
rect 78476 217382 78536 217410
rect 79304 217382 79640 217410
rect 80132 217382 80468 217410
rect 80960 217382 81296 217410
rect 81880 217382 82216 217410
rect 82708 217382 82768 217410
rect 83536 217382 83872 217410
rect 84364 217382 84700 217410
rect 85192 217382 85528 217410
rect 86020 217382 86356 217410
rect 86848 217382 86908 217410
rect 87768 217382 88196 217410
rect 88596 217382 88932 217410
rect 89424 217382 89576 217410
rect 90252 217382 90588 217410
rect 91080 217382 91416 217410
rect 91908 217382 92336 217410
rect 92736 217382 93072 217410
rect 93656 217382 93808 217410
rect 94484 217382 94820 217410
rect 95312 217382 95648 217410
rect 96140 217382 96568 217410
rect 96968 217382 97304 217410
rect 97796 217382 97856 217410
rect 98624 217382 99052 217410
rect 99544 217382 99880 217410
rect 100372 217382 100708 217410
rect 101200 217382 101536 217410
rect 101968 217410 101996 223246
rect 103256 217410 103284 225966
rect 103992 217410 104020 228686
rect 106556 226092 106608 226098
rect 106556 226034 106608 226040
rect 105728 223372 105780 223378
rect 105728 223314 105780 223320
rect 104716 220312 104768 220318
rect 104716 220254 104768 220260
rect 104728 217410 104756 220254
rect 105740 217410 105768 223314
rect 106568 217410 106596 226034
rect 107488 217410 107516 228754
rect 108212 227520 108264 227526
rect 108212 227462 108264 227468
rect 108224 217410 108252 227462
rect 109868 226160 109920 226166
rect 109868 226102 109920 226108
rect 108856 223440 108908 223446
rect 108856 223382 108908 223388
rect 108868 217410 108896 223382
rect 109880 217410 109908 226102
rect 110708 217410 110736 228822
rect 112996 226228 113048 226234
rect 112996 226170 113048 226176
rect 112444 221944 112496 221950
rect 112444 221886 112496 221892
rect 111616 220448 111668 220454
rect 111616 220390 111668 220396
rect 111628 217410 111656 220390
rect 112456 217410 112484 221886
rect 113008 217410 113036 226170
rect 114204 217410 114232 228890
rect 116584 226296 116636 226302
rect 116584 226238 116636 226244
rect 114928 224732 114980 224738
rect 114928 224674 114980 224680
rect 114940 217410 114968 224674
rect 115756 223508 115808 223514
rect 115756 223450 115808 223456
rect 115768 217410 115796 223450
rect 116596 217410 116624 226238
rect 117240 217410 117268 228958
rect 119896 225548 119948 225554
rect 119896 225490 119948 225496
rect 119160 222080 119212 222086
rect 119160 222022 119212 222028
rect 118332 220584 118384 220590
rect 118332 220526 118384 220532
rect 118344 217410 118372 220526
rect 119172 217410 119200 222022
rect 119908 217410 119936 225490
rect 120828 217410 120856 229026
rect 127532 228336 127584 228342
rect 127532 228278 127584 228284
rect 124128 227044 124180 227050
rect 124128 226986 124180 226992
rect 123392 225480 123444 225486
rect 123392 225422 123444 225428
rect 122472 222148 122524 222154
rect 122472 222090 122524 222096
rect 121276 220516 121328 220522
rect 121276 220458 121328 220464
rect 101968 217382 102028 217410
rect 102856 217382 103284 217410
rect 103684 217382 104020 217410
rect 104512 217382 104756 217410
rect 105432 217382 105768 217410
rect 106260 217382 106596 217410
rect 107088 217382 107516 217410
rect 107916 217382 108252 217410
rect 108744 217382 108896 217410
rect 109572 217382 109908 217410
rect 110400 217382 110736 217410
rect 111320 217382 111656 217410
rect 112148 217382 112484 217410
rect 112976 217382 113036 217410
rect 113804 217382 114232 217410
rect 114632 217382 114968 217410
rect 115460 217382 115796 217410
rect 116288 217382 116624 217410
rect 117208 217382 117268 217410
rect 118036 217382 118372 217410
rect 118864 217382 119200 217410
rect 119692 217382 119936 217410
rect 120520 217382 120856 217410
rect 121288 217410 121316 220458
rect 122484 217410 122512 222090
rect 123404 217410 123432 225422
rect 124140 217410 124168 226986
rect 125048 226976 125100 226982
rect 125048 226918 125100 226924
rect 125060 217410 125088 226918
rect 126796 225412 126848 225418
rect 126796 225354 126848 225360
rect 125876 223576 125928 223582
rect 125876 223518 125928 223524
rect 125888 217410 125916 223518
rect 126808 217410 126836 225354
rect 127544 217410 127572 228278
rect 131028 228268 131080 228274
rect 131028 228210 131080 228216
rect 130108 225344 130160 225350
rect 130108 225286 130160 225292
rect 129280 221400 129332 221406
rect 129280 221342 129332 221348
rect 128176 220652 128228 220658
rect 128176 220594 128228 220600
rect 128188 217410 128216 220594
rect 129292 217410 129320 221342
rect 130120 217410 130148 225286
rect 131040 217410 131068 228210
rect 132316 222828 132368 222834
rect 132316 222770 132368 222776
rect 131764 220788 131816 220794
rect 131764 220730 131816 220736
rect 131776 217410 131804 220730
rect 132328 217410 132356 222770
rect 132420 220794 132448 229910
rect 134248 227112 134300 227118
rect 134248 227054 134300 227060
rect 133512 225276 133564 225282
rect 133512 225218 133564 225224
rect 132408 220788 132460 220794
rect 132408 220730 132460 220736
rect 133524 217410 133552 225218
rect 134260 217410 134288 227054
rect 135996 224392 136048 224398
rect 135996 224334 136048 224340
rect 134984 220720 135036 220726
rect 134984 220662 135036 220668
rect 134996 217410 135024 220662
rect 136008 217410 136036 224334
rect 136376 224330 136404 230182
rect 155868 230172 155920 230178
rect 155868 230114 155920 230120
rect 146208 230104 146260 230110
rect 146208 230046 146260 230052
rect 139308 230036 139360 230042
rect 139308 229978 139360 229984
rect 137744 228200 137796 228206
rect 137744 228142 137796 228148
rect 136364 224324 136416 224330
rect 136364 224266 136416 224272
rect 136456 224324 136508 224330
rect 136456 224266 136508 224272
rect 121288 217382 121348 217410
rect 122176 217382 122512 217410
rect 123096 217382 123432 217410
rect 123924 217382 124168 217410
rect 124752 217382 125088 217410
rect 125580 217382 125916 217410
rect 126408 217382 126836 217410
rect 127236 217382 127572 217410
rect 128064 217382 128216 217410
rect 128984 217382 129320 217410
rect 129812 217382 130148 217410
rect 130640 217382 131068 217410
rect 131468 217382 131804 217410
rect 132296 217382 132356 217410
rect 133124 217382 133552 217410
rect 133952 217382 134288 217410
rect 134872 217382 135024 217410
rect 135700 217382 136036 217410
rect 136468 217410 136496 224266
rect 137756 217410 137784 228142
rect 139216 224460 139268 224466
rect 139216 224402 139268 224408
rect 138480 220788 138532 220794
rect 138480 220730 138532 220736
rect 138492 217410 138520 220730
rect 139228 217410 139256 224402
rect 139320 220794 139348 229978
rect 140044 229696 140096 229702
rect 140044 229638 140096 229644
rect 140056 227186 140084 229638
rect 144368 228132 144420 228138
rect 144368 228074 144420 228080
rect 141056 227316 141108 227322
rect 141056 227258 141108 227264
rect 140044 227180 140096 227186
rect 140044 227122 140096 227128
rect 140136 227180 140188 227186
rect 140136 227122 140188 227128
rect 139308 220788 139360 220794
rect 139308 220730 139360 220736
rect 140148 217410 140176 227122
rect 141068 217410 141096 227258
rect 143448 227248 143500 227254
rect 143448 227190 143500 227196
rect 142712 224528 142764 224534
rect 142712 224470 142764 224476
rect 141884 220788 141936 220794
rect 141884 220730 141936 220736
rect 141896 217410 141924 220730
rect 142724 217410 142752 224470
rect 143460 217410 143488 227190
rect 144380 217410 144408 228074
rect 146116 224596 146168 224602
rect 146116 224538 146168 224544
rect 145196 220380 145248 220386
rect 145196 220322 145248 220328
rect 145208 217410 145236 220322
rect 146128 217410 146156 224538
rect 146220 220386 146248 230046
rect 151820 229628 151872 229634
rect 151820 229570 151872 229576
rect 149704 229560 149756 229566
rect 149704 229502 149756 229508
rect 146392 229492 146444 229498
rect 146392 229434 146444 229440
rect 146404 227390 146432 229434
rect 149716 227526 149744 229502
rect 149704 227520 149756 227526
rect 149704 227462 149756 227468
rect 150348 227520 150400 227526
rect 150348 227462 150400 227468
rect 147496 227452 147548 227458
rect 147496 227394 147548 227400
rect 146392 227384 146444 227390
rect 146392 227326 146444 227332
rect 146944 227384 146996 227390
rect 146944 227326 146996 227332
rect 146208 220380 146260 220386
rect 146208 220322 146260 220328
rect 146956 217410 146984 227326
rect 147508 217410 147536 227394
rect 149428 224664 149480 224670
rect 149428 224606 149480 224612
rect 148600 220040 148652 220046
rect 148600 219982 148652 219988
rect 148612 217410 148640 219982
rect 149440 217410 149468 224606
rect 150360 217410 150388 227462
rect 151832 224738 151860 229570
rect 154488 228064 154540 228070
rect 154488 228006 154540 228012
rect 153660 227588 153712 227594
rect 153660 227530 153712 227536
rect 151820 224732 151872 224738
rect 151820 224674 151872 224680
rect 152924 224732 152976 224738
rect 152924 224674 152976 224680
rect 151084 221332 151136 221338
rect 151084 221274 151136 221280
rect 151096 217410 151124 221274
rect 151728 219972 151780 219978
rect 151728 219914 151780 219920
rect 151740 217410 151768 219914
rect 152936 217410 152964 224674
rect 153672 217410 153700 227530
rect 154500 217410 154528 228006
rect 155776 224800 155828 224806
rect 155776 224742 155828 224748
rect 155316 220380 155368 220386
rect 155316 220322 155368 220328
rect 155328 217410 155356 220322
rect 136468 217382 136528 217410
rect 137356 217382 137784 217410
rect 138184 217382 138520 217410
rect 139012 217382 139256 217410
rect 139840 217382 140176 217410
rect 140760 217382 141096 217410
rect 141588 217382 141924 217410
rect 142416 217382 142752 217410
rect 143244 217382 143488 217410
rect 144072 217382 144408 217410
rect 144900 217382 145236 217410
rect 145728 217382 146156 217410
rect 146648 217382 146984 217410
rect 147476 217382 147536 217410
rect 148304 217382 148640 217410
rect 149132 217382 149468 217410
rect 149960 217382 150388 217410
rect 150788 217382 151124 217410
rect 151616 217382 151768 217410
rect 152536 217382 152964 217410
rect 153364 217382 153700 217410
rect 154192 217382 154528 217410
rect 155020 217382 155356 217410
rect 155788 217410 155816 224742
rect 155880 220386 155908 230114
rect 162860 229356 162912 229362
rect 162860 229298 162912 229304
rect 161296 227996 161348 228002
rect 161296 227938 161348 227944
rect 160376 227724 160428 227730
rect 160376 227666 160428 227672
rect 157064 227656 157116 227662
rect 157064 227598 157116 227604
rect 155868 220380 155920 220386
rect 155868 220322 155920 220328
rect 157076 217410 157104 227598
rect 159548 224868 159600 224874
rect 159548 224810 159600 224816
rect 157800 221264 157852 221270
rect 157800 221206 157852 221212
rect 157812 217410 157840 221206
rect 158628 219904 158680 219910
rect 158628 219846 158680 219852
rect 158640 217410 158668 219846
rect 159560 217410 159588 224810
rect 160388 217410 160416 227666
rect 161308 217410 161336 227938
rect 162872 226982 162900 229298
rect 162860 226976 162912 226982
rect 162860 226918 162912 226924
rect 163688 226976 163740 226982
rect 163688 226918 163740 226924
rect 162768 224936 162820 224942
rect 162768 224878 162820 224884
rect 162032 222692 162084 222698
rect 162032 222634 162084 222640
rect 162044 217410 162072 222634
rect 162780 217410 162808 224878
rect 163700 217410 163728 226918
rect 164608 226840 164660 226846
rect 164608 226782 164660 226788
rect 164620 217410 164648 226782
rect 155788 217382 155848 217410
rect 156676 217382 157104 217410
rect 157504 217382 157840 217410
rect 158424 217382 158668 217410
rect 159252 217382 159588 217410
rect 160080 217382 160416 217410
rect 160908 217382 161336 217410
rect 161736 217382 162072 217410
rect 162564 217382 162808 217410
rect 163392 217382 163728 217410
rect 164312 217382 164648 217410
rect 164896 217326 164924 241402
rect 185584 237448 185636 237454
rect 189080 237448 189132 237454
rect 185584 237390 185636 237396
rect 189078 237416 189080 237425
rect 189132 237416 189134 237425
rect 185596 235006 185624 237390
rect 189078 237351 189134 237360
rect 182916 235000 182968 235006
rect 182916 234942 182968 234948
rect 185584 235000 185636 235006
rect 185584 234942 185636 234948
rect 182928 233510 182956 234942
rect 178040 233504 178092 233510
rect 178040 233446 178092 233452
rect 182916 233504 182968 233510
rect 182916 233446 182968 233452
rect 178052 231674 178080 233446
rect 190380 231742 190408 247959
rect 415306 246392 415362 246401
rect 415306 246327 415362 246336
rect 415320 245682 415348 246327
rect 191104 245676 191156 245682
rect 191104 245618 191156 245624
rect 415308 245676 415360 245682
rect 415308 245618 415360 245624
rect 565084 245676 565136 245682
rect 565084 245618 565136 245624
rect 190368 231736 190420 231742
rect 190368 231678 190420 231684
rect 191116 231674 191144 245618
rect 414386 243128 414442 243137
rect 414386 243063 414442 243072
rect 414400 242962 414428 243063
rect 414388 242956 414440 242962
rect 414388 242898 414440 242904
rect 414294 240000 414350 240009
rect 414294 239935 414350 239944
rect 414202 233608 414258 233617
rect 414202 233543 414258 233552
rect 414216 232558 414244 233543
rect 414204 232552 414256 232558
rect 414204 232494 414256 232500
rect 414308 232422 414336 239935
rect 414938 236736 414994 236745
rect 414938 236671 414994 236680
rect 414952 232490 414980 236671
rect 414940 232484 414992 232490
rect 414940 232426 414992 232432
rect 414296 232416 414348 232422
rect 414296 232358 414348 232364
rect 178040 231668 178092 231674
rect 178040 231610 178092 231616
rect 191104 231668 191156 231674
rect 191104 231610 191156 231616
rect 179328 230444 179380 230450
rect 179328 230386 179380 230392
rect 175188 230376 175240 230382
rect 175188 230318 175240 230324
rect 169668 230308 169720 230314
rect 169668 230250 169720 230256
rect 166908 226908 166960 226914
rect 166908 226850 166960 226856
rect 166264 224188 166316 224194
rect 166264 224130 166316 224136
rect 165436 219836 165488 219842
rect 165436 219778 165488 219784
rect 165448 217410 165476 219778
rect 166276 217410 166304 224130
rect 166920 217410 166948 226850
rect 169576 224120 169628 224126
rect 169576 224062 169628 224068
rect 167920 221196 167972 221202
rect 167920 221138 167972 221144
rect 167932 217410 167960 221138
rect 168748 220380 168800 220386
rect 168748 220322 168800 220328
rect 168760 217410 168788 220322
rect 169588 217410 169616 224062
rect 169680 220386 169708 230250
rect 171048 227928 171100 227934
rect 171048 227870 171100 227876
rect 170496 225208 170548 225214
rect 170496 225150 170548 225156
rect 169668 220380 169720 220386
rect 169668 220322 169720 220328
rect 170508 217410 170536 225150
rect 171060 217410 171088 227870
rect 173808 226772 173860 226778
rect 173808 226714 173860 226720
rect 172980 224052 173032 224058
rect 172980 223994 173032 224000
rect 172152 219768 172204 219774
rect 172152 219710 172204 219716
rect 172164 217410 172192 219710
rect 172992 217410 173020 223994
rect 173820 217410 173848 226714
rect 174636 226704 174688 226710
rect 174636 226646 174688 226652
rect 174648 217410 174676 226646
rect 175200 217410 175228 230318
rect 177212 226636 177264 226642
rect 177212 226578 177264 226584
rect 176476 223984 176528 223990
rect 176476 223926 176528 223932
rect 176488 217410 176516 223926
rect 177224 217410 177252 226578
rect 177856 222760 177908 222766
rect 177856 222702 177908 222708
rect 177868 217410 177896 222702
rect 179340 220386 179368 230386
rect 186964 229424 187016 229430
rect 186964 229366 187016 229372
rect 180800 229288 180852 229294
rect 180800 229230 180852 229236
rect 180616 225140 180668 225146
rect 180616 225082 180668 225088
rect 179696 223916 179748 223922
rect 179696 223858 179748 223864
rect 178868 220380 178920 220386
rect 178868 220322 178920 220328
rect 179328 220380 179380 220386
rect 179328 220322 179380 220328
rect 178880 217410 178908 220322
rect 179708 217410 179736 223858
rect 180628 217410 180656 225082
rect 180812 222698 180840 229230
rect 183192 223848 183244 223854
rect 183192 223790 183244 223796
rect 180800 222692 180852 222698
rect 180800 222634 180852 222640
rect 181352 222692 181404 222698
rect 181352 222634 181404 222640
rect 181364 217410 181392 222634
rect 181996 219632 182048 219638
rect 181996 219574 182048 219580
rect 182008 217410 182036 219574
rect 183204 217410 183232 223790
rect 186228 223780 186280 223786
rect 186228 223722 186280 223728
rect 184756 222556 184808 222562
rect 184756 222498 184808 222504
rect 183928 221128 183980 221134
rect 183928 221070 183980 221076
rect 183940 217410 183968 221070
rect 184768 217410 184796 222498
rect 185584 219700 185636 219706
rect 185584 219642 185636 219648
rect 185596 217410 185624 219642
rect 186240 217410 186268 223722
rect 186976 219706 187004 229366
rect 192312 228410 192340 231676
rect 192404 231662 192602 231690
rect 192680 231662 192970 231690
rect 192300 228404 192352 228410
rect 192300 228346 192352 228352
rect 190276 226568 190328 226574
rect 190276 226510 190328 226516
rect 187332 222624 187384 222630
rect 187332 222566 187384 222572
rect 186964 219700 187016 219706
rect 186964 219642 187016 219648
rect 187344 217410 187372 222566
rect 188160 222488 188212 222494
rect 188160 222430 188212 222436
rect 188172 217410 188200 222430
rect 189816 221060 189868 221066
rect 189816 221002 189868 221008
rect 188896 219632 188948 219638
rect 188896 219574 188948 219580
rect 188908 217410 188936 219574
rect 189828 217410 189856 221002
rect 165140 217382 165476 217410
rect 165968 217382 166304 217410
rect 166796 217382 166948 217410
rect 167624 217382 167960 217410
rect 168452 217382 168788 217410
rect 169280 217382 169616 217410
rect 170200 217382 170536 217410
rect 171028 217382 171088 217410
rect 171856 217382 172192 217410
rect 172684 217382 173020 217410
rect 173512 217382 173848 217410
rect 174340 217382 174676 217410
rect 175168 217382 175228 217410
rect 176088 217382 176516 217410
rect 176916 217382 177252 217410
rect 177744 217382 177896 217410
rect 178572 217382 178908 217410
rect 179400 217382 179736 217410
rect 180228 217382 180656 217410
rect 181056 217382 181392 217410
rect 181976 217382 182036 217410
rect 182804 217382 183232 217410
rect 183632 217382 183968 217410
rect 184460 217382 184796 217410
rect 185288 217382 185624 217410
rect 186116 217382 186268 217410
rect 186944 217382 187372 217410
rect 187864 217382 188200 217410
rect 188692 217382 188936 217410
rect 189520 217382 189856 217410
rect 190288 217410 190316 226510
rect 192404 222873 192432 231662
rect 192680 225622 192708 231662
rect 193324 228478 193352 231676
rect 193416 231662 193706 231690
rect 193312 228472 193364 228478
rect 193312 228414 193364 228420
rect 192668 225616 192720 225622
rect 192668 225558 192720 225564
rect 192852 225004 192904 225010
rect 192852 224946 192904 224952
rect 192390 222864 192446 222873
rect 192390 222799 192446 222808
rect 191564 222420 191616 222426
rect 191564 222362 191616 222368
rect 191576 217410 191604 222362
rect 192300 220380 192352 220386
rect 192300 220322 192352 220328
rect 192312 217410 192340 220322
rect 192864 220114 192892 224946
rect 193416 221513 193444 231662
rect 194060 223009 194088 231676
rect 194140 228404 194192 228410
rect 194140 228346 194192 228352
rect 194046 223000 194102 223009
rect 194046 222935 194102 222944
rect 193402 221504 193458 221513
rect 193402 221439 193458 221448
rect 192944 220992 192996 220998
rect 192944 220934 192996 220940
rect 192852 220108 192904 220114
rect 192852 220050 192904 220056
rect 192956 217410 192984 220934
rect 194152 219434 194180 228346
rect 194428 225690 194456 231676
rect 194796 229809 194824 231676
rect 194888 231662 195178 231690
rect 194782 229800 194838 229809
rect 194782 229735 194838 229744
rect 194416 225684 194468 225690
rect 194416 225626 194468 225632
rect 194888 221474 194916 231662
rect 194968 228472 195020 228478
rect 194968 228414 195020 228420
rect 194876 221468 194928 221474
rect 194876 221410 194928 221416
rect 194980 219434 195008 228414
rect 195440 224233 195468 231676
rect 195808 226953 195836 231676
rect 196176 229945 196204 231676
rect 196268 231662 196558 231690
rect 196162 229936 196218 229945
rect 196162 229871 196218 229880
rect 195794 226944 195850 226953
rect 195794 226879 195850 226888
rect 195426 224224 195482 224233
rect 195426 224159 195482 224168
rect 196268 221542 196296 231662
rect 196622 230344 196678 230353
rect 196622 230279 196678 230288
rect 196532 222352 196584 222358
rect 196532 222294 196584 222300
rect 196256 221536 196308 221542
rect 196256 221478 196308 221484
rect 195152 220924 195204 220930
rect 195152 220866 195204 220872
rect 195164 219502 195192 220866
rect 195704 219564 195756 219570
rect 195704 219506 195756 219512
rect 195152 219496 195204 219502
rect 195152 219438 195204 219444
rect 194060 219406 194180 219434
rect 194888 219406 195008 219434
rect 194060 217410 194088 219406
rect 194888 217410 194916 219406
rect 195716 217410 195744 219506
rect 196544 217410 196572 222294
rect 196636 220153 196664 230279
rect 196912 222970 196940 231676
rect 197280 227089 197308 231676
rect 197266 227080 197322 227089
rect 197266 227015 197322 227024
rect 197648 225010 197676 231676
rect 197740 231662 198030 231690
rect 197636 225004 197688 225010
rect 197636 224946 197688 224952
rect 196900 222964 196952 222970
rect 196900 222906 196952 222912
rect 197740 221649 197768 231662
rect 198188 223032 198240 223038
rect 198188 222974 198240 222980
rect 197726 221640 197782 221649
rect 197726 221575 197782 221584
rect 197268 221536 197320 221542
rect 197268 221478 197320 221484
rect 196622 220144 196678 220153
rect 196622 220079 196678 220088
rect 197280 217410 197308 221478
rect 198200 217410 198228 222974
rect 198292 222970 198320 231676
rect 198384 231662 198674 231690
rect 198280 222964 198332 222970
rect 198280 222906 198332 222912
rect 198384 222902 198412 231662
rect 199028 230353 199056 231676
rect 199120 231662 199410 231690
rect 199014 230344 199070 230353
rect 199014 230279 199070 230288
rect 199016 225684 199068 225690
rect 199016 225626 199068 225632
rect 198372 222896 198424 222902
rect 198372 222838 198424 222844
rect 199028 217410 199056 225626
rect 199120 221785 199148 231662
rect 199764 224505 199792 231676
rect 199750 224496 199806 224505
rect 199750 224431 199806 224440
rect 200132 224369 200160 231676
rect 200500 229770 200528 231676
rect 200592 231662 200882 231690
rect 200488 229764 200540 229770
rect 200488 229706 200540 229712
rect 200118 224360 200174 224369
rect 200118 224295 200174 224304
rect 199936 222964 199988 222970
rect 199936 222906 199988 222912
rect 199106 221776 199162 221785
rect 199106 221711 199162 221720
rect 199948 217410 199976 222906
rect 200592 221921 200620 231662
rect 200672 229764 200724 229770
rect 200672 229706 200724 229712
rect 200684 225690 200712 229706
rect 200672 225684 200724 225690
rect 200672 225626 200724 225632
rect 201144 223106 201172 231676
rect 201512 227225 201540 231676
rect 201604 231662 201894 231690
rect 201972 231662 202262 231690
rect 201498 227216 201554 227225
rect 201498 227151 201554 227160
rect 201408 225616 201460 225622
rect 201408 225558 201460 225564
rect 201132 223100 201184 223106
rect 201132 223042 201184 223048
rect 200764 222896 200816 222902
rect 200764 222838 200816 222844
rect 200578 221912 200634 221921
rect 200578 221847 200634 221856
rect 200776 217410 200804 222838
rect 201420 217410 201448 225558
rect 201604 220289 201632 231662
rect 201972 221610 202000 231662
rect 202616 224641 202644 231676
rect 202984 225758 203012 231676
rect 203352 229906 203380 231676
rect 203444 231662 203734 231690
rect 203340 229900 203392 229906
rect 203340 229842 203392 229848
rect 202972 225752 203024 225758
rect 202972 225694 203024 225700
rect 203248 225684 203300 225690
rect 203248 225626 203300 225632
rect 202602 224632 202658 224641
rect 202602 224567 202658 224576
rect 201960 221604 202012 221610
rect 201960 221546 202012 221552
rect 202420 221604 202472 221610
rect 202420 221546 202472 221552
rect 201590 220280 201646 220289
rect 202432 220250 202460 221546
rect 201590 220215 201646 220224
rect 202420 220244 202472 220250
rect 202420 220186 202472 220192
rect 202420 219496 202472 219502
rect 202420 219438 202472 219444
rect 202432 217410 202460 219438
rect 203260 217410 203288 225626
rect 203444 221678 203472 231662
rect 203996 223174 204024 231676
rect 204378 231662 204484 231690
rect 203984 223168 204036 223174
rect 203984 223110 204036 223116
rect 204456 222018 204484 231662
rect 204548 231662 204746 231690
rect 204824 231662 205114 231690
rect 205192 231662 205482 231690
rect 204444 222012 204496 222018
rect 204444 221954 204496 221960
rect 203432 221672 203484 221678
rect 203432 221614 203484 221620
rect 203708 221672 203760 221678
rect 203708 221614 203760 221620
rect 203720 220318 203748 221614
rect 203708 220312 203760 220318
rect 203708 220254 203760 220260
rect 204548 220250 204576 231662
rect 204824 221746 204852 231662
rect 204904 223100 204956 223106
rect 204904 223042 204956 223048
rect 204812 221740 204864 221746
rect 204812 221682 204864 221688
rect 204536 220244 204588 220250
rect 204536 220186 204588 220192
rect 204076 220176 204128 220182
rect 204076 220118 204128 220124
rect 204088 217410 204116 220118
rect 204916 217410 204944 223042
rect 205192 221814 205220 231662
rect 205836 229702 205864 231676
rect 206204 229838 206232 231676
rect 206192 229832 206244 229838
rect 206192 229774 206244 229780
rect 205824 229696 205876 229702
rect 205824 229638 205876 229644
rect 206572 228313 206600 231676
rect 206664 231662 206862 231690
rect 206558 228304 206614 228313
rect 206558 228239 206614 228248
rect 205548 221876 205600 221882
rect 205548 221818 205600 221824
rect 205180 221808 205232 221814
rect 205180 221750 205232 221756
rect 205560 217410 205588 221818
rect 206664 221814 206692 231662
rect 206744 229832 206796 229838
rect 206744 229774 206796 229780
rect 206756 221882 206784 229774
rect 207216 225826 207244 231676
rect 207204 225820 207256 225826
rect 207204 225762 207256 225768
rect 206836 225752 206888 225758
rect 206836 225694 206888 225700
rect 206744 221876 206796 221882
rect 206744 221818 206796 221824
rect 206652 221808 206704 221814
rect 206652 221750 206704 221756
rect 206192 220516 206244 220522
rect 206192 220458 206244 220464
rect 206204 220318 206232 220458
rect 206192 220312 206244 220318
rect 206192 220254 206244 220260
rect 206848 217410 206876 225694
rect 207584 224262 207612 231676
rect 207952 228449 207980 231676
rect 208044 231662 208334 231690
rect 207938 228440 207994 228449
rect 207938 228375 207994 228384
rect 207572 224256 207624 224262
rect 207572 224198 207624 224204
rect 208044 223145 208072 231662
rect 208308 225820 208360 225826
rect 208308 225762 208360 225768
rect 208030 223136 208086 223145
rect 208030 223071 208086 223080
rect 208216 221808 208268 221814
rect 208216 221750 208268 221756
rect 206928 221740 206980 221746
rect 206928 221682 206980 221688
rect 206940 220454 206968 221682
rect 208228 220522 208256 221750
rect 208216 220516 208268 220522
rect 208216 220458 208268 220464
rect 206928 220448 206980 220454
rect 206928 220390 206980 220396
rect 207480 220244 207532 220250
rect 207480 220186 207532 220192
rect 207492 217410 207520 220186
rect 208320 217410 208348 225762
rect 208688 225593 208716 231676
rect 209056 229498 209084 231676
rect 209044 229492 209096 229498
rect 209044 229434 209096 229440
rect 209424 228546 209452 231676
rect 209412 228540 209464 228546
rect 209412 228482 209464 228488
rect 208674 225584 208730 225593
rect 208674 225519 208730 225528
rect 209700 223174 209728 231676
rect 209872 228540 209924 228546
rect 209872 228482 209924 228488
rect 209688 223168 209740 223174
rect 209688 223110 209740 223116
rect 209688 221468 209740 221474
rect 209688 221410 209740 221416
rect 209136 220108 209188 220114
rect 209136 220050 209188 220056
rect 209148 217410 209176 220050
rect 209700 217410 209728 221410
rect 209884 220182 209912 228482
rect 210068 225729 210096 231676
rect 210160 231662 210450 231690
rect 210054 225720 210110 225729
rect 210054 225655 210110 225664
rect 210160 221610 210188 231662
rect 210804 228614 210832 231676
rect 210792 228608 210844 228614
rect 210792 228550 210844 228556
rect 210424 223508 210476 223514
rect 210424 223450 210476 223456
rect 210436 223310 210464 223450
rect 210424 223304 210476 223310
rect 211172 223281 211200 231676
rect 211540 225894 211568 231676
rect 211632 231662 211922 231690
rect 211528 225888 211580 225894
rect 211528 225830 211580 225836
rect 210424 223246 210476 223252
rect 211158 223272 211214 223281
rect 211158 223207 211214 223216
rect 210148 221604 210200 221610
rect 210148 221546 210200 221552
rect 211632 220930 211660 231662
rect 212276 228682 212304 231676
rect 212448 229900 212500 229906
rect 212448 229842 212500 229848
rect 212264 228676 212316 228682
rect 212264 228618 212316 228624
rect 211712 225888 211764 225894
rect 211712 225830 211764 225836
rect 211620 220924 211672 220930
rect 211620 220866 211672 220872
rect 209872 220176 209924 220182
rect 209872 220118 209924 220124
rect 210792 220176 210844 220182
rect 210792 220118 210844 220124
rect 210804 217410 210832 220118
rect 211724 217410 211752 225830
rect 212460 217410 212488 229842
rect 212552 223242 212580 231676
rect 212920 225962 212948 231676
rect 213288 230246 213316 231676
rect 213276 230240 213328 230246
rect 213276 230182 213328 230188
rect 213656 228750 213684 231676
rect 213644 228744 213696 228750
rect 213644 228686 213696 228692
rect 213828 228608 213880 228614
rect 213828 228550 213880 228556
rect 212908 225956 212960 225962
rect 212908 225898 212960 225904
rect 212540 223236 212592 223242
rect 212540 223178 212592 223184
rect 213368 221604 213420 221610
rect 213368 221546 213420 221552
rect 213380 217410 213408 221546
rect 213840 220250 213868 228550
rect 213920 223508 213972 223514
rect 213920 223450 213972 223456
rect 213932 220318 213960 223450
rect 214024 223378 214052 231676
rect 214392 226030 214420 231676
rect 214484 231662 214774 231690
rect 214380 226024 214432 226030
rect 214380 225966 214432 225972
rect 214012 223372 214064 223378
rect 214012 223314 214064 223320
rect 214484 221678 214512 231662
rect 215128 228818 215156 231676
rect 215116 228812 215168 228818
rect 215116 228754 215168 228760
rect 215116 228676 215168 228682
rect 215116 228618 215168 228624
rect 214472 221672 214524 221678
rect 214472 221614 214524 221620
rect 214196 220720 214248 220726
rect 214196 220662 214248 220668
rect 213920 220312 213972 220318
rect 213920 220254 213972 220260
rect 213828 220244 213880 220250
rect 213828 220186 213880 220192
rect 214208 217410 214236 220662
rect 215128 217410 215156 228618
rect 215300 225956 215352 225962
rect 215300 225898 215352 225904
rect 215312 220726 215340 225898
rect 215404 223446 215432 231676
rect 215772 226098 215800 231676
rect 216140 229566 216168 231676
rect 216128 229560 216180 229566
rect 216128 229502 216180 229508
rect 216508 228886 216536 231676
rect 216784 231662 216890 231690
rect 216496 228880 216548 228886
rect 216496 228822 216548 228828
rect 216680 228812 216732 228818
rect 216680 228754 216732 228760
rect 215760 226092 215812 226098
rect 215760 226034 215812 226040
rect 215392 223440 215444 223446
rect 215392 223382 215444 223388
rect 216588 221672 216640 221678
rect 216588 221614 216640 221620
rect 215300 220720 215352 220726
rect 215300 220662 215352 220668
rect 215852 220244 215904 220250
rect 215852 220186 215904 220192
rect 215864 217410 215892 220186
rect 216600 217410 216628 221614
rect 216692 220590 216720 228754
rect 216784 221950 216812 231662
rect 217244 226166 217272 231676
rect 217336 231662 217626 231690
rect 217232 226160 217284 226166
rect 217232 226102 217284 226108
rect 216772 221944 216824 221950
rect 216772 221886 216824 221892
rect 217336 221746 217364 231662
rect 217980 228954 218008 231676
rect 217968 228948 218020 228954
rect 217968 228890 218020 228896
rect 218060 226160 218112 226166
rect 218060 226102 218112 226108
rect 217324 221740 217376 221746
rect 217324 221682 217376 221688
rect 218072 220658 218100 226102
rect 218256 223310 218284 231676
rect 218624 226234 218652 231676
rect 218992 229634 219020 231676
rect 219256 230240 219308 230246
rect 219256 230182 219308 230188
rect 218980 229628 219032 229634
rect 218980 229570 219032 229576
rect 218612 226228 218664 226234
rect 218612 226170 218664 226176
rect 218244 223304 218296 223310
rect 218244 223246 218296 223252
rect 218428 221740 218480 221746
rect 218428 221682 218480 221688
rect 218060 220652 218112 220658
rect 218060 220594 218112 220600
rect 216680 220584 216732 220590
rect 216680 220526 216732 220532
rect 217600 220312 217652 220318
rect 217600 220254 217652 220260
rect 217612 217410 217640 220254
rect 218440 217410 218468 221682
rect 219268 217410 219296 230182
rect 219360 229022 219388 231676
rect 219544 231662 219742 231690
rect 219348 229016 219400 229022
rect 219348 228958 219400 228964
rect 219544 222086 219572 231662
rect 220096 226302 220124 231676
rect 220188 231662 220478 231690
rect 220084 226296 220136 226302
rect 220084 226238 220136 226244
rect 219532 222080 219584 222086
rect 219532 222022 219584 222028
rect 220084 221876 220136 221882
rect 220084 221818 220136 221824
rect 220096 217410 220124 221818
rect 220188 221814 220216 231662
rect 220832 229090 220860 231676
rect 221016 231662 221122 231690
rect 221200 231662 221490 231690
rect 220820 229084 220872 229090
rect 220820 229026 220872 229032
rect 220636 226024 220688 226030
rect 220636 225966 220688 225972
rect 220176 221808 220228 221814
rect 220176 221750 220228 221756
rect 220648 217410 220676 225966
rect 221016 222154 221044 231662
rect 221200 225554 221228 231662
rect 221188 225548 221240 225554
rect 221188 225490 221240 225496
rect 221844 223514 221872 231676
rect 222108 228744 222160 228750
rect 222108 228686 222160 228692
rect 221832 223508 221884 223514
rect 221832 223450 221884 223456
rect 221004 222148 221056 222154
rect 221004 222090 221056 222096
rect 221740 221808 221792 221814
rect 221740 221750 221792 221756
rect 221752 217410 221780 221750
rect 222120 220794 222148 228686
rect 222212 227050 222240 231676
rect 222200 227044 222252 227050
rect 222200 226986 222252 226992
rect 222580 223582 222608 231676
rect 222948 225486 222976 231676
rect 223316 229362 223344 231676
rect 223304 229356 223356 229362
rect 223304 229298 223356 229304
rect 223684 228342 223712 231676
rect 223776 231662 223974 231690
rect 223672 228336 223724 228342
rect 223672 228278 223724 228284
rect 223120 226228 223172 226234
rect 223120 226170 223172 226176
rect 222936 225480 222988 225486
rect 222936 225422 222988 225428
rect 222568 223576 222620 223582
rect 222568 223518 222620 223524
rect 222108 220788 222160 220794
rect 222108 220730 222160 220736
rect 222568 220448 222620 220454
rect 222568 220390 222620 220396
rect 222580 217410 222608 220390
rect 223132 220046 223160 226170
rect 223488 221944 223540 221950
rect 223488 221886 223540 221892
rect 223120 220040 223172 220046
rect 223120 219982 223172 219988
rect 223500 217410 223528 221886
rect 223776 221406 223804 231662
rect 224040 228948 224092 228954
rect 224040 228890 224092 228896
rect 223764 221400 223816 221406
rect 223764 221342 223816 221348
rect 224052 219978 224080 228890
rect 224328 225418 224356 231676
rect 224696 228818 224724 231676
rect 224684 228812 224736 228818
rect 224684 228754 224736 228760
rect 225064 228274 225092 231676
rect 225052 228268 225104 228274
rect 225052 228210 225104 228216
rect 224960 226092 225012 226098
rect 224960 226034 225012 226040
rect 224316 225412 224368 225418
rect 224316 225354 224368 225360
rect 224868 222012 224920 222018
rect 224868 221954 224920 221960
rect 224316 220380 224368 220386
rect 224316 220322 224368 220328
rect 224040 219972 224092 219978
rect 224040 219914 224092 219920
rect 224328 217410 224356 220322
rect 224880 217410 224908 221954
rect 224972 220522 225000 226034
rect 225432 222834 225460 231676
rect 225800 225350 225828 231676
rect 226168 229974 226196 231676
rect 226156 229968 226208 229974
rect 226156 229910 226208 229916
rect 226248 229968 226300 229974
rect 226248 229910 226300 229916
rect 225788 225344 225840 225350
rect 225788 225286 225840 225292
rect 225420 222828 225472 222834
rect 225420 222770 225472 222776
rect 224960 220516 225012 220522
rect 224960 220458 225012 220464
rect 226260 219434 226288 229910
rect 226536 227118 226564 231676
rect 226524 227112 226576 227118
rect 226524 227054 226576 227060
rect 226812 224398 226840 231676
rect 227180 225282 227208 231676
rect 227272 231662 227562 231690
rect 227272 226166 227300 231662
rect 227536 229696 227588 229702
rect 227536 229638 227588 229644
rect 227260 226160 227312 226166
rect 227260 226102 227312 226108
rect 227352 226160 227404 226166
rect 227352 226102 227404 226108
rect 227168 225276 227220 225282
rect 227168 225218 227220 225224
rect 226800 224392 226852 224398
rect 226800 224334 226852 224340
rect 226800 222080 226852 222086
rect 226800 222022 226852 222028
rect 226076 219406 226288 219434
rect 226076 217410 226104 219406
rect 226812 217410 226840 222022
rect 227364 219910 227392 226102
rect 227352 219904 227404 219910
rect 227352 219846 227404 219852
rect 227548 217410 227576 229638
rect 227720 228880 227772 228886
rect 227720 228822 227772 228828
rect 227732 219842 227760 228822
rect 227916 228206 227944 231676
rect 227904 228200 227956 228206
rect 227904 228142 227956 228148
rect 228284 224466 228312 231676
rect 228272 224460 228324 224466
rect 228272 224402 228324 224408
rect 228652 224330 228680 231676
rect 229020 230042 229048 231676
rect 229008 230036 229060 230042
rect 229008 229978 229060 229984
rect 229388 227322 229416 231676
rect 229376 227316 229428 227322
rect 229376 227258 229428 227264
rect 229664 224534 229692 231676
rect 230032 227186 230060 231676
rect 230296 228812 230348 228818
rect 230296 228754 230348 228760
rect 230020 227180 230072 227186
rect 230020 227122 230072 227128
rect 229652 224528 229704 224534
rect 229652 224470 229704 224476
rect 228640 224324 228692 224330
rect 228640 224266 228692 224272
rect 228456 222148 228508 222154
rect 228456 222090 228508 222096
rect 227720 219836 227772 219842
rect 227720 219778 227772 219784
rect 228468 217410 228496 222090
rect 229376 220516 229428 220522
rect 229376 220458 229428 220464
rect 229388 217410 229416 220458
rect 230308 217410 230336 228754
rect 230400 228750 230428 231676
rect 230388 228744 230440 228750
rect 230388 228686 230440 228692
rect 230768 228138 230796 231676
rect 230756 228132 230808 228138
rect 230756 228074 230808 228080
rect 231136 224602 231164 231676
rect 231504 227254 231532 231676
rect 231872 230110 231900 231676
rect 231860 230104 231912 230110
rect 231860 230046 231912 230052
rect 232240 227458 232268 231676
rect 232332 231662 232530 231690
rect 232228 227452 232280 227458
rect 232228 227394 232280 227400
rect 231492 227248 231544 227254
rect 231492 227190 231544 227196
rect 232332 224670 232360 231662
rect 232884 227390 232912 231676
rect 233148 230036 233200 230042
rect 233148 229978 233200 229984
rect 232872 227384 232924 227390
rect 232872 227326 232924 227332
rect 232780 227248 232832 227254
rect 232780 227190 232832 227196
rect 232320 224664 232372 224670
rect 232320 224606 232372 224612
rect 231124 224596 231176 224602
rect 231124 224538 231176 224544
rect 232412 224324 232464 224330
rect 232412 224266 232464 224272
rect 231676 221400 231728 221406
rect 231676 221342 231728 221348
rect 231032 220584 231084 220590
rect 231032 220526 231084 220532
rect 231044 217410 231072 220526
rect 231688 217410 231716 221342
rect 232424 219774 232452 224266
rect 232688 220788 232740 220794
rect 232688 220730 232740 220736
rect 232412 219768 232464 219774
rect 232412 219710 232464 219716
rect 232700 217410 232728 220730
rect 232792 219706 232820 227190
rect 233160 220794 233188 229978
rect 233252 226234 233280 231676
rect 233528 231662 233634 231690
rect 233528 229094 233556 231662
rect 233436 229066 233556 229094
rect 233240 226228 233292 226234
rect 233240 226170 233292 226176
rect 233436 221338 233464 229066
rect 233516 228812 233568 228818
rect 233516 228754 233568 228760
rect 233424 221332 233476 221338
rect 233424 221274 233476 221280
rect 233148 220788 233200 220794
rect 233148 220730 233200 220736
rect 232780 219700 232832 219706
rect 232780 219642 232832 219648
rect 233528 217410 233556 228754
rect 233988 224738 234016 231676
rect 234356 227526 234384 231676
rect 234528 230104 234580 230110
rect 234528 230046 234580 230052
rect 234344 227520 234396 227526
rect 234344 227462 234396 227468
rect 233976 224732 234028 224738
rect 233976 224674 234028 224680
rect 234540 219434 234568 230046
rect 234724 228954 234752 231676
rect 234712 228948 234764 228954
rect 234712 228890 234764 228896
rect 235092 228070 235120 231676
rect 235080 228064 235132 228070
rect 235080 228006 235132 228012
rect 234712 227112 234764 227118
rect 234712 227054 234764 227060
rect 234620 224460 234672 224466
rect 234620 224402 234672 224408
rect 234632 219638 234660 224402
rect 234620 219632 234672 219638
rect 234620 219574 234672 219580
rect 234724 219570 234752 227054
rect 235368 224806 235396 231676
rect 235736 227594 235764 231676
rect 236104 230178 236132 231676
rect 236196 231662 236486 231690
rect 236092 230172 236144 230178
rect 236092 230114 236144 230120
rect 235724 227588 235776 227594
rect 235724 227530 235776 227536
rect 235356 224800 235408 224806
rect 235356 224742 235408 224748
rect 235264 221332 235316 221338
rect 235264 221274 235316 221280
rect 234712 219564 234764 219570
rect 234712 219506 234764 219512
rect 234448 219406 234568 219434
rect 234448 217410 234476 219406
rect 235276 217410 235304 221274
rect 236196 221270 236224 231662
rect 236840 224874 236868 231676
rect 237208 227662 237236 231676
rect 237196 227656 237248 227662
rect 237196 227598 237248 227604
rect 237380 227180 237432 227186
rect 237380 227122 237432 227128
rect 237012 227044 237064 227050
rect 237012 226986 237064 226992
rect 236828 224868 236880 224874
rect 236828 224810 236880 224816
rect 236184 221264 236236 221270
rect 236184 221206 236236 221212
rect 235908 220652 235960 220658
rect 235908 220594 235960 220600
rect 235920 217410 235948 220594
rect 237024 217410 237052 226986
rect 237392 219502 237420 227122
rect 237576 226166 237604 231676
rect 237944 228002 237972 231676
rect 237932 227996 237984 228002
rect 237932 227938 237984 227944
rect 237564 226160 237616 226166
rect 237564 226102 237616 226108
rect 238220 224942 238248 231676
rect 238588 227730 238616 231676
rect 238956 229294 238984 231676
rect 238944 229288 238996 229294
rect 238944 229230 238996 229236
rect 238576 227724 238628 227730
rect 238576 227666 238628 227672
rect 239324 226846 239352 231676
rect 239312 226840 239364 226846
rect 239312 226782 239364 226788
rect 238208 224936 238260 224942
rect 238208 224878 238260 224884
rect 239692 224194 239720 231676
rect 239784 231662 240074 231690
rect 239784 226982 239812 231662
rect 240048 230172 240100 230178
rect 240048 230114 240100 230120
rect 239772 226976 239824 226982
rect 239772 226918 239824 226924
rect 239956 224256 240008 224262
rect 239956 224198 240008 224204
rect 239680 224188 239732 224194
rect 239680 224130 239732 224136
rect 238576 221264 238628 221270
rect 238576 221206 238628 221212
rect 237748 220720 237800 220726
rect 237748 220662 237800 220668
rect 237380 219496 237432 219502
rect 237380 219438 237432 219444
rect 237760 217410 237788 220662
rect 238588 217410 238616 221206
rect 239404 220788 239456 220794
rect 239404 220730 239456 220736
rect 239416 217410 239444 220730
rect 239968 217410 239996 224198
rect 240060 220794 240088 230114
rect 240428 228886 240456 231676
rect 240520 231662 240810 231690
rect 240416 228880 240468 228886
rect 240416 228822 240468 228828
rect 240520 221202 240548 231662
rect 241072 224126 241100 231676
rect 241440 226914 241468 231676
rect 241808 230314 241836 231676
rect 241796 230308 241848 230314
rect 241796 230250 241848 230256
rect 242176 227934 242204 231676
rect 242164 227928 242216 227934
rect 242164 227870 242216 227876
rect 241428 226908 241480 226914
rect 241428 226850 241480 226856
rect 241060 224120 241112 224126
rect 241060 224062 241112 224068
rect 242544 224058 242572 231676
rect 242912 225214 242940 231676
rect 242900 225208 242952 225214
rect 242900 225150 242952 225156
rect 243280 224330 243308 231676
rect 243648 226710 243676 231676
rect 243636 226704 243688 226710
rect 243636 226646 243688 226652
rect 243268 224324 243320 224330
rect 243268 224266 243320 224272
rect 243636 224324 243688 224330
rect 243636 224266 243688 224272
rect 242532 224052 242584 224058
rect 242532 223994 242584 224000
rect 240508 221196 240560 221202
rect 240508 221138 240560 221144
rect 241980 221196 242032 221202
rect 241980 221138 242032 221144
rect 240048 220788 240100 220794
rect 240048 220730 240100 220736
rect 241152 220788 241204 220794
rect 241152 220730 241204 220736
rect 241164 217410 241192 220730
rect 241992 217410 242020 221138
rect 242808 219904 242860 219910
rect 242808 219846 242860 219852
rect 242820 217410 242848 219846
rect 243648 217410 243676 224266
rect 243924 223990 243952 231676
rect 244188 230308 244240 230314
rect 244188 230250 244240 230256
rect 243912 223984 243964 223990
rect 243912 223926 243964 223932
rect 244200 217410 244228 230250
rect 244292 226778 244320 231676
rect 244660 230382 244688 231676
rect 244648 230376 244700 230382
rect 244648 230318 244700 230324
rect 244924 229560 244976 229566
rect 244924 229502 244976 229508
rect 244280 226772 244332 226778
rect 244280 226714 244332 226720
rect 244936 221542 244964 229502
rect 245028 222766 245056 231676
rect 245396 223922 245424 231676
rect 245764 226642 245792 231676
rect 246132 230450 246160 231676
rect 246120 230444 246172 230450
rect 246120 230386 246172 230392
rect 245752 226636 245804 226642
rect 245752 226578 245804 226584
rect 245384 223916 245436 223922
rect 245384 223858 245436 223864
rect 245016 222760 245068 222766
rect 245016 222702 245068 222708
rect 246500 222698 246528 231676
rect 246776 223854 246804 231676
rect 246948 230376 247000 230382
rect 246948 230318 247000 230324
rect 246856 224392 246908 224398
rect 246856 224334 246908 224340
rect 246764 223848 246816 223854
rect 246764 223790 246816 223796
rect 246488 222692 246540 222698
rect 246488 222634 246540 222640
rect 244924 221536 244976 221542
rect 244924 221478 244976 221484
rect 245292 221536 245344 221542
rect 245292 221478 245344 221484
rect 245304 217410 245332 221478
rect 246120 219972 246172 219978
rect 246120 219914 246172 219920
rect 246132 217410 246160 219914
rect 246868 217410 246896 224334
rect 246960 219978 246988 230318
rect 247144 225146 247172 231676
rect 247512 227254 247540 231676
rect 247500 227248 247552 227254
rect 247500 227190 247552 227196
rect 247132 225140 247184 225146
rect 247132 225082 247184 225088
rect 247880 222562 247908 231676
rect 248248 223786 248276 231676
rect 248524 231662 248630 231690
rect 248328 229628 248380 229634
rect 248328 229570 248380 229576
rect 248236 223780 248288 223786
rect 248236 223722 248288 223728
rect 247868 222556 247920 222562
rect 247868 222498 247920 222504
rect 248340 220046 248368 229570
rect 248524 221134 248552 231662
rect 248984 229430 249012 231676
rect 248972 229424 249024 229430
rect 248972 229366 249024 229372
rect 249352 222494 249380 231676
rect 249444 231662 249642 231690
rect 249340 222488 249392 222494
rect 249340 222430 249392 222436
rect 248512 221128 248564 221134
rect 248512 221070 248564 221076
rect 248696 221128 248748 221134
rect 248696 221070 248748 221076
rect 247868 220040 247920 220046
rect 247868 219982 247920 219988
rect 248328 220040 248380 220046
rect 248328 219982 248380 219988
rect 246948 219972 247000 219978
rect 246948 219914 247000 219920
rect 247880 217410 247908 219982
rect 248708 217410 248736 221070
rect 249444 221066 249472 231662
rect 249996 222630 250024 231676
rect 250364 224466 250392 231676
rect 250352 224460 250404 224466
rect 250352 224402 250404 224408
rect 250352 223168 250404 223174
rect 250352 223110 250404 223116
rect 249984 222624 250036 222630
rect 249984 222566 250036 222572
rect 249432 221060 249484 221066
rect 249432 221002 249484 221008
rect 249524 219904 249576 219910
rect 249524 219846 249576 219852
rect 249536 217410 249564 219846
rect 250364 217410 250392 223110
rect 250732 222426 250760 231676
rect 250824 231662 251114 231690
rect 250720 222420 250772 222426
rect 250720 222362 250772 222368
rect 250824 220998 250852 231662
rect 251468 226574 251496 231676
rect 251456 226568 251508 226574
rect 251456 226510 251508 226516
rect 251836 226098 251864 231676
rect 252204 228478 252232 231676
rect 252296 231662 252494 231690
rect 252192 228472 252244 228478
rect 252192 228414 252244 228420
rect 252008 228336 252060 228342
rect 252008 228278 252060 228284
rect 251824 226092 251876 226098
rect 251824 226034 251876 226040
rect 250812 220992 250864 220998
rect 250812 220934 250864 220940
rect 250996 219768 251048 219774
rect 250996 219710 251048 219716
rect 251008 217410 251036 219710
rect 252020 217410 252048 228278
rect 252296 222358 252324 231662
rect 252848 228410 252876 231676
rect 252836 228404 252888 228410
rect 252836 228346 252888 228352
rect 253216 227118 253244 231676
rect 253204 227112 253256 227118
rect 253204 227054 253256 227060
rect 253584 223038 253612 231676
rect 253848 226092 253900 226098
rect 253848 226034 253900 226040
rect 253572 223032 253624 223038
rect 253572 222974 253624 222980
rect 252284 222352 252336 222358
rect 252284 222294 252336 222300
rect 252100 220108 252152 220114
rect 252100 220050 252152 220056
rect 252112 219706 252140 220050
rect 252928 219904 252980 219910
rect 252928 219846 252980 219852
rect 252100 219700 252152 219706
rect 252100 219642 252152 219648
rect 252940 217410 252968 219846
rect 253860 217410 253888 226034
rect 253952 222970 253980 231676
rect 254320 229566 254348 231676
rect 254688 229770 254716 231676
rect 254676 229764 254728 229770
rect 254676 229706 254728 229712
rect 254308 229560 254360 229566
rect 254308 229502 254360 229508
rect 255056 225622 255084 231676
rect 255228 229764 255280 229770
rect 255228 229706 255280 229712
rect 255136 227112 255188 227118
rect 255136 227054 255188 227060
rect 255044 225616 255096 225622
rect 255044 225558 255096 225564
rect 253940 222964 253992 222970
rect 253940 222906 253992 222912
rect 254584 220176 254636 220182
rect 254584 220118 254636 220124
rect 254596 217410 254624 220118
rect 255148 217410 255176 227054
rect 255240 220182 255268 229706
rect 255332 225690 255360 231676
rect 255320 225684 255372 225690
rect 255320 225626 255372 225632
rect 255700 222902 255728 231676
rect 255964 229220 256016 229226
rect 255964 229162 256016 229168
rect 255688 222896 255740 222902
rect 255688 222838 255740 222844
rect 255228 220176 255280 220182
rect 255228 220118 255280 220124
rect 255976 220114 256004 229162
rect 256068 227186 256096 231676
rect 256056 227180 256108 227186
rect 256056 227122 256108 227128
rect 256436 223106 256464 231676
rect 256804 225758 256832 231676
rect 257172 228546 257200 231676
rect 257540 229838 257568 231676
rect 257528 229832 257580 229838
rect 257528 229774 257580 229780
rect 257344 229152 257396 229158
rect 257344 229094 257396 229100
rect 257160 228540 257212 228546
rect 257160 228482 257212 228488
rect 256792 225752 256844 225758
rect 256792 225694 256844 225700
rect 257068 225616 257120 225622
rect 257068 225558 257120 225564
rect 256424 223100 256476 223106
rect 256424 223042 256476 223048
rect 255964 220108 256016 220114
rect 255964 220050 256016 220056
rect 256240 219836 256292 219842
rect 256240 219778 256292 219784
rect 256252 217410 256280 219778
rect 257080 217410 257108 225558
rect 257356 219706 257384 229094
rect 257908 225826 257936 231676
rect 258198 231662 258304 231690
rect 257896 225820 257948 225826
rect 257896 225762 257948 225768
rect 258276 221474 258304 231662
rect 258552 228614 258580 231676
rect 258920 229158 258948 231676
rect 259012 231662 259302 231690
rect 258908 229152 258960 229158
rect 258908 229094 258960 229100
rect 258540 228608 258592 228614
rect 258540 228550 258592 228556
rect 258816 227180 258868 227186
rect 258816 227122 258868 227128
rect 258264 221468 258316 221474
rect 258264 221410 258316 221416
rect 257896 220176 257948 220182
rect 257896 220118 257948 220124
rect 257344 219700 257396 219706
rect 257344 219642 257396 219648
rect 257908 217410 257936 220118
rect 258828 217410 258856 227122
rect 259012 225894 259040 231662
rect 259368 229832 259420 229838
rect 259368 229774 259420 229780
rect 259000 225888 259052 225894
rect 259000 225830 259052 225836
rect 259380 217410 259408 229774
rect 259656 221610 259684 231676
rect 260024 229226 260052 231676
rect 260392 229906 260420 231676
rect 260380 229900 260432 229906
rect 260380 229842 260432 229848
rect 260104 229628 260156 229634
rect 260104 229570 260156 229576
rect 260012 229220 260064 229226
rect 260012 229162 260064 229168
rect 259644 221604 259696 221610
rect 259644 221546 259696 221552
rect 260116 220318 260144 229570
rect 260760 228682 260788 231676
rect 260748 228676 260800 228682
rect 260748 228618 260800 228624
rect 260564 228404 260616 228410
rect 260564 228346 260616 228352
rect 260104 220312 260156 220318
rect 260104 220254 260156 220260
rect 260576 217410 260604 228346
rect 261036 221678 261064 231676
rect 261404 225962 261432 231676
rect 261496 231662 261786 231690
rect 261864 231662 262154 231690
rect 262324 231662 262522 231690
rect 262600 231662 262890 231690
rect 261392 225956 261444 225962
rect 261392 225898 261444 225904
rect 261024 221672 261076 221678
rect 261024 221614 261076 221620
rect 261496 220250 261524 231662
rect 261864 221746 261892 231662
rect 262128 222896 262180 222902
rect 262128 222838 262180 222844
rect 261852 221740 261904 221746
rect 261852 221682 261904 221688
rect 261484 220244 261536 220250
rect 261484 220186 261536 220192
rect 261300 219632 261352 219638
rect 261300 219574 261352 219580
rect 261312 217410 261340 219574
rect 262140 217410 262168 222838
rect 262324 221882 262352 231662
rect 262600 229634 262628 231662
rect 262864 230444 262916 230450
rect 262864 230386 262916 230392
rect 262876 230110 262904 230386
rect 263244 230246 263272 231676
rect 263626 231662 263732 231690
rect 263232 230240 263284 230246
rect 263232 230182 263284 230188
rect 262864 230104 262916 230110
rect 262864 230046 262916 230052
rect 263508 229900 263560 229906
rect 263508 229842 263560 229848
rect 262588 229628 262640 229634
rect 262588 229570 262640 229576
rect 263416 225684 263468 225690
rect 263416 225626 263468 225632
rect 262312 221876 262364 221882
rect 262312 221818 262364 221824
rect 262588 220516 262640 220522
rect 262588 220458 262640 220464
rect 262956 220516 263008 220522
rect 262956 220458 263008 220464
rect 262600 220250 262628 220458
rect 262588 220244 262640 220250
rect 262588 220186 262640 220192
rect 262968 217410 262996 220458
rect 190288 217382 190348 217410
rect 191176 217382 191604 217410
rect 192004 217382 192340 217410
rect 192832 217382 192984 217410
rect 193752 217382 194088 217410
rect 194580 217382 194916 217410
rect 195408 217382 195744 217410
rect 196236 217382 196572 217410
rect 197064 217382 197308 217410
rect 197892 217382 198228 217410
rect 198720 217382 199056 217410
rect 199640 217382 199976 217410
rect 200468 217382 200804 217410
rect 201296 217382 201448 217410
rect 202124 217382 202460 217410
rect 202952 217382 203288 217410
rect 203780 217382 204116 217410
rect 204608 217382 204944 217410
rect 205528 217382 205588 217410
rect 206356 217382 206876 217410
rect 207184 217382 207520 217410
rect 208012 217382 208348 217410
rect 208840 217382 209176 217410
rect 209668 217382 209728 217410
rect 210496 217382 210832 217410
rect 211416 217382 211752 217410
rect 212244 217382 212488 217410
rect 213072 217382 213408 217410
rect 213900 217382 214236 217410
rect 214728 217382 215156 217410
rect 215556 217382 215892 217410
rect 216384 217382 216628 217410
rect 217304 217382 217640 217410
rect 218132 217382 218468 217410
rect 218960 217382 219296 217410
rect 219788 217382 220124 217410
rect 220616 217382 220676 217410
rect 221444 217382 221780 217410
rect 222272 217382 222608 217410
rect 223192 217382 223528 217410
rect 224020 217382 224356 217410
rect 224848 217382 224908 217410
rect 225676 217382 226104 217410
rect 226504 217382 226840 217410
rect 227332 217382 227576 217410
rect 228160 217382 228496 217410
rect 229080 217382 229416 217410
rect 229908 217382 230336 217410
rect 230736 217382 231072 217410
rect 231564 217382 231716 217410
rect 232392 217382 232728 217410
rect 233220 217382 233556 217410
rect 234048 217382 234476 217410
rect 234968 217382 235304 217410
rect 235796 217382 235948 217410
rect 236624 217382 237052 217410
rect 237452 217382 237788 217410
rect 238280 217382 238616 217410
rect 239108 217382 239444 217410
rect 239936 217382 239996 217410
rect 240856 217382 241192 217410
rect 241684 217382 242020 217410
rect 242512 217382 242848 217410
rect 243340 217382 243676 217410
rect 244168 217382 244228 217410
rect 244996 217382 245332 217410
rect 245824 217382 246160 217410
rect 246744 217382 246896 217410
rect 247572 217382 247908 217410
rect 248400 217382 248736 217410
rect 249228 217382 249564 217410
rect 250056 217382 250392 217410
rect 250884 217382 251036 217410
rect 251712 217382 252048 217410
rect 252632 217382 252968 217410
rect 253460 217382 253888 217410
rect 254288 217382 254624 217410
rect 255116 217382 255176 217410
rect 255944 217382 256280 217410
rect 256772 217382 257108 217410
rect 257600 217382 257936 217410
rect 258520 217382 258856 217410
rect 259348 217382 259408 217410
rect 260176 217382 260604 217410
rect 261004 217382 261340 217410
rect 261832 217382 262168 217410
rect 262660 217382 262996 217410
rect 263428 217410 263456 225626
rect 263520 220522 263548 229842
rect 263704 221814 263732 231662
rect 263796 231662 263902 231690
rect 263796 221950 263824 231662
rect 264256 226030 264284 231676
rect 264348 231662 264638 231690
rect 265006 231662 265112 231690
rect 264244 226024 264296 226030
rect 264244 225966 264296 225972
rect 263784 221944 263836 221950
rect 263784 221886 263836 221892
rect 263692 221808 263744 221814
rect 263692 221750 263744 221756
rect 263508 220516 263560 220522
rect 263508 220458 263560 220464
rect 264348 220454 264376 231662
rect 265084 222018 265112 231662
rect 265176 231662 265374 231690
rect 265452 231662 265742 231690
rect 265176 222086 265204 231662
rect 265164 222080 265216 222086
rect 265164 222022 265216 222028
rect 265072 222012 265124 222018
rect 265072 221954 265124 221960
rect 264336 220448 264388 220454
rect 264336 220390 264388 220396
rect 265452 220386 265480 231662
rect 266096 229974 266124 231676
rect 266084 229968 266136 229974
rect 266084 229910 266136 229916
rect 265532 222964 265584 222970
rect 265532 222906 265584 222912
rect 265440 220380 265492 220386
rect 265440 220322 265492 220328
rect 264704 220312 264756 220318
rect 264704 220254 264756 220260
rect 264716 217410 264744 220254
rect 265544 217410 265572 222906
rect 266464 222154 266492 231676
rect 266740 228750 266768 231676
rect 267108 229702 267136 231676
rect 267200 231662 267490 231690
rect 267096 229696 267148 229702
rect 267096 229638 267148 229644
rect 266728 228744 266780 228750
rect 266728 228686 266780 228692
rect 266452 222148 266504 222154
rect 266452 222090 266504 222096
rect 267200 220250 267228 231662
rect 267844 221406 267872 231676
rect 268212 228818 268240 231676
rect 268304 231662 268594 231690
rect 268200 228812 268252 228818
rect 268200 228754 268252 228760
rect 267832 221400 267884 221406
rect 267832 221342 267884 221348
rect 268304 220590 268332 231662
rect 268948 230110 268976 231676
rect 269224 231662 269330 231690
rect 268936 230104 268988 230110
rect 268936 230046 268988 230052
rect 268384 229696 268436 229702
rect 268384 229638 268436 229644
rect 268292 220584 268344 220590
rect 268292 220526 268344 220532
rect 267188 220244 267240 220250
rect 267188 220186 267240 220192
rect 266176 220108 266228 220114
rect 266176 220050 266228 220056
rect 266188 217410 266216 220050
rect 268016 219700 268068 219706
rect 268016 219642 268068 219648
rect 267188 219496 267240 219502
rect 267188 219438 267240 219444
rect 267200 217410 267228 219438
rect 268028 217410 268056 219642
rect 268396 219502 268424 229638
rect 268936 224460 268988 224466
rect 268936 224402 268988 224408
rect 268384 219496 268436 219502
rect 268384 219438 268436 219444
rect 268948 217410 268976 224402
rect 269224 221338 269252 231662
rect 269592 227050 269620 231676
rect 269960 230450 269988 231676
rect 270052 231662 270342 231690
rect 269948 230444 270000 230450
rect 269948 230386 270000 230392
rect 269580 227044 269632 227050
rect 269580 226986 269632 226992
rect 269212 221332 269264 221338
rect 269212 221274 269264 221280
rect 269672 220788 269724 220794
rect 269672 220730 269724 220736
rect 269684 217410 269712 220730
rect 270052 220658 270080 231662
rect 270316 230036 270368 230042
rect 270316 229978 270368 229984
rect 270132 229628 270184 229634
rect 270132 229570 270184 229576
rect 270144 220726 270172 229570
rect 270132 220720 270184 220726
rect 270132 220662 270184 220668
rect 270040 220652 270092 220658
rect 270040 220594 270092 220600
rect 270328 217410 270356 229978
rect 270408 229968 270460 229974
rect 270408 229910 270460 229916
rect 270420 220794 270448 229910
rect 270696 221270 270724 231676
rect 271064 224262 271092 231676
rect 271144 230376 271196 230382
rect 271144 230318 271196 230324
rect 271052 224256 271104 224262
rect 271052 224198 271104 224204
rect 270684 221264 270736 221270
rect 270684 221206 270736 221212
rect 271156 220794 271184 230318
rect 271328 230104 271380 230110
rect 271328 230046 271380 230052
rect 271236 229288 271288 229294
rect 271236 229230 271288 229236
rect 270408 220788 270460 220794
rect 270408 220730 270460 220736
rect 271144 220788 271196 220794
rect 271144 220730 271196 220736
rect 271248 220182 271276 229230
rect 271236 220176 271288 220182
rect 271236 220118 271288 220124
rect 271340 219774 271368 230046
rect 271432 229634 271460 231676
rect 271800 230178 271828 231676
rect 271984 231662 272182 231690
rect 272260 231662 272458 231690
rect 271788 230172 271840 230178
rect 271788 230114 271840 230120
rect 271420 229628 271472 229634
rect 271420 229570 271472 229576
rect 271984 221202 272012 231662
rect 272260 224330 272288 231662
rect 272812 230382 272840 231676
rect 272904 231662 273194 231690
rect 273456 231662 273562 231690
rect 273640 231662 273930 231690
rect 272800 230376 272852 230382
rect 272800 230318 272852 230324
rect 272248 224324 272300 224330
rect 272248 224266 272300 224272
rect 272248 221468 272300 221474
rect 272248 221410 272300 221416
rect 271972 221196 272024 221202
rect 271972 221138 272024 221144
rect 271420 220652 271472 220658
rect 271420 220594 271472 220600
rect 271328 219768 271380 219774
rect 271328 219710 271380 219716
rect 271432 217410 271460 220594
rect 272260 217410 272288 221410
rect 272904 220046 272932 231662
rect 272984 229560 273036 229566
rect 272984 229502 273036 229508
rect 272892 220040 272944 220046
rect 272892 219982 272944 219988
rect 272996 219638 273024 229502
rect 273456 221542 273484 231662
rect 273640 224398 273668 231662
rect 274284 230314 274312 231676
rect 274652 230450 274680 231676
rect 274836 231662 275034 231690
rect 275112 231662 275310 231690
rect 274640 230444 274692 230450
rect 274640 230386 274692 230392
rect 274272 230308 274324 230314
rect 274272 230250 274324 230256
rect 274548 230308 274600 230314
rect 274548 230250 274600 230256
rect 273904 229424 273956 229430
rect 273904 229366 273956 229372
rect 273916 229094 273944 229366
rect 273824 229066 273944 229094
rect 273628 224392 273680 224398
rect 273628 224334 273680 224340
rect 273444 221536 273496 221542
rect 273444 221478 273496 221484
rect 273076 220584 273128 220590
rect 273076 220526 273128 220532
rect 272984 219632 273036 219638
rect 272984 219574 273036 219580
rect 273088 217410 273116 220526
rect 273824 220318 273852 229066
rect 274560 220794 274588 230250
rect 274836 221134 274864 231662
rect 275112 223174 275140 231662
rect 275376 230172 275428 230178
rect 275376 230114 275428 230120
rect 275284 229492 275336 229498
rect 275284 229434 275336 229440
rect 275100 223168 275152 223174
rect 275100 223110 275152 223116
rect 274824 221128 274876 221134
rect 274824 221070 274876 221076
rect 273904 220788 273956 220794
rect 273904 220730 273956 220736
rect 274548 220788 274600 220794
rect 274548 220730 274600 220736
rect 273812 220312 273864 220318
rect 273812 220254 273864 220260
rect 273916 217410 273944 220730
rect 274456 220720 274508 220726
rect 274456 220662 274508 220668
rect 274468 217410 274496 220662
rect 275296 219706 275324 229434
rect 275388 220658 275416 230114
rect 275664 229634 275692 231676
rect 276046 231662 276244 231690
rect 275652 229628 275704 229634
rect 275652 229570 275704 229576
rect 275560 221536 275612 221542
rect 275560 221478 275612 221484
rect 275376 220652 275428 220658
rect 275376 220594 275428 220600
rect 275284 219700 275336 219706
rect 275284 219642 275336 219648
rect 275572 217410 275600 221478
rect 276216 219978 276244 231662
rect 276400 228478 276428 231676
rect 276492 231662 276782 231690
rect 276388 228472 276440 228478
rect 276388 228414 276440 228420
rect 276492 226098 276520 231662
rect 276664 230444 276716 230450
rect 276664 230386 276716 230392
rect 276480 226092 276532 226098
rect 276480 226034 276532 226040
rect 276676 220590 276704 230386
rect 276756 230240 276808 230246
rect 276756 230182 276808 230188
rect 276768 220726 276796 230182
rect 277136 230110 277164 231676
rect 277518 231662 277624 231690
rect 277124 230104 277176 230110
rect 277124 230046 277176 230052
rect 277308 230036 277360 230042
rect 277308 229978 277360 229984
rect 277320 229786 277348 229978
rect 277228 229758 277348 229786
rect 277228 229702 277256 229758
rect 277216 229696 277268 229702
rect 277216 229638 277268 229644
rect 277308 229696 277360 229702
rect 277308 229638 277360 229644
rect 277492 229696 277544 229702
rect 277492 229638 277544 229644
rect 276756 220720 276808 220726
rect 276756 220662 276808 220668
rect 276664 220584 276716 220590
rect 276664 220526 276716 220532
rect 276204 219972 276256 219978
rect 276204 219914 276256 219920
rect 276480 219496 276532 219502
rect 276480 219438 276532 219444
rect 276492 217410 276520 219438
rect 277320 217410 277348 229638
rect 277504 229362 277532 229638
rect 277492 229356 277544 229362
rect 277492 229298 277544 229304
rect 277596 219910 277624 231662
rect 277768 230444 277820 230450
rect 277768 230386 277820 230392
rect 277780 230178 277808 230386
rect 277676 230172 277728 230178
rect 277676 230114 277728 230120
rect 277768 230172 277820 230178
rect 277768 230114 277820 230120
rect 277688 229702 277716 230114
rect 277676 229696 277728 229702
rect 277676 229638 277728 229644
rect 277872 227118 277900 231676
rect 278044 230308 278096 230314
rect 278044 230250 278096 230256
rect 277860 227112 277912 227118
rect 277860 227054 277912 227060
rect 277584 219904 277636 219910
rect 277584 219846 277636 219852
rect 278056 219502 278084 230250
rect 278148 225622 278176 231676
rect 278516 229770 278544 231676
rect 278898 231662 279004 231690
rect 278504 229764 278556 229770
rect 278504 229706 278556 229712
rect 278688 229764 278740 229770
rect 278688 229706 278740 229712
rect 278136 225616 278188 225622
rect 278136 225558 278188 225564
rect 278700 220794 278728 229706
rect 278136 220788 278188 220794
rect 278136 220730 278188 220736
rect 278688 220788 278740 220794
rect 278688 220730 278740 220736
rect 278044 219496 278096 219502
rect 278044 219438 278096 219444
rect 278148 217410 278176 220730
rect 278596 220108 278648 220114
rect 278596 220050 278648 220056
rect 263428 217382 263488 217410
rect 264408 217382 264744 217410
rect 265236 217382 265572 217410
rect 266064 217382 266216 217410
rect 266892 217382 267228 217410
rect 267720 217382 268056 217410
rect 268548 217382 268976 217410
rect 269376 217382 269712 217410
rect 270296 217382 270356 217410
rect 271124 217382 271460 217410
rect 271952 217382 272288 217410
rect 272780 217382 273116 217410
rect 273608 217382 273944 217410
rect 274436 217382 274496 217410
rect 275264 217382 275600 217410
rect 276184 217382 276520 217410
rect 277012 217382 277348 217410
rect 277840 217382 278176 217410
rect 278608 217410 278636 220050
rect 278976 219842 279004 231662
rect 279252 227186 279280 231676
rect 279424 230376 279476 230382
rect 279424 230318 279476 230324
rect 279240 227180 279292 227186
rect 279240 227122 279292 227128
rect 279436 220182 279464 230318
rect 279620 228410 279648 231676
rect 279988 229294 280016 231676
rect 280356 229838 280384 231676
rect 280344 229832 280396 229838
rect 280344 229774 280396 229780
rect 280068 229628 280120 229634
rect 280068 229570 280120 229576
rect 279976 229288 280028 229294
rect 279976 229230 280028 229236
rect 279608 228404 279660 228410
rect 279608 228346 279660 228352
rect 279424 220176 279476 220182
rect 279424 220118 279476 220124
rect 278964 219836 279016 219842
rect 278964 219778 279016 219784
rect 280080 219434 280108 229570
rect 280724 222902 280752 231676
rect 281000 225690 281028 231676
rect 281092 231662 281382 231690
rect 281092 229566 281120 231662
rect 281736 229906 281764 231676
rect 281724 229900 281776 229906
rect 281724 229842 281776 229848
rect 281356 229832 281408 229838
rect 281356 229774 281408 229780
rect 281080 229560 281132 229566
rect 281080 229502 281132 229508
rect 280988 225684 281040 225690
rect 280988 225626 281040 225632
rect 280712 222896 280764 222902
rect 280712 222838 280764 222844
rect 280620 220176 280672 220182
rect 280620 220118 280672 220124
rect 279896 219406 280108 219434
rect 279896 217410 279924 219406
rect 280632 217410 280660 220118
rect 281368 217410 281396 229774
rect 281448 229288 281500 229294
rect 281448 229230 281500 229236
rect 281460 220182 281488 229230
rect 282104 222970 282132 231676
rect 282472 230042 282500 231676
rect 282460 230036 282512 230042
rect 282460 229978 282512 229984
rect 282840 229430 282868 231676
rect 283208 230382 283236 231676
rect 283196 230376 283248 230382
rect 283196 230318 283248 230324
rect 282828 229424 282880 229430
rect 282828 229366 282880 229372
rect 282828 229220 282880 229226
rect 282828 229162 282880 229168
rect 282092 222964 282144 222970
rect 282092 222906 282144 222912
rect 282840 220794 282868 229162
rect 283576 224466 283604 231676
rect 283852 230110 283880 231676
rect 283944 231662 284234 231690
rect 283840 230104 283892 230110
rect 283840 230046 283892 230052
rect 283944 229498 283972 231662
rect 284208 230036 284260 230042
rect 284208 229978 284260 229984
rect 283932 229492 283984 229498
rect 283932 229434 283984 229440
rect 284116 229152 284168 229158
rect 284116 229094 284168 229100
rect 283564 224460 283616 224466
rect 283564 224402 283616 224408
rect 282368 220788 282420 220794
rect 282368 220730 282420 220736
rect 282828 220788 282880 220794
rect 282828 220730 282880 220736
rect 281448 220176 281500 220182
rect 281448 220118 281500 220124
rect 282380 217410 282408 220730
rect 283196 220312 283248 220318
rect 283196 220254 283248 220260
rect 283208 217410 283236 220254
rect 284128 217410 284156 229094
rect 284220 220318 284248 229978
rect 284588 229974 284616 231676
rect 284680 231662 284970 231690
rect 284576 229968 284628 229974
rect 284576 229910 284628 229916
rect 284680 221474 284708 231662
rect 285324 230450 285352 231676
rect 285312 230444 285364 230450
rect 285312 230386 285364 230392
rect 285588 230308 285640 230314
rect 285588 230250 285640 230256
rect 285496 229968 285548 229974
rect 285496 229910 285548 229916
rect 284668 221468 284720 221474
rect 284668 221410 284720 221416
rect 284208 220312 284260 220318
rect 284208 220254 284260 220260
rect 285508 220114 285536 229910
rect 284852 220108 284904 220114
rect 284852 220050 284904 220056
rect 285496 220108 285548 220114
rect 285496 220050 285548 220056
rect 284864 217410 284892 220050
rect 285600 217410 285628 230250
rect 285692 229702 285720 231676
rect 286060 230178 286088 231676
rect 286152 231662 286442 231690
rect 286048 230172 286100 230178
rect 286048 230114 286100 230120
rect 285680 229696 285732 229702
rect 285680 229638 285732 229644
rect 286152 221542 286180 231662
rect 286704 229362 286732 231676
rect 286968 230444 287020 230450
rect 286968 230386 287020 230392
rect 286692 229356 286744 229362
rect 286692 229298 286744 229304
rect 286140 221536 286192 221542
rect 286140 221478 286192 221484
rect 286980 220794 287008 230386
rect 287072 230246 287100 231676
rect 287440 230382 287468 231676
rect 287532 231662 287822 231690
rect 287428 230376 287480 230382
rect 287428 230318 287480 230324
rect 287060 230240 287112 230246
rect 287060 230182 287112 230188
rect 286508 220788 286560 220794
rect 286508 220730 286560 220736
rect 286968 220788 287020 220794
rect 286968 220730 287020 220736
rect 287336 220788 287388 220794
rect 287336 220730 287388 220736
rect 286520 217410 286548 220730
rect 287348 217410 287376 220730
rect 287532 220182 287560 231662
rect 288176 229294 288204 231676
rect 288348 230444 288400 230450
rect 288348 230386 288400 230392
rect 288164 229288 288216 229294
rect 288164 229230 288216 229236
rect 287520 220176 287572 220182
rect 287520 220118 287572 220124
rect 288360 217410 288388 230386
rect 288544 229770 288572 231676
rect 288532 229764 288584 229770
rect 288532 229706 288584 229712
rect 288912 229634 288940 231676
rect 288900 229628 288952 229634
rect 288900 229570 288952 229576
rect 289280 229226 289308 231676
rect 289268 229220 289320 229226
rect 289268 229162 289320 229168
rect 289556 229158 289584 231676
rect 289924 229838 289952 231676
rect 290292 230042 290320 231676
rect 290660 230314 290688 231676
rect 290752 231662 291042 231690
rect 290648 230308 290700 230314
rect 290648 230250 290700 230256
rect 290280 230036 290332 230042
rect 290280 229978 290332 229984
rect 289912 229832 289964 229838
rect 289912 229774 289964 229780
rect 289544 229152 289596 229158
rect 289544 229094 289596 229100
rect 290752 229094 290780 231662
rect 291396 229974 291424 231676
rect 291764 230382 291792 231676
rect 291856 231662 292146 231690
rect 292224 231662 292422 231690
rect 291752 230376 291804 230382
rect 291752 230318 291804 230324
rect 291384 229968 291436 229974
rect 291384 229910 291436 229916
rect 290660 229066 290780 229094
rect 290660 220794 290688 229066
rect 290648 220788 290700 220794
rect 290648 220730 290700 220736
rect 290740 220788 290792 220794
rect 290740 220730 290792 220736
rect 289084 220720 289136 220726
rect 289084 220662 289136 220668
rect 289096 217410 289124 220662
rect 289636 220040 289688 220046
rect 289636 219982 289688 219988
rect 289648 217410 289676 219982
rect 290752 217410 290780 220730
rect 291856 220726 291884 231662
rect 292224 220794 292252 231662
rect 292776 230450 292804 231676
rect 292868 231662 293158 231690
rect 293236 231662 293526 231690
rect 292764 230444 292816 230450
rect 292764 230386 292816 230392
rect 292580 230376 292632 230382
rect 292580 230318 292632 230324
rect 292592 224262 292620 230318
rect 292580 224256 292632 224262
rect 292580 224198 292632 224204
rect 292212 220788 292264 220794
rect 292212 220730 292264 220736
rect 292488 220788 292540 220794
rect 292488 220730 292540 220736
rect 291844 220720 291896 220726
rect 291844 220662 291896 220668
rect 291568 220312 291620 220318
rect 291568 220254 291620 220260
rect 291580 217410 291608 220254
rect 292500 217410 292528 220730
rect 292868 220046 292896 231662
rect 293236 220794 293264 231662
rect 293880 230382 293908 231676
rect 293972 231662 294262 231690
rect 294340 231662 294630 231690
rect 294998 231662 295196 231690
rect 293868 230376 293920 230382
rect 293868 230318 293920 230324
rect 293500 224256 293552 224262
rect 293500 224198 293552 224204
rect 293224 220788 293276 220794
rect 293224 220730 293276 220736
rect 293224 220584 293276 220590
rect 293224 220526 293276 220532
rect 292856 220040 292908 220046
rect 292856 219982 292908 219988
rect 293236 217410 293264 220526
rect 278608 217382 278668 217410
rect 279496 217382 279924 217410
rect 280324 217382 280660 217410
rect 281152 217382 281396 217410
rect 282072 217382 282408 217410
rect 282900 217382 283236 217410
rect 283728 217382 284156 217410
rect 284556 217382 284892 217410
rect 285384 217382 285628 217410
rect 286212 217382 286548 217410
rect 287040 217382 287376 217410
rect 287960 217382 288388 217410
rect 288788 217382 289124 217410
rect 289616 217382 289676 217410
rect 290444 217382 290780 217410
rect 291272 217382 291608 217410
rect 292100 217382 292528 217410
rect 292928 217382 293264 217410
rect 293512 217410 293540 224198
rect 293972 220318 294000 231662
rect 294340 220590 294368 231662
rect 295168 229094 295196 231662
rect 295260 229362 295288 231676
rect 295536 231662 295642 231690
rect 295720 231662 296010 231690
rect 295248 229356 295300 229362
rect 295248 229298 295300 229304
rect 295168 229066 295380 229094
rect 294972 220788 295024 220794
rect 294972 220730 295024 220736
rect 294328 220584 294380 220590
rect 294328 220526 294380 220532
rect 293960 220312 294012 220318
rect 293960 220254 294012 220260
rect 294984 217410 295012 220730
rect 293512 217382 293848 217410
rect 294676 217382 295012 217410
rect 295352 217410 295380 229066
rect 295536 220794 295564 231662
rect 295720 229094 295748 231662
rect 296364 229226 296392 231676
rect 296732 229906 296760 231676
rect 296824 231662 297114 231690
rect 296720 229900 296772 229906
rect 296720 229842 296772 229848
rect 296352 229220 296404 229226
rect 296352 229162 296404 229168
rect 296824 229094 296852 231662
rect 297468 230450 297496 231676
rect 297850 231662 298048 231690
rect 297456 230444 297508 230450
rect 297456 230386 297508 230392
rect 296904 229356 296956 229362
rect 296904 229298 296956 229304
rect 295720 229066 295932 229094
rect 295524 220788 295576 220794
rect 295524 220730 295576 220736
rect 295904 217410 295932 229066
rect 296732 229066 296852 229094
rect 296732 217870 296760 229066
rect 296916 219434 296944 229298
rect 298020 220794 298048 231662
rect 298112 230382 298140 231676
rect 298100 230376 298152 230382
rect 298100 230318 298152 230324
rect 298480 229430 298508 231676
rect 298848 230246 298876 231676
rect 299230 231662 299428 231690
rect 299296 230376 299348 230382
rect 299296 230318 299348 230324
rect 298836 230240 298888 230246
rect 298836 230182 298888 230188
rect 298468 229424 298520 229430
rect 298468 229366 298520 229372
rect 298468 229220 298520 229226
rect 298468 229162 298520 229168
rect 298008 220788 298060 220794
rect 298008 220730 298060 220736
rect 296824 219406 296944 219434
rect 296720 217864 296772 217870
rect 296720 217806 296772 217812
rect 296824 217410 296852 219406
rect 297640 217864 297692 217870
rect 297640 217806 297692 217812
rect 297652 217410 297680 217806
rect 298480 217410 298508 229162
rect 299308 220590 299336 230318
rect 299296 220584 299348 220590
rect 299296 220526 299348 220532
rect 299400 220454 299428 231662
rect 299584 230382 299612 231676
rect 299966 231662 300256 231690
rect 300334 231662 300624 231690
rect 300228 230450 300256 231662
rect 299940 230444 299992 230450
rect 299940 230386 299992 230392
rect 300216 230444 300268 230450
rect 300216 230386 300268 230392
rect 299572 230376 299624 230382
rect 299572 230318 299624 230324
rect 299572 229900 299624 229906
rect 299572 229842 299624 229848
rect 299388 220448 299440 220454
rect 299388 220390 299440 220396
rect 299584 217870 299612 229842
rect 299572 217864 299624 217870
rect 299572 217806 299624 217812
rect 299952 217410 299980 230386
rect 300492 230376 300544 230382
rect 300492 230318 300544 230324
rect 300504 219638 300532 230318
rect 300492 219632 300544 219638
rect 300492 219574 300544 219580
rect 300596 219502 300624 231662
rect 300688 229566 300716 231676
rect 300978 231662 301268 231690
rect 301346 231662 301636 231690
rect 301714 231662 302004 231690
rect 300676 229560 300728 229566
rect 300676 229502 300728 229508
rect 301136 229424 301188 229430
rect 301136 229366 301188 229372
rect 300584 219496 300636 219502
rect 300584 219438 300636 219444
rect 301148 219434 301176 229366
rect 301240 221474 301268 231662
rect 301228 221468 301280 221474
rect 301228 221410 301280 221416
rect 301608 219570 301636 231662
rect 301976 220114 302004 231662
rect 302068 229838 302096 231676
rect 302450 231662 302740 231690
rect 302818 231662 303108 231690
rect 303186 231662 303476 231690
rect 302424 230240 302476 230246
rect 302424 230182 302476 230188
rect 302056 229832 302108 229838
rect 302056 229774 302108 229780
rect 302436 229094 302464 230182
rect 302436 229066 302648 229094
rect 302240 220788 302292 220794
rect 302240 220730 302292 220736
rect 301964 220108 302016 220114
rect 301964 220050 302016 220056
rect 301596 219564 301648 219570
rect 301596 219506 301648 219512
rect 301148 219406 301268 219434
rect 300216 217864 300268 217870
rect 300216 217806 300268 217812
rect 295352 217382 295504 217410
rect 295904 217382 296332 217410
rect 296824 217382 297160 217410
rect 297652 217382 297988 217410
rect 298480 217382 298816 217410
rect 299736 217382 299980 217410
rect 300228 217410 300256 217806
rect 301240 217410 301268 219406
rect 302252 217410 302280 220730
rect 300228 217382 300564 217410
rect 301240 217382 301392 217410
rect 302220 217382 302280 217410
rect 302620 217410 302648 229066
rect 302712 225690 302740 231662
rect 302700 225684 302752 225690
rect 302700 225626 302752 225632
rect 303080 220726 303108 231662
rect 303068 220720 303120 220726
rect 303068 220662 303120 220668
rect 303448 220658 303476 231662
rect 303540 229974 303568 231676
rect 303528 229968 303580 229974
rect 303528 229910 303580 229916
rect 303816 225758 303844 231676
rect 303988 230444 304040 230450
rect 303988 230386 304040 230392
rect 304000 229094 304028 230386
rect 304184 230382 304212 231676
rect 304566 231662 304856 231690
rect 304172 230376 304224 230382
rect 304172 230318 304224 230324
rect 304000 229066 304304 229094
rect 303804 225752 303856 225758
rect 303804 225694 303856 225700
rect 303436 220652 303488 220658
rect 303436 220594 303488 220600
rect 303620 220584 303672 220590
rect 303620 220526 303672 220532
rect 303632 217410 303660 220526
rect 304276 217410 304304 229066
rect 304828 220522 304856 231662
rect 304920 230466 304948 231676
rect 304920 230438 305040 230466
rect 304908 230376 304960 230382
rect 304908 230318 304960 230324
rect 304816 220516 304868 220522
rect 304816 220458 304868 220464
rect 304920 220250 304948 230318
rect 305012 229906 305040 230438
rect 305000 229900 305052 229906
rect 305000 229842 305052 229848
rect 305288 227050 305316 231676
rect 305656 230382 305684 231676
rect 306038 231662 306144 231690
rect 305644 230376 305696 230382
rect 305644 230318 305696 230324
rect 305552 229560 305604 229566
rect 305552 229502 305604 229508
rect 305276 227044 305328 227050
rect 305276 226986 305328 226992
rect 305564 220862 305592 229502
rect 305552 220856 305604 220862
rect 305552 220798 305604 220804
rect 306116 220454 306144 231662
rect 306196 230376 306248 230382
rect 306196 230318 306248 230324
rect 306208 220590 306236 230318
rect 306392 222970 306420 231676
rect 306668 228546 306696 231676
rect 307036 230382 307064 231676
rect 307024 230376 307076 230382
rect 307024 230318 307076 230324
rect 306656 228540 306708 228546
rect 306656 228482 306708 228488
rect 306380 222964 306432 222970
rect 306380 222906 306432 222912
rect 306196 220584 306248 220590
rect 306196 220526 306248 220532
rect 305276 220448 305328 220454
rect 305276 220390 305328 220396
rect 306104 220448 306156 220454
rect 306104 220390 306156 220396
rect 304908 220244 304960 220250
rect 304908 220186 304960 220192
rect 305288 217410 305316 220390
rect 307404 220318 307432 231676
rect 307576 230376 307628 230382
rect 307576 230318 307628 230324
rect 307588 220386 307616 230318
rect 307772 224398 307800 231676
rect 308140 228410 308168 231676
rect 308128 228404 308180 228410
rect 308128 228346 308180 228352
rect 307760 224392 307812 224398
rect 307760 224334 307812 224340
rect 308508 222902 308536 231676
rect 308784 231662 308890 231690
rect 308496 222896 308548 222902
rect 308496 222838 308548 222844
rect 308588 220856 308640 220862
rect 308588 220798 308640 220804
rect 307576 220380 307628 220386
rect 307576 220322 307628 220328
rect 307392 220312 307444 220318
rect 307392 220254 307444 220260
rect 306932 219632 306984 219638
rect 306932 219574 306984 219580
rect 306380 219496 306432 219502
rect 306380 219438 306432 219444
rect 306392 217410 306420 219438
rect 306944 217410 306972 219574
rect 307760 219564 307812 219570
rect 307760 219506 307812 219512
rect 307772 217410 307800 219506
rect 308600 217410 308628 220798
rect 308784 220182 308812 231662
rect 309244 224330 309272 231676
rect 309520 227458 309548 231676
rect 309888 228478 309916 231676
rect 309876 228472 309928 228478
rect 309876 228414 309928 228420
rect 309508 227452 309560 227458
rect 309508 227394 309560 227400
rect 309232 224324 309284 224330
rect 309232 224266 309284 224272
rect 308772 220176 308824 220182
rect 308772 220118 308824 220124
rect 310256 220114 310284 231676
rect 310624 230314 310652 231676
rect 310612 230308 310664 230314
rect 310612 230250 310664 230256
rect 310992 225622 311020 231676
rect 311164 229832 311216 229838
rect 311164 229774 311216 229780
rect 310980 225616 311032 225622
rect 310980 225558 311032 225564
rect 311176 222154 311204 229774
rect 311360 224262 311388 231676
rect 311728 230450 311756 231676
rect 311716 230444 311768 230450
rect 311716 230386 311768 230392
rect 312096 230382 312124 231676
rect 312084 230376 312136 230382
rect 312084 230318 312136 230324
rect 312372 230042 312400 231676
rect 312360 230036 312412 230042
rect 312360 229978 312412 229984
rect 312544 229968 312596 229974
rect 312544 229910 312596 229916
rect 311440 229900 311492 229906
rect 311440 229842 311492 229848
rect 311348 224256 311400 224262
rect 311348 224198 311400 224204
rect 311452 223038 311480 229842
rect 311440 223032 311492 223038
rect 311440 222974 311492 222980
rect 312556 222154 312584 229910
rect 312740 227322 312768 231676
rect 313108 229294 313136 231676
rect 313188 230376 313240 230382
rect 313188 230318 313240 230324
rect 313096 229288 313148 229294
rect 313096 229230 313148 229236
rect 312728 227316 312780 227322
rect 312728 227258 312780 227264
rect 311164 222148 311216 222154
rect 311164 222090 311216 222096
rect 311992 222148 312044 222154
rect 311992 222090 312044 222096
rect 312544 222148 312596 222154
rect 312544 222090 312596 222096
rect 310520 221468 310572 221474
rect 310520 221410 310572 221416
rect 309416 220108 309468 220114
rect 309416 220050 309468 220056
rect 310244 220108 310296 220114
rect 310244 220050 310296 220056
rect 309428 217410 309456 220050
rect 310532 217410 310560 221410
rect 311164 220720 311216 220726
rect 311164 220662 311216 220668
rect 311176 217410 311204 220662
rect 312004 217410 312032 222090
rect 313200 221202 313228 230318
rect 313476 229634 313504 231676
rect 313844 229974 313872 231676
rect 313832 229968 313884 229974
rect 313832 229910 313884 229916
rect 313464 229628 313516 229634
rect 313464 229570 313516 229576
rect 313556 225684 313608 225690
rect 313556 225626 313608 225632
rect 313188 221196 313240 221202
rect 313188 221138 313240 221144
rect 312820 220652 312872 220658
rect 312820 220594 312872 220600
rect 312832 217410 312860 220594
rect 313568 217410 313596 225626
rect 314212 223242 314240 231676
rect 314476 230308 314528 230314
rect 314476 230250 314528 230256
rect 314488 225690 314516 230250
rect 314580 230246 314608 231676
rect 314948 230382 314976 231676
rect 314936 230376 314988 230382
rect 314936 230318 314988 230324
rect 314568 230240 314620 230246
rect 314568 230182 314620 230188
rect 315224 229770 315252 231676
rect 315304 230444 315356 230450
rect 315304 230386 315356 230392
rect 315212 229764 315264 229770
rect 315212 229706 315264 229712
rect 314568 229628 314620 229634
rect 314568 229570 314620 229576
rect 314476 225684 314528 225690
rect 314476 225626 314528 225632
rect 314200 223236 314252 223242
rect 314200 223178 314252 223184
rect 314580 221270 314608 229570
rect 315316 229094 315344 230386
rect 315316 229066 315436 229094
rect 315304 222148 315356 222154
rect 315304 222090 315356 222096
rect 314568 221264 314620 221270
rect 314568 221206 314620 221212
rect 314660 220244 314712 220250
rect 314660 220186 314712 220192
rect 314672 217410 314700 220186
rect 315316 217410 315344 222090
rect 315408 220250 315436 229066
rect 315592 227390 315620 231676
rect 315868 231662 315974 231690
rect 315868 230110 315896 231662
rect 316328 230382 316356 231676
rect 315948 230376 316000 230382
rect 315948 230318 316000 230324
rect 316316 230376 316368 230382
rect 316316 230318 316368 230324
rect 315856 230104 315908 230110
rect 315856 230046 315908 230052
rect 315580 227384 315632 227390
rect 315580 227326 315632 227332
rect 315960 221338 315988 230318
rect 316696 229906 316724 231676
rect 316684 229900 316736 229906
rect 316684 229842 316736 229848
rect 317064 223174 317092 231676
rect 317328 230376 317380 230382
rect 317328 230318 317380 230324
rect 317052 223168 317104 223174
rect 317052 223110 317104 223116
rect 317340 221406 317368 230318
rect 317432 230314 317460 231676
rect 317420 230308 317472 230314
rect 317420 230250 317472 230256
rect 317800 230246 317828 231676
rect 317788 230240 317840 230246
rect 317788 230182 317840 230188
rect 318076 229838 318104 231676
rect 318064 229832 318116 229838
rect 318064 229774 318116 229780
rect 318064 229288 318116 229294
rect 318064 229230 318116 229236
rect 317420 225752 317472 225758
rect 317420 225694 317472 225700
rect 317328 221400 317380 221406
rect 317328 221342 317380 221348
rect 315948 221332 316000 221338
rect 315948 221274 316000 221280
rect 316132 220516 316184 220522
rect 316132 220458 316184 220464
rect 315396 220244 315448 220250
rect 315396 220186 315448 220192
rect 316144 217410 316172 220458
rect 317432 217410 317460 225694
rect 317880 220584 317932 220590
rect 317880 220526 317932 220532
rect 302620 217382 303048 217410
rect 303632 217382 303876 217410
rect 304276 217382 304704 217410
rect 305288 217382 305624 217410
rect 306392 217382 306452 217410
rect 306944 217382 307280 217410
rect 307772 217382 308108 217410
rect 308600 217382 308936 217410
rect 309428 217382 309764 217410
rect 310532 217382 310592 217410
rect 311176 217382 311512 217410
rect 312004 217382 312340 217410
rect 312832 217382 313168 217410
rect 313568 217382 313996 217410
rect 314672 217382 314824 217410
rect 315316 217382 315652 217410
rect 316144 217382 316480 217410
rect 317400 217382 317460 217410
rect 317892 217410 317920 220526
rect 318076 219978 318104 229230
rect 318444 227254 318472 231676
rect 318708 230240 318760 230246
rect 318708 230182 318760 230188
rect 318432 227248 318484 227254
rect 318432 227190 318484 227196
rect 318720 222154 318748 230182
rect 318812 229702 318840 231676
rect 319194 231662 319484 231690
rect 319562 231662 319852 231690
rect 319260 230376 319312 230382
rect 319260 230318 319312 230324
rect 318800 229696 318852 229702
rect 318800 229638 318852 229644
rect 319272 223106 319300 230318
rect 319352 230172 319404 230178
rect 319352 230114 319404 230120
rect 319260 223100 319312 223106
rect 319260 223042 319312 223048
rect 318892 223032 318944 223038
rect 318892 222974 318944 222980
rect 318708 222148 318760 222154
rect 318708 222090 318760 222096
rect 318064 219972 318116 219978
rect 318064 219914 318116 219920
rect 318904 217410 318932 222974
rect 319364 220046 319392 230114
rect 319456 221542 319484 231662
rect 319444 221536 319496 221542
rect 319444 221478 319496 221484
rect 319824 221474 319852 231662
rect 319916 230382 319944 231676
rect 319904 230376 319956 230382
rect 319904 230318 319956 230324
rect 320284 230314 320312 231676
rect 320666 231662 320864 231690
rect 320942 231662 321232 231690
rect 320272 230308 320324 230314
rect 320272 230250 320324 230256
rect 320272 227044 320324 227050
rect 320272 226986 320324 226992
rect 319812 221468 319864 221474
rect 319812 221410 319864 221416
rect 319536 220448 319588 220454
rect 319536 220390 319588 220396
rect 319352 220040 319404 220046
rect 319352 219982 319404 219988
rect 319548 217410 319576 220390
rect 320284 217410 320312 226986
rect 320836 222086 320864 231662
rect 320824 222080 320876 222086
rect 320824 222022 320876 222028
rect 321204 221950 321232 231662
rect 321296 227186 321324 231676
rect 321664 230246 321692 231676
rect 322046 231662 322336 231690
rect 322414 231662 322704 231690
rect 321652 230240 321704 230246
rect 321652 230182 321704 230188
rect 322204 230104 322256 230110
rect 322204 230046 322256 230052
rect 321284 227180 321336 227186
rect 321284 227122 321336 227128
rect 321928 222964 321980 222970
rect 321928 222906 321980 222912
rect 321192 221944 321244 221950
rect 321192 221886 321244 221892
rect 321560 220380 321612 220386
rect 321560 220322 321612 220328
rect 321572 217410 321600 220322
rect 317892 217382 318228 217410
rect 318904 217382 319056 217410
rect 319548 217382 319884 217410
rect 320284 217382 320712 217410
rect 321540 217382 321600 217410
rect 321940 217410 321968 222906
rect 322216 220522 322244 230046
rect 322308 222018 322336 231662
rect 322296 222012 322348 222018
rect 322296 221954 322348 221960
rect 322676 221882 322704 231662
rect 322768 225962 322796 231676
rect 323136 230450 323164 231676
rect 323124 230444 323176 230450
rect 323124 230386 323176 230392
rect 323504 230382 323532 231676
rect 323492 230376 323544 230382
rect 323492 230318 323544 230324
rect 323780 230110 323808 231676
rect 323768 230104 323820 230110
rect 323768 230046 323820 230052
rect 323676 228540 323728 228546
rect 323676 228482 323728 228488
rect 322756 225956 322808 225962
rect 322756 225898 322808 225904
rect 322664 221876 322716 221882
rect 322664 221818 322716 221824
rect 322204 220516 322256 220522
rect 322204 220458 322256 220464
rect 322940 220312 322992 220318
rect 322940 220254 322992 220260
rect 322952 217410 322980 220254
rect 323688 217410 323716 228482
rect 324148 225826 324176 231676
rect 324530 231662 324820 231690
rect 324898 231662 325188 231690
rect 325266 231662 325556 231690
rect 324228 230376 324280 230382
rect 324228 230318 324280 230324
rect 324136 225820 324188 225826
rect 324136 225762 324188 225768
rect 324240 221814 324268 230318
rect 324504 222896 324556 222902
rect 324504 222838 324556 222844
rect 324228 221808 324280 221814
rect 324228 221750 324280 221756
rect 324516 217410 324544 222838
rect 324792 220794 324820 231662
rect 325160 221746 325188 231662
rect 325148 221740 325200 221746
rect 325148 221682 325200 221688
rect 325528 221610 325556 231662
rect 325620 227118 325648 231676
rect 326002 231662 326292 231690
rect 326370 231662 326568 231690
rect 325608 227112 325660 227118
rect 325608 227054 325660 227060
rect 325700 224392 325752 224398
rect 325700 224334 325752 224340
rect 325516 221604 325568 221610
rect 325516 221546 325568 221552
rect 324780 220788 324832 220794
rect 324780 220730 324832 220736
rect 325712 217410 325740 224334
rect 326264 220726 326292 231662
rect 326540 221678 326568 231662
rect 326632 222970 326660 231676
rect 327000 225894 327028 231676
rect 327368 229566 327396 231676
rect 327356 229560 327408 229566
rect 327356 229502 327408 229508
rect 327736 228886 327764 231676
rect 327724 228880 327776 228886
rect 327724 228822 327776 228828
rect 328104 228750 328132 231676
rect 328472 230450 328500 231676
rect 328460 230444 328512 230450
rect 328460 230386 328512 230392
rect 328840 229634 328868 231676
rect 328828 229628 328880 229634
rect 328828 229570 328880 229576
rect 329208 228954 329236 231676
rect 329196 228948 329248 228954
rect 329196 228890 329248 228896
rect 328092 228744 328144 228750
rect 328092 228686 328144 228692
rect 327816 228472 327868 228478
rect 327816 228414 327868 228420
rect 327080 228404 327132 228410
rect 327080 228346 327132 228352
rect 326988 225888 327040 225894
rect 326988 225830 327040 225836
rect 326620 222964 326672 222970
rect 326620 222906 326672 222912
rect 326528 221672 326580 221678
rect 326528 221614 326580 221620
rect 326252 220720 326304 220726
rect 326252 220662 326304 220668
rect 326252 220176 326304 220182
rect 326252 220118 326304 220124
rect 326264 217410 326292 220118
rect 327092 217410 327120 228346
rect 327828 217410 327856 228414
rect 329484 227050 329512 231676
rect 329852 230450 329880 231676
rect 329564 230444 329616 230450
rect 329564 230386 329616 230392
rect 329840 230444 329892 230450
rect 329840 230386 329892 230392
rect 329472 227044 329524 227050
rect 329472 226986 329524 226992
rect 328736 224324 328788 224330
rect 328736 224266 328788 224272
rect 328748 217410 328776 224266
rect 329576 220658 329604 230386
rect 330220 230178 330248 231676
rect 330116 230172 330168 230178
rect 330116 230114 330168 230120
rect 330208 230172 330260 230178
rect 330208 230114 330260 230120
rect 330128 229634 330156 230114
rect 329656 229628 329708 229634
rect 329656 229570 329708 229576
rect 330116 229628 330168 229634
rect 330116 229570 330168 229576
rect 329564 220652 329616 220658
rect 329564 220594 329616 220600
rect 329668 220590 329696 229570
rect 330588 228818 330616 231676
rect 330852 230444 330904 230450
rect 330852 230386 330904 230392
rect 330576 228812 330628 228818
rect 330576 228754 330628 228760
rect 330392 227452 330444 227458
rect 330392 227394 330444 227400
rect 329656 220584 329708 220590
rect 329656 220526 329708 220532
rect 329840 220108 329892 220114
rect 329840 220050 329892 220056
rect 329852 217410 329880 220050
rect 330404 217410 330432 227394
rect 330864 220454 330892 230386
rect 330956 223038 330984 231676
rect 331036 230172 331088 230178
rect 331036 230114 331088 230120
rect 330944 223032 330996 223038
rect 330944 222974 330996 222980
rect 330852 220448 330904 220454
rect 330852 220390 330904 220396
rect 331048 220318 331076 230114
rect 331324 229362 331352 231676
rect 331692 230450 331720 231676
rect 331680 230444 331732 230450
rect 331680 230386 331732 230392
rect 331312 229356 331364 229362
rect 331312 229298 331364 229304
rect 332060 229022 332088 231676
rect 332232 229356 332284 229362
rect 332232 229298 332284 229304
rect 332048 229016 332100 229022
rect 332048 228958 332100 228964
rect 331220 225684 331272 225690
rect 331220 225626 331272 225632
rect 331036 220312 331088 220318
rect 331036 220254 331088 220260
rect 331232 217870 331260 225626
rect 331312 224256 331364 224262
rect 331312 224198 331364 224204
rect 331220 217864 331272 217870
rect 331220 217806 331272 217812
rect 331324 217410 331352 224198
rect 332244 220386 332272 229298
rect 332336 224738 332364 231676
rect 332416 230444 332468 230450
rect 332416 230386 332468 230392
rect 332324 224732 332376 224738
rect 332324 224674 332376 224680
rect 332232 220380 332284 220386
rect 332232 220322 332284 220328
rect 332428 220182 332456 230386
rect 332704 229430 332732 231676
rect 333072 230450 333100 231676
rect 333454 231662 333652 231690
rect 333624 230518 333652 231662
rect 333716 231662 333822 231690
rect 333612 230512 333664 230518
rect 333612 230454 333664 230460
rect 333060 230444 333112 230450
rect 333060 230386 333112 230392
rect 332692 229424 332744 229430
rect 332692 229366 332744 229372
rect 333716 224466 333744 231662
rect 333796 230444 333848 230450
rect 333796 230386 333848 230392
rect 333704 224460 333756 224466
rect 333704 224402 333756 224408
rect 332968 220244 333020 220250
rect 332968 220186 333020 220192
rect 332416 220176 332468 220182
rect 332416 220118 332468 220124
rect 332140 217864 332192 217870
rect 332140 217806 332192 217812
rect 332152 217410 332180 217806
rect 332980 217410 333008 220186
rect 333808 220114 333836 230386
rect 333888 229424 333940 229430
rect 333888 229366 333940 229372
rect 333900 220250 333928 229366
rect 334176 228206 334204 231676
rect 334544 229430 334572 231676
rect 334716 229696 334768 229702
rect 334716 229638 334768 229644
rect 334624 229628 334676 229634
rect 334624 229570 334676 229576
rect 334532 229424 334584 229430
rect 334532 229366 334584 229372
rect 334164 228200 334216 228206
rect 334164 228142 334216 228148
rect 333980 227316 334032 227322
rect 333980 227258 334032 227264
rect 333888 220244 333940 220250
rect 333888 220186 333940 220192
rect 333796 220108 333848 220114
rect 333796 220050 333848 220056
rect 333992 217870 334020 227258
rect 334072 225616 334124 225622
rect 334072 225558 334124 225564
rect 333980 217864 334032 217870
rect 333980 217806 334032 217812
rect 334084 217410 334112 225558
rect 334636 219706 334664 229570
rect 334728 219774 334756 229638
rect 334912 228682 334940 231676
rect 334900 228676 334952 228682
rect 334900 228618 334952 228624
rect 335188 227322 335216 231676
rect 335176 227316 335228 227322
rect 335176 227258 335228 227264
rect 335556 224126 335584 231676
rect 335924 226098 335952 231676
rect 336292 228614 336320 231676
rect 336660 230178 336688 231676
rect 336648 230172 336700 230178
rect 336648 230114 336700 230120
rect 336924 230036 336976 230042
rect 336924 229978 336976 229984
rect 336280 228608 336332 228614
rect 336280 228550 336332 228556
rect 335912 226092 335964 226098
rect 335912 226034 335964 226040
rect 335544 224120 335596 224126
rect 335544 224062 335596 224068
rect 335544 221196 335596 221202
rect 335544 221138 335596 221144
rect 334716 219768 334768 219774
rect 334716 219710 334768 219716
rect 334624 219700 334676 219706
rect 334624 219642 334676 219648
rect 334716 217864 334768 217870
rect 334716 217806 334768 217812
rect 334728 217410 334756 217806
rect 335556 217410 335584 221138
rect 336740 219972 336792 219978
rect 336740 219914 336792 219920
rect 336752 217410 336780 219914
rect 336936 219434 336964 229978
rect 337028 224602 337056 231676
rect 337410 231662 337700 231690
rect 337384 230308 337436 230314
rect 337384 230250 337436 230256
rect 337016 224596 337068 224602
rect 337016 224538 337068 224544
rect 337396 219842 337424 230250
rect 337672 222902 337700 231662
rect 337764 228546 337792 231676
rect 338040 229634 338068 231676
rect 338028 229628 338080 229634
rect 338028 229570 338080 229576
rect 337752 228540 337804 228546
rect 337752 228482 337804 228488
rect 338408 224670 338436 231676
rect 338790 231662 339080 231690
rect 338764 230240 338816 230246
rect 338764 230182 338816 230188
rect 338396 224664 338448 224670
rect 338396 224606 338448 224612
rect 338120 223236 338172 223242
rect 338120 223178 338172 223184
rect 337660 222896 337712 222902
rect 337660 222838 337712 222844
rect 337384 219836 337436 219842
rect 337384 219778 337436 219784
rect 336936 219406 337148 219434
rect 321940 217382 322368 217410
rect 322952 217382 323288 217410
rect 323688 217382 324116 217410
rect 324516 217382 324944 217410
rect 325712 217382 325772 217410
rect 326264 217382 326600 217410
rect 327092 217382 327428 217410
rect 327828 217382 328256 217410
rect 328748 217382 329176 217410
rect 329852 217382 330004 217410
rect 330404 217382 330832 217410
rect 331324 217382 331660 217410
rect 332152 217382 332488 217410
rect 332980 217382 333316 217410
rect 334084 217382 334144 217410
rect 334728 217382 335064 217410
rect 335556 217382 335892 217410
rect 336720 217382 336780 217410
rect 337120 217410 337148 219406
rect 338132 217410 338160 223178
rect 338776 219910 338804 230182
rect 339052 225214 339080 231662
rect 339144 230314 339172 231676
rect 339132 230308 339184 230314
rect 339132 230250 339184 230256
rect 339512 229498 339540 231676
rect 339500 229492 339552 229498
rect 339500 229434 339552 229440
rect 339040 225208 339092 225214
rect 339040 225150 339092 225156
rect 339880 224398 339908 231676
rect 340144 230376 340196 230382
rect 340144 230318 340196 230324
rect 339868 224392 339920 224398
rect 339868 224334 339920 224340
rect 338856 221264 338908 221270
rect 338856 221206 338908 221212
rect 338764 219904 338816 219910
rect 338764 219846 338816 219852
rect 338868 217410 338896 221206
rect 339684 220040 339736 220046
rect 339684 219982 339736 219988
rect 339696 217410 339724 219982
rect 340156 219978 340184 230318
rect 340248 225146 340276 231676
rect 340616 228478 340644 231676
rect 340892 229702 340920 231676
rect 341274 231662 341472 231690
rect 341248 229968 341300 229974
rect 341248 229910 341300 229916
rect 340880 229696 340932 229702
rect 340880 229638 340932 229644
rect 340604 228472 340656 228478
rect 340604 228414 340656 228420
rect 340236 225140 340288 225146
rect 340236 225082 340288 225088
rect 340144 219972 340196 219978
rect 340144 219914 340196 219920
rect 341260 217410 341288 229910
rect 341340 227384 341392 227390
rect 341340 227326 341392 227332
rect 337120 217382 337548 217410
rect 338132 217382 338376 217410
rect 338868 217382 339204 217410
rect 339696 217382 340032 217410
rect 340952 217382 341288 217410
rect 341352 217410 341380 227326
rect 341444 224330 341472 231662
rect 341524 229560 341576 229566
rect 341524 229502 341576 229508
rect 341432 224324 341484 224330
rect 341432 224266 341484 224272
rect 341536 220046 341564 229502
rect 341628 225690 341656 231676
rect 341996 230382 342024 231676
rect 341984 230376 342036 230382
rect 341984 230318 342036 230324
rect 342364 229362 342392 231676
rect 342352 229356 342404 229362
rect 342352 229298 342404 229304
rect 341616 225684 341668 225690
rect 341616 225626 341668 225632
rect 342732 224534 342760 231676
rect 342904 229424 342956 229430
rect 342904 229366 342956 229372
rect 342916 224754 342944 229366
rect 343100 225758 343128 231676
rect 343272 229356 343324 229362
rect 343272 229298 343324 229304
rect 343088 225752 343140 225758
rect 343088 225694 343140 225700
rect 342916 224726 343128 224754
rect 342720 224528 342772 224534
rect 342720 224470 342772 224476
rect 342260 221332 342312 221338
rect 342260 221274 342312 221280
rect 341524 220040 341576 220046
rect 341524 219982 341576 219988
rect 342272 217410 342300 221274
rect 343100 220522 343128 224726
rect 343284 221066 343312 229298
rect 343468 228070 343496 231676
rect 343744 230042 343772 231676
rect 343732 230036 343784 230042
rect 343732 229978 343784 229984
rect 343732 229764 343784 229770
rect 343732 229706 343784 229712
rect 343744 229094 343772 229706
rect 343744 229066 343864 229094
rect 343456 228064 343508 228070
rect 343456 228006 343508 228012
rect 343272 221060 343324 221066
rect 343272 221002 343324 221008
rect 342996 220516 343048 220522
rect 342996 220458 343048 220464
rect 343088 220516 343140 220522
rect 343088 220458 343140 220464
rect 343008 217410 343036 220458
rect 343836 217410 343864 229066
rect 344112 224262 344140 231676
rect 344480 225622 344508 231676
rect 344848 229770 344876 231676
rect 344836 229764 344888 229770
rect 344836 229706 344888 229712
rect 345216 228410 345244 231676
rect 345204 228404 345256 228410
rect 345204 228346 345256 228352
rect 344468 225616 344520 225622
rect 344468 225558 344520 225564
rect 344100 224256 344152 224262
rect 344100 224198 344152 224204
rect 345584 224194 345612 231676
rect 345952 225282 345980 231676
rect 346320 228138 346348 231676
rect 346492 229900 346544 229906
rect 346492 229842 346544 229848
rect 346308 228132 346360 228138
rect 346308 228074 346360 228080
rect 345940 225276 345992 225282
rect 345940 225218 345992 225224
rect 346504 224210 346532 229842
rect 346596 229094 346624 231676
rect 346596 229066 346716 229094
rect 345572 224188 345624 224194
rect 346504 224182 346624 224210
rect 345572 224130 345624 224136
rect 345020 223168 345072 223174
rect 345020 223110 345072 223116
rect 345032 217410 345060 223110
rect 345572 221400 345624 221406
rect 345572 221342 345624 221348
rect 345584 217410 345612 221342
rect 346492 219700 346544 219706
rect 346492 219642 346544 219648
rect 346504 217410 346532 219642
rect 346596 219434 346624 224182
rect 346688 222426 346716 229066
rect 346964 223786 346992 231676
rect 347332 223922 347360 231676
rect 347700 230246 347728 231676
rect 347688 230240 347740 230246
rect 347688 230182 347740 230188
rect 348068 229094 348096 231676
rect 348068 229066 348188 229094
rect 348056 227248 348108 227254
rect 348056 227190 348108 227196
rect 347320 223916 347372 223922
rect 347320 223858 347372 223864
rect 346952 223780 347004 223786
rect 346952 223722 347004 223728
rect 346676 222420 346728 222426
rect 346676 222362 346728 222368
rect 346596 219406 347268 219434
rect 347240 217410 347268 219406
rect 348068 217410 348096 227190
rect 348160 222494 348188 229066
rect 348436 223854 348464 231676
rect 348804 225350 348832 231676
rect 349172 228274 349200 231676
rect 349160 228268 349212 228274
rect 349160 228210 349212 228216
rect 348792 225344 348844 225350
rect 348792 225286 348844 225292
rect 348424 223848 348476 223854
rect 348424 223790 348476 223796
rect 349448 222562 349476 231676
rect 349816 223990 349844 231676
rect 350184 230654 350212 231676
rect 350172 230648 350224 230654
rect 350172 230590 350224 230596
rect 350552 229634 350580 231676
rect 350934 231662 351224 231690
rect 351302 231662 351592 231690
rect 350908 229832 350960 229838
rect 350908 229774 350960 229780
rect 350540 229628 350592 229634
rect 350540 229570 350592 229576
rect 349804 223984 349856 223990
rect 349804 223926 349856 223932
rect 350632 223100 350684 223106
rect 350632 223042 350684 223048
rect 349436 222556 349488 222562
rect 349436 222498 349488 222504
rect 348148 222488 348200 222494
rect 348148 222430 348200 222436
rect 349160 222148 349212 222154
rect 349160 222090 349212 222096
rect 349172 217410 349200 222090
rect 349804 219768 349856 219774
rect 349804 219710 349856 219716
rect 349816 217410 349844 219710
rect 350644 217870 350672 223042
rect 350632 217864 350684 217870
rect 350632 217806 350684 217812
rect 350920 217410 350948 229774
rect 351196 222630 351224 231662
rect 351184 222624 351236 222630
rect 351184 222566 351236 222572
rect 351564 221202 351592 231662
rect 351656 226574 351684 231676
rect 352024 229906 352052 231676
rect 352012 229900 352064 229906
rect 352012 229842 352064 229848
rect 351644 226568 351696 226574
rect 351644 226510 351696 226516
rect 352300 223378 352328 231676
rect 352564 229560 352616 229566
rect 352564 229502 352616 229508
rect 352288 223372 352340 223378
rect 352288 223314 352340 223320
rect 352576 221542 352604 229502
rect 352668 222698 352696 231676
rect 353050 231662 353248 231690
rect 352656 222692 352708 222698
rect 352656 222634 352708 222640
rect 352380 221536 352432 221542
rect 352380 221478 352432 221484
rect 352564 221536 352616 221542
rect 352564 221478 352616 221484
rect 351552 221196 351604 221202
rect 351552 221138 351604 221144
rect 351460 217864 351512 217870
rect 351460 217806 351512 217812
rect 351472 217410 351500 217806
rect 352392 217410 352420 221478
rect 353220 219366 353248 231662
rect 353404 228342 353432 231676
rect 353392 228336 353444 228342
rect 353392 228278 353444 228284
rect 353772 223242 353800 231676
rect 354154 231662 354444 231690
rect 353944 229492 353996 229498
rect 353944 229434 353996 229440
rect 353760 223236 353812 223242
rect 353760 223178 353812 223184
rect 353956 221338 353984 229434
rect 354036 221468 354088 221474
rect 354036 221410 354088 221416
rect 353944 221332 353996 221338
rect 353944 221274 353996 221280
rect 353300 219836 353352 219842
rect 353300 219778 353352 219784
rect 353208 219360 353260 219366
rect 353208 219302 353260 219308
rect 353312 217410 353340 219778
rect 354048 217410 354076 221410
rect 354416 219434 354444 231662
rect 354508 226642 354536 231676
rect 354876 229838 354904 231676
rect 354864 229832 354916 229838
rect 354864 229774 354916 229780
rect 354772 227180 354824 227186
rect 354772 227122 354824 227128
rect 354496 226636 354548 226642
rect 354496 226578 354548 226584
rect 354404 219428 354456 219434
rect 354404 219370 354456 219376
rect 354784 217410 354812 227122
rect 355152 222766 355180 231676
rect 355520 229498 355548 231676
rect 355508 229492 355560 229498
rect 355508 229434 355560 229440
rect 355888 226710 355916 231676
rect 356256 229974 356284 231676
rect 356244 229968 356296 229974
rect 356244 229910 356296 229916
rect 355876 226704 355928 226710
rect 355876 226646 355928 226652
rect 356624 222834 356652 231676
rect 356992 225418 357020 231676
rect 357072 229968 357124 229974
rect 357072 229910 357124 229916
rect 356980 225412 357032 225418
rect 356980 225354 357032 225360
rect 356612 222828 356664 222834
rect 356612 222770 356664 222776
rect 355140 222760 355192 222766
rect 355140 222702 355192 222708
rect 356060 222080 356112 222086
rect 356060 222022 356112 222028
rect 356072 217410 356100 222022
rect 357084 221270 357112 229910
rect 357360 226778 357388 231676
rect 357728 229294 357756 231676
rect 357716 229288 357768 229294
rect 357716 229230 357768 229236
rect 357348 226772 357400 226778
rect 357348 226714 357400 226720
rect 358004 223582 358032 231676
rect 358372 226030 358400 231676
rect 358740 226846 358768 231676
rect 359108 229974 359136 231676
rect 359096 229968 359148 229974
rect 359096 229910 359148 229916
rect 358728 226840 358780 226846
rect 358728 226782 358780 226788
rect 358360 226024 358412 226030
rect 358360 225966 358412 225972
rect 358176 225956 358228 225962
rect 358176 225898 358228 225904
rect 357992 223576 358044 223582
rect 357992 223518 358044 223524
rect 357532 221944 357584 221950
rect 357532 221886 357584 221892
rect 357072 221264 357124 221270
rect 357072 221206 357124 221212
rect 356520 219904 356572 219910
rect 356520 219846 356572 219852
rect 341352 217382 341780 217410
rect 342272 217382 342608 217410
rect 343008 217382 343436 217410
rect 343836 217382 344264 217410
rect 345032 217382 345092 217410
rect 345584 217382 345920 217410
rect 346504 217382 346840 217410
rect 347240 217382 347668 217410
rect 348068 217382 348496 217410
rect 349172 217382 349324 217410
rect 349816 217382 350152 217410
rect 350920 217382 350980 217410
rect 351472 217382 351808 217410
rect 352392 217382 352728 217410
rect 353312 217382 353556 217410
rect 354048 217382 354384 217410
rect 354784 217382 355212 217410
rect 356040 217382 356100 217410
rect 356532 217410 356560 219846
rect 357544 217410 357572 221886
rect 358188 217410 358216 225898
rect 359476 223514 359504 231676
rect 359844 225486 359872 231676
rect 360108 229968 360160 229974
rect 360108 229910 360160 229916
rect 359832 225480 359884 225486
rect 359832 225422 359884 225428
rect 359464 223508 359516 223514
rect 359464 223450 359516 223456
rect 359096 222012 359148 222018
rect 359096 221954 359148 221960
rect 359108 217410 359136 221954
rect 360120 221338 360148 229910
rect 360212 227662 360240 231676
rect 360580 229974 360608 231676
rect 360870 231662 361160 231690
rect 360568 229968 360620 229974
rect 360568 229910 360620 229916
rect 360200 227656 360252 227662
rect 360200 227598 360252 227604
rect 360292 227112 360344 227118
rect 360292 227054 360344 227060
rect 360108 221332 360160 221338
rect 360108 221274 360160 221280
rect 360200 219972 360252 219978
rect 360200 219914 360252 219920
rect 360212 217410 360240 219914
rect 360304 219502 360332 227054
rect 361132 223446 361160 231662
rect 361224 229430 361252 231676
rect 361304 229968 361356 229974
rect 361304 229910 361356 229916
rect 361212 229424 361264 229430
rect 361212 229366 361264 229372
rect 361120 223440 361172 223446
rect 361120 223382 361172 223388
rect 360752 221876 360804 221882
rect 360752 221818 360804 221824
rect 360292 219496 360344 219502
rect 360292 219438 360344 219444
rect 360764 217410 360792 221818
rect 361316 221406 361344 229910
rect 361592 226914 361620 231676
rect 361960 229974 361988 231676
rect 362342 231662 362632 231690
rect 362710 231662 362908 231690
rect 362604 230058 362632 231662
rect 362604 230030 362816 230058
rect 362788 229974 362816 230030
rect 361948 229968 362000 229974
rect 361948 229910 362000 229916
rect 362684 229968 362736 229974
rect 362684 229910 362736 229916
rect 362776 229968 362828 229974
rect 362776 229910 362828 229916
rect 361580 226908 361632 226914
rect 361580 226850 361632 226856
rect 361580 225820 361632 225826
rect 361580 225762 361632 225768
rect 361304 221400 361356 221406
rect 361304 221342 361356 221348
rect 361592 217410 361620 225762
rect 362696 222154 362724 229910
rect 362880 225554 362908 231662
rect 363064 226982 363092 231676
rect 363446 231662 363644 231690
rect 363722 231662 364012 231690
rect 364090 231662 364288 231690
rect 363144 227316 363196 227322
rect 363144 227258 363196 227264
rect 363052 226976 363104 226982
rect 363052 226918 363104 226924
rect 362960 225888 363012 225894
rect 362960 225830 363012 225836
rect 362868 225548 362920 225554
rect 362868 225490 362920 225496
rect 362684 222148 362736 222154
rect 362684 222090 362736 222096
rect 362408 221808 362460 221814
rect 362408 221750 362460 221756
rect 362420 217410 362448 221750
rect 362972 219842 363000 225830
rect 363156 219978 363184 227258
rect 363616 222086 363644 231662
rect 363604 222080 363656 222086
rect 363604 222022 363656 222028
rect 363984 221950 364012 231662
rect 364260 226302 364288 231662
rect 364444 227730 364472 231676
rect 364826 231662 365116 231690
rect 364524 230104 364576 230110
rect 364524 230046 364576 230052
rect 364432 227724 364484 227730
rect 364432 227666 364484 227672
rect 364248 226296 364300 226302
rect 364248 226238 364300 226244
rect 363972 221944 364024 221950
rect 363972 221886 364024 221892
rect 363236 220788 363288 220794
rect 363236 220730 363288 220736
rect 363144 219972 363196 219978
rect 363144 219914 363196 219920
rect 362960 219836 363012 219842
rect 362960 219778 363012 219784
rect 363248 217410 363276 220730
rect 364536 217410 364564 230046
rect 365088 222018 365116 231662
rect 365180 229090 365208 231676
rect 365168 229084 365220 229090
rect 365168 229026 365220 229032
rect 365352 227044 365404 227050
rect 365352 226986 365404 226992
rect 365076 222012 365128 222018
rect 365076 221954 365128 221960
rect 365364 219910 365392 226986
rect 365548 226234 365576 231676
rect 365916 227594 365944 231676
rect 366298 231662 366496 231690
rect 365904 227588 365956 227594
rect 365904 227530 365956 227536
rect 365536 226228 365588 226234
rect 365536 226170 365588 226176
rect 365996 223032 366048 223038
rect 365996 222974 366048 222980
rect 365812 221740 365864 221746
rect 365812 221682 365864 221688
rect 365352 219904 365404 219910
rect 365352 219846 365404 219852
rect 364984 219496 365036 219502
rect 364984 219438 365036 219444
rect 356532 217382 356868 217410
rect 357544 217382 357696 217410
rect 358188 217382 358616 217410
rect 359108 217382 359444 217410
rect 360212 217382 360272 217410
rect 360764 217382 361100 217410
rect 361592 217382 361928 217410
rect 362420 217382 362756 217410
rect 363248 217382 363584 217410
rect 364504 217382 364564 217410
rect 364996 217410 365024 219438
rect 365824 217410 365852 221682
rect 366008 220794 366036 222974
rect 366468 221882 366496 231662
rect 366560 229566 366588 231676
rect 366548 229560 366600 229566
rect 366548 229502 366600 229508
rect 366928 226166 366956 231676
rect 367296 227526 367324 231676
rect 367678 231662 367968 231690
rect 367284 227520 367336 227526
rect 367284 227462 367336 227468
rect 366916 226160 366968 226166
rect 366916 226102 366968 226108
rect 367744 226092 367796 226098
rect 367744 226034 367796 226040
rect 366456 221876 366508 221882
rect 366456 221818 366508 221824
rect 367468 221604 367520 221610
rect 367468 221546 367520 221552
rect 365996 220788 366048 220794
rect 365996 220730 366048 220736
rect 366640 220720 366692 220726
rect 366640 220662 366692 220668
rect 366652 217410 366680 220662
rect 367480 217410 367508 221546
rect 367756 220726 367784 226034
rect 367940 221814 367968 231662
rect 368032 230110 368060 231676
rect 368020 230104 368072 230110
rect 368020 230046 368072 230052
rect 368400 226098 368428 231676
rect 368768 227458 368796 231676
rect 369150 231662 369348 231690
rect 368756 227452 368808 227458
rect 368756 227394 368808 227400
rect 368388 226092 368440 226098
rect 368388 226034 368440 226040
rect 367928 221808 367980 221814
rect 367928 221750 367980 221756
rect 369320 221746 369348 231662
rect 369412 229226 369440 231676
rect 369400 229220 369452 229226
rect 369400 229162 369452 229168
rect 369780 225962 369808 231676
rect 370148 227390 370176 231676
rect 370530 231662 370820 231690
rect 370228 229016 370280 229022
rect 370228 228958 370280 228964
rect 370136 227384 370188 227390
rect 370136 227326 370188 227332
rect 369768 225956 369820 225962
rect 369768 225898 369820 225904
rect 369308 221740 369360 221746
rect 369308 221682 369360 221688
rect 369124 221672 369176 221678
rect 369124 221614 369176 221620
rect 367744 220720 367796 220726
rect 367744 220662 367796 220668
rect 368480 219836 368532 219842
rect 368480 219778 368532 219784
rect 368492 217410 368520 219778
rect 369136 217410 369164 221614
rect 370240 220046 370268 228958
rect 370792 221678 370820 231662
rect 370884 224874 370912 231676
rect 371252 225894 371280 231676
rect 371332 228948 371384 228954
rect 371332 228890 371384 228896
rect 371240 225888 371292 225894
rect 371240 225830 371292 225836
rect 370872 224868 370924 224874
rect 370872 224810 370924 224816
rect 371240 222964 371292 222970
rect 371240 222906 371292 222912
rect 370780 221672 370832 221678
rect 370780 221614 370832 221620
rect 370044 220040 370096 220046
rect 370044 219982 370096 219988
rect 370228 220040 370280 220046
rect 370228 219982 370280 219988
rect 370056 217410 370084 219982
rect 371252 217410 371280 222906
rect 371344 219502 371372 228890
rect 371620 227322 371648 231676
rect 371884 230444 371936 230450
rect 371884 230386 371936 230392
rect 371608 227316 371660 227322
rect 371608 227258 371660 227264
rect 371896 220658 371924 230386
rect 371988 229362 372016 231676
rect 371976 229356 372028 229362
rect 371976 229298 372028 229304
rect 372264 224806 372292 231676
rect 372632 225826 372660 231676
rect 372712 228880 372764 228886
rect 372712 228822 372764 228828
rect 372620 225820 372672 225826
rect 372620 225762 372672 225768
rect 372252 224800 372304 224806
rect 372252 224742 372304 224748
rect 372620 224732 372672 224738
rect 372620 224674 372672 224680
rect 371700 220652 371752 220658
rect 371700 220594 371752 220600
rect 371884 220652 371936 220658
rect 371884 220594 371936 220600
rect 371332 219496 371384 219502
rect 371332 219438 371384 219444
rect 364996 217382 365332 217410
rect 365824 217382 366160 217410
rect 366652 217382 366988 217410
rect 367480 217382 367816 217410
rect 368492 217382 368644 217410
rect 369136 217382 369472 217410
rect 370056 217382 370392 217410
rect 371220 217382 371280 217410
rect 371712 217410 371740 220594
rect 372632 219774 372660 224674
rect 372620 219768 372672 219774
rect 372620 219710 372672 219716
rect 372724 217410 372752 228822
rect 373000 227254 373028 231676
rect 373368 229022 373396 231676
rect 373356 229016 373408 229022
rect 373356 228958 373408 228964
rect 372988 227248 373040 227254
rect 372988 227190 373040 227196
rect 373736 224738 373764 231676
rect 374000 228744 374052 228750
rect 374000 228686 374052 228692
rect 373724 224732 373776 224738
rect 373724 224674 373776 224680
rect 373356 220584 373408 220590
rect 373356 220526 373408 220532
rect 373368 217410 373396 220526
rect 374012 219434 374040 228686
rect 374104 224942 374132 231676
rect 374472 227186 374500 231676
rect 374460 227180 374512 227186
rect 374460 227122 374512 227128
rect 374840 227118 374868 231676
rect 375116 228954 375144 231676
rect 375104 228948 375156 228954
rect 375104 228890 375156 228896
rect 375288 228812 375340 228818
rect 375288 228754 375340 228760
rect 374828 227112 374880 227118
rect 374828 227054 374880 227060
rect 374092 224936 374144 224942
rect 374092 224878 374144 224884
rect 375300 220590 375328 228754
rect 375484 227798 375512 231676
rect 375852 230081 375880 231676
rect 376024 230172 376076 230178
rect 376024 230114 376076 230120
rect 375838 230072 375894 230081
rect 375838 230007 375894 230016
rect 375472 227792 375524 227798
rect 375472 227734 375524 227740
rect 375288 220584 375340 220590
rect 375288 220526 375340 220532
rect 376036 220454 376064 230114
rect 376116 229288 376168 229294
rect 376116 229230 376168 229236
rect 376128 221134 376156 229230
rect 376220 223417 376248 231676
rect 376588 228886 376616 231676
rect 376956 230353 376984 231676
rect 376942 230344 376998 230353
rect 376942 230279 376998 230288
rect 377324 230217 377352 231676
rect 377310 230208 377366 230217
rect 377310 230143 377366 230152
rect 376576 228880 376628 228886
rect 376576 228822 376628 228828
rect 377692 224641 377720 231676
rect 377968 228818 377996 231676
rect 378336 230178 378364 231676
rect 378324 230172 378376 230178
rect 378324 230114 378376 230120
rect 378704 229945 378732 231676
rect 378968 230308 379020 230314
rect 378968 230250 379020 230256
rect 378690 229936 378746 229945
rect 378690 229871 378746 229880
rect 378600 229220 378652 229226
rect 378600 229162 378652 229168
rect 377956 228812 378008 228818
rect 377956 228754 378008 228760
rect 378508 228200 378560 228206
rect 378508 228142 378560 228148
rect 377678 224632 377734 224641
rect 377678 224567 377734 224576
rect 378048 224460 378100 224466
rect 378048 224402 378100 224408
rect 377312 224120 377364 224126
rect 377312 224062 377364 224068
rect 376206 223408 376262 223417
rect 376206 223343 376262 223352
rect 376116 221128 376168 221134
rect 376116 221070 376168 221076
rect 377324 220454 377352 224062
rect 375380 220448 375432 220454
rect 375380 220390 375432 220396
rect 376024 220448 376076 220454
rect 376024 220390 376076 220396
rect 377312 220448 377364 220454
rect 377312 220390 377364 220396
rect 374012 219406 374132 219434
rect 374104 217410 374132 219406
rect 375392 217410 375420 220390
rect 376208 220380 376260 220386
rect 376208 220322 376260 220328
rect 376220 219842 376248 220322
rect 376944 220312 376996 220318
rect 376944 220254 376996 220260
rect 376208 219836 376260 219842
rect 376208 219778 376260 219784
rect 375932 219496 375984 219502
rect 375932 219438 375984 219444
rect 371712 217382 372048 217410
rect 372724 217382 372876 217410
rect 373368 217382 373704 217410
rect 374104 217382 374532 217410
rect 375360 217382 375420 217410
rect 375944 217410 375972 219438
rect 376956 217410 376984 220254
rect 377588 219904 377640 219910
rect 377588 219846 377640 219852
rect 377600 217410 377628 219846
rect 378060 219706 378088 224402
rect 378416 219836 378468 219842
rect 378416 219778 378468 219784
rect 378048 219700 378100 219706
rect 378048 219642 378100 219648
rect 378428 217410 378456 219778
rect 378520 219502 378548 228142
rect 378612 224126 378640 229162
rect 378980 228206 379008 230250
rect 378968 228200 379020 228206
rect 378968 228142 379020 228148
rect 378692 224596 378744 224602
rect 378692 224538 378744 224544
rect 378600 224120 378652 224126
rect 378600 224062 378652 224068
rect 378704 220318 378732 224538
rect 379072 223281 379100 231676
rect 379058 223272 379114 223281
rect 379058 223207 379114 223216
rect 378692 220312 378744 220318
rect 378692 220254 378744 220260
rect 378508 219496 378560 219502
rect 378508 219438 378560 219444
rect 379440 219298 379468 231676
rect 379704 227792 379756 227798
rect 379704 227734 379756 227740
rect 379520 220584 379572 220590
rect 379520 220526 379572 220532
rect 379612 220584 379664 220590
rect 379612 220526 379664 220532
rect 379428 219292 379480 219298
rect 379428 219234 379480 219240
rect 379532 217410 379560 220526
rect 379624 220386 379652 220526
rect 379612 220380 379664 220386
rect 379612 220322 379664 220328
rect 379716 219842 379744 227734
rect 379808 222970 379836 231676
rect 380176 229809 380204 231676
rect 380440 230376 380492 230382
rect 380440 230318 380492 230324
rect 380162 229800 380218 229809
rect 380162 229735 380218 229744
rect 380256 229696 380308 229702
rect 380256 229638 380308 229644
rect 380164 224664 380216 224670
rect 380164 224606 380216 224612
rect 379796 222964 379848 222970
rect 379796 222906 379848 222912
rect 380176 220182 380204 224606
rect 380268 220930 380296 229638
rect 380452 227798 380480 230318
rect 380440 227792 380492 227798
rect 380440 227734 380492 227740
rect 380544 227361 380572 231676
rect 380530 227352 380586 227361
rect 380530 227287 380586 227296
rect 380256 220924 380308 220930
rect 380256 220866 380308 220872
rect 380072 220176 380124 220182
rect 380072 220118 380124 220124
rect 380164 220176 380216 220182
rect 380164 220118 380216 220124
rect 379704 219836 379756 219842
rect 379704 219778 379756 219784
rect 380084 217410 380112 220118
rect 380820 219230 380848 231676
rect 381188 230382 381216 231676
rect 381570 231662 381860 231690
rect 381176 230376 381228 230382
rect 381176 230318 381228 230324
rect 381832 224346 381860 231662
rect 381924 224505 381952 231676
rect 382292 230450 382320 231676
rect 382280 230444 382332 230450
rect 382280 230386 382332 230392
rect 382660 230382 382688 231676
rect 382188 230376 382240 230382
rect 382188 230318 382240 230324
rect 382648 230376 382700 230382
rect 382648 230318 382700 230324
rect 381910 224496 381966 224505
rect 381910 224431 381966 224440
rect 381832 224318 381952 224346
rect 380900 220788 380952 220794
rect 380900 220730 380952 220736
rect 380808 219224 380860 219230
rect 380808 219166 380860 219172
rect 380912 217410 380940 220730
rect 381924 220289 381952 224318
rect 382200 220425 382228 230318
rect 383028 227225 383056 231676
rect 383410 231662 383516 231690
rect 383384 230376 383436 230382
rect 383384 230318 383436 230324
rect 383108 229424 383160 229430
rect 383108 229366 383160 229372
rect 383014 227216 383070 227225
rect 383014 227151 383070 227160
rect 383120 225214 383148 229366
rect 382280 225208 382332 225214
rect 382280 225150 382332 225156
rect 383108 225208 383160 225214
rect 383108 225150 383160 225156
rect 382186 220416 382242 220425
rect 382186 220351 382242 220360
rect 381910 220280 381966 220289
rect 381820 220244 381872 220250
rect 382292 220250 382320 225150
rect 383396 220794 383424 230318
rect 383384 220788 383436 220794
rect 383384 220730 383436 220736
rect 381910 220215 381966 220224
rect 382280 220244 382332 220250
rect 381820 220186 381872 220192
rect 382280 220186 382332 220192
rect 381832 217410 381860 220186
rect 382648 220040 382700 220046
rect 382648 219982 382700 219988
rect 382660 217410 382688 219982
rect 383488 219094 383516 231662
rect 383568 230444 383620 230450
rect 383568 230386 383620 230392
rect 383580 219162 383608 230386
rect 383672 230382 383700 231676
rect 383660 230376 383712 230382
rect 383660 230318 383712 230324
rect 384040 224369 384068 231676
rect 384408 229294 384436 231676
rect 384790 231662 384896 231690
rect 384396 229288 384448 229294
rect 384396 229230 384448 229236
rect 384026 224360 384082 224369
rect 384026 224295 384082 224304
rect 384868 220153 384896 231662
rect 385144 230586 385172 231676
rect 385132 230580 385184 230586
rect 385132 230522 385184 230528
rect 385512 230382 385540 231676
rect 384948 230376 385000 230382
rect 384948 230318 385000 230324
rect 385500 230376 385552 230382
rect 385500 230318 385552 230324
rect 384854 220144 384910 220153
rect 383660 220108 383712 220114
rect 384854 220079 384910 220088
rect 383660 220050 383712 220056
rect 383568 219156 383620 219162
rect 383568 219098 383620 219104
rect 383476 219088 383528 219094
rect 383476 219030 383528 219036
rect 383672 217410 383700 220050
rect 384960 220046 384988 230318
rect 385880 230314 385908 231676
rect 386248 230518 386276 231676
rect 386236 230512 386288 230518
rect 386236 230454 386288 230460
rect 386524 230382 386552 231676
rect 386892 230450 386920 231676
rect 386880 230444 386932 230450
rect 386880 230386 386932 230392
rect 386328 230376 386380 230382
rect 386328 230318 386380 230324
rect 386512 230376 386564 230382
rect 386512 230318 386564 230324
rect 385868 230308 385920 230314
rect 385868 230250 385920 230256
rect 385684 230036 385736 230042
rect 385684 229978 385736 229984
rect 385696 229094 385724 229978
rect 385696 229066 385816 229094
rect 385684 225140 385736 225146
rect 385684 225082 385736 225088
rect 385696 220114 385724 225082
rect 385788 220998 385816 229066
rect 385776 220992 385828 220998
rect 385776 220934 385828 220940
rect 385960 220652 386012 220658
rect 385960 220594 386012 220600
rect 385684 220108 385736 220114
rect 385684 220050 385736 220056
rect 384948 220040 385000 220046
rect 384948 219982 385000 219988
rect 384304 219768 384356 219774
rect 384304 219710 384356 219716
rect 384316 217410 384344 219710
rect 385132 219496 385184 219502
rect 385132 219438 385184 219444
rect 385144 217410 385172 219438
rect 385972 217410 386000 220594
rect 386340 219026 386368 230318
rect 386972 229492 387024 229498
rect 386972 229434 387024 229440
rect 386984 225146 387012 229434
rect 387260 228721 387288 231676
rect 387642 231662 387748 231690
rect 387720 230466 387748 231662
rect 387720 230438 387840 230466
rect 387812 230382 387840 230438
rect 387708 230376 387760 230382
rect 387708 230318 387760 230324
rect 387800 230376 387852 230382
rect 387800 230318 387852 230324
rect 387616 230240 387668 230246
rect 387616 230182 387668 230188
rect 387524 230104 387576 230110
rect 387524 230046 387576 230052
rect 387246 228712 387302 228721
rect 387246 228647 387302 228656
rect 387248 228064 387300 228070
rect 387248 228006 387300 228012
rect 386972 225140 387024 225146
rect 386972 225082 387024 225088
rect 386972 224392 387024 224398
rect 386972 224334 387024 224340
rect 386788 220516 386840 220522
rect 386788 220458 386840 220464
rect 386328 219020 386380 219026
rect 386328 218962 386380 218968
rect 386800 217410 386828 220458
rect 386984 219910 387012 224334
rect 386972 219904 387024 219910
rect 386972 219846 387024 219852
rect 387260 219774 387288 228006
rect 387536 224058 387564 230046
rect 387628 227934 387656 230182
rect 387616 227928 387668 227934
rect 387616 227870 387668 227876
rect 387524 224052 387576 224058
rect 387524 223994 387576 224000
rect 387248 219768 387300 219774
rect 387248 219710 387300 219716
rect 387720 218958 387748 230318
rect 387996 230110 388024 231676
rect 387984 230104 388036 230110
rect 387984 230046 388036 230052
rect 388076 229628 388128 229634
rect 388076 229570 388128 229576
rect 388088 228002 388116 229570
rect 388076 227996 388128 228002
rect 388076 227938 388128 227944
rect 388364 227089 388392 231676
rect 388444 230444 388496 230450
rect 388444 230386 388496 230392
rect 388350 227080 388406 227089
rect 388350 227015 388406 227024
rect 388456 220658 388484 230386
rect 388732 224670 388760 231676
rect 389100 230246 389128 231676
rect 389088 230240 389140 230246
rect 389088 230182 389140 230188
rect 389272 228676 389324 228682
rect 389272 228618 389324 228624
rect 388720 224664 388772 224670
rect 388720 224606 388772 224612
rect 389180 222964 389232 222970
rect 389180 222906 389232 222912
rect 388444 220652 388496 220658
rect 388444 220594 388496 220600
rect 389192 220561 389220 222906
rect 389178 220552 389234 220561
rect 389178 220487 389234 220496
rect 388536 220448 388588 220454
rect 388536 220390 388588 220396
rect 387800 219700 387852 219706
rect 387800 219642 387852 219648
rect 387708 218952 387760 218958
rect 387708 218894 387760 218900
rect 387812 217410 387840 219642
rect 388548 217410 388576 220390
rect 389284 217410 389312 228618
rect 389376 223145 389404 231676
rect 389744 224602 389772 231676
rect 389732 224596 389784 224602
rect 389732 224538 389784 224544
rect 390112 223310 390140 231676
rect 390100 223304 390152 223310
rect 390100 223246 390152 223252
rect 389362 223136 389418 223145
rect 389362 223071 389418 223080
rect 390480 223009 390508 231676
rect 390848 226001 390876 231676
rect 391112 230308 391164 230314
rect 391112 230250 391164 230256
rect 390834 225992 390890 226001
rect 390834 225927 390890 225936
rect 390466 223000 390522 223009
rect 390466 222935 390522 222944
rect 390652 222896 390704 222902
rect 390652 222838 390704 222844
rect 390560 220720 390612 220726
rect 390560 220662 390612 220668
rect 390572 217410 390600 220662
rect 390664 219502 390692 222838
rect 391124 219978 391152 230250
rect 391216 229702 391244 231676
rect 391204 229696 391256 229702
rect 391204 229638 391256 229644
rect 391584 223106 391612 231676
rect 391952 228750 391980 231676
rect 392228 229430 392256 231676
rect 392610 231662 392900 231690
rect 392584 229696 392636 229702
rect 392584 229638 392636 229644
rect 392216 229424 392268 229430
rect 392216 229366 392268 229372
rect 391940 228744 391992 228750
rect 391940 228686 391992 228692
rect 392492 228608 392544 228614
rect 392492 228550 392544 228556
rect 391572 223100 391624 223106
rect 391572 223042 391624 223048
rect 391940 220312 391992 220318
rect 391940 220254 391992 220260
rect 391020 219972 391072 219978
rect 391020 219914 391072 219920
rect 391112 219972 391164 219978
rect 391112 219914 391164 219920
rect 390652 219496 390704 219502
rect 390652 219438 390704 219444
rect 375944 217382 376280 217410
rect 376956 217382 377108 217410
rect 377600 217382 377936 217410
rect 378428 217382 378764 217410
rect 379532 217382 379592 217410
rect 380084 217382 380420 217410
rect 380912 217382 381248 217410
rect 381832 217382 382168 217410
rect 382660 217382 382996 217410
rect 383672 217382 383824 217410
rect 384316 217382 384652 217410
rect 385144 217382 385480 217410
rect 385972 217382 386308 217410
rect 386800 217382 387136 217410
rect 387812 217382 388056 217410
rect 388548 217382 388884 217410
rect 389284 217382 389712 217410
rect 390540 217382 390600 217410
rect 391032 217410 391060 219914
rect 391952 217410 391980 220254
rect 392504 219434 392532 228550
rect 392596 220522 392624 229638
rect 392872 221785 392900 231662
rect 392964 228682 392992 231676
rect 393332 230450 393360 231676
rect 393320 230444 393372 230450
rect 393320 230386 393372 230392
rect 393700 229498 393728 231676
rect 393688 229492 393740 229498
rect 393688 229434 393740 229440
rect 392952 228676 393004 228682
rect 392952 228618 393004 228624
rect 394068 225865 394096 231676
rect 394450 231662 394556 231690
rect 394054 225856 394110 225865
rect 394054 225791 394110 225800
rect 392858 221776 392914 221785
rect 392858 221711 392914 221720
rect 392584 220516 392636 220522
rect 392584 220458 392636 220464
rect 394528 219502 394556 231662
rect 394608 230444 394660 230450
rect 394608 230386 394660 230392
rect 394620 220454 394648 230386
rect 394804 222970 394832 231676
rect 395080 229226 395108 231676
rect 395462 231662 395752 231690
rect 395068 229220 395120 229226
rect 395068 229162 395120 229168
rect 395724 229094 395752 231662
rect 395632 229066 395752 229094
rect 394792 222964 394844 222970
rect 394792 222906 394844 222912
rect 394700 220584 394752 220590
rect 394700 220526 394752 220532
rect 394608 220448 394660 220454
rect 394608 220390 394660 220396
rect 393596 219496 393648 219502
rect 393596 219438 393648 219444
rect 394516 219496 394568 219502
rect 394516 219438 394568 219444
rect 392504 219406 392624 219434
rect 392596 217410 392624 219406
rect 393608 217410 393636 219438
rect 394712 217410 394740 220526
rect 395632 220386 395660 229066
rect 395712 223304 395764 223310
rect 395712 223246 395764 223252
rect 395724 220590 395752 223246
rect 395816 223174 395844 231676
rect 396198 231662 396488 231690
rect 396566 231662 396856 231690
rect 396934 231662 397224 231690
rect 396172 228540 396224 228546
rect 396172 228482 396224 228488
rect 395804 223168 395856 223174
rect 395804 223110 395856 223116
rect 395712 220584 395764 220590
rect 395712 220526 395764 220532
rect 395620 220380 395672 220386
rect 395620 220322 395672 220328
rect 395252 220176 395304 220182
rect 395252 220118 395304 220124
rect 395264 217410 395292 220118
rect 396184 217410 396212 228482
rect 396460 225729 396488 231662
rect 396724 230240 396776 230246
rect 396724 230182 396776 230188
rect 396446 225720 396502 225729
rect 396446 225655 396502 225664
rect 396356 223304 396408 223310
rect 396356 223246 396408 223252
rect 396368 223106 396396 223246
rect 396356 223100 396408 223106
rect 396356 223042 396408 223048
rect 396736 220726 396764 230182
rect 396724 220720 396776 220726
rect 396724 220662 396776 220668
rect 396828 220318 396856 231662
rect 397196 221649 397224 231662
rect 397288 228546 397316 231676
rect 397656 229634 397684 231676
rect 397644 229628 397696 229634
rect 397644 229570 397696 229576
rect 397276 228540 397328 228546
rect 397276 228482 397328 228488
rect 397932 223038 397960 231676
rect 398104 230240 398156 230246
rect 398104 230182 398156 230188
rect 398116 229906 398144 230182
rect 398104 229900 398156 229906
rect 398104 229842 398156 229848
rect 398300 228614 398328 231676
rect 398668 230314 398696 231676
rect 398656 230308 398708 230314
rect 398656 230250 398708 230256
rect 399036 230042 399064 231676
rect 399024 230036 399076 230042
rect 399024 229978 399076 229984
rect 398564 229628 398616 229634
rect 398564 229570 398616 229576
rect 398656 229628 398708 229634
rect 398656 229570 398708 229576
rect 398288 228608 398340 228614
rect 398288 228550 398340 228556
rect 397920 223032 397972 223038
rect 397920 222974 397972 222980
rect 397182 221640 397238 221649
rect 397182 221575 397238 221584
rect 397736 221536 397788 221542
rect 397736 221478 397788 221484
rect 396816 220312 396868 220318
rect 396816 220254 396868 220260
rect 396908 220244 396960 220250
rect 396908 220186 396960 220192
rect 396920 217410 396948 220186
rect 397748 217410 397776 221478
rect 398576 220182 398604 229570
rect 398668 229362 398696 229570
rect 398656 229356 398708 229362
rect 398656 229298 398708 229304
rect 399404 228585 399432 231676
rect 399772 229906 399800 231676
rect 400048 231662 400154 231690
rect 399760 229900 399812 229906
rect 399760 229842 399812 229848
rect 399390 228576 399446 228585
rect 399390 228511 399446 228520
rect 399392 228200 399444 228206
rect 399392 228142 399444 228148
rect 398840 223168 398892 223174
rect 398840 223110 398892 223116
rect 398852 222970 398880 223110
rect 398840 222964 398892 222970
rect 398840 222906 398892 222912
rect 398564 220176 398616 220182
rect 398564 220118 398616 220124
rect 398840 219904 398892 219910
rect 398840 219846 398892 219852
rect 398852 217410 398880 219846
rect 399404 217410 399432 228142
rect 400048 224466 400076 231662
rect 400128 230036 400180 230042
rect 400128 229978 400180 229984
rect 400036 224460 400088 224466
rect 400036 224402 400088 224408
rect 400140 221610 400168 229978
rect 400508 225593 400536 231676
rect 400680 230376 400732 230382
rect 400680 230318 400732 230324
rect 400494 225584 400550 225593
rect 400494 225519 400550 225528
rect 400128 221604 400180 221610
rect 400128 221546 400180 221552
rect 400312 220108 400364 220114
rect 400312 220050 400364 220056
rect 400324 217410 400352 220050
rect 400692 219910 400720 230318
rect 400784 229702 400812 231676
rect 401152 230042 401180 231676
rect 401140 230036 401192 230042
rect 401140 229978 401192 229984
rect 400772 229696 400824 229702
rect 400772 229638 400824 229644
rect 401520 229498 401548 231676
rect 401888 230450 401916 231676
rect 401876 230444 401928 230450
rect 401876 230386 401928 230392
rect 400956 229492 401008 229498
rect 400956 229434 401008 229440
rect 401508 229492 401560 229498
rect 401508 229434 401560 229440
rect 400968 221921 400996 229434
rect 402256 224398 402284 231676
rect 402624 228449 402652 231676
rect 402992 229362 403020 231676
rect 403360 230382 403388 231676
rect 403348 230376 403400 230382
rect 403348 230318 403400 230324
rect 403072 230240 403124 230246
rect 403072 230182 403124 230188
rect 402980 229356 403032 229362
rect 402980 229298 403032 229304
rect 402980 228472 403032 228478
rect 402610 228440 402666 228449
rect 402980 228414 403032 228420
rect 402610 228375 402666 228384
rect 402244 224392 402296 224398
rect 402244 224334 402296 224340
rect 401876 224324 401928 224330
rect 401876 224266 401928 224272
rect 400954 221912 401010 221921
rect 400954 221847 401010 221856
rect 401140 221468 401192 221474
rect 401140 221410 401192 221416
rect 400680 219904 400732 219910
rect 400680 219846 400732 219852
rect 401152 217410 401180 221410
rect 401888 217410 401916 224266
rect 402992 217410 403020 228414
rect 403084 227866 403112 230182
rect 403072 227860 403124 227866
rect 403072 227802 403124 227808
rect 403636 225690 403664 231676
rect 404004 230246 404032 231676
rect 404386 231662 404676 231690
rect 404176 230376 404228 230382
rect 404176 230318 404228 230324
rect 403992 230240 404044 230246
rect 403992 230182 404044 230188
rect 403532 225684 403584 225690
rect 403532 225626 403584 225632
rect 403624 225684 403676 225690
rect 403624 225626 403676 225632
rect 403544 217410 403572 225626
rect 404188 221542 404216 230318
rect 404360 229628 404412 229634
rect 404360 229570 404412 229576
rect 404268 229356 404320 229362
rect 404268 229298 404320 229304
rect 404176 221536 404228 221542
rect 404176 221478 404228 221484
rect 404280 220114 404308 229298
rect 404372 228206 404400 229570
rect 404360 228200 404412 228206
rect 404360 228142 404412 228148
rect 404648 222970 404676 231662
rect 404740 229362 404768 231676
rect 405004 229492 405056 229498
rect 405004 229434 405056 229440
rect 404728 229356 404780 229362
rect 404728 229298 404780 229304
rect 404636 222964 404688 222970
rect 404636 222906 404688 222912
rect 405016 221513 405044 229434
rect 405108 229158 405136 231676
rect 405096 229152 405148 229158
rect 405096 229094 405148 229100
rect 405476 223718 405504 231676
rect 405844 230314 405872 231676
rect 406212 230382 406240 231676
rect 406304 231662 406502 231690
rect 406200 230376 406252 230382
rect 406200 230318 406252 230324
rect 405740 230308 405792 230314
rect 405740 230250 405792 230256
rect 405832 230308 405884 230314
rect 405832 230250 405884 230256
rect 405752 229498 405780 230250
rect 405740 229492 405792 229498
rect 405740 229434 405792 229440
rect 406108 227792 406160 227798
rect 406108 227734 406160 227740
rect 405924 224528 405976 224534
rect 405924 224470 405976 224476
rect 405464 223712 405516 223718
rect 405464 223654 405516 223660
rect 405002 221504 405058 221513
rect 405002 221439 405058 221448
rect 404452 220924 404504 220930
rect 404452 220866 404504 220872
rect 404268 220108 404320 220114
rect 404268 220050 404320 220056
rect 404464 217410 404492 220866
rect 405936 217410 405964 224470
rect 391032 217382 391368 217410
rect 391952 217382 392196 217410
rect 392596 217382 393024 217410
rect 393608 217382 393944 217410
rect 394712 217382 394772 217410
rect 395264 217382 395600 217410
rect 396184 217382 396428 217410
rect 396920 217382 397256 217410
rect 397748 217382 398084 217410
rect 398852 217382 398912 217410
rect 399404 217382 399832 217410
rect 400324 217382 400660 217410
rect 401152 217382 401488 217410
rect 401888 217382 402316 217410
rect 402992 217382 403144 217410
rect 403544 217382 403972 217410
rect 404464 217382 404800 217410
rect 405720 217382 405964 217410
rect 406120 217410 406148 227734
rect 406304 221474 406332 231662
rect 406856 230246 406884 231676
rect 407028 230376 407080 230382
rect 407028 230318 407080 230324
rect 406660 230240 406712 230246
rect 406660 230182 406712 230188
rect 406844 230240 406896 230246
rect 406844 230182 406896 230188
rect 406476 229968 406528 229974
rect 406476 229910 406528 229916
rect 406384 229764 406436 229770
rect 406384 229706 406436 229712
rect 406292 221468 406344 221474
rect 406292 221410 406344 221416
rect 406396 219638 406424 229706
rect 406488 228070 406516 229910
rect 406672 229770 406700 230182
rect 407040 230042 407068 230318
rect 406752 230036 406804 230042
rect 406752 229978 406804 229984
rect 407028 230036 407080 230042
rect 407028 229978 407080 229984
rect 406660 229764 406712 229770
rect 406660 229706 406712 229712
rect 406476 228064 406528 228070
rect 406476 228006 406528 228012
rect 406764 224534 406792 229978
rect 407224 229974 407252 231676
rect 407212 229968 407264 229974
rect 407212 229910 407264 229916
rect 407120 229832 407172 229838
rect 407120 229774 407172 229780
rect 407132 229634 407160 229774
rect 407120 229628 407172 229634
rect 407120 229570 407172 229576
rect 407120 225752 407172 225758
rect 407120 225694 407172 225700
rect 406752 224528 406804 224534
rect 406752 224470 406804 224476
rect 406384 219632 406436 219638
rect 406384 219574 406436 219580
rect 407132 217410 407160 225694
rect 407592 222902 407620 231676
rect 407764 229900 407816 229906
rect 407764 229842 407816 229848
rect 407776 229634 407804 229842
rect 407672 229628 407724 229634
rect 407672 229570 407724 229576
rect 407764 229628 407816 229634
rect 407764 229570 407816 229576
rect 407580 222896 407632 222902
rect 407580 222838 407632 222844
rect 407684 220930 407712 229570
rect 407960 226953 407988 231676
rect 408328 229770 408356 231676
rect 408316 229764 408368 229770
rect 408316 229706 408368 229712
rect 408408 229220 408460 229226
rect 408408 229162 408460 229168
rect 407946 226944 408002 226953
rect 407946 226879 408002 226888
rect 408420 225758 408448 229162
rect 408500 228404 408552 228410
rect 408500 228346 408552 228352
rect 408408 225752 408460 225758
rect 408408 225694 408460 225700
rect 407856 221060 407908 221066
rect 407856 221002 407908 221008
rect 407672 220924 407724 220930
rect 407672 220866 407724 220872
rect 407868 217410 407896 221002
rect 408512 219570 408540 228346
rect 408696 224330 408724 231676
rect 409064 230382 409092 231676
rect 409052 230376 409104 230382
rect 409052 230318 409104 230324
rect 409340 229226 409368 231676
rect 409604 230308 409656 230314
rect 409604 230250 409656 230256
rect 409328 229220 409380 229226
rect 409328 229162 409380 229168
rect 408684 224324 408736 224330
rect 408684 224266 408736 224272
rect 408592 224256 408644 224262
rect 409616 224233 409644 230250
rect 409708 227050 409736 231676
rect 409788 230308 409840 230314
rect 409788 230250 409840 230256
rect 409800 230042 409828 230250
rect 409788 230036 409840 230042
rect 409788 229978 409840 229984
rect 410076 229362 410104 231676
rect 410444 229838 410472 231676
rect 410432 229832 410484 229838
rect 410432 229774 410484 229780
rect 409788 229356 409840 229362
rect 409788 229298 409840 229304
rect 410064 229356 410116 229362
rect 410064 229298 410116 229304
rect 409800 228478 409828 229298
rect 409788 228472 409840 228478
rect 409788 228414 409840 228420
rect 410812 228410 410840 231676
rect 410996 231662 411194 231690
rect 410800 228404 410852 228410
rect 410800 228346 410852 228352
rect 409972 228132 410024 228138
rect 409972 228074 410024 228080
rect 409696 227044 409748 227050
rect 409696 226986 409748 226992
rect 408592 224198 408644 224204
rect 409602 224224 409658 224233
rect 408500 219564 408552 219570
rect 408500 219506 408552 219512
rect 408604 217410 408632 224198
rect 409602 224159 409658 224168
rect 409984 219774 410012 228074
rect 410248 225616 410300 225622
rect 410248 225558 410300 225564
rect 409880 219768 409932 219774
rect 409880 219710 409932 219716
rect 409972 219768 410024 219774
rect 409972 219710 410024 219716
rect 409892 217410 409920 219710
rect 406120 217382 406548 217410
rect 407132 217382 407376 217410
rect 407868 217382 408204 217410
rect 408604 217382 409032 217410
rect 409860 217382 409920 217410
rect 410260 217410 410288 225558
rect 410996 222873 411024 231662
rect 411168 230376 411220 230382
rect 411168 230318 411220 230324
rect 411352 230376 411404 230382
rect 411352 230318 411404 230324
rect 411076 230240 411128 230246
rect 411076 230182 411128 230188
rect 411088 225622 411116 230182
rect 411180 228313 411208 230318
rect 411260 230240 411312 230246
rect 411260 230182 411312 230188
rect 411272 229158 411300 230182
rect 411364 229974 411392 230318
rect 411352 229968 411404 229974
rect 411352 229910 411404 229916
rect 411548 229770 411576 231676
rect 411536 229764 411588 229770
rect 411536 229706 411588 229712
rect 411352 229288 411404 229294
rect 411352 229230 411404 229236
rect 411260 229152 411312 229158
rect 411260 229094 411312 229100
rect 411166 228304 411222 228313
rect 411166 228239 411222 228248
rect 411076 225616 411128 225622
rect 411076 225558 411128 225564
rect 411364 224262 411392 229230
rect 411916 229226 411944 231676
rect 423680 230648 423732 230654
rect 423680 230590 423732 230596
rect 416688 229560 416740 229566
rect 416688 229502 416740 229508
rect 411904 229220 411956 229226
rect 411904 229162 411956 229168
rect 414020 225276 414072 225282
rect 414020 225218 414072 225224
rect 412272 224324 412324 224330
rect 412272 224266 412324 224272
rect 411352 224256 411404 224262
rect 411352 224198 411404 224204
rect 411996 224188 412048 224194
rect 411996 224130 412048 224136
rect 410982 222864 411038 222873
rect 410982 222799 411038 222808
rect 411260 220992 411312 220998
rect 411260 220934 411312 220940
rect 411272 217410 411300 220934
rect 412008 217410 412036 224130
rect 412284 223718 412312 224266
rect 412272 223712 412324 223718
rect 412272 223654 412324 223660
rect 412916 219632 412968 219638
rect 412916 219574 412968 219580
rect 412928 217410 412956 219574
rect 414032 217410 414060 225218
rect 416700 223786 416728 229502
rect 420184 229220 420236 229226
rect 420184 229162 420236 229168
rect 420196 228138 420224 229162
rect 423692 229094 423720 230590
rect 507860 230580 507912 230586
rect 507860 230522 507912 230528
rect 456156 230444 456208 230450
rect 456156 230386 456208 230392
rect 428646 230344 428702 230353
rect 428646 230279 428702 230288
rect 423692 229066 423812 229094
rect 423036 228268 423088 228274
rect 423036 228210 423088 228216
rect 420184 228132 420236 228138
rect 420184 228074 420236 228080
rect 419540 227928 419592 227934
rect 419540 227870 419592 227876
rect 417056 223916 417108 223922
rect 417056 223858 417108 223864
rect 415492 223780 415544 223786
rect 415492 223722 415544 223728
rect 416688 223780 416740 223786
rect 416688 223722 416740 223728
rect 415308 222420 415360 222426
rect 415308 222362 415360 222368
rect 415320 220386 415348 222362
rect 415308 220380 415360 220386
rect 415308 220322 415360 220328
rect 414572 219564 414624 219570
rect 414572 219506 414624 219512
rect 414584 217410 414612 219506
rect 415504 217410 415532 223722
rect 416228 219768 416280 219774
rect 416228 219710 416280 219716
rect 416240 217410 416268 219710
rect 417068 217410 417096 223858
rect 418712 223848 418764 223854
rect 418712 223790 418764 223796
rect 418160 220380 418212 220386
rect 418160 220322 418212 220328
rect 418172 217410 418200 220322
rect 418724 217410 418752 223790
rect 419552 217410 419580 227870
rect 420368 225344 420420 225350
rect 420368 225286 420420 225292
rect 420380 217410 420408 225286
rect 422392 223984 422444 223990
rect 422392 223926 422444 223932
rect 421196 222488 421248 222494
rect 421196 222430 421248 222436
rect 421208 217410 421236 222430
rect 422404 217410 422432 223926
rect 423048 217410 423076 228210
rect 423784 217410 423812 229066
rect 426440 227996 426492 228002
rect 426440 227938 426492 227944
rect 425060 222556 425112 222562
rect 425060 222498 425112 222504
rect 425072 217410 425100 222498
rect 425520 221196 425572 221202
rect 425520 221138 425572 221144
rect 410260 217382 410688 217410
rect 411272 217382 411608 217410
rect 412008 217382 412436 217410
rect 412928 217382 413264 217410
rect 414032 217382 414092 217410
rect 414584 217382 414920 217410
rect 415504 217382 415748 217410
rect 416240 217382 416576 217410
rect 417068 217382 417496 217410
rect 418172 217382 418324 217410
rect 418724 217382 419152 217410
rect 419552 217382 419980 217410
rect 420380 217382 420808 217410
rect 421208 217382 421636 217410
rect 422404 217382 422464 217410
rect 423048 217382 423384 217410
rect 423784 217382 424212 217410
rect 425040 217382 425100 217410
rect 425532 217410 425560 221138
rect 426452 217410 426480 227938
rect 427084 226568 427136 226574
rect 427084 226510 427136 226516
rect 427096 217410 427124 226510
rect 428660 222630 428688 230279
rect 443644 230172 443696 230178
rect 443644 230114 443696 230120
rect 441712 229492 441764 229498
rect 441712 229434 441764 229440
rect 430764 229424 430816 229430
rect 430764 229366 430816 229372
rect 430776 229094 430804 229366
rect 435548 229356 435600 229362
rect 435548 229298 435600 229304
rect 430776 229066 431448 229094
rect 429660 227860 429712 227866
rect 429660 227802 429712 227808
rect 429292 222692 429344 222698
rect 429292 222634 429344 222640
rect 427912 222624 427964 222630
rect 427912 222566 427964 222572
rect 428648 222624 428700 222630
rect 428648 222566 428700 222572
rect 427924 217410 427952 222566
rect 429304 217410 429332 222634
rect 425532 217382 425868 217410
rect 426452 217382 426696 217410
rect 427096 217382 427524 217410
rect 427924 217382 428352 217410
rect 429272 217382 429332 217410
rect 429672 217410 429700 227802
rect 431420 223378 431448 229066
rect 433340 228336 433392 228342
rect 433340 228278 433392 228284
rect 431316 223372 431368 223378
rect 431316 223314 431368 223320
rect 431408 223372 431460 223378
rect 431408 223314 431460 223320
rect 430580 219360 430632 219366
rect 430580 219302 430632 219308
rect 430592 217410 430620 219302
rect 431328 217410 431356 223314
rect 432236 219428 432288 219434
rect 432236 219370 432288 219376
rect 432248 217410 432276 219370
rect 433352 217410 433380 228278
rect 433800 226636 433852 226642
rect 433800 226578 433852 226584
rect 433812 217410 433840 226578
rect 434720 225140 434772 225146
rect 434720 225082 434772 225088
rect 434732 217870 434760 225082
rect 435560 223242 435588 229298
rect 440608 226772 440660 226778
rect 440608 226714 440660 226720
rect 437480 226704 437532 226710
rect 437480 226646 437532 226652
rect 434812 223236 434864 223242
rect 434812 223178 434864 223184
rect 435548 223236 435600 223242
rect 435548 223178 435600 223184
rect 434720 217864 434772 217870
rect 434720 217806 434772 217812
rect 434824 217410 434852 223178
rect 436468 221060 436520 221066
rect 436468 221002 436520 221008
rect 435640 217864 435692 217870
rect 435640 217806 435692 217812
rect 435652 217410 435680 217806
rect 436480 217410 436508 221002
rect 437492 217410 437520 226646
rect 438860 225412 438912 225418
rect 438860 225354 438912 225360
rect 438032 222760 438084 222766
rect 438032 222702 438084 222708
rect 438044 217410 438072 222702
rect 438872 217410 438900 225354
rect 439780 221264 439832 221270
rect 439780 221206 439832 221212
rect 439792 217410 439820 221206
rect 440620 217410 440648 226714
rect 441724 226030 441752 229434
rect 441620 226024 441672 226030
rect 441620 225966 441672 225972
rect 441712 226024 441764 226030
rect 441712 225966 441764 225972
rect 441632 217870 441660 225966
rect 441712 222828 441764 222834
rect 441712 222770 441764 222776
rect 441620 217864 441672 217870
rect 441620 217806 441672 217812
rect 441724 217410 441752 222770
rect 443656 221270 443684 230114
rect 453304 229696 453356 229702
rect 453304 229638 453356 229644
rect 449164 229628 449216 229634
rect 449164 229570 449216 229576
rect 449176 227662 449204 229570
rect 447324 227656 447376 227662
rect 447324 227598 447376 227604
rect 449164 227656 449216 227662
rect 449164 227598 449216 227604
rect 444380 226840 444432 226846
rect 444380 226782 444432 226788
rect 443644 221264 443696 221270
rect 443644 221206 443696 221212
rect 443184 221128 443236 221134
rect 443184 221070 443236 221076
rect 442356 217864 442408 217870
rect 442356 217806 442408 217812
rect 442368 217410 442396 217806
rect 443196 217410 443224 221070
rect 444392 217410 444420 226782
rect 445760 225480 445812 225486
rect 445760 225422 445812 225428
rect 444748 223576 444800 223582
rect 444748 223518 444800 223524
rect 429672 217382 430100 217410
rect 430592 217382 430928 217410
rect 431328 217382 431756 217410
rect 432248 217382 432584 217410
rect 433352 217382 433412 217410
rect 433812 217382 434240 217410
rect 434824 217382 435160 217410
rect 435652 217382 435988 217410
rect 436480 217382 436816 217410
rect 437492 217382 437644 217410
rect 438044 217382 438472 217410
rect 438872 217382 439300 217410
rect 439792 217382 440128 217410
rect 440620 217382 441048 217410
rect 441724 217382 441876 217410
rect 442368 217382 442704 217410
rect 443196 217382 443532 217410
rect 444360 217382 444420 217410
rect 444760 217410 444788 223518
rect 445772 217410 445800 225422
rect 446588 221332 446640 221338
rect 446588 221274 446640 221280
rect 446600 217410 446628 221274
rect 447336 217410 447364 227598
rect 450636 226908 450688 226914
rect 450636 226850 450688 226856
rect 448980 225208 449032 225214
rect 448980 225150 449032 225156
rect 448612 223508 448664 223514
rect 448612 223450 448664 223456
rect 448624 217410 448652 223450
rect 444760 217382 445188 217410
rect 445772 217382 446016 217410
rect 446600 217382 446936 217410
rect 447336 217382 447764 217410
rect 448592 217382 448652 217410
rect 448992 217410 449020 225150
rect 449900 221400 449952 221406
rect 449900 221342 449952 221348
rect 449912 217410 449940 221342
rect 450648 217410 450676 226850
rect 452660 225548 452712 225554
rect 452660 225490 452712 225496
rect 451464 223440 451516 223446
rect 451464 223382 451516 223388
rect 451476 217410 451504 223382
rect 452672 217410 452700 225490
rect 453316 222154 453344 229638
rect 454040 228064 454092 228070
rect 454040 228006 454092 228012
rect 453212 222148 453264 222154
rect 453212 222090 453264 222096
rect 453304 222148 453356 222154
rect 453304 222090 453356 222096
rect 453224 217410 453252 222090
rect 454052 217870 454080 228006
rect 454132 226976 454184 226982
rect 454132 226918 454184 226924
rect 454040 217864 454092 217870
rect 454040 217806 454092 217812
rect 454144 217410 454172 226918
rect 456168 226302 456196 230386
rect 461584 230376 461636 230382
rect 461584 230318 461636 230324
rect 460940 229084 460992 229090
rect 460940 229026 460992 229032
rect 457352 227724 457404 227730
rect 457352 227666 457404 227672
rect 455696 226296 455748 226302
rect 455696 226238 455748 226244
rect 456156 226296 456208 226302
rect 456156 226238 456208 226244
rect 454960 217864 455012 217870
rect 454960 217806 455012 217812
rect 454972 217410 455000 217806
rect 455708 217410 455736 226238
rect 456800 222080 456852 222086
rect 456800 222022 456852 222028
rect 456812 217410 456840 222022
rect 457364 217410 457392 227666
rect 459560 226228 459612 226234
rect 459560 226170 459612 226176
rect 458364 221944 458416 221950
rect 458364 221886 458416 221892
rect 458376 217410 458404 221886
rect 459572 217410 459600 226170
rect 460020 222012 460072 222018
rect 460020 221954 460072 221960
rect 448992 217382 449420 217410
rect 449912 217382 450248 217410
rect 450648 217382 451076 217410
rect 451476 217382 451904 217410
rect 452672 217382 452824 217410
rect 453224 217382 453652 217410
rect 454144 217382 454480 217410
rect 454972 217382 455308 217410
rect 455708 217382 456136 217410
rect 456812 217382 456964 217410
rect 457364 217382 457792 217410
rect 458376 217382 458712 217410
rect 459540 217382 459600 217410
rect 460032 217410 460060 221954
rect 460952 217870 460980 229026
rect 461596 227594 461624 230318
rect 467104 230308 467156 230314
rect 467104 230250 467156 230256
rect 461216 227588 461268 227594
rect 461216 227530 461268 227536
rect 461584 227588 461636 227594
rect 461584 227530 461636 227536
rect 461228 219434 461256 227530
rect 464160 227520 464212 227526
rect 464160 227462 464212 227468
rect 462412 226160 462464 226166
rect 462412 226102 462464 226108
rect 461044 219406 461256 219434
rect 460940 217864 460992 217870
rect 460940 217806 460992 217812
rect 461044 217410 461072 219406
rect 461676 217864 461728 217870
rect 461676 217806 461728 217812
rect 461688 217410 461716 217806
rect 462424 217410 462452 226102
rect 463700 221876 463752 221882
rect 463700 221818 463752 221824
rect 463712 217410 463740 221818
rect 460032 217382 460368 217410
rect 461044 217382 461196 217410
rect 461688 217382 462024 217410
rect 462424 217382 462852 217410
rect 463680 217382 463740 217410
rect 464172 217410 464200 227462
rect 465080 226092 465132 226098
rect 465080 226034 465132 226040
rect 465092 217870 465120 226034
rect 465172 223780 465224 223786
rect 465172 223722 465224 223728
rect 465080 217864 465132 217870
rect 465080 217806 465132 217812
rect 465184 217410 465212 223722
rect 467116 221814 467144 230250
rect 468484 230240 468536 230246
rect 468484 230182 468536 230188
rect 478142 230208 478198 230217
rect 468496 227458 468524 230182
rect 478142 230143 478198 230152
rect 476120 228200 476172 228206
rect 476120 228142 476172 228148
rect 467840 227452 467892 227458
rect 467840 227394 467892 227400
rect 468484 227452 468536 227458
rect 468484 227394 468536 227400
rect 466736 221808 466788 221814
rect 466736 221750 466788 221756
rect 467104 221808 467156 221814
rect 467104 221750 467156 221756
rect 465908 217864 465960 217870
rect 465908 217806 465960 217812
rect 465920 217410 465948 217806
rect 466748 217410 466776 221750
rect 467852 217410 467880 227394
rect 470876 227384 470928 227390
rect 470876 227326 470928 227332
rect 469220 225956 469272 225962
rect 469220 225898 469272 225904
rect 468300 224052 468352 224058
rect 468300 223994 468352 224000
rect 468312 217410 468340 223994
rect 469232 217410 469260 225898
rect 470140 221740 470192 221746
rect 470140 221682 470192 221688
rect 470152 217410 470180 221682
rect 470888 217410 470916 227326
rect 474188 227316 474240 227322
rect 474188 227258 474240 227264
rect 471980 225888 472032 225894
rect 471980 225830 472032 225836
rect 471992 217870 472020 225830
rect 472072 224120 472124 224126
rect 472072 224062 472124 224068
rect 471980 217864 472032 217870
rect 471980 217806 472032 217812
rect 472084 217410 472112 224062
rect 473544 221672 473596 221678
rect 473544 221614 473596 221620
rect 472624 217864 472676 217870
rect 472624 217806 472676 217812
rect 472636 217410 472664 217806
rect 473556 217410 473584 221614
rect 474200 217410 474228 227258
rect 475016 224868 475068 224874
rect 475016 224810 475068 224816
rect 475028 217410 475056 224810
rect 476132 217870 476160 228142
rect 478156 227254 478184 230143
rect 486422 230072 486478 230081
rect 486422 230007 486478 230016
rect 480260 229016 480312 229022
rect 480260 228958 480312 228964
rect 477592 227248 477644 227254
rect 477592 227190 477644 227196
rect 478144 227248 478196 227254
rect 478144 227190 478196 227196
rect 476212 225820 476264 225826
rect 476212 225762 476264 225768
rect 476120 217864 476172 217870
rect 476120 217806 476172 217812
rect 476224 217410 476252 225762
rect 476856 217864 476908 217870
rect 476856 217806 476908 217812
rect 476868 217410 476896 217806
rect 477604 217410 477632 227190
rect 479248 224936 479300 224942
rect 479248 224878 479300 224884
rect 478972 224800 479024 224806
rect 478972 224742 479024 224748
rect 478984 217410 479012 224742
rect 464172 217382 464600 217410
rect 465184 217382 465428 217410
rect 465920 217382 466256 217410
rect 466748 217382 467084 217410
rect 467852 217382 467912 217410
rect 468312 217382 468740 217410
rect 469232 217382 469568 217410
rect 470152 217382 470488 217410
rect 470888 217382 471316 217410
rect 472084 217382 472144 217410
rect 472636 217382 472972 217410
rect 473556 217382 473800 217410
rect 474200 217382 474628 217410
rect 475028 217382 475456 217410
rect 476224 217382 476376 217410
rect 476868 217382 477204 217410
rect 477604 217382 478032 217410
rect 478860 217382 479012 217410
rect 479260 217410 479288 224878
rect 480272 217410 480300 228958
rect 483480 228948 483532 228954
rect 483480 228890 483532 228896
rect 480904 227180 480956 227186
rect 480904 227122 480956 227128
rect 480916 217410 480944 227122
rect 483112 227112 483164 227118
rect 483112 227054 483164 227060
rect 481824 224732 481876 224738
rect 481824 224674 481876 224680
rect 481836 217410 481864 224674
rect 483124 217410 483152 227054
rect 479260 217382 479688 217410
rect 480272 217382 480516 217410
rect 480916 217382 481344 217410
rect 481836 217382 482264 217410
rect 483092 217382 483152 217410
rect 483492 217410 483520 228890
rect 485136 228132 485188 228138
rect 485136 228074 485188 228080
rect 484400 219836 484452 219842
rect 484400 219778 484452 219784
rect 484412 217410 484440 219778
rect 485148 217410 485176 228074
rect 486436 218142 486464 230007
rect 493322 229936 493378 229945
rect 493322 229871 493378 229880
rect 493336 229094 493364 229871
rect 496082 229800 496138 229809
rect 496082 229735 496138 229744
rect 493336 229066 493456 229094
rect 487712 228880 487764 228886
rect 487712 228822 487764 228828
rect 486424 218136 486476 218142
rect 486424 218078 486476 218084
rect 486436 217410 486464 218078
rect 487528 218068 487580 218074
rect 487528 218010 487580 218016
rect 487540 217410 487568 218010
rect 483492 217382 483920 217410
rect 484412 217382 484748 217410
rect 485148 217382 485576 217410
rect 486404 217382 486464 217410
rect 487232 217382 487568 217410
rect 487724 217410 487752 228822
rect 491300 228812 491352 228818
rect 491300 228754 491352 228760
rect 489368 227248 489420 227254
rect 489368 227190 489420 227196
rect 487802 223408 487858 223417
rect 487802 223343 487858 223352
rect 487816 218414 487844 223343
rect 488540 222624 488592 222630
rect 488540 222566 488592 222572
rect 487804 218408 487856 218414
rect 487804 218350 487856 218356
rect 487816 218074 487844 218350
rect 487804 218068 487856 218074
rect 487804 218010 487856 218016
rect 488552 217410 488580 222566
rect 489380 218346 489408 227190
rect 490194 224632 490250 224641
rect 490194 224567 490250 224576
rect 489368 218340 489420 218346
rect 489368 218282 489420 218288
rect 489828 218340 489880 218346
rect 489828 218282 489880 218288
rect 489840 217410 489868 218282
rect 487724 217382 488152 217410
rect 488552 217396 488980 217410
rect 488552 217382 488994 217396
rect 489808 217382 489868 217410
rect 164884 217320 164936 217326
rect 164884 217262 164936 217268
rect 488966 216866 488994 217382
rect 489090 216880 489146 216889
rect 488966 216852 489090 216866
rect 488980 216838 489090 216852
rect 489090 216815 489146 216824
rect 490208 216458 490236 224567
rect 491312 217410 491340 228754
rect 491392 221264 491444 221270
rect 491392 221206 491444 221212
rect 491404 217870 491432 221206
rect 493428 218210 493456 229066
rect 494058 223272 494114 223281
rect 494058 223207 494114 223216
rect 493416 218204 493468 218210
rect 493416 218146 493468 218152
rect 491392 217864 491444 217870
rect 491392 217806 491444 217812
rect 492588 217864 492640 217870
rect 492588 217806 492640 217812
rect 492600 217410 492628 217806
rect 493428 217410 493456 218146
rect 491312 217382 491464 217410
rect 492292 217382 492628 217410
rect 493120 217382 493456 217410
rect 494072 216866 494100 223207
rect 495622 220552 495678 220561
rect 495622 220487 495678 220496
rect 494520 219292 494572 219298
rect 494520 219234 494572 219240
rect 494532 217410 494560 219234
rect 495636 217546 495664 220487
rect 496096 218142 496124 229735
rect 496910 227352 496966 227361
rect 496910 227287 496966 227296
rect 496084 218136 496136 218142
rect 496084 218078 496136 218084
rect 495636 217518 495710 217546
rect 494532 217382 494868 217410
rect 495682 216866 495710 217518
rect 496096 217410 496124 218078
rect 496924 217410 496952 227287
rect 502522 227216 502578 227225
rect 502522 227151 502578 227160
rect 499578 224496 499634 224505
rect 499578 224431 499634 224440
rect 498658 220416 498714 220425
rect 498658 220351 498714 220360
rect 498200 219224 498252 219230
rect 498200 219166 498252 219172
rect 498212 217410 498240 219166
rect 496096 217382 496524 217410
rect 496924 217382 497688 217410
rect 498180 217382 498240 217410
rect 498672 217410 498700 220351
rect 498672 217382 499160 217410
rect 499592 217394 499620 224431
rect 502432 220788 502484 220794
rect 502432 220730 502484 220736
rect 499670 220280 499726 220289
rect 499670 220215 499726 220224
rect 499684 218278 499712 220215
rect 502444 219570 502472 220730
rect 502432 219564 502484 219570
rect 502432 219506 502484 219512
rect 501236 219156 501288 219162
rect 501236 219098 501288 219104
rect 499672 218272 499724 218278
rect 499672 218214 499724 218220
rect 500224 218272 500276 218278
rect 500224 218214 500276 218220
rect 500236 217410 500264 218214
rect 501248 217410 501276 219098
rect 502444 217410 502472 219506
rect 497660 217258 497688 217382
rect 497648 217252 497700 217258
rect 497648 217194 497700 217200
rect 494040 216850 494376 216866
rect 495682 216852 496032 216866
rect 494040 216844 494388 216850
rect 494040 216838 494336 216844
rect 495696 216838 496032 216852
rect 494336 216786 494388 216792
rect 496004 216753 496032 216838
rect 499132 216782 499160 217382
rect 499580 217388 499632 217394
rect 499928 217382 500264 217410
rect 500756 217394 500908 217410
rect 500756 217388 500920 217394
rect 500756 217382 500868 217388
rect 499580 217330 499632 217336
rect 501248 217382 501584 217410
rect 502412 217382 502472 217410
rect 500868 217330 500920 217336
rect 502536 216918 502564 227151
rect 505374 224360 505430 224369
rect 505374 224295 505430 224304
rect 505008 220788 505060 220794
rect 505008 220730 505060 220736
rect 505020 220046 505048 220730
rect 505008 220040 505060 220046
rect 505008 219982 505060 219988
rect 503720 219088 503772 219094
rect 503720 219030 503772 219036
rect 503732 217410 503760 219030
rect 505020 217410 505048 219982
rect 503732 217382 504068 217410
rect 504896 217382 505048 217410
rect 505388 217410 505416 224295
rect 506480 224188 506532 224194
rect 506480 224130 506532 224136
rect 506492 217410 506520 224130
rect 507214 220144 507270 220153
rect 507214 220079 507270 220088
rect 507228 219473 507256 220079
rect 507214 219464 507270 219473
rect 507214 219399 507270 219408
rect 507228 217410 507256 219399
rect 507872 217410 507900 230522
rect 511264 230512 511316 230518
rect 511264 230454 511316 230460
rect 509884 219972 509936 219978
rect 509884 219914 509936 219920
rect 509896 219638 509924 219914
rect 509884 219632 509936 219638
rect 509884 219574 509936 219580
rect 508780 219020 508832 219026
rect 508780 218962 508832 218968
rect 508412 217796 508464 217802
rect 508412 217738 508464 217744
rect 508424 217410 508452 217738
rect 505388 217382 506152 217410
rect 506492 217382 506644 217410
rect 507228 217382 507472 217410
rect 507872 217382 508452 217410
rect 508792 217410 508820 218962
rect 509896 217410 509924 219574
rect 511276 218482 511304 230454
rect 515404 230104 515456 230110
rect 515404 230046 515456 230052
rect 513378 228712 513434 228721
rect 513378 228647 513434 228656
rect 512828 220652 512880 220658
rect 512828 220594 512880 220600
rect 512840 219706 512868 220594
rect 512828 219700 512880 219706
rect 512828 219642 512880 219648
rect 511356 218952 511408 218958
rect 511356 218894 511408 218900
rect 511264 218476 511316 218482
rect 511264 218418 511316 218424
rect 511276 217546 511304 218418
rect 511184 217518 511304 217546
rect 511184 217410 511212 217518
rect 508792 217382 509128 217410
rect 509896 217382 509956 217410
rect 510784 217382 511212 217410
rect 511368 217410 511396 218894
rect 512840 217410 512868 219642
rect 511368 217382 511704 217410
rect 512532 217382 512868 217410
rect 506124 216986 506152 217382
rect 513392 217002 513420 228647
rect 513840 219904 513892 219910
rect 513840 219846 513892 219852
rect 513852 217410 513880 219846
rect 515416 219774 515444 230046
rect 539600 230036 539652 230042
rect 539600 229978 539652 229984
rect 523040 228744 523092 228750
rect 523040 228686 523092 228692
rect 515494 227080 515550 227089
rect 515494 227015 515550 227024
rect 515404 219768 515456 219774
rect 515404 219710 515456 219716
rect 515416 217410 515444 219710
rect 515508 218550 515536 227015
rect 521658 225992 521714 226001
rect 521658 225927 521714 225936
rect 516232 224664 516284 224670
rect 516232 224606 516284 224612
rect 515496 218544 515548 218550
rect 515496 218486 515548 218492
rect 516048 218544 516100 218550
rect 516048 218486 516100 218492
rect 516060 217410 516088 218486
rect 513852 217382 514188 217410
rect 515016 217382 515444 217410
rect 515844 217382 516088 217410
rect 516244 217410 516272 224606
rect 518900 224596 518952 224602
rect 518900 224538 518952 224544
rect 518162 223136 518218 223145
rect 518162 223071 518218 223080
rect 517520 220720 517572 220726
rect 517520 220662 517572 220668
rect 517532 219910 517560 220662
rect 517520 219904 517572 219910
rect 517520 219846 517572 219852
rect 517532 217410 517560 219846
rect 518176 218618 518204 223071
rect 518164 218612 518216 218618
rect 518164 218554 518216 218560
rect 518440 218612 518492 218618
rect 518440 218554 518492 218560
rect 518452 217410 518480 218554
rect 516244 217382 516672 217410
rect 517532 217382 517592 217410
rect 518420 217382 518480 217410
rect 518912 217410 518940 224538
rect 520462 223000 520518 223009
rect 520462 222935 520518 222944
rect 520004 220584 520056 220590
rect 520004 220526 520056 220532
rect 520016 217410 520044 220526
rect 518912 217382 519248 217410
rect 520016 217382 520076 217410
rect 513656 217048 513708 217054
rect 513360 216996 513656 217002
rect 513360 216990 513708 216996
rect 506112 216980 506164 216986
rect 513360 216974 513696 216990
rect 506112 216922 506164 216928
rect 502524 216912 502576 216918
rect 503536 216912 503588 216918
rect 502524 216854 502576 216860
rect 503240 216860 503536 216866
rect 503240 216854 503588 216860
rect 503240 216838 503576 216854
rect 499120 216776 499172 216782
rect 495990 216744 496046 216753
rect 499120 216718 499172 216724
rect 495990 216679 496046 216688
rect 520476 216458 520504 222935
rect 521672 217410 521700 225927
rect 522580 220516 522632 220522
rect 522580 220458 522632 220464
rect 522592 217410 522620 220458
rect 523052 217938 523080 228686
rect 526352 228676 526404 228682
rect 526352 228618 526404 228624
rect 525064 223372 525116 223378
rect 525064 223314 525116 223320
rect 523132 223304 523184 223310
rect 523132 223246 523184 223252
rect 523040 217932 523092 217938
rect 523040 217874 523092 217880
rect 521672 217382 521732 217410
rect 522560 217382 522620 217410
rect 523144 216458 523172 223246
rect 525076 220726 525104 223314
rect 525890 221776 525946 221785
rect 525890 221711 525946 221720
rect 525064 220720 525116 220726
rect 525064 220662 525116 220668
rect 523960 217932 524012 217938
rect 523960 217874 524012 217880
rect 523972 217410 524000 217874
rect 525076 217410 525104 220662
rect 525904 217546 525932 221711
rect 525904 217518 525978 217546
rect 523972 217382 524308 217410
rect 525076 217382 525136 217410
rect 525950 216594 525978 217518
rect 526364 217410 526392 228618
rect 538220 228608 538272 228614
rect 538220 228550 538272 228556
rect 536840 228540 536892 228546
rect 536840 228482 536892 228488
rect 528926 225856 528982 225865
rect 528926 225791 528982 225800
rect 528098 221912 528154 221921
rect 528098 221847 528154 221856
rect 527272 220448 527324 220454
rect 527272 220390 527324 220396
rect 527284 217410 527312 220390
rect 528112 217410 528140 221847
rect 528940 217410 528968 225791
rect 531412 225752 531464 225758
rect 531412 225694 531464 225700
rect 534078 225720 534134 225729
rect 530584 223168 530636 223174
rect 530584 223110 530636 223116
rect 529940 219836 529992 219842
rect 529940 219778 529992 219784
rect 529952 219502 529980 219778
rect 529940 219496 529992 219502
rect 529940 219438 529992 219444
rect 529952 217410 529980 219438
rect 526364 217382 526792 217410
rect 527284 217382 527620 217410
rect 528112 217396 528448 217410
rect 528112 217382 528462 217396
rect 528940 217382 529368 217410
rect 529952 217382 530196 217410
rect 525950 216580 526300 216594
rect 525964 216566 526300 216580
rect 490208 216442 490972 216458
rect 520476 216442 521240 216458
rect 523144 216442 523816 216458
rect 526272 216442 526300 216566
rect 528434 216458 528462 217382
rect 530596 216458 530624 223110
rect 531424 217410 531452 225694
rect 534078 225655 534134 225664
rect 533068 223100 533120 223106
rect 533068 223042 533120 223048
rect 532700 220312 532752 220318
rect 532700 220254 532752 220260
rect 531424 217382 531852 217410
rect 532712 217138 532740 220254
rect 532680 217122 533016 217138
rect 532680 217116 533028 217122
rect 532680 217110 532976 217116
rect 532976 217058 533028 217064
rect 533080 216458 533108 223042
rect 534092 217410 534120 225655
rect 536010 221640 536066 221649
rect 536010 221575 536066 221584
rect 535368 220244 535420 220250
rect 535368 220186 535420 220192
rect 535380 217410 535408 220186
rect 534092 217382 534336 217410
rect 535256 217382 535408 217410
rect 536024 217410 536052 221575
rect 536852 217410 536880 228482
rect 537392 220176 537444 220182
rect 537392 220118 537444 220124
rect 537404 217410 537432 220118
rect 538232 217938 538260 228550
rect 539612 225758 539640 229978
rect 547144 229968 547196 229974
rect 547144 229910 547196 229916
rect 541530 228576 541586 228585
rect 541530 228511 541586 228520
rect 540428 226024 540480 226030
rect 540428 225966 540480 225972
rect 539600 225752 539652 225758
rect 539600 225694 539652 225700
rect 538312 223032 538364 223038
rect 538312 222974 538364 222980
rect 538220 217932 538272 217938
rect 538220 217874 538272 217880
rect 536024 217382 536420 217410
rect 536852 217382 536912 217410
rect 537404 217382 537892 217410
rect 528434 216444 528600 216458
rect 528448 216442 528600 216444
rect 530596 216442 531268 216458
rect 533080 216442 533844 216458
rect 536392 216442 536420 217382
rect 537864 217190 537892 217382
rect 537852 217184 537904 217190
rect 537852 217126 537904 217132
rect 538324 216458 538352 222974
rect 540440 219978 540468 225966
rect 541440 221604 541492 221610
rect 541440 221546 541492 221552
rect 540428 219972 540480 219978
rect 540428 219914 540480 219920
rect 539048 217932 539100 217938
rect 539048 217874 539100 217880
rect 539060 217410 539088 217874
rect 540440 217410 540468 219914
rect 541452 219026 541480 221546
rect 541440 219020 541492 219026
rect 541440 218962 541492 218968
rect 541452 217410 541480 218962
rect 539060 217382 539396 217410
rect 540224 217382 540468 217410
rect 541144 217382 541480 217410
rect 541544 217410 541572 228511
rect 543004 227656 543056 227662
rect 543004 227598 543056 227604
rect 543016 220046 543044 227598
rect 544014 225584 544070 225593
rect 544014 225519 544070 225528
rect 543188 224460 543240 224466
rect 543188 224402 543240 224408
rect 543004 220040 543056 220046
rect 543004 219982 543056 219988
rect 543016 217410 543044 219982
rect 543200 219094 543228 224402
rect 543188 219088 543240 219094
rect 543188 219030 543240 219036
rect 543648 219088 543700 219094
rect 543648 219030 543700 219036
rect 543660 217410 543688 219030
rect 541544 217382 541972 217410
rect 542800 217382 543044 217410
rect 543628 217382 543688 217410
rect 544028 217410 544056 225519
rect 545764 224528 545816 224534
rect 545764 224470 545816 224476
rect 545212 222148 545264 222154
rect 545212 222090 545264 222096
rect 545224 217530 545252 222090
rect 545776 219162 545804 224470
rect 547156 221610 547184 229910
rect 563704 229832 563756 229838
rect 563704 229774 563756 229780
rect 551284 229152 551336 229158
rect 551284 229094 551336 229100
rect 549258 228440 549314 228449
rect 549258 228375 549314 228384
rect 548156 226296 548208 226302
rect 548156 226238 548208 226244
rect 547144 221604 547196 221610
rect 547144 221546 547196 221552
rect 546682 221504 546738 221513
rect 546682 221439 546738 221448
rect 545764 219156 545816 219162
rect 545764 219098 545816 219104
rect 545212 217524 545264 217530
rect 545212 217466 545264 217472
rect 545224 217410 545252 217466
rect 545776 217410 545804 219098
rect 546696 217410 546724 221439
rect 548168 220182 548196 226238
rect 548248 224392 548300 224398
rect 548248 224334 548300 224340
rect 548156 220176 548208 220182
rect 548156 220118 548208 220124
rect 548168 217410 548196 220118
rect 544028 217382 544456 217410
rect 545224 217382 545284 217410
rect 545776 217382 546112 217410
rect 546696 217382 547032 217410
rect 547860 217382 548196 217410
rect 548260 216458 548288 224334
rect 549272 217410 549300 228375
rect 551296 221678 551324 229094
rect 553952 228472 554004 228478
rect 553952 228414 554004 228420
rect 552664 227588 552716 227594
rect 552664 227530 552716 227536
rect 552020 225684 552072 225690
rect 552020 225626 552072 225632
rect 551284 221672 551336 221678
rect 551284 221614 551336 221620
rect 551284 221536 551336 221542
rect 551284 221478 551336 221484
rect 551296 220114 551324 221478
rect 549996 220108 550048 220114
rect 549996 220050 550048 220056
rect 551284 220108 551336 220114
rect 551284 220050 551336 220056
rect 549272 217382 549516 217410
rect 550008 217274 550036 220050
rect 551296 217410 551324 220050
rect 552032 217410 552060 225626
rect 552676 220658 552704 227530
rect 553964 224954 553992 228414
rect 554964 227452 555016 227458
rect 554964 227394 555016 227400
rect 553964 224926 554176 224954
rect 553676 222964 553728 222970
rect 553676 222906 553728 222912
rect 552664 220652 552716 220658
rect 552664 220594 552716 220600
rect 551172 217382 551324 217410
rect 552000 217382 552060 217410
rect 552676 217410 552704 220594
rect 553688 218686 553716 222906
rect 553676 218680 553728 218686
rect 553676 218622 553728 218628
rect 553688 217410 553716 218622
rect 554148 217410 554176 224926
rect 554976 217410 555004 227394
rect 561678 226944 561734 226953
rect 561678 226879 561734 226888
rect 560300 225752 560352 225758
rect 560300 225694 560352 225700
rect 559196 225616 559248 225622
rect 559196 225558 559248 225564
rect 556160 224324 556212 224330
rect 556160 224266 556212 224272
rect 555700 217456 555752 217462
rect 552676 217382 552920 217410
rect 553688 217382 553748 217410
rect 554148 217382 554576 217410
rect 554976 217404 555700 217410
rect 554976 217398 555752 217404
rect 556172 217410 556200 224266
rect 556710 224224 556766 224233
rect 556710 224159 556766 224168
rect 556724 217410 556752 224159
rect 557816 221808 557868 221814
rect 557816 221750 557868 221756
rect 557828 217598 557856 221750
rect 558460 221468 558512 221474
rect 558460 221410 558512 221416
rect 558472 220862 558500 221410
rect 558460 220856 558512 220862
rect 558460 220798 558512 220804
rect 557816 217592 557868 217598
rect 557816 217534 557868 217540
rect 557828 217410 557856 217534
rect 558472 217410 558500 220798
rect 559208 217410 559236 225558
rect 560312 217666 560340 225694
rect 560944 222896 560996 222902
rect 560944 222838 560996 222844
rect 560576 220516 560628 220522
rect 560576 220458 560628 220464
rect 560588 220318 560616 220458
rect 560576 220312 560628 220318
rect 560576 220254 560628 220260
rect 560300 217660 560352 217666
rect 560300 217602 560352 217608
rect 560312 217410 560340 217602
rect 554976 217382 555740 217398
rect 556172 217382 556568 217410
rect 556724 217382 557060 217410
rect 557828 217382 557888 217410
rect 558472 217382 558808 217410
rect 559208 217382 559636 217410
rect 560312 217382 560464 217410
rect 550548 217320 550600 217326
rect 550008 217268 550548 217274
rect 550008 217262 550600 217268
rect 550008 217246 550588 217262
rect 538324 216442 538904 216458
rect 548260 216442 549024 216458
rect 556540 216442 556568 217382
rect 560956 216458 560984 222838
rect 561692 217410 561720 226879
rect 563612 224256 563664 224262
rect 563612 224198 563664 224204
rect 561772 221604 561824 221610
rect 561772 221546 561824 221552
rect 561784 217734 561812 221546
rect 563624 220998 563652 224198
rect 563612 220992 563664 220998
rect 563612 220934 563664 220940
rect 561772 217728 561824 217734
rect 561772 217670 561824 217676
rect 562876 217728 562928 217734
rect 562876 217670 562928 217676
rect 562888 217410 562916 217670
rect 563624 217410 563652 220934
rect 563716 220930 563744 229774
rect 564438 228304 564494 228313
rect 564438 228239 564494 228248
rect 563704 220924 563756 220930
rect 563704 220866 563756 220872
rect 564452 217410 564480 228239
rect 565096 221474 565124 245618
rect 570604 229764 570656 229770
rect 570604 229706 570656 229712
rect 569132 228404 569184 228410
rect 569132 228346 569184 228352
rect 565912 227044 565964 227050
rect 565912 226986 565964 226992
rect 565452 221672 565504 221678
rect 565452 221614 565504 221620
rect 565084 221468 565136 221474
rect 565084 221410 565136 221416
rect 565464 219502 565492 221614
rect 565452 219496 565504 219502
rect 565452 219438 565504 219444
rect 565464 217410 565492 219438
rect 565924 217410 565952 226986
rect 567200 223236 567252 223242
rect 567200 223178 567252 223184
rect 567212 217410 567240 223178
rect 569144 220998 569172 228346
rect 569314 222864 569370 222873
rect 569314 222799 569370 222808
rect 569132 220992 569184 220998
rect 569132 220934 569184 220940
rect 567936 220924 567988 220930
rect 567936 220866 567988 220872
rect 567948 219230 567976 220866
rect 567936 219224 567988 219230
rect 567936 219166 567988 219172
rect 561692 217382 562120 217410
rect 562888 217382 562948 217410
rect 563624 217382 563776 217410
rect 564452 217382 564696 217410
rect 565464 217382 565524 217410
rect 565924 217382 566688 217410
rect 567180 217382 567240 217410
rect 567948 217410 567976 219166
rect 569144 217410 569172 220934
rect 567948 217382 568008 217410
rect 568836 217382 569172 217410
rect 569328 217410 569356 222799
rect 570616 218958 570644 229706
rect 570604 218952 570656 218958
rect 570604 218894 570656 218900
rect 570616 217410 570644 218894
rect 571444 217410 571472 255274
rect 571536 229094 571564 258062
rect 571536 229066 571840 229094
rect 569328 217382 569664 217410
rect 570584 217382 570644 217410
rect 571412 217382 571472 217410
rect 571812 217410 571840 229066
rect 572732 217410 572760 262210
rect 574744 252612 574796 252618
rect 574744 252554 574796 252560
rect 574100 248464 574152 248470
rect 574100 248406 574152 248412
rect 574112 229094 574140 248406
rect 574112 229066 574324 229094
rect 573548 221468 573600 221474
rect 573548 221410 573600 221416
rect 573560 217410 573588 221410
rect 574192 220380 574244 220386
rect 574192 220322 574244 220328
rect 571812 217382 572240 217410
rect 572732 217382 573068 217410
rect 573560 217382 573896 217410
rect 566660 216714 566688 217382
rect 566648 216708 566700 216714
rect 566648 216650 566700 216656
rect 560956 216442 561628 216458
rect 574204 216442 574232 220322
rect 574296 217410 574324 229066
rect 574756 220590 574784 252554
rect 623044 242956 623096 242962
rect 623044 242898 623096 242904
rect 577504 232416 577556 232422
rect 577504 232358 577556 232364
rect 577228 220720 577280 220726
rect 577228 220662 577280 220668
rect 574744 220584 574796 220590
rect 574744 220526 574796 220532
rect 575480 220584 575532 220590
rect 575480 220526 575532 220532
rect 574836 219904 574888 219910
rect 574836 219846 574888 219852
rect 574296 217382 574724 217410
rect 574848 216442 574876 219846
rect 575492 217410 575520 220526
rect 576400 220516 576452 220522
rect 576400 220458 576452 220464
rect 577136 220516 577188 220522
rect 577136 220458 577188 220464
rect 576308 219156 576360 219162
rect 576308 219098 576360 219104
rect 576216 219088 576268 219094
rect 576216 219030 576268 219036
rect 576124 219020 576176 219026
rect 576124 218962 576176 218968
rect 576032 218680 576084 218686
rect 576032 218622 576084 218628
rect 575940 218612 575992 218618
rect 575940 218554 575992 218560
rect 575848 217796 575900 217802
rect 575848 217738 575900 217744
rect 575492 217382 575552 217410
rect 575756 217252 575808 217258
rect 575756 217194 575808 217200
rect 575664 216708 575716 216714
rect 575664 216650 575716 216656
rect 490208 216436 490984 216442
rect 490208 216430 490932 216436
rect 520476 216436 521252 216442
rect 520476 216430 521200 216436
rect 490932 216378 490984 216384
rect 523144 216436 523828 216442
rect 523144 216430 523776 216436
rect 521200 216378 521252 216384
rect 523776 216378 523828 216384
rect 526260 216436 526312 216442
rect 528448 216436 528612 216442
rect 528448 216430 528560 216436
rect 526260 216378 526312 216384
rect 530596 216436 531280 216442
rect 530596 216430 531228 216436
rect 528560 216378 528612 216384
rect 533080 216436 533856 216442
rect 533080 216430 533804 216436
rect 531228 216378 531280 216384
rect 533804 216378 533856 216384
rect 536380 216436 536432 216442
rect 538324 216436 538916 216442
rect 538324 216430 538864 216436
rect 536380 216378 536432 216384
rect 548260 216436 549036 216442
rect 548260 216430 548984 216436
rect 538864 216378 538916 216384
rect 548984 216378 549036 216384
rect 556528 216436 556580 216442
rect 560956 216436 561640 216442
rect 560956 216430 561588 216436
rect 556528 216378 556580 216384
rect 561588 216378 561640 216384
rect 574192 216436 574244 216442
rect 574192 216378 574244 216384
rect 574836 216436 574888 216442
rect 574836 216378 574888 216384
rect 575676 213314 575704 216650
rect 575768 213858 575796 217194
rect 575756 213852 575808 213858
rect 575756 213794 575808 213800
rect 575860 213790 575888 217738
rect 575848 213784 575900 213790
rect 575848 213726 575900 213732
rect 575952 213722 575980 218554
rect 575940 213716 575992 213722
rect 575940 213658 575992 213664
rect 576044 213382 576072 218622
rect 576136 213586 576164 218962
rect 576124 213580 576176 213586
rect 576124 213522 576176 213528
rect 576228 213518 576256 219030
rect 576216 213512 576268 213518
rect 576216 213454 576268 213460
rect 576320 213450 576348 219098
rect 576412 214674 576440 220458
rect 577044 219496 577096 219502
rect 577044 219438 577096 219444
rect 576952 217388 577004 217394
rect 576952 217330 577004 217336
rect 576400 214668 576452 214674
rect 576400 214610 576452 214616
rect 576964 213926 576992 217330
rect 577056 214606 577084 219438
rect 577148 214878 577176 220458
rect 577136 214872 577188 214878
rect 577136 214814 577188 214820
rect 577240 214742 577268 220662
rect 577228 214736 577280 214742
rect 577228 214678 577280 214684
rect 577044 214600 577096 214606
rect 577044 214542 577096 214548
rect 576952 213920 577004 213926
rect 576952 213862 577004 213868
rect 576308 213444 576360 213450
rect 576308 213386 576360 213392
rect 576032 213376 576084 213382
rect 576032 213318 576084 213324
rect 575664 213308 575716 213314
rect 575664 213250 575716 213256
rect 577516 213246 577544 232358
rect 604460 231736 604512 231742
rect 604460 231678 604512 231684
rect 604472 230518 604500 231678
rect 604460 230512 604512 230518
rect 604460 230454 604512 230460
rect 605748 230512 605800 230518
rect 605748 230454 605800 230460
rect 578882 216200 578938 216209
rect 578882 216135 578938 216144
rect 577872 216096 577924 216102
rect 577872 216038 577924 216044
rect 577884 213654 577912 216038
rect 577872 213648 577924 213654
rect 577872 213590 577924 213596
rect 577504 213240 577556 213246
rect 577504 213182 577556 213188
rect 578422 211712 578478 211721
rect 578422 211647 578478 211656
rect 578436 206990 578464 211647
rect 578514 210216 578570 210225
rect 578514 210151 578570 210160
rect 578424 206984 578476 206990
rect 578424 206926 578476 206932
rect 578528 205630 578556 210151
rect 578896 209710 578924 216135
rect 579066 214704 579122 214713
rect 579066 214639 579122 214648
rect 578974 213208 579030 213217
rect 578974 213143 579030 213152
rect 578884 209704 578936 209710
rect 578884 209646 578936 209652
rect 578988 208350 579016 213143
rect 579080 209778 579108 214639
rect 580264 209840 580316 209846
rect 580264 209782 580316 209788
rect 579068 209772 579120 209778
rect 579068 209714 579120 209720
rect 579526 208720 579582 208729
rect 579526 208655 579582 208664
rect 578976 208344 579028 208350
rect 578976 208286 579028 208292
rect 578790 207224 578846 207233
rect 578790 207159 578846 207168
rect 578516 205624 578568 205630
rect 578516 205566 578568 205572
rect 578804 204270 578832 207159
rect 579434 205728 579490 205737
rect 579434 205663 579490 205672
rect 578792 204264 578844 204270
rect 578792 204206 578844 204212
rect 578882 204232 578938 204241
rect 578882 204167 578938 204176
rect 578896 201414 578924 204167
rect 579448 202842 579476 205663
rect 579540 205562 579568 208655
rect 579528 205556 579580 205562
rect 579528 205498 579580 205504
rect 579436 202836 579488 202842
rect 579436 202778 579488 202784
rect 579250 202736 579306 202745
rect 579250 202671 579306 202680
rect 579264 201482 579292 202671
rect 579252 201476 579304 201482
rect 579252 201418 579304 201424
rect 578884 201408 578936 201414
rect 578884 201350 578936 201356
rect 578238 201240 578294 201249
rect 578238 201175 578294 201184
rect 578252 200122 578280 201175
rect 578240 200116 578292 200122
rect 578240 200058 578292 200064
rect 578422 199744 578478 199753
rect 578422 199679 578478 199688
rect 578436 198694 578464 199679
rect 578424 198688 578476 198694
rect 578424 198630 578476 198636
rect 579066 198248 579122 198257
rect 579066 198183 579122 198192
rect 579080 197334 579108 198183
rect 579068 197328 579120 197334
rect 579068 197270 579120 197276
rect 579526 196752 579582 196761
rect 579526 196687 579582 196696
rect 579540 196654 579568 196687
rect 579528 196648 579580 196654
rect 579528 196590 579580 196596
rect 579528 195288 579580 195294
rect 579526 195256 579528 195265
rect 579580 195256 579582 195265
rect 579526 195191 579582 195200
rect 579528 193860 579580 193866
rect 579528 193802 579580 193808
rect 579540 193633 579568 193802
rect 579526 193624 579582 193633
rect 579526 193559 579582 193568
rect 579528 192500 579580 192506
rect 579528 192442 579580 192448
rect 579540 192137 579568 192442
rect 579526 192128 579582 192137
rect 579526 192063 579582 192072
rect 579252 191888 579304 191894
rect 579252 191830 579304 191836
rect 579264 190641 579292 191830
rect 579250 190632 579306 190641
rect 579250 190567 579306 190576
rect 578240 190528 578292 190534
rect 578240 190470 578292 190476
rect 578252 189145 578280 190470
rect 579528 189168 579580 189174
rect 578238 189136 578294 189145
rect 579528 189110 579580 189116
rect 578238 189071 578294 189080
rect 579252 189100 579304 189106
rect 579252 189042 579304 189048
rect 578792 187740 578844 187746
rect 578792 187682 578844 187688
rect 578804 184657 578832 187682
rect 579264 187649 579292 189042
rect 579250 187640 579306 187649
rect 579250 187575 579306 187584
rect 579344 186380 579396 186386
rect 579344 186322 579396 186328
rect 578976 185020 579028 185026
rect 578976 184962 579028 184968
rect 578790 184648 578846 184657
rect 578790 184583 578846 184592
rect 578240 182232 578292 182238
rect 578240 182174 578292 182180
rect 578252 177177 578280 182174
rect 578332 180940 578384 180946
rect 578332 180882 578384 180888
rect 578238 177168 578294 177177
rect 578238 177103 578294 177112
rect 578344 175681 578372 180882
rect 578424 180872 578476 180878
rect 578424 180814 578476 180820
rect 578330 175672 578386 175681
rect 578330 175607 578386 175616
rect 578436 174185 578464 180814
rect 578988 180169 579016 184962
rect 579068 184952 579120 184958
rect 579068 184894 579120 184900
rect 579080 181665 579108 184894
rect 579252 183592 579304 183598
rect 579252 183534 579304 183540
rect 579066 181656 579122 181665
rect 579066 181591 579122 181600
rect 578974 180160 579030 180169
rect 578974 180095 579030 180104
rect 578792 179444 578844 179450
rect 578792 179386 578844 179392
rect 578700 178084 578752 178090
rect 578700 178026 578752 178032
rect 578422 174176 578478 174185
rect 578422 174111 578478 174120
rect 578712 171193 578740 178026
rect 578804 172689 578832 179386
rect 579264 178673 579292 183534
rect 579356 183161 579384 186322
rect 579540 186153 579568 189110
rect 579526 186144 579582 186153
rect 579526 186079 579582 186088
rect 579342 183152 579398 183161
rect 579342 183087 579398 183096
rect 579250 178664 579306 178673
rect 579250 178599 579306 178608
rect 579436 176792 579488 176798
rect 579436 176734 579488 176740
rect 579252 176724 579304 176730
rect 579252 176666 579304 176672
rect 578790 172680 578846 172689
rect 578790 172615 578846 172624
rect 579160 172576 579212 172582
rect 579160 172518 579212 172524
rect 578698 171184 578754 171193
rect 578698 171119 578754 171128
rect 578976 169856 579028 169862
rect 578976 169798 579028 169804
rect 578884 168428 578936 168434
rect 578884 168370 578936 168376
rect 578700 166728 578752 166734
rect 578700 166670 578752 166676
rect 578712 166569 578740 166670
rect 578698 166560 578754 166569
rect 578698 166495 578754 166504
rect 578240 164620 578292 164626
rect 578240 164562 578292 164568
rect 578252 164393 578280 164562
rect 578238 164384 578294 164393
rect 578238 164319 578294 164328
rect 578896 156097 578924 168370
rect 578988 157593 579016 169798
rect 579068 169788 579120 169794
rect 579068 169730 579120 169736
rect 579080 159089 579108 169730
rect 579172 162081 579200 172518
rect 579264 168065 579292 176666
rect 579344 171148 579396 171154
rect 579344 171090 579396 171096
rect 579250 168056 579306 168065
rect 579250 167991 579306 168000
rect 579158 162072 579214 162081
rect 579158 162007 579214 162016
rect 579356 160585 579384 171090
rect 579448 169561 579476 176734
rect 579434 169552 579490 169561
rect 579434 169487 579490 169496
rect 579528 164212 579580 164218
rect 579528 164154 579580 164160
rect 579540 163577 579568 164154
rect 579526 163568 579582 163577
rect 579526 163503 579582 163512
rect 579342 160576 579398 160585
rect 579342 160511 579398 160520
rect 579436 160132 579488 160138
rect 579436 160074 579488 160080
rect 579066 159080 579122 159089
rect 579066 159015 579122 159024
rect 579344 158772 579396 158778
rect 579344 158714 579396 158720
rect 578974 157584 579030 157593
rect 578974 157519 579030 157528
rect 578882 156088 578938 156097
rect 578882 156023 578938 156032
rect 578516 154692 578568 154698
rect 578516 154634 578568 154640
rect 578528 154601 578556 154634
rect 579160 154624 579212 154630
rect 578514 154592 578570 154601
rect 579160 154566 579212 154572
rect 578514 154527 578570 154536
rect 579068 153332 579120 153338
rect 579068 153274 579120 153280
rect 578976 153264 579028 153270
rect 578976 153206 579028 153212
rect 578884 150476 578936 150482
rect 578884 150418 578936 150424
rect 578516 148708 578568 148714
rect 578516 148650 578568 148656
rect 578528 148617 578556 148650
rect 578514 148608 578570 148617
rect 578514 148543 578570 148552
rect 578516 147348 578568 147354
rect 578516 147290 578568 147296
rect 578528 146985 578556 147290
rect 578514 146976 578570 146985
rect 578514 146911 578570 146920
rect 578608 144900 578660 144906
rect 578608 144842 578660 144848
rect 578620 143993 578648 144842
rect 578606 143984 578662 143993
rect 578606 143919 578662 143928
rect 578896 129033 578924 150418
rect 578988 132025 579016 153206
rect 579080 133521 579108 153274
rect 579172 135017 579200 154566
rect 579252 153128 579304 153134
rect 579250 153096 579252 153105
rect 579304 153096 579306 153105
rect 579250 153031 579306 153040
rect 579252 152992 579304 152998
rect 579252 152934 579304 152940
rect 579264 139505 579292 152934
rect 579356 141001 579384 158714
rect 579448 152998 579476 160074
rect 579436 152992 579488 152998
rect 579436 152934 579488 152940
rect 579528 151768 579580 151774
rect 579528 151710 579580 151716
rect 579540 151609 579568 151710
rect 579526 151600 579582 151609
rect 579526 151535 579582 151544
rect 579436 150272 579488 150278
rect 579436 150214 579488 150220
rect 579448 150113 579476 150214
rect 579434 150104 579490 150113
rect 579434 150039 579490 150048
rect 580276 147354 580304 209782
rect 603172 209772 603224 209778
rect 603172 209714 603224 209720
rect 603080 209704 603132 209710
rect 603080 209646 603132 209652
rect 603092 209545 603120 209646
rect 603078 209536 603134 209545
rect 603078 209471 603134 209480
rect 603184 208593 603212 209714
rect 603170 208584 603226 208593
rect 603170 208519 603226 208528
rect 603080 208344 603132 208350
rect 603080 208286 603132 208292
rect 603092 207505 603120 208286
rect 603078 207496 603134 207505
rect 603078 207431 603134 207440
rect 603080 206984 603132 206990
rect 603080 206926 603132 206932
rect 603092 206553 603120 206926
rect 603078 206544 603134 206553
rect 603078 206479 603134 206488
rect 603080 205624 603132 205630
rect 603080 205566 603132 205572
rect 603092 205465 603120 205566
rect 603172 205556 603224 205562
rect 603172 205498 603224 205504
rect 603078 205456 603134 205465
rect 603078 205391 603134 205400
rect 603184 204513 603212 205498
rect 603170 204504 603226 204513
rect 603170 204439 603226 204448
rect 603080 204264 603132 204270
rect 603080 204206 603132 204212
rect 603092 203425 603120 204206
rect 603078 203416 603134 203425
rect 603078 203351 603134 203360
rect 603080 202836 603132 202842
rect 603080 202778 603132 202784
rect 603092 202473 603120 202778
rect 603078 202464 603134 202473
rect 603078 202399 603134 202408
rect 603172 201476 603224 201482
rect 603172 201418 603224 201424
rect 603080 201408 603132 201414
rect 603078 201376 603080 201385
rect 603132 201376 603134 201385
rect 603078 201311 603134 201320
rect 603184 200433 603212 201418
rect 603170 200424 603226 200433
rect 603170 200359 603226 200368
rect 603080 200116 603132 200122
rect 603080 200058 603132 200064
rect 603092 199345 603120 200058
rect 603078 199336 603134 199345
rect 603078 199271 603134 199280
rect 603080 198688 603132 198694
rect 603080 198630 603132 198636
rect 603092 198393 603120 198630
rect 603078 198384 603134 198393
rect 603078 198319 603134 198328
rect 603172 197328 603224 197334
rect 603078 197296 603134 197305
rect 603172 197270 603224 197276
rect 603078 197231 603134 197240
rect 603092 196654 603120 197231
rect 603080 196648 603132 196654
rect 603080 196590 603132 196596
rect 603184 196353 603212 197270
rect 603170 196344 603226 196353
rect 603170 196279 603226 196288
rect 603080 195288 603132 195294
rect 603078 195256 603080 195265
rect 603132 195256 603134 195265
rect 603078 195191 603134 195200
rect 603078 194304 603134 194313
rect 603078 194239 603134 194248
rect 603092 193866 603120 194239
rect 603080 193860 603132 193866
rect 603080 193802 603132 193808
rect 603078 193216 603134 193225
rect 603078 193151 603134 193160
rect 603092 192506 603120 193151
rect 603080 192500 603132 192506
rect 603080 192442 603132 192448
rect 603078 192264 603134 192273
rect 603078 192199 603134 192208
rect 603092 191894 603120 192199
rect 603080 191888 603132 191894
rect 603080 191830 603132 191836
rect 603078 191176 603134 191185
rect 603078 191111 603134 191120
rect 603092 190534 603120 191111
rect 603080 190528 603132 190534
rect 603080 190470 603132 190476
rect 603170 190224 603226 190233
rect 603170 190159 603226 190168
rect 603080 189168 603132 189174
rect 603078 189136 603080 189145
rect 603132 189136 603134 189145
rect 603184 189106 603212 190159
rect 603078 189071 603134 189080
rect 603172 189100 603224 189106
rect 603172 189042 603224 189048
rect 603078 188184 603134 188193
rect 603078 188119 603134 188128
rect 603092 187746 603120 188119
rect 603080 187740 603132 187746
rect 603080 187682 603132 187688
rect 603078 187096 603134 187105
rect 603078 187031 603134 187040
rect 603092 186386 603120 187031
rect 603080 186380 603132 186386
rect 603080 186322 603132 186328
rect 603170 186144 603226 186153
rect 603170 186079 603226 186088
rect 603078 185056 603134 185065
rect 603078 184991 603080 185000
rect 603132 184991 603134 185000
rect 603080 184962 603132 184968
rect 603184 184958 603212 186079
rect 603172 184952 603224 184958
rect 603172 184894 603224 184900
rect 603078 184104 603134 184113
rect 603078 184039 603134 184048
rect 603092 183598 603120 184039
rect 603080 183592 603132 183598
rect 603080 183534 603132 183540
rect 603078 183016 603134 183025
rect 603078 182951 603134 182960
rect 603092 182238 603120 182951
rect 603080 182232 603132 182238
rect 603080 182174 603132 182180
rect 603170 182064 603226 182073
rect 603170 181999 603226 182008
rect 603078 180976 603134 180985
rect 603184 180946 603212 181999
rect 603078 180911 603134 180920
rect 603172 180940 603224 180946
rect 603092 180878 603120 180911
rect 603172 180882 603224 180888
rect 603080 180872 603132 180878
rect 603080 180814 603132 180820
rect 603078 180024 603134 180033
rect 603078 179959 603134 179968
rect 603092 179450 603120 179959
rect 603080 179444 603132 179450
rect 603080 179386 603132 179392
rect 603078 178936 603134 178945
rect 603078 178871 603134 178880
rect 603092 178090 603120 178871
rect 603080 178084 603132 178090
rect 603080 178026 603132 178032
rect 603170 177984 603226 177993
rect 603170 177919 603226 177928
rect 603078 176896 603134 176905
rect 603078 176831 603134 176840
rect 603092 176730 603120 176831
rect 603184 176798 603212 177919
rect 603172 176792 603224 176798
rect 603172 176734 603224 176740
rect 603080 176724 603132 176730
rect 603080 176666 603132 176672
rect 603078 175944 603134 175953
rect 603078 175879 603134 175888
rect 603092 175302 603120 175879
rect 581644 175296 581696 175302
rect 581644 175238 581696 175244
rect 603080 175296 603132 175302
rect 603080 175238 603132 175244
rect 580356 173936 580408 173942
rect 580356 173878 580408 173884
rect 580368 164626 580396 173878
rect 581656 166734 581684 175238
rect 603078 174856 603134 174865
rect 603078 174791 603134 174800
rect 603092 173942 603120 174791
rect 603080 173936 603132 173942
rect 603080 173878 603132 173884
rect 603722 173904 603778 173913
rect 603722 173839 603778 173848
rect 603078 172816 603134 172825
rect 603078 172751 603134 172760
rect 603092 172582 603120 172751
rect 603080 172576 603132 172582
rect 603080 172518 603132 172524
rect 603078 171864 603134 171873
rect 603078 171799 603134 171808
rect 603092 171154 603120 171799
rect 603080 171148 603132 171154
rect 603080 171090 603132 171096
rect 603170 170776 603226 170785
rect 603170 170711 603226 170720
rect 603080 169856 603132 169862
rect 603078 169824 603080 169833
rect 603132 169824 603134 169833
rect 603184 169794 603212 170711
rect 603078 169759 603134 169768
rect 603172 169788 603224 169794
rect 603172 169730 603224 169736
rect 603078 168736 603134 168745
rect 603078 168671 603134 168680
rect 603092 168434 603120 168671
rect 603080 168428 603132 168434
rect 603080 168370 603132 168376
rect 603078 167784 603134 167793
rect 603078 167719 603134 167728
rect 603092 167074 603120 167719
rect 583116 167068 583168 167074
rect 583116 167010 583168 167016
rect 603080 167068 603132 167074
rect 603080 167010 603132 167016
rect 581644 166728 581696 166734
rect 581644 166670 581696 166676
rect 581736 165640 581788 165646
rect 581736 165582 581788 165588
rect 580356 164620 580408 164626
rect 580356 164562 580408 164568
rect 581644 164280 581696 164286
rect 581644 164222 581696 164228
rect 580356 162920 580408 162926
rect 580356 162862 580408 162868
rect 580368 148714 580396 162862
rect 581656 150278 581684 164222
rect 581748 153134 581776 165582
rect 583024 161492 583076 161498
rect 583024 161434 583076 161440
rect 581736 153128 581788 153134
rect 581736 153070 581788 153076
rect 581644 150272 581696 150278
rect 581644 150214 581696 150220
rect 580356 148708 580408 148714
rect 580356 148650 580408 148656
rect 580264 147348 580316 147354
rect 580264 147290 580316 147296
rect 583036 146130 583064 161434
rect 583128 154698 583156 167010
rect 603078 166696 603134 166705
rect 603078 166631 603134 166640
rect 603092 165646 603120 166631
rect 603080 165640 603132 165646
rect 603080 165582 603132 165588
rect 603078 164656 603134 164665
rect 603078 164591 603134 164600
rect 603092 164286 603120 164591
rect 603080 164280 603132 164286
rect 603080 164222 603132 164228
rect 603736 164218 603764 173839
rect 603814 165744 603870 165753
rect 603814 165679 603870 165688
rect 603724 164212 603776 164218
rect 603724 164154 603776 164160
rect 603078 163704 603134 163713
rect 603078 163639 603134 163648
rect 603092 162926 603120 163639
rect 603080 162920 603132 162926
rect 603080 162862 603132 162868
rect 603078 162616 603134 162625
rect 603078 162551 603134 162560
rect 603092 161498 603120 162551
rect 603722 161664 603778 161673
rect 603722 161599 603778 161608
rect 603080 161492 603132 161498
rect 603080 161434 603132 161440
rect 603078 160576 603134 160585
rect 603078 160511 603134 160520
rect 603092 160138 603120 160511
rect 603080 160132 603132 160138
rect 603080 160074 603132 160080
rect 603078 159624 603134 159633
rect 603078 159559 603134 159568
rect 603092 158778 603120 159559
rect 603080 158772 603132 158778
rect 603080 158714 603132 158720
rect 603170 158536 603226 158545
rect 603170 158471 603226 158480
rect 603078 157584 603134 157593
rect 603078 157519 603134 157528
rect 603092 157486 603120 157519
rect 585876 157480 585928 157486
rect 585876 157422 585928 157428
rect 603080 157480 603132 157486
rect 603080 157422 603132 157428
rect 584404 157412 584456 157418
rect 584404 157354 584456 157360
rect 583116 154692 583168 154698
rect 583116 154634 583168 154640
rect 579528 146124 579580 146130
rect 579528 146066 579580 146072
rect 583024 146124 583076 146130
rect 583024 146066 583076 146072
rect 579540 145489 579568 146066
rect 579526 145480 579582 145489
rect 579526 145415 579582 145424
rect 583116 144968 583168 144974
rect 583116 144910 583168 144916
rect 580356 143608 580408 143614
rect 580356 143550 580408 143556
rect 579528 142656 579580 142662
rect 579528 142598 579580 142604
rect 579540 142497 579568 142598
rect 579526 142488 579582 142497
rect 579526 142423 579582 142432
rect 579342 140992 579398 141001
rect 579342 140927 579398 140936
rect 579250 139496 579306 139505
rect 579250 139431 579306 139440
rect 579526 138000 579582 138009
rect 579526 137935 579528 137944
rect 579580 137935 579582 137944
rect 579528 137906 579580 137912
rect 579528 136536 579580 136542
rect 579526 136504 579528 136513
rect 579580 136504 579582 136513
rect 579526 136439 579582 136448
rect 579158 135008 579214 135017
rect 579158 134943 579214 134952
rect 580264 133952 580316 133958
rect 580264 133894 580316 133900
rect 579066 133512 579122 133521
rect 579066 133447 579122 133456
rect 578974 132016 579030 132025
rect 578974 131951 579030 131960
rect 579252 131096 579304 131102
rect 579252 131038 579304 131044
rect 579264 130529 579292 131038
rect 579250 130520 579306 130529
rect 579250 130455 579306 130464
rect 578882 129024 578938 129033
rect 578882 128959 578938 128968
rect 578884 128308 578936 128314
rect 578884 128250 578936 128256
rect 578896 127537 578924 128250
rect 578882 127528 578938 127537
rect 578882 127463 578938 127472
rect 579068 126948 579120 126954
rect 579068 126890 579120 126896
rect 579080 126041 579108 126890
rect 579066 126032 579122 126041
rect 579066 125967 579122 125976
rect 578424 125588 578476 125594
rect 578424 125530 578476 125536
rect 578436 124545 578464 125530
rect 578422 124536 578478 124545
rect 578422 124471 578478 124480
rect 579252 124160 579304 124166
rect 579252 124102 579304 124108
rect 579264 122913 579292 124102
rect 579250 122904 579306 122913
rect 579250 122839 579306 122848
rect 579528 121440 579580 121446
rect 579526 121408 579528 121417
rect 579580 121408 579582 121417
rect 579526 121343 579582 121352
rect 579252 120080 579304 120086
rect 579252 120022 579304 120028
rect 579264 119921 579292 120022
rect 579250 119912 579306 119921
rect 579250 119847 579306 119856
rect 579160 118720 579212 118726
rect 579160 118662 579212 118668
rect 578608 118448 578660 118454
rect 578606 118416 578608 118425
rect 578660 118416 578662 118425
rect 578606 118351 578662 118360
rect 579068 117360 579120 117366
rect 579068 117302 579120 117308
rect 578976 114572 579028 114578
rect 578976 114514 579028 114520
rect 578884 113212 578936 113218
rect 578884 113154 578936 113160
rect 578424 112668 578476 112674
rect 578424 112610 578476 112616
rect 578436 112441 578464 112610
rect 578422 112432 578478 112441
rect 578422 112367 578478 112376
rect 578700 111784 578752 111790
rect 578700 111726 578752 111732
rect 578712 110945 578740 111726
rect 578698 110936 578754 110945
rect 578698 110871 578754 110880
rect 578516 103488 578568 103494
rect 578514 103456 578516 103465
rect 578568 103456 578570 103465
rect 578514 103391 578570 103400
rect 578332 102128 578384 102134
rect 578332 102070 578384 102076
rect 578344 101969 578372 102070
rect 578330 101960 578386 101969
rect 578330 101895 578386 101904
rect 578700 100700 578752 100706
rect 578700 100642 578752 100648
rect 578712 100337 578740 100642
rect 578698 100328 578754 100337
rect 578698 100263 578754 100272
rect 578608 96620 578660 96626
rect 578608 96562 578660 96568
rect 578620 95849 578648 96562
rect 578606 95840 578662 95849
rect 578606 95775 578662 95784
rect 578700 95192 578752 95198
rect 578700 95134 578752 95140
rect 578712 94353 578740 95134
rect 578698 94344 578754 94353
rect 578698 94279 578754 94288
rect 578516 81388 578568 81394
rect 578516 81330 578568 81336
rect 578528 80889 578556 81330
rect 578514 80880 578570 80889
rect 578514 80815 578570 80824
rect 576124 77308 576176 77314
rect 576124 77250 576176 77256
rect 52276 53168 52328 53174
rect 52276 53110 52328 53116
rect 346308 53168 346360 53174
rect 346308 53110 346360 53116
rect 145380 53100 145432 53106
rect 145380 53042 145432 53048
rect 84824 52686 85160 52714
rect 52184 51740 52236 51746
rect 52184 51682 52236 51688
rect 60740 51740 60792 51746
rect 60740 51682 60792 51688
rect 60752 51066 60780 51682
rect 60740 51060 60792 51066
rect 60740 51002 60792 51008
rect 85132 50289 85160 52686
rect 145392 50810 145420 53042
rect 150328 52822 150388 52850
rect 150360 51066 150388 52822
rect 346320 52714 346348 53110
rect 215832 52686 216168 52714
rect 281336 52686 281488 52714
rect 346320 52686 347176 52714
rect 412344 52686 412496 52714
rect 477848 52686 478184 52714
rect 189078 51776 189134 51785
rect 189078 51711 189134 51720
rect 189092 51066 189120 51711
rect 150348 51060 150400 51066
rect 150348 51002 150400 51008
rect 189080 51060 189132 51066
rect 189080 51002 189132 51008
rect 145084 50782 145420 50810
rect 216140 50425 216168 52686
rect 281460 50561 281488 52686
rect 347148 52426 347176 52686
rect 347136 52420 347188 52426
rect 347136 52362 347188 52368
rect 281446 50552 281502 50561
rect 281446 50487 281502 50496
rect 216126 50416 216182 50425
rect 216126 50351 216182 50360
rect 85118 50280 85174 50289
rect 85118 50215 85174 50224
rect 142356 44305 142384 46716
rect 412468 46617 412496 52686
rect 478156 49774 478184 52686
rect 543016 52686 543352 52714
rect 543016 50289 543044 52686
rect 543002 50280 543058 50289
rect 543002 50215 543058 50224
rect 478144 49768 478196 49774
rect 478144 49710 478196 49716
rect 478788 49768 478840 49774
rect 478788 49710 478840 49716
rect 412454 46608 412510 46617
rect 412454 46543 412510 46552
rect 473174 46336 473230 46345
rect 473174 46271 473230 46280
rect 470138 46200 470194 46209
rect 470138 46135 470194 46144
rect 419722 45520 419778 45529
rect 419722 45455 419778 45464
rect 415398 45384 415454 45393
rect 415398 45319 415454 45328
rect 241520 45008 241572 45014
rect 241518 44976 241520 44985
rect 246120 45008 246172 45014
rect 241572 44976 241574 44985
rect 241518 44911 241574 44920
rect 246118 44976 246120 44985
rect 246172 44976 246174 44985
rect 246118 44911 246174 44920
rect 251086 44976 251142 44985
rect 251086 44911 251088 44920
rect 251140 44911 251142 44920
rect 255870 44976 255926 44985
rect 255870 44911 255872 44920
rect 251088 44882 251140 44888
rect 255924 44911 255926 44920
rect 255872 44882 255924 44888
rect 241520 44872 241572 44878
rect 241518 44840 241520 44849
rect 246120 44872 246172 44878
rect 241572 44840 241574 44849
rect 241518 44775 241574 44784
rect 246118 44840 246120 44849
rect 405556 44872 405608 44878
rect 246172 44840 246174 44849
rect 246118 44775 246174 44784
rect 251086 44840 251142 44849
rect 251086 44775 251088 44784
rect 251140 44775 251142 44784
rect 255870 44840 255926 44849
rect 405556 44814 405608 44820
rect 255870 44775 255872 44784
rect 251088 44746 251140 44752
rect 255924 44775 255926 44784
rect 255872 44746 255924 44752
rect 142342 44296 142398 44305
rect 142342 44231 142398 44240
rect 361762 43616 361818 43625
rect 361762 43551 361818 43560
rect 307298 43480 307354 43489
rect 307298 43415 307354 43424
rect 187514 42120 187570 42129
rect 187358 42078 187514 42106
rect 194322 42120 194378 42129
rect 194074 42078 194322 42106
rect 187514 42055 187570 42064
rect 307312 42106 307340 43415
rect 310104 42392 310160 42401
rect 310104 42327 310160 42336
rect 307004 42078 307340 42106
rect 310118 42092 310146 42327
rect 361776 42092 361804 43551
rect 365074 42120 365130 42129
rect 364918 42078 365074 42106
rect 194322 42055 194378 42064
rect 405568 42092 405596 44814
rect 415412 42364 415440 45319
rect 419736 42772 419764 45455
rect 365074 42055 365130 42064
rect 416686 41848 416742 41857
rect 416622 41806 416686 41834
rect 460570 41848 460626 41857
rect 460368 41806 460570 41834
rect 416686 41783 416742 41792
rect 470152 41820 470180 46135
rect 473188 42534 473216 46271
rect 478800 44713 478828 49710
rect 576136 44985 576164 77250
rect 578896 73273 578924 113154
rect 578988 76265 579016 114514
rect 579080 79393 579108 117302
rect 579172 82385 579200 118662
rect 579528 117292 579580 117298
rect 579528 117234 579580 117240
rect 579540 116929 579568 117234
rect 579526 116920 579582 116929
rect 579526 116855 579582 116864
rect 579528 115592 579580 115598
rect 579528 115534 579580 115540
rect 579540 115433 579568 115534
rect 579526 115424 579582 115433
rect 579526 115359 579582 115368
rect 579252 114504 579304 114510
rect 579252 114446 579304 114452
rect 579264 113937 579292 114446
rect 579250 113928 579306 113937
rect 579250 113863 579306 113872
rect 579436 109608 579488 109614
rect 579436 109550 579488 109556
rect 579448 109449 579476 109550
rect 579434 109440 579490 109449
rect 579434 109375 579490 109384
rect 579252 108792 579304 108798
rect 579252 108734 579304 108740
rect 579264 107953 579292 108734
rect 579250 107944 579306 107953
rect 579250 107879 579306 107888
rect 579528 107636 579580 107642
rect 579528 107578 579580 107584
rect 579540 106457 579568 107578
rect 579526 106448 579582 106457
rect 579526 106383 579582 106392
rect 579528 106276 579580 106282
rect 579528 106218 579580 106224
rect 579540 104961 579568 106218
rect 579526 104952 579582 104961
rect 579526 104887 579582 104896
rect 580276 103494 580304 133894
rect 580368 118454 580396 143550
rect 583024 138032 583076 138038
rect 583024 137974 583076 137980
rect 581644 136672 581696 136678
rect 581644 136614 581696 136620
rect 580356 118448 580408 118454
rect 580356 118390 580408 118396
rect 581656 108798 581684 136614
rect 581736 129056 581788 129062
rect 581736 128998 581788 129004
rect 581748 120086 581776 128998
rect 581736 120080 581788 120086
rect 581736 120022 581788 120028
rect 583036 109614 583064 137974
rect 583128 121446 583156 144910
rect 584416 142662 584444 157354
rect 584588 147688 584640 147694
rect 584588 147630 584640 147636
rect 584404 142656 584456 142662
rect 584404 142598 584456 142604
rect 584404 139460 584456 139466
rect 584404 139402 584456 139408
rect 583116 121440 583168 121446
rect 583116 121382 583168 121388
rect 584416 112674 584444 139402
rect 584600 128314 584628 147630
rect 585784 142180 585836 142186
rect 585784 142122 585836 142128
rect 584588 128308 584640 128314
rect 584588 128250 584640 128256
rect 584496 127016 584548 127022
rect 584496 126958 584548 126964
rect 584404 112668 584456 112674
rect 584404 112610 584456 112616
rect 583116 112464 583168 112470
rect 583116 112406 583168 112412
rect 583024 109608 583076 109614
rect 583024 109550 583076 109556
rect 581644 108792 581696 108798
rect 581644 108734 581696 108740
rect 581736 107704 581788 107710
rect 581736 107646 581788 107652
rect 580264 103488 580316 103494
rect 580264 103430 580316 103436
rect 581644 102196 581696 102202
rect 581644 102138 581696 102144
rect 580264 100768 580316 100774
rect 580264 100710 580316 100716
rect 579528 98932 579580 98938
rect 579528 98874 579580 98880
rect 579540 98841 579568 98874
rect 579526 98832 579582 98841
rect 579526 98767 579582 98776
rect 579528 97640 579580 97646
rect 579528 97582 579580 97588
rect 579540 97345 579568 97582
rect 579526 97336 579582 97345
rect 579526 97271 579582 97280
rect 579528 93832 579580 93838
rect 579528 93774 579580 93780
rect 579540 92857 579568 93774
rect 579526 92848 579582 92857
rect 579526 92783 579582 92792
rect 579528 92472 579580 92478
rect 579528 92414 579580 92420
rect 579540 91361 579568 92414
rect 579526 91352 579582 91361
rect 579526 91287 579582 91296
rect 579528 91044 579580 91050
rect 579528 90986 579580 90992
rect 579540 89865 579568 90986
rect 579526 89856 579582 89865
rect 579526 89791 579582 89800
rect 579528 89684 579580 89690
rect 579528 89626 579580 89632
rect 579540 88369 579568 89626
rect 579526 88360 579582 88369
rect 579526 88295 579582 88304
rect 579528 86964 579580 86970
rect 579528 86906 579580 86912
rect 579540 86873 579568 86906
rect 579526 86864 579582 86873
rect 579526 86799 579582 86808
rect 579528 85536 579580 85542
rect 579528 85478 579580 85484
rect 579540 85377 579568 85478
rect 579526 85368 579582 85377
rect 579526 85303 579582 85312
rect 579528 84176 579580 84182
rect 579528 84118 579580 84124
rect 579540 83881 579568 84118
rect 579526 83872 579582 83881
rect 579526 83807 579582 83816
rect 579158 82376 579214 82385
rect 579158 82311 579214 82320
rect 579066 79384 579122 79393
rect 579066 79319 579122 79328
rect 579528 78668 579580 78674
rect 579528 78610 579580 78616
rect 579540 77897 579568 78610
rect 579526 77888 579582 77897
rect 579526 77823 579582 77832
rect 579068 77376 579120 77382
rect 579068 77318 579120 77324
rect 578974 76256 579030 76265
rect 578974 76191 579030 76200
rect 578882 73264 578938 73273
rect 578882 73199 578938 73208
rect 578332 68944 578384 68950
rect 578332 68886 578384 68892
rect 578344 68785 578372 68886
rect 578330 68776 578386 68785
rect 578330 68711 578386 68720
rect 578700 61396 578752 61402
rect 578700 61338 578752 61344
rect 578712 61305 578740 61338
rect 578698 61296 578754 61305
rect 578698 61231 578754 61240
rect 578976 60716 579028 60722
rect 578976 60658 579028 60664
rect 578988 59809 579016 60658
rect 578974 59800 579030 59809
rect 578974 59735 579030 59744
rect 578884 58812 578936 58818
rect 578884 58754 578936 58760
rect 578896 58313 578924 58754
rect 578882 58304 578938 58313
rect 578882 58239 578938 58248
rect 578884 57928 578936 57934
rect 578884 57870 578936 57876
rect 578332 57248 578384 57254
rect 578332 57190 578384 57196
rect 578240 55684 578292 55690
rect 578240 55626 578292 55632
rect 578252 55321 578280 55626
rect 578238 55312 578294 55321
rect 578238 55247 578294 55256
rect 578344 53825 578372 57190
rect 578896 56817 578924 57870
rect 578882 56808 578938 56817
rect 578882 56743 578938 56752
rect 578330 53816 578386 53825
rect 578330 53751 578386 53760
rect 579080 53106 579108 77318
rect 579528 75880 579580 75886
rect 579528 75822 579580 75828
rect 579540 74769 579568 75822
rect 579526 74760 579582 74769
rect 579526 74695 579582 74704
rect 579526 71768 579582 71777
rect 579526 71703 579528 71712
rect 579580 71703 579582 71712
rect 579528 71674 579580 71680
rect 579528 70372 579580 70378
rect 579528 70314 579580 70320
rect 579540 70281 579568 70314
rect 579526 70272 579582 70281
rect 579526 70207 579582 70216
rect 579528 67584 579580 67590
rect 579528 67526 579580 67532
rect 579540 67289 579568 67526
rect 579526 67280 579582 67289
rect 579526 67215 579582 67224
rect 579252 65816 579304 65822
rect 579250 65784 579252 65793
rect 579304 65784 579306 65793
rect 579250 65719 579306 65728
rect 579528 64320 579580 64326
rect 579526 64288 579528 64297
rect 579580 64288 579582 64297
rect 579526 64223 579582 64232
rect 579528 63504 579580 63510
rect 579528 63446 579580 63452
rect 579540 62801 579568 63446
rect 579526 62792 579582 62801
rect 579526 62727 579582 62736
rect 580276 55690 580304 100710
rect 580356 98660 580408 98666
rect 580356 98602 580408 98608
rect 580368 68950 580396 98602
rect 580356 68944 580408 68950
rect 580356 68886 580408 68892
rect 581656 57934 581684 102138
rect 581748 65822 581776 107646
rect 583024 102264 583076 102270
rect 583024 102206 583076 102212
rect 581736 65816 581788 65822
rect 581736 65758 581788 65764
rect 583036 58818 583064 102206
rect 583128 97646 583156 112406
rect 584404 104916 584456 104922
rect 584404 104858 584456 104864
rect 583116 97640 583168 97646
rect 583116 97582 583168 97588
rect 584416 61402 584444 104858
rect 584508 95198 584536 126958
rect 585796 115598 585824 142122
rect 585888 136542 585916 157422
rect 603184 157418 603212 158471
rect 603172 157412 603224 157418
rect 603172 157354 603224 157360
rect 603078 156496 603134 156505
rect 603078 156431 603134 156440
rect 603092 155990 603120 156431
rect 587256 155984 587308 155990
rect 587256 155926 587308 155932
rect 603080 155984 603132 155990
rect 603080 155926 603132 155932
rect 587164 151836 587216 151842
rect 587164 151778 587216 151784
rect 585876 136536 585928 136542
rect 585876 136478 585928 136484
rect 587176 131102 587204 151778
rect 587268 137970 587296 155926
rect 603078 155544 603134 155553
rect 603078 155479 603134 155488
rect 603092 154630 603120 155479
rect 603080 154624 603132 154630
rect 603080 154566 603132 154572
rect 603170 154456 603226 154465
rect 603170 154391 603226 154400
rect 603078 153504 603134 153513
rect 603078 153439 603134 153448
rect 603092 153270 603120 153439
rect 603184 153338 603212 154391
rect 603172 153332 603224 153338
rect 603172 153274 603224 153280
rect 603080 153264 603132 153270
rect 603080 153206 603132 153212
rect 603078 152416 603134 152425
rect 603078 152351 603134 152360
rect 603092 151842 603120 152351
rect 603080 151836 603132 151842
rect 603080 151778 603132 151784
rect 603078 151464 603134 151473
rect 603078 151399 603134 151408
rect 603092 150482 603120 151399
rect 603080 150476 603132 150482
rect 603080 150418 603132 150424
rect 603170 150376 603226 150385
rect 603170 150311 603226 150320
rect 603078 149424 603134 149433
rect 603078 149359 603134 149368
rect 603092 149190 603120 149359
rect 592776 149184 592828 149190
rect 592776 149126 592828 149132
rect 603080 149184 603132 149190
rect 603080 149126 603132 149132
rect 589924 149116 589976 149122
rect 589924 149058 589976 149064
rect 588544 146328 588596 146334
rect 588544 146270 588596 146276
rect 587256 137964 587308 137970
rect 587256 137906 587308 137912
rect 587348 135312 587400 135318
rect 587348 135254 587400 135260
rect 587164 131096 587216 131102
rect 587164 131038 587216 131044
rect 585876 129804 585928 129810
rect 585876 129746 585928 129752
rect 585784 115592 585836 115598
rect 585784 115534 585836 115540
rect 585784 106344 585836 106350
rect 585784 106286 585836 106292
rect 584496 95192 584548 95198
rect 584496 95134 584548 95140
rect 585796 64326 585824 106286
rect 585888 98938 585916 129746
rect 587256 121508 587308 121514
rect 587256 121450 587308 121456
rect 587164 109064 587216 109070
rect 587164 109006 587216 109012
rect 585876 98932 585928 98938
rect 585876 98874 585928 98880
rect 587176 67590 587204 109006
rect 587268 85542 587296 121450
rect 587360 107642 587388 135254
rect 588556 124166 588584 146270
rect 588636 131776 588688 131782
rect 588636 131718 588688 131724
rect 588544 124160 588596 124166
rect 588544 124102 588596 124108
rect 588544 120148 588596 120154
rect 588544 120090 588596 120096
rect 587348 107636 587400 107642
rect 587348 107578 587400 107584
rect 587256 85536 587308 85542
rect 587256 85478 587308 85484
rect 588556 84182 588584 120090
rect 588648 106282 588676 131718
rect 589936 125594 589964 149058
rect 591304 140820 591356 140826
rect 591304 140762 591356 140768
rect 590016 132524 590068 132530
rect 590016 132466 590068 132472
rect 589924 125588 589976 125594
rect 589924 125530 589976 125536
rect 589924 122868 589976 122874
rect 589924 122810 589976 122816
rect 588636 106276 588688 106282
rect 588636 106218 588688 106224
rect 589936 86970 589964 122810
rect 590028 102134 590056 132466
rect 591316 114510 591344 140762
rect 592788 126954 592816 149126
rect 603184 149122 603212 150311
rect 603172 149116 603224 149122
rect 603172 149058 603224 149064
rect 603078 148336 603134 148345
rect 603078 148271 603134 148280
rect 603092 147694 603120 148271
rect 603080 147688 603132 147694
rect 603080 147630 603132 147636
rect 603078 147384 603134 147393
rect 603078 147319 603134 147328
rect 603092 146334 603120 147319
rect 603080 146328 603132 146334
rect 603080 146270 603132 146276
rect 603170 146296 603226 146305
rect 603170 146231 603226 146240
rect 603184 144974 603212 146231
rect 603172 144968 603224 144974
rect 603172 144910 603224 144916
rect 603736 144906 603764 161599
rect 603828 151774 603856 165679
rect 603816 151768 603868 151774
rect 603816 151710 603868 151716
rect 603906 145344 603962 145353
rect 603906 145279 603962 145288
rect 603724 144900 603776 144906
rect 603724 144842 603776 144848
rect 603078 144256 603134 144265
rect 603078 144191 603134 144200
rect 603092 143614 603120 144191
rect 603080 143608 603132 143614
rect 603080 143550 603132 143556
rect 603722 143304 603778 143313
rect 603722 143239 603778 143248
rect 603078 142216 603134 142225
rect 603078 142151 603080 142160
rect 603132 142151 603134 142160
rect 603080 142122 603132 142128
rect 603078 141264 603134 141273
rect 603078 141199 603134 141208
rect 603092 140826 603120 141199
rect 603080 140820 603132 140826
rect 603080 140762 603132 140768
rect 603078 140176 603134 140185
rect 603078 140111 603134 140120
rect 603092 139466 603120 140111
rect 603080 139460 603132 139466
rect 603080 139402 603132 139408
rect 603170 139224 603226 139233
rect 603170 139159 603226 139168
rect 603078 138136 603134 138145
rect 598296 138100 598348 138106
rect 603184 138106 603212 139159
rect 603078 138071 603134 138080
rect 603172 138100 603224 138106
rect 598296 138042 598348 138048
rect 596916 131164 596968 131170
rect 596916 131106 596968 131112
rect 594064 128376 594116 128382
rect 594064 128318 594116 128324
rect 592776 126948 592828 126954
rect 592776 126890 592828 126896
rect 592684 125656 592736 125662
rect 592684 125598 592736 125604
rect 591396 124228 591448 124234
rect 591396 124170 591448 124176
rect 591304 114504 591356 114510
rect 591304 114446 591356 114452
rect 590016 102128 590068 102134
rect 590016 102070 590068 102076
rect 591304 99408 591356 99414
rect 591304 99350 591356 99356
rect 589924 86964 589976 86970
rect 589924 86906 589976 86912
rect 588544 84176 588596 84182
rect 588544 84118 588596 84124
rect 587164 67584 587216 67590
rect 587164 67526 587216 67532
rect 585784 64320 585836 64326
rect 585784 64262 585836 64268
rect 584404 61396 584456 61402
rect 584404 61338 584456 61344
rect 583024 58812 583076 58818
rect 583024 58754 583076 58760
rect 581644 57928 581696 57934
rect 581644 57870 581696 57876
rect 591316 57254 591344 99350
rect 591408 91050 591436 124170
rect 592696 93838 592724 125598
rect 594076 96626 594104 128318
rect 595444 110492 595496 110498
rect 595444 110434 595496 110440
rect 594064 96620 594116 96626
rect 594064 96562 594116 96568
rect 592684 93832 592736 93838
rect 592684 93774 592736 93780
rect 591396 91044 591448 91050
rect 591396 90986 591448 90992
rect 595456 70378 595484 110434
rect 596824 103964 596876 103970
rect 596824 103906 596876 103912
rect 595444 70372 595496 70378
rect 595444 70314 595496 70320
rect 596836 63510 596864 103906
rect 596928 100706 596956 131106
rect 598204 111852 598256 111858
rect 598204 111794 598256 111800
rect 596916 100700 596968 100706
rect 596916 100642 596968 100648
rect 598216 71738 598244 111794
rect 598308 111790 598336 138042
rect 603092 138038 603120 138071
rect 603172 138042 603224 138048
rect 603080 138032 603132 138038
rect 603080 137974 603132 137980
rect 603078 137184 603134 137193
rect 603078 137119 603134 137128
rect 603092 136678 603120 137119
rect 603080 136672 603132 136678
rect 603080 136614 603132 136620
rect 603078 136096 603134 136105
rect 603078 136031 603134 136040
rect 603092 135318 603120 136031
rect 603080 135312 603132 135318
rect 603080 135254 603132 135260
rect 603170 135144 603226 135153
rect 603170 135079 603226 135088
rect 603078 134056 603134 134065
rect 603078 133991 603134 134000
rect 603092 133958 603120 133991
rect 603080 133952 603132 133958
rect 603080 133894 603132 133900
rect 603078 133104 603134 133113
rect 603078 133039 603134 133048
rect 603092 132530 603120 133039
rect 603080 132524 603132 132530
rect 603080 132466 603132 132472
rect 603078 132016 603134 132025
rect 603078 131951 603134 131960
rect 603092 131170 603120 131951
rect 603184 131782 603212 135079
rect 603172 131776 603224 131782
rect 603172 131718 603224 131724
rect 603080 131164 603132 131170
rect 603080 131106 603132 131112
rect 603078 131064 603134 131073
rect 603078 130999 603134 131008
rect 603092 129810 603120 130999
rect 603080 129804 603132 129810
rect 603080 129746 603132 129752
rect 603078 129024 603134 129033
rect 603078 128959 603134 128968
rect 603092 128382 603120 128959
rect 603080 128376 603132 128382
rect 603080 128318 603132 128324
rect 603078 127936 603134 127945
rect 603078 127871 603134 127880
rect 603092 127022 603120 127871
rect 603080 127016 603132 127022
rect 603080 126958 603132 126964
rect 603170 126984 603226 126993
rect 603170 126919 603226 126928
rect 603078 125896 603134 125905
rect 603078 125831 603134 125840
rect 603092 125730 603120 125831
rect 601056 125724 601108 125730
rect 601056 125666 601108 125672
rect 603080 125724 603132 125730
rect 603080 125666 603132 125672
rect 600964 116000 601016 116006
rect 600964 115942 601016 115948
rect 599584 114640 599636 114646
rect 599584 114582 599636 114588
rect 598296 111784 598348 111790
rect 598296 111726 598348 111732
rect 599596 75886 599624 114582
rect 600976 78674 601004 115942
rect 601068 92478 601096 125666
rect 603184 125662 603212 126919
rect 603172 125656 603224 125662
rect 603172 125598 603224 125604
rect 603078 124944 603134 124953
rect 603078 124879 603134 124888
rect 603092 124234 603120 124879
rect 603080 124228 603132 124234
rect 603080 124170 603132 124176
rect 602434 123856 602490 123865
rect 602434 123791 602490 123800
rect 602342 118824 602398 118833
rect 602342 118759 602398 118768
rect 601056 92472 601108 92478
rect 601056 92414 601108 92420
rect 602356 81394 602384 118759
rect 602448 89690 602476 123791
rect 603078 122904 603134 122913
rect 603078 122839 603080 122848
rect 603132 122839 603134 122848
rect 603080 122810 603132 122816
rect 603078 121816 603134 121825
rect 603078 121751 603134 121760
rect 603092 121514 603120 121751
rect 603080 121508 603132 121514
rect 603080 121450 603132 121456
rect 603078 120864 603134 120873
rect 603078 120799 603134 120808
rect 603092 120154 603120 120799
rect 603080 120148 603132 120154
rect 603080 120090 603132 120096
rect 603078 119776 603134 119785
rect 603078 119711 603134 119720
rect 603092 118726 603120 119711
rect 603080 118720 603132 118726
rect 603080 118662 603132 118668
rect 603078 117736 603134 117745
rect 603078 117671 603134 117680
rect 603092 117366 603120 117671
rect 603080 117360 603132 117366
rect 603080 117302 603132 117308
rect 603736 117298 603764 143239
rect 603814 129976 603870 129985
rect 603814 129911 603870 129920
rect 603724 117292 603776 117298
rect 603724 117234 603776 117240
rect 603446 116784 603502 116793
rect 603446 116719 603502 116728
rect 603460 116006 603488 116719
rect 603448 116000 603500 116006
rect 603448 115942 603500 115948
rect 603078 115696 603134 115705
rect 603078 115631 603134 115640
rect 603092 114578 603120 115631
rect 603170 114744 603226 114753
rect 603170 114679 603226 114688
rect 603184 114646 603212 114679
rect 603172 114640 603224 114646
rect 603172 114582 603224 114588
rect 603080 114572 603132 114578
rect 603080 114514 603132 114520
rect 603078 113656 603134 113665
rect 603078 113591 603134 113600
rect 603092 113218 603120 113591
rect 603080 113212 603132 113218
rect 603080 113154 603132 113160
rect 603078 112704 603134 112713
rect 603078 112639 603134 112648
rect 603092 111858 603120 112639
rect 603828 112470 603856 129911
rect 603920 129062 603948 145279
rect 603908 129056 603960 129062
rect 603908 128998 603960 129004
rect 603816 112464 603868 112470
rect 603816 112406 603868 112412
rect 603080 111852 603132 111858
rect 603080 111794 603132 111800
rect 603078 111616 603134 111625
rect 603078 111551 603134 111560
rect 603092 110498 603120 111551
rect 603814 110664 603870 110673
rect 603814 110599 603870 110608
rect 603080 110492 603132 110498
rect 603080 110434 603132 110440
rect 603078 109576 603134 109585
rect 603078 109511 603134 109520
rect 603092 109070 603120 109511
rect 603080 109064 603132 109070
rect 603080 109006 603132 109012
rect 603078 108624 603134 108633
rect 603078 108559 603134 108568
rect 603092 107710 603120 108559
rect 603080 107704 603132 107710
rect 603080 107646 603132 107652
rect 603078 107536 603134 107545
rect 603078 107471 603134 107480
rect 603092 106350 603120 107471
rect 603170 106584 603226 106593
rect 603170 106519 603226 106528
rect 603080 106344 603132 106350
rect 603080 106286 603132 106292
rect 603078 105496 603134 105505
rect 603078 105431 603134 105440
rect 603092 104922 603120 105431
rect 603080 104916 603132 104922
rect 603080 104858 603132 104864
rect 603184 103970 603212 106519
rect 603722 104544 603778 104553
rect 603722 104479 603778 104488
rect 603172 103964 603224 103970
rect 603172 103906 603224 103912
rect 603170 103456 603226 103465
rect 603170 103391 603226 103400
rect 603078 102504 603134 102513
rect 603078 102439 603134 102448
rect 603092 102202 603120 102439
rect 603184 102270 603212 103391
rect 603172 102264 603224 102270
rect 603172 102206 603224 102212
rect 603080 102196 603132 102202
rect 603080 102138 603132 102144
rect 603078 101416 603134 101425
rect 603078 101351 603134 101360
rect 603092 100774 603120 101351
rect 603080 100768 603132 100774
rect 603080 100710 603132 100716
rect 603078 100464 603134 100473
rect 603078 100399 603134 100408
rect 603092 99414 603120 100399
rect 603080 99408 603132 99414
rect 603080 99350 603132 99356
rect 602436 89684 602488 89690
rect 602436 89626 602488 89632
rect 602344 81388 602396 81394
rect 602344 81330 602396 81336
rect 600964 78668 601016 78674
rect 600964 78610 601016 78616
rect 599584 75880 599636 75886
rect 599584 75822 599636 75828
rect 598204 71732 598256 71738
rect 598204 71674 598256 71680
rect 596824 63504 596876 63510
rect 596824 63446 596876 63452
rect 603736 60722 603764 104479
rect 603828 98666 603856 110599
rect 603816 98660 603868 98666
rect 603816 98602 603868 98608
rect 605760 77994 605788 230454
rect 621204 220992 621256 220998
rect 621204 220934 621256 220940
rect 619824 220924 619876 220930
rect 619824 220866 619876 220872
rect 618812 220856 618864 220862
rect 618812 220798 618864 220804
rect 605932 220244 605984 220250
rect 605932 220186 605984 220192
rect 605944 216102 605972 220186
rect 615500 220176 615552 220182
rect 615500 220118 615552 220124
rect 609612 220108 609664 220114
rect 609612 220050 609664 220056
rect 608416 218544 608468 218550
rect 608416 218486 608468 218492
rect 606668 218408 606720 218414
rect 606668 218350 606720 218356
rect 605932 216096 605984 216102
rect 605932 216038 605984 216044
rect 606680 210202 606708 218350
rect 607496 216980 607548 216986
rect 607496 216922 607548 216928
rect 607128 215348 607180 215354
rect 607128 215290 607180 215296
rect 607140 210202 607168 215290
rect 607508 213178 607536 216922
rect 607588 216844 607640 216850
rect 607588 216786 607640 216792
rect 607496 213172 607548 213178
rect 607496 213114 607548 213120
rect 607600 210202 607628 216786
rect 608048 213852 608100 213858
rect 608048 213794 608100 213800
rect 608060 210202 608088 213794
rect 608428 213110 608456 218486
rect 608508 216912 608560 216918
rect 608508 216854 608560 216860
rect 608520 214010 608548 216854
rect 608520 213982 608640 214010
rect 608508 213920 608560 213926
rect 608508 213862 608560 213868
rect 608416 213104 608468 213110
rect 608416 213046 608468 213052
rect 608520 210202 608548 213862
rect 606648 210174 606708 210202
rect 607108 210174 607168 210202
rect 607568 210174 607628 210202
rect 608028 210174 608088 210202
rect 608488 210174 608548 210202
rect 608612 210066 608640 213982
rect 609624 213858 609652 220050
rect 614120 220040 614172 220046
rect 614120 219982 614172 219988
rect 613384 219972 613436 219978
rect 613384 219914 613436 219920
rect 612004 219836 612056 219842
rect 612004 219778 612056 219784
rect 609888 218476 609940 218482
rect 609888 218418 609940 218424
rect 609900 213874 609928 218418
rect 610808 217048 610860 217054
rect 610808 216990 610860 216996
rect 610346 216880 610402 216889
rect 610346 216815 610402 216824
rect 609612 213852 609664 213858
rect 609900 213846 610020 213874
rect 609612 213794 609664 213800
rect 609888 213784 609940 213790
rect 609888 213726 609940 213732
rect 609428 213172 609480 213178
rect 609428 213114 609480 213120
rect 609440 210202 609468 213114
rect 609900 210202 609928 213726
rect 609408 210174 609468 210202
rect 609868 210174 609928 210202
rect 609992 210066 610020 213846
rect 610360 213790 610388 216815
rect 610348 213784 610400 213790
rect 610348 213726 610400 213732
rect 610820 210202 610848 216990
rect 612016 216374 612044 219778
rect 613396 216442 613424 219914
rect 613384 216436 613436 216442
rect 613384 216378 613436 216384
rect 612004 216368 612056 216374
rect 612004 216310 612056 216316
rect 614132 216306 614160 219982
rect 615512 216510 615540 220118
rect 616788 219224 616840 219230
rect 616788 219166 616840 219172
rect 615500 216504 615552 216510
rect 615500 216446 615552 216452
rect 614120 216300 614172 216306
rect 614120 216242 614172 216248
rect 615500 215892 615552 215898
rect 615500 215834 615552 215840
rect 615040 215824 615092 215830
rect 615040 215766 615092 215772
rect 614580 215756 614632 215762
rect 614580 215698 614632 215704
rect 614028 215688 614080 215694
rect 614028 215630 614080 215636
rect 613568 215620 613620 215626
rect 613568 215562 613620 215568
rect 613108 215552 613160 215558
rect 613108 215494 613160 215500
rect 612648 215484 612700 215490
rect 612648 215426 612700 215432
rect 612188 215416 612240 215422
rect 612188 215358 612240 215364
rect 611728 213716 611780 213722
rect 611728 213658 611780 213664
rect 611268 213104 611320 213110
rect 611268 213046 611320 213052
rect 611280 210202 611308 213046
rect 611740 210202 611768 213658
rect 612200 210202 612228 215358
rect 612660 210202 612688 215426
rect 613120 210202 613148 215494
rect 613580 210202 613608 215562
rect 614040 210202 614068 215630
rect 614592 210202 614620 215698
rect 615052 210202 615080 215766
rect 615512 210202 615540 215834
rect 615960 213580 616012 213586
rect 615960 213522 616012 213528
rect 615972 210202 616000 213522
rect 616800 213518 616828 219166
rect 617524 218952 617576 218958
rect 617524 218894 617576 218900
rect 617340 213648 617392 213654
rect 617340 213590 617392 213596
rect 616420 213512 616472 213518
rect 616420 213454 616472 213460
rect 616788 213512 616840 213518
rect 616788 213454 616840 213460
rect 616432 210202 616460 213454
rect 616880 213444 616932 213450
rect 616880 213386 616932 213392
rect 616892 210202 616920 213386
rect 617352 210202 617380 213590
rect 617536 213450 617564 218894
rect 618168 217116 618220 217122
rect 618168 217058 618220 217064
rect 617800 213852 617852 213858
rect 617800 213794 617852 213800
rect 617524 213444 617576 213450
rect 617524 213386 617576 213392
rect 617812 210202 617840 213794
rect 618180 213654 618208 217058
rect 618720 215960 618772 215966
rect 618720 215902 618772 215908
rect 618168 213648 618220 213654
rect 618168 213590 618220 213596
rect 618260 213376 618312 213382
rect 618260 213318 618312 213324
rect 618272 210202 618300 213318
rect 618732 210202 618760 215902
rect 610788 210174 610848 210202
rect 611248 210174 611308 210202
rect 611708 210174 611768 210202
rect 612168 210174 612228 210202
rect 612628 210174 612688 210202
rect 613088 210174 613148 210202
rect 613548 210174 613608 210202
rect 614008 210174 614068 210202
rect 614560 210174 614620 210202
rect 615020 210174 615080 210202
rect 615480 210174 615540 210202
rect 615940 210174 616000 210202
rect 616400 210174 616460 210202
rect 616860 210174 616920 210202
rect 617320 210174 617380 210202
rect 617780 210174 617840 210202
rect 618240 210174 618300 210202
rect 618700 210174 618760 210202
rect 618824 210066 618852 220798
rect 618996 217184 619048 217190
rect 618996 217126 619048 217132
rect 619008 213586 619036 217126
rect 619640 216028 619692 216034
rect 619640 215970 619692 215976
rect 618996 213580 619048 213586
rect 618996 213522 619048 213528
rect 619652 210202 619680 215970
rect 619620 210174 619680 210202
rect 619836 210066 619864 220866
rect 620284 218340 620336 218346
rect 620284 218282 620336 218288
rect 619916 217864 619968 217870
rect 619916 217806 619968 217812
rect 619928 213858 619956 217806
rect 619916 213852 619968 213858
rect 619916 213794 619968 213800
rect 620296 213382 620324 218282
rect 621020 217524 621072 217530
rect 621020 217466 621072 217472
rect 621032 213722 621060 217466
rect 621020 213716 621072 213722
rect 621020 213658 621072 213664
rect 620284 213376 620336 213382
rect 620284 213318 620336 213324
rect 620560 213308 620612 213314
rect 620560 213250 620612 213256
rect 620572 210202 620600 213250
rect 621216 210202 621244 220934
rect 622952 219564 623004 219570
rect 622952 219506 623004 219512
rect 622584 216776 622636 216782
rect 622490 216744 622546 216753
rect 622584 216718 622636 216724
rect 622490 216679 622546 216688
rect 622032 213852 622084 213858
rect 622032 213794 622084 213800
rect 621480 213784 621532 213790
rect 621480 213726 621532 213732
rect 621492 210202 621520 213726
rect 622044 210202 622072 213794
rect 622504 210202 622532 216679
rect 620540 210174 620600 210202
rect 621000 210174 621244 210202
rect 621460 210174 621520 210202
rect 622012 210174 622072 210202
rect 622472 210174 622532 210202
rect 622596 210066 622624 216718
rect 622964 210338 622992 219506
rect 623056 213314 623084 242898
rect 639144 232552 639196 232558
rect 639144 232494 639196 232500
rect 638224 232484 638276 232490
rect 638224 232426 638276 232432
rect 636844 230512 636896 230518
rect 636844 230454 636896 230460
rect 623872 220788 623924 220794
rect 623872 220730 623924 220736
rect 623780 219632 623832 219638
rect 623780 219574 623832 219580
rect 623044 213308 623096 213314
rect 623044 213250 623096 213256
rect 623792 212430 623820 219574
rect 623780 212424 623832 212430
rect 623780 212366 623832 212372
rect 622964 210310 623084 210338
rect 623056 210066 623084 210310
rect 623884 210202 623912 220730
rect 632336 220652 632388 220658
rect 632336 220594 632388 220600
rect 625252 219768 625304 219774
rect 625252 219710 625304 219716
rect 623962 219464 624018 219473
rect 623962 219399 624018 219408
rect 623852 210174 623912 210202
rect 623976 210066 624004 219399
rect 625264 212430 625292 219710
rect 625528 219700 625580 219706
rect 625528 219642 625580 219648
rect 624424 212424 624476 212430
rect 624424 212366 624476 212372
rect 625252 212424 625304 212430
rect 625252 212366 625304 212372
rect 624436 210066 624464 212366
rect 625540 210202 625568 219642
rect 629944 218204 629996 218210
rect 629944 218146 629996 218152
rect 629208 217320 629260 217326
rect 629208 217262 629260 217268
rect 628472 216368 628524 216374
rect 628472 216310 628524 216316
rect 626172 216232 626224 216238
rect 626172 216174 626224 216180
rect 625712 212424 625764 212430
rect 625712 212366 625764 212372
rect 625724 210202 625752 212366
rect 626184 210202 626212 216174
rect 628012 216164 628064 216170
rect 628012 216106 628064 216112
rect 627092 214872 627144 214878
rect 627092 214814 627144 214820
rect 626632 214668 626684 214674
rect 626632 214610 626684 214616
rect 626644 210202 626672 214610
rect 627104 210202 627132 214814
rect 627552 214736 627604 214742
rect 627552 214678 627604 214684
rect 627564 210202 627592 214678
rect 628024 210202 628052 216106
rect 628484 210202 628512 216310
rect 629220 213654 629248 217262
rect 629484 216096 629536 216102
rect 629484 216038 629536 216044
rect 628932 213648 628984 213654
rect 628932 213590 628984 213596
rect 629208 213648 629260 213654
rect 629208 213590 629260 213596
rect 628944 210202 628972 213590
rect 629496 210202 629524 216038
rect 629956 213858 629984 218146
rect 631784 216504 631836 216510
rect 631784 216446 631836 216452
rect 630404 216436 630456 216442
rect 630404 216378 630456 216384
rect 629944 213852 629996 213858
rect 629944 213794 629996 213800
rect 629944 213580 629996 213586
rect 629944 213522 629996 213528
rect 629956 210202 629984 213522
rect 630416 210202 630444 216378
rect 630864 216300 630916 216306
rect 630864 216242 630916 216248
rect 630876 210202 630904 216242
rect 631324 213716 631376 213722
rect 631324 213658 631376 213664
rect 631336 210202 631364 213658
rect 631796 210202 631824 216446
rect 632244 213648 632296 213654
rect 632244 213590 632296 213596
rect 632256 210202 632284 213590
rect 625448 210174 625568 210202
rect 625692 210174 625752 210202
rect 626152 210174 626212 210202
rect 626612 210174 626672 210202
rect 627072 210174 627132 210202
rect 627532 210174 627592 210202
rect 627992 210174 628052 210202
rect 628452 210174 628512 210202
rect 628912 210174 628972 210202
rect 629464 210174 629524 210202
rect 629924 210174 629984 210202
rect 630384 210174 630444 210202
rect 630844 210174 630904 210202
rect 631304 210174 631364 210202
rect 631764 210174 631824 210202
rect 632224 210174 632284 210202
rect 625448 210066 625476 210174
rect 608612 210038 608948 210066
rect 609992 210038 610328 210066
rect 618824 210038 619160 210066
rect 619836 210038 620080 210066
rect 622596 210038 622932 210066
rect 623056 210038 623392 210066
rect 623976 210038 624312 210066
rect 624436 210038 624772 210066
rect 625232 210038 625476 210066
rect 632348 210066 632376 220594
rect 636016 218272 636068 218278
rect 636016 218214 636068 218220
rect 634544 217728 634596 217734
rect 634544 217670 634596 217676
rect 634084 217660 634136 217666
rect 634084 217602 634136 217608
rect 633624 217592 633676 217598
rect 633624 217534 633676 217540
rect 633164 217456 633216 217462
rect 633164 217398 633216 217404
rect 633176 210202 633204 217398
rect 633636 210202 633664 217534
rect 634096 210202 634124 217602
rect 634556 210202 634584 217670
rect 635004 214600 635056 214606
rect 635004 214542 635056 214548
rect 635016 210202 635044 214542
rect 636028 213790 636056 218214
rect 636108 218136 636160 218142
rect 636108 218078 636160 218084
rect 636120 213926 636148 218078
rect 636108 213920 636160 213926
rect 636108 213862 636160 213868
rect 636856 213858 636884 230454
rect 638236 213926 638264 232426
rect 639156 229094 639184 232494
rect 647344 230489 647372 278122
rect 648724 277394 648752 277780
rect 648632 277366 648752 277394
rect 648632 267073 648660 277366
rect 648618 267064 648674 267073
rect 648618 266999 648674 267008
rect 649356 231396 649408 231402
rect 649356 231338 649408 231344
rect 647330 230480 647386 230489
rect 647330 230415 647386 230424
rect 649368 229094 649396 231338
rect 639156 229066 639368 229094
rect 649368 229066 649580 229094
rect 638316 218068 638368 218074
rect 638316 218010 638368 218016
rect 637396 213920 637448 213926
rect 637396 213862 637448 213868
rect 638224 213920 638276 213926
rect 638224 213862 638276 213868
rect 636568 213852 636620 213858
rect 636568 213794 636620 213800
rect 636844 213852 636896 213858
rect 636844 213794 636896 213800
rect 636016 213784 636068 213790
rect 636016 213726 636068 213732
rect 635464 213512 635516 213518
rect 635464 213454 635516 213460
rect 635476 210202 635504 213454
rect 635924 213444 635976 213450
rect 635924 213386 635976 213392
rect 635936 210202 635964 213386
rect 636384 213376 636436 213382
rect 636384 213318 636436 213324
rect 636396 210202 636424 213318
rect 633144 210174 633204 210202
rect 633604 210174 633664 210202
rect 634064 210174 634124 210202
rect 634524 210174 634584 210202
rect 634984 210174 635044 210202
rect 635444 210174 635504 210202
rect 635904 210174 635964 210202
rect 636364 210174 636424 210202
rect 636580 210066 636608 213794
rect 637408 210202 637436 213862
rect 637856 213784 637908 213790
rect 637856 213726 637908 213732
rect 637868 210202 637896 213726
rect 638328 210202 638356 218010
rect 639236 213852 639288 213858
rect 639236 213794 639288 213800
rect 639248 210202 639276 213794
rect 637376 210174 637436 210202
rect 637836 210174 637896 210202
rect 638296 210174 638356 210202
rect 639216 210174 639276 210202
rect 639340 210066 639368 229066
rect 647148 218884 647200 218890
rect 647148 218826 647200 218832
rect 640616 213920 640668 213926
rect 640616 213862 640668 213868
rect 640156 213240 640208 213246
rect 640156 213182 640208 213188
rect 640168 210202 640196 213182
rect 640628 210202 640656 213862
rect 641076 213308 641128 213314
rect 641076 213250 641128 213256
rect 642732 213308 642784 213314
rect 642732 213250 642784 213256
rect 641088 210202 641116 213250
rect 641824 210310 642128 210338
rect 641824 210202 641852 210310
rect 640136 210174 640196 210202
rect 640596 210174 640656 210202
rect 641056 210174 641116 210202
rect 641516 210174 641852 210202
rect 642100 210066 642128 210310
rect 642744 210202 642772 213250
rect 643836 213240 643888 213246
rect 643836 213182 643888 213188
rect 643204 210310 643508 210338
rect 643204 210202 643232 210310
rect 642436 210188 642772 210202
rect 642422 210174 642772 210188
rect 642896 210174 643232 210202
rect 642422 210066 642450 210174
rect 632348 210038 632684 210066
rect 636580 210038 636916 210066
rect 639340 210038 639676 210066
rect 642100 210052 642450 210066
rect 643480 210066 643508 210310
rect 643848 210202 643876 213182
rect 646964 213036 647016 213042
rect 646964 212978 647016 212984
rect 645584 212628 645636 212634
rect 645584 212570 645636 212576
rect 644584 210310 644980 210338
rect 644584 210202 644612 210310
rect 643816 210188 643876 210202
rect 643802 210174 643876 210188
rect 644368 210174 644612 210202
rect 643802 210066 643830 210174
rect 643480 210052 643830 210066
rect 644952 210066 644980 210310
rect 645596 210202 645624 212570
rect 646056 210310 646360 210338
rect 646056 210202 646084 210310
rect 645288 210188 645624 210202
rect 645274 210174 645624 210188
rect 645748 210174 646084 210202
rect 645274 210066 645302 210174
rect 644952 210052 645302 210066
rect 646332 210066 646360 210310
rect 646976 210202 647004 212978
rect 647160 210202 647188 218826
rect 648526 213072 648582 213081
rect 648526 213007 648582 213016
rect 647436 210310 647740 210338
rect 647436 210202 647464 210310
rect 646668 210188 647004 210202
rect 646654 210174 647004 210188
rect 647128 210174 647464 210202
rect 646654 210066 646682 210174
rect 646332 210052 646682 210066
rect 647712 210066 647740 210310
rect 648540 210202 648568 213007
rect 648816 210310 649120 210338
rect 648816 210202 648844 210310
rect 648508 210174 648844 210202
rect 649092 210066 649120 210310
rect 649552 210066 649580 229066
rect 650012 213314 650040 984778
rect 651380 984768 651432 984774
rect 651380 984710 651432 984716
rect 650092 984700 650144 984706
rect 650092 984642 650144 984648
rect 650000 213308 650052 213314
rect 650000 213250 650052 213256
rect 650104 212634 650132 984642
rect 650644 231464 650696 231470
rect 650644 231406 650696 231412
rect 650656 229094 650684 231406
rect 650656 229066 650960 229094
rect 650092 212628 650144 212634
rect 650092 212570 650144 212576
rect 650196 210310 650500 210338
rect 650196 210066 650224 210310
rect 642100 210038 642436 210052
rect 643480 210038 643816 210052
rect 644952 210038 645288 210052
rect 646332 210038 646668 210052
rect 647712 210038 648048 210066
rect 649092 210038 649428 210066
rect 649552 210038 650224 210066
rect 650472 210066 650500 210310
rect 650932 210066 650960 229066
rect 651392 213246 651420 984710
rect 651472 984632 651524 984638
rect 651472 984574 651524 984580
rect 651380 213240 651432 213246
rect 651380 213182 651432 213188
rect 651484 213042 651512 984574
rect 651654 975896 651710 975905
rect 651654 975831 651710 975840
rect 651668 975730 651696 975831
rect 651656 975724 651708 975730
rect 651656 975666 651708 975672
rect 652022 962568 652078 962577
rect 652022 962503 652078 962512
rect 651562 949376 651618 949385
rect 651562 949311 651618 949320
rect 651576 948122 651604 949311
rect 651564 948116 651616 948122
rect 651564 948058 651616 948064
rect 652036 939826 652064 962503
rect 652024 939820 652076 939826
rect 652024 939762 652076 939768
rect 658936 937242 658964 991646
rect 659016 957840 659068 957846
rect 659016 957782 659068 957788
rect 658924 937236 658976 937242
rect 658924 937178 658976 937184
rect 659028 937038 659056 957782
rect 660316 938602 660344 993006
rect 660304 938596 660356 938602
rect 660304 938538 660356 938544
rect 651564 937032 651616 937038
rect 651564 936974 651616 936980
rect 659016 937032 659068 937038
rect 659016 936974 659068 936980
rect 651576 936193 651604 936974
rect 651562 936184 651618 936193
rect 651562 936119 651618 936128
rect 661696 935678 661724 995590
rect 666652 992996 666704 993002
rect 666652 992938 666704 992944
rect 666560 991636 666612 991642
rect 666560 991578 666612 991584
rect 665456 991500 665508 991506
rect 665456 991442 665508 991448
rect 663064 990140 663116 990146
rect 663064 990082 663116 990088
rect 663076 937378 663104 990082
rect 663064 937372 663116 937378
rect 663064 937314 663116 937320
rect 661684 935672 661736 935678
rect 661684 935614 661736 935620
rect 651562 922720 651618 922729
rect 651562 922655 651618 922664
rect 651576 921874 651604 922655
rect 651564 921868 651616 921874
rect 651564 921810 651616 921816
rect 651562 909528 651618 909537
rect 651562 909463 651564 909472
rect 651616 909463 651618 909472
rect 661684 909492 661736 909498
rect 651564 909434 651616 909440
rect 661684 909434 661736 909440
rect 651562 896200 651618 896209
rect 651562 896135 651618 896144
rect 651576 895694 651604 896135
rect 651564 895688 651616 895694
rect 651564 895630 651616 895636
rect 660304 895688 660356 895694
rect 660304 895630 660356 895636
rect 652022 882872 652078 882881
rect 652022 882807 652078 882816
rect 651562 869680 651618 869689
rect 651562 869615 651618 869624
rect 651576 869446 651604 869615
rect 651564 869440 651616 869446
rect 651564 869382 651616 869388
rect 652036 868698 652064 882807
rect 652024 868692 652076 868698
rect 652024 868634 652076 868640
rect 651562 856352 651618 856361
rect 651562 856287 651618 856296
rect 651576 855642 651604 856287
rect 651564 855636 651616 855642
rect 651564 855578 651616 855584
rect 651562 843024 651618 843033
rect 651562 842959 651618 842968
rect 651576 841838 651604 842959
rect 651564 841832 651616 841838
rect 651564 841774 651616 841780
rect 651562 829832 651618 829841
rect 651562 829767 651618 829776
rect 651576 829462 651604 829767
rect 651564 829456 651616 829462
rect 651564 829398 651616 829404
rect 658924 829456 658976 829462
rect 658924 829398 658976 829404
rect 651562 816504 651618 816513
rect 651562 816439 651618 816448
rect 651576 815658 651604 816439
rect 651564 815652 651616 815658
rect 651564 815594 651616 815600
rect 651562 803312 651618 803321
rect 651562 803247 651618 803256
rect 651576 803214 651604 803247
rect 651564 803208 651616 803214
rect 651564 803150 651616 803156
rect 651654 789984 651710 789993
rect 651654 789919 651710 789928
rect 651668 789410 651696 789919
rect 651656 789404 651708 789410
rect 651656 789346 651708 789352
rect 658936 779006 658964 829398
rect 658924 779000 658976 779006
rect 658924 778942 658976 778948
rect 651562 776656 651618 776665
rect 651562 776591 651618 776600
rect 651576 775606 651604 776591
rect 651564 775600 651616 775606
rect 651564 775542 651616 775548
rect 658924 775600 658976 775606
rect 658924 775542 658976 775548
rect 651562 763328 651618 763337
rect 651562 763263 651618 763272
rect 651576 763230 651604 763263
rect 651564 763224 651616 763230
rect 651564 763166 651616 763172
rect 651562 750136 651618 750145
rect 651562 750071 651618 750080
rect 651576 749494 651604 750071
rect 651564 749488 651616 749494
rect 651564 749430 651616 749436
rect 651562 736808 651618 736817
rect 651562 736743 651618 736752
rect 651576 735622 651604 736743
rect 651564 735616 651616 735622
rect 651564 735558 651616 735564
rect 658936 734874 658964 775542
rect 660316 760578 660344 895630
rect 661696 760714 661724 909434
rect 664444 855636 664496 855642
rect 664444 855578 664496 855584
rect 663064 841832 663116 841838
rect 663064 841774 663116 841780
rect 661776 789404 661828 789410
rect 661776 789346 661828 789352
rect 661684 760708 661736 760714
rect 661684 760650 661736 760656
rect 660304 760572 660356 760578
rect 660304 760514 660356 760520
rect 660304 735616 660356 735622
rect 660304 735558 660356 735564
rect 658924 734868 658976 734874
rect 658924 734810 658976 734816
rect 652022 723480 652078 723489
rect 652022 723415 652078 723424
rect 652036 723178 652064 723415
rect 652024 723172 652076 723178
rect 652024 723114 652076 723120
rect 658924 723172 658976 723178
rect 658924 723114 658976 723120
rect 651562 710288 651618 710297
rect 651562 710223 651618 710232
rect 651576 709374 651604 710223
rect 651564 709368 651616 709374
rect 651564 709310 651616 709316
rect 652022 696960 652078 696969
rect 652022 696895 652078 696904
rect 651838 683632 651894 683641
rect 651838 683567 651894 683576
rect 651852 683194 651880 683567
rect 651840 683188 651892 683194
rect 651840 683130 651892 683136
rect 651562 670440 651618 670449
rect 651562 670375 651618 670384
rect 651576 669390 651604 670375
rect 651564 669384 651616 669390
rect 651564 669326 651616 669332
rect 651562 657112 651618 657121
rect 651562 657047 651618 657056
rect 651576 656946 651604 657047
rect 651564 656940 651616 656946
rect 651564 656882 651616 656888
rect 651562 643784 651618 643793
rect 651562 643719 651618 643728
rect 651576 643142 651604 643719
rect 651564 643136 651616 643142
rect 651564 643078 651616 643084
rect 651562 630592 651618 630601
rect 651562 630527 651618 630536
rect 651576 629338 651604 630527
rect 651564 629332 651616 629338
rect 651564 629274 651616 629280
rect 651562 603936 651618 603945
rect 651562 603871 651618 603880
rect 651576 603158 651604 603871
rect 651564 603152 651616 603158
rect 651564 603094 651616 603100
rect 651562 590744 651618 590753
rect 651562 590679 651564 590688
rect 651616 590679 651618 590688
rect 651564 590650 651616 590656
rect 652036 581058 652064 696895
rect 658936 689314 658964 723114
rect 658924 689308 658976 689314
rect 658924 689250 658976 689256
rect 658924 683188 658976 683194
rect 658924 683130 658976 683136
rect 652390 617264 652446 617273
rect 652390 617199 652446 617208
rect 652404 616894 652432 617199
rect 652392 616888 652444 616894
rect 652392 616830 652444 616836
rect 652024 581052 652076 581058
rect 652024 580994 652076 581000
rect 658936 579834 658964 683130
rect 659016 669384 659068 669390
rect 659016 669326 659068 669332
rect 659028 643754 659056 669326
rect 659016 643748 659068 643754
rect 659016 643690 659068 643696
rect 660316 625190 660344 735558
rect 661788 669458 661816 789346
rect 663076 715018 663104 841774
rect 664456 716310 664484 855578
rect 664536 763224 664588 763230
rect 664536 763166 664588 763172
rect 664444 716304 664496 716310
rect 664444 716246 664496 716252
rect 663064 715012 663116 715018
rect 663064 714954 663116 714960
rect 661776 669452 661828 669458
rect 661776 669394 661828 669400
rect 663064 656940 663116 656946
rect 663064 656882 663116 656888
rect 661776 629332 661828 629338
rect 661776 629274 661828 629280
rect 660304 625184 660356 625190
rect 660304 625126 660356 625132
rect 659016 616888 659068 616894
rect 659016 616830 659068 616836
rect 659028 599622 659056 616830
rect 660304 603152 660356 603158
rect 660304 603094 660356 603100
rect 659016 599616 659068 599622
rect 659016 599558 659068 599564
rect 658924 579828 658976 579834
rect 658924 579770 658976 579776
rect 651562 577416 651618 577425
rect 651562 577351 651618 577360
rect 651576 576910 651604 577351
rect 651564 576904 651616 576910
rect 651564 576846 651616 576852
rect 659016 576904 659068 576910
rect 659016 576846 659068 576852
rect 652114 564088 652170 564097
rect 652114 564023 652170 564032
rect 652128 563106 652156 564023
rect 652116 563100 652168 563106
rect 652116 563042 652168 563048
rect 658924 563100 658976 563106
rect 658924 563042 658976 563048
rect 658936 554062 658964 563042
rect 658924 554056 658976 554062
rect 658924 553998 658976 554004
rect 651562 550896 651618 550905
rect 651562 550831 651618 550840
rect 651576 550662 651604 550831
rect 651564 550656 651616 550662
rect 651564 550598 651616 550604
rect 651562 537568 651618 537577
rect 651562 537503 651618 537512
rect 651576 536858 651604 537503
rect 651564 536852 651616 536858
rect 651564 536794 651616 536800
rect 651562 524240 651618 524249
rect 651562 524175 651618 524184
rect 651576 523054 651604 524175
rect 651564 523048 651616 523054
rect 651564 522990 651616 522996
rect 651562 511048 651618 511057
rect 651562 510983 651618 510992
rect 651576 510678 651604 510983
rect 651564 510672 651616 510678
rect 651564 510614 651616 510620
rect 651562 497720 651618 497729
rect 651562 497655 651618 497664
rect 651576 496874 651604 497655
rect 651564 496868 651616 496874
rect 651564 496810 651616 496816
rect 658924 496868 658976 496874
rect 658924 496810 658976 496816
rect 651562 484528 651618 484537
rect 651562 484463 651618 484472
rect 651576 484430 651604 484463
rect 651564 484424 651616 484430
rect 651564 484366 651616 484372
rect 651654 471200 651710 471209
rect 651654 471135 651710 471144
rect 651668 470626 651696 471135
rect 651656 470620 651708 470626
rect 651656 470562 651708 470568
rect 651562 457872 651618 457881
rect 651562 457807 651618 457816
rect 651576 456822 651604 457807
rect 651564 456816 651616 456822
rect 651564 456758 651616 456764
rect 651562 444544 651618 444553
rect 651562 444479 651618 444488
rect 651576 444446 651604 444479
rect 651564 444440 651616 444446
rect 651564 444382 651616 444388
rect 651562 431352 651618 431361
rect 651562 431287 651618 431296
rect 651576 430642 651604 431287
rect 651564 430636 651616 430642
rect 651564 430578 651616 430584
rect 651562 418024 651618 418033
rect 651562 417959 651618 417968
rect 651576 416838 651604 417959
rect 651564 416832 651616 416838
rect 651564 416774 651616 416780
rect 652022 404696 652078 404705
rect 652022 404631 652078 404640
rect 652036 404394 652064 404631
rect 652024 404388 652076 404394
rect 652024 404330 652076 404336
rect 651562 391504 651618 391513
rect 651562 391439 651618 391448
rect 651576 390590 651604 391439
rect 651564 390584 651616 390590
rect 651564 390526 651616 390532
rect 651564 378208 651616 378214
rect 651562 378176 651564 378185
rect 651616 378176 651618 378185
rect 651562 378111 651618 378120
rect 652022 364848 652078 364857
rect 652022 364783 652078 364792
rect 652036 364410 652064 364783
rect 652024 364404 652076 364410
rect 652024 364346 652076 364352
rect 658936 357610 658964 496810
rect 659028 491434 659056 576846
rect 660316 491570 660344 603094
rect 661684 550656 661736 550662
rect 661684 550598 661736 550604
rect 660304 491564 660356 491570
rect 660304 491506 660356 491512
rect 659016 491428 659068 491434
rect 659016 491370 659068 491376
rect 660396 484424 660448 484430
rect 660396 484366 660448 484372
rect 659016 444440 659068 444446
rect 659016 444382 659068 444388
rect 658924 357604 658976 357610
rect 658924 357546 658976 357552
rect 651562 351656 651618 351665
rect 651562 351591 651618 351600
rect 651576 350606 651604 351591
rect 651564 350600 651616 350606
rect 651564 350542 651616 350548
rect 651654 338328 651710 338337
rect 651654 338263 651710 338272
rect 651668 338162 651696 338263
rect 651656 338156 651708 338162
rect 651656 338098 651708 338104
rect 651562 325000 651618 325009
rect 651562 324935 651618 324944
rect 651576 324358 651604 324935
rect 651564 324352 651616 324358
rect 651564 324294 651616 324300
rect 659028 312050 659056 444382
rect 660304 430636 660356 430642
rect 660304 430578 660356 430584
rect 659016 312044 659068 312050
rect 659016 311986 659068 311992
rect 652390 311808 652446 311817
rect 652390 311743 652446 311752
rect 652404 310554 652432 311743
rect 652392 310548 652444 310554
rect 652392 310490 652444 310496
rect 652022 298480 652078 298489
rect 652022 298415 652078 298424
rect 651562 285288 651618 285297
rect 651562 285223 651618 285232
rect 651576 284374 651604 285223
rect 651564 284368 651616 284374
rect 651564 284310 651616 284316
rect 651472 213036 651524 213042
rect 651472 212978 651524 212984
rect 652036 210458 652064 298415
rect 659660 278112 659712 278118
rect 659660 278054 659712 278060
rect 658280 278044 658332 278050
rect 658280 277986 658332 277992
rect 655520 231328 655572 231334
rect 655520 231270 655572 231276
rect 652760 231260 652812 231266
rect 652760 231202 652812 231208
rect 652024 210452 652076 210458
rect 652024 210394 652076 210400
rect 651668 210310 651972 210338
rect 651668 210066 651696 210310
rect 650472 210038 650808 210066
rect 650932 210038 651696 210066
rect 651944 210066 651972 210310
rect 652772 210202 652800 231202
rect 654138 218512 654194 218521
rect 654138 218447 654194 218456
rect 653048 210310 653352 210338
rect 653048 210202 653076 210310
rect 652740 210174 653076 210202
rect 653324 210066 653352 210310
rect 654152 210202 654180 218447
rect 654428 210310 654732 210338
rect 654428 210202 654456 210310
rect 654120 210174 654456 210202
rect 654704 210066 654732 210310
rect 655532 210202 655560 231270
rect 656900 218816 656952 218822
rect 656900 218758 656952 218764
rect 655808 210310 656112 210338
rect 655808 210202 655836 210310
rect 655500 210174 655836 210202
rect 656084 210066 656112 210310
rect 656912 210202 656940 218758
rect 657188 210310 657492 210338
rect 657188 210202 657216 210310
rect 656880 210174 657216 210202
rect 657464 210066 657492 210310
rect 658292 210202 658320 277986
rect 659672 229094 659700 278054
rect 660316 267782 660344 430578
rect 660408 357746 660436 484366
rect 661696 403170 661724 550598
rect 661788 534274 661816 629274
rect 663076 535634 663104 656882
rect 664548 625394 664576 763166
rect 664536 625388 664588 625394
rect 664536 625330 664588 625336
rect 664444 590708 664496 590714
rect 664444 590650 664496 590656
rect 663064 535628 663116 535634
rect 663064 535570 663116 535576
rect 661776 534268 661828 534274
rect 661776 534210 661828 534216
rect 663156 523048 663208 523054
rect 663156 522990 663208 522996
rect 663064 416832 663116 416838
rect 663064 416774 663116 416780
rect 661776 404388 661828 404394
rect 661776 404330 661828 404336
rect 661684 403164 661736 403170
rect 661684 403106 661736 403112
rect 660396 357740 660448 357746
rect 660396 357682 660448 357688
rect 661788 267986 661816 404330
rect 663076 268122 663104 416774
rect 663168 403306 663196 522990
rect 664456 491706 664484 590650
rect 664536 536852 664588 536858
rect 664536 536794 664588 536800
rect 664444 491700 664496 491706
rect 664444 491642 664496 491648
rect 664444 470620 664496 470626
rect 664444 470562 664496 470568
rect 663156 403300 663208 403306
rect 663156 403242 663208 403248
rect 664456 313410 664484 470562
rect 664548 403442 664576 536794
rect 664536 403436 664588 403442
rect 664536 403378 664588 403384
rect 664536 378208 664588 378214
rect 664536 378150 664588 378156
rect 664444 313404 664496 313410
rect 664444 313346 664496 313352
rect 663064 268116 663116 268122
rect 663064 268058 663116 268064
rect 661776 267980 661828 267986
rect 661776 267922 661828 267928
rect 660304 267776 660356 267782
rect 660304 267718 660356 267724
rect 662420 264240 662472 264246
rect 662420 264182 662472 264188
rect 661040 231192 661092 231198
rect 661040 231134 661092 231140
rect 661052 229094 661080 231134
rect 659672 229066 659792 229094
rect 661052 229066 661172 229094
rect 658568 210310 658872 210338
rect 658568 210202 658596 210310
rect 658260 210174 658596 210202
rect 658844 210066 658872 210310
rect 659764 210202 659792 229066
rect 660040 210310 660344 210338
rect 660040 210202 660068 210310
rect 659732 210174 660068 210202
rect 660316 210066 660344 210310
rect 661144 210202 661172 229066
rect 662432 210594 662460 264182
rect 663984 231668 664036 231674
rect 663984 231610 664036 231616
rect 663800 231600 663852 231606
rect 663800 231542 663852 231548
rect 662512 231124 662564 231130
rect 662512 231066 662564 231072
rect 662524 229094 662552 231066
rect 662524 229066 662644 229094
rect 662512 218748 662564 218754
rect 662512 218690 662564 218696
rect 662420 210588 662472 210594
rect 662420 210530 662472 210536
rect 661420 210310 661724 210338
rect 661420 210202 661448 210310
rect 661112 210174 661448 210202
rect 661696 210066 661724 210310
rect 662524 210202 662552 218690
rect 662492 210174 662552 210202
rect 662616 210066 662644 229066
rect 663812 212430 663840 231542
rect 663892 231532 663944 231538
rect 663892 231474 663944 231480
rect 663800 212424 663852 212430
rect 663800 212366 663852 212372
rect 663904 212362 663932 231474
rect 663996 229094 664024 231610
rect 663996 229066 664208 229094
rect 663892 212356 663944 212362
rect 663892 212298 663944 212304
rect 663064 210588 663116 210594
rect 663064 210530 663116 210536
rect 663076 210066 663104 210530
rect 664180 210202 664208 229066
rect 664548 222222 664576 378150
rect 664536 222216 664588 222222
rect 664536 222158 664588 222164
rect 665272 214396 665324 214402
rect 665272 214338 665324 214344
rect 664444 212424 664496 212430
rect 664444 212366 664496 212372
rect 664352 212356 664404 212362
rect 664352 212298 664404 212304
rect 664364 210202 664392 212298
rect 664088 210174 664208 210202
rect 664332 210174 664392 210202
rect 664088 210066 664116 210174
rect 651944 210038 652280 210066
rect 653324 210038 653660 210066
rect 654704 210038 655040 210066
rect 656084 210038 656420 210066
rect 657464 210038 657800 210066
rect 658844 210038 659272 210066
rect 660316 210038 660652 210066
rect 661696 210038 662032 210066
rect 662616 210038 662952 210066
rect 663076 210038 663412 210066
rect 663872 210038 664116 210066
rect 664456 210066 664484 212366
rect 665284 210202 665312 214338
rect 665252 210174 665312 210202
rect 664456 210038 664792 210066
rect 638408 209840 638460 209846
rect 638460 209788 638756 209794
rect 638408 209782 638756 209788
rect 638420 209766 638756 209782
rect 665468 209710 665496 991442
rect 665824 815652 665876 815658
rect 665824 815594 665876 815600
rect 665836 670818 665864 815594
rect 665824 670812 665876 670818
rect 665824 670754 665876 670760
rect 665824 510672 665876 510678
rect 665824 510614 665876 510620
rect 665836 357882 665864 510614
rect 665824 357876 665876 357882
rect 665824 357818 665876 357824
rect 666192 214260 666244 214266
rect 666192 214202 666244 214208
rect 665732 214124 665784 214130
rect 665732 214066 665784 214072
rect 665744 210202 665772 214066
rect 666204 210202 666232 214202
rect 665712 210174 665772 210202
rect 666172 210174 666232 210202
rect 665456 209704 665508 209710
rect 665456 209646 665508 209652
rect 666572 189009 666600 991578
rect 666664 194041 666692 992938
rect 666836 992928 666888 992934
rect 666836 992870 666888 992876
rect 666744 991568 666796 991574
rect 666744 991510 666796 991516
rect 666756 199073 666784 991510
rect 666848 204241 666876 992870
rect 672724 975724 672776 975730
rect 672724 975666 672776 975672
rect 669964 961920 670016 961926
rect 669964 961862 670016 961868
rect 668676 643136 668728 643142
rect 668676 643078 668728 643084
rect 668584 568608 668636 568614
rect 668584 568550 668636 568556
rect 668124 214192 668176 214198
rect 668124 214134 668176 214140
rect 667204 210452 667256 210458
rect 667204 210394 667256 210400
rect 666928 209704 666980 209710
rect 666928 209646 666980 209652
rect 666940 209273 666968 209646
rect 666926 209264 666982 209273
rect 666926 209199 666982 209208
rect 666834 204232 666890 204241
rect 666834 204167 666890 204176
rect 666848 200841 666876 204167
rect 666834 200832 666890 200841
rect 666834 200767 666890 200776
rect 666742 199064 666798 199073
rect 666742 198999 666798 199008
rect 666650 194032 666706 194041
rect 666650 193967 666706 193976
rect 666664 190641 666692 193967
rect 666650 190632 666706 190641
rect 666650 190567 666706 190576
rect 666558 189000 666614 189009
rect 666558 188935 666614 188944
rect 666572 185609 666600 188935
rect 666558 185600 666614 185609
rect 666558 185535 666614 185544
rect 666558 163568 666614 163577
rect 666558 163503 666614 163512
rect 666572 161537 666600 163503
rect 666558 161528 666614 161537
rect 666558 161463 666614 161472
rect 666558 153368 666614 153377
rect 666558 153303 666614 153312
rect 666572 151881 666600 153303
rect 666558 151872 666614 151881
rect 666558 151807 666614 151816
rect 666558 151600 666614 151609
rect 666558 151535 666614 151544
rect 666572 149977 666600 151535
rect 666558 149968 666614 149977
rect 666558 149903 666614 149912
rect 666558 142080 666614 142089
rect 666558 142015 666614 142024
rect 666572 139777 666600 142015
rect 666558 139768 666614 139777
rect 666558 139703 666614 139712
rect 667216 132666 667244 210394
rect 667938 209264 667994 209273
rect 667938 209199 667994 209208
rect 667952 205873 667980 209199
rect 667938 205864 667994 205873
rect 667938 205799 667994 205808
rect 667938 199064 667994 199073
rect 667938 198999 667994 199008
rect 667952 195673 667980 198999
rect 667938 195664 667994 195673
rect 667938 195599 667994 195608
rect 668030 183832 668086 183841
rect 668030 183767 668086 183776
rect 668044 180441 668072 183767
rect 668030 180432 668086 180441
rect 668030 180367 668086 180376
rect 667940 178832 667992 178838
rect 667938 178800 667940 178809
rect 667992 178800 667994 178809
rect 667938 178735 667994 178744
rect 667952 175409 667980 178735
rect 667938 175400 667994 175409
rect 667938 175335 667994 175344
rect 667940 173664 667992 173670
rect 667938 173632 667940 173641
rect 667992 173632 667994 173641
rect 667938 173567 667994 173576
rect 667952 171193 667980 173567
rect 667938 171184 667994 171193
rect 667938 171119 667994 171128
rect 667938 168600 667994 168609
rect 667938 168535 667994 168544
rect 667952 165209 667980 168535
rect 667938 165200 667994 165209
rect 667938 165135 667994 165144
rect 667938 158400 667994 158409
rect 667938 158335 667994 158344
rect 667952 155009 667980 158335
rect 667938 155000 667994 155009
rect 667938 154935 667994 154944
rect 667940 143336 667992 143342
rect 667940 143278 667992 143284
rect 667952 143177 667980 143278
rect 667938 143168 667994 143177
rect 667938 143103 667994 143112
rect 668032 138236 668084 138242
rect 668032 138178 668084 138184
rect 668044 138145 668072 138178
rect 668030 138136 668086 138145
rect 668030 138071 668086 138080
rect 668044 134745 668072 138071
rect 668030 134736 668086 134745
rect 668030 134671 668086 134680
rect 667204 132660 667256 132666
rect 667204 132602 667256 132608
rect 666558 132424 666614 132433
rect 666558 132359 666614 132368
rect 666572 129577 666600 132359
rect 666558 129568 666614 129577
rect 666558 129503 666614 129512
rect 668032 128172 668084 128178
rect 668032 128114 668084 128120
rect 668044 127945 668072 128114
rect 668030 127936 668086 127945
rect 668030 127871 668086 127880
rect 668044 124545 668072 127871
rect 668030 124536 668086 124545
rect 668030 124471 668086 124480
rect 667940 123888 667992 123894
rect 667940 123830 667992 123836
rect 667952 122913 667980 123830
rect 667938 122904 667994 122913
rect 667938 122839 667994 122848
rect 666558 122768 666614 122777
rect 666558 122703 666614 122712
rect 666572 119513 666600 122703
rect 666558 119504 666614 119513
rect 666558 119439 666614 119448
rect 667940 111308 667992 111314
rect 667940 111250 667992 111256
rect 667952 110945 667980 111250
rect 667938 110936 667994 110945
rect 667938 110871 667994 110880
rect 667940 110356 667992 110362
rect 667940 110298 667992 110304
rect 667952 109313 667980 110298
rect 667938 109304 667994 109313
rect 667938 109239 667994 109248
rect 668136 107545 668164 214134
rect 668308 184204 668360 184210
rect 668308 184146 668360 184152
rect 668320 183841 668348 184146
rect 668306 183832 668362 183841
rect 668306 183767 668362 183776
rect 668400 164008 668452 164014
rect 668400 163950 668452 163956
rect 668412 163577 668440 163950
rect 668398 163568 668454 163577
rect 668398 163503 668454 163512
rect 668596 158409 668624 568550
rect 668688 535770 668716 643078
rect 668676 535764 668728 535770
rect 668676 535706 668728 535712
rect 668676 524476 668728 524482
rect 668676 524418 668728 524424
rect 668582 158400 668638 158409
rect 668582 158335 668638 158344
rect 668688 153377 668716 524418
rect 668952 214328 669004 214334
rect 668952 214270 669004 214276
rect 668860 214056 668912 214062
rect 668860 213998 668912 214004
rect 668768 213988 668820 213994
rect 668768 213930 668820 213936
rect 668674 153368 668730 153377
rect 668674 153303 668730 153312
rect 668308 148572 668360 148578
rect 668308 148514 668360 148520
rect 668320 148209 668348 148514
rect 668306 148200 668362 148209
rect 668306 148135 668362 148144
rect 668320 144945 668348 148135
rect 668306 144936 668362 144945
rect 668306 144871 668362 144880
rect 668584 133000 668636 133006
rect 668582 132968 668584 132977
rect 668636 132968 668638 132977
rect 668582 132903 668638 132912
rect 668676 131164 668728 131170
rect 668676 131106 668728 131112
rect 668584 129804 668636 129810
rect 668584 129746 668636 129752
rect 668492 117292 668544 117298
rect 668492 117234 668544 117240
rect 668504 116113 668532 117234
rect 668490 116104 668546 116113
rect 668490 116039 668546 116048
rect 668492 114368 668544 114374
rect 668490 114336 668492 114345
rect 668544 114336 668546 114345
rect 668490 114271 668546 114280
rect 668122 107536 668178 107545
rect 668122 107471 668178 107480
rect 668596 100881 668624 129746
rect 668688 104145 668716 131106
rect 668780 128382 668808 213930
rect 668872 129810 668900 213998
rect 668964 131170 668992 214270
rect 668952 131164 669004 131170
rect 668952 131106 669004 131112
rect 668860 129804 668912 129810
rect 668860 129746 668912 129752
rect 668768 128376 668820 128382
rect 668768 128318 668820 128324
rect 668674 104136 668730 104145
rect 668674 104071 668730 104080
rect 668780 102513 668808 128318
rect 668860 122868 668912 122874
rect 668860 122810 668912 122816
rect 668872 112713 668900 122810
rect 669228 117836 669280 117842
rect 669228 117778 669280 117784
rect 669240 117745 669268 117778
rect 669226 117736 669282 117745
rect 669226 117671 669282 117680
rect 668858 112704 668914 112713
rect 668858 112639 668914 112648
rect 669228 106140 669280 106146
rect 669228 106082 669280 106088
rect 669240 105913 669268 106082
rect 669226 105904 669282 105913
rect 669226 105839 669282 105848
rect 668766 102504 668822 102513
rect 668766 102439 668822 102448
rect 668582 100872 668638 100881
rect 668582 100807 668638 100816
rect 605852 100014 606740 100042
rect 605748 77988 605800 77994
rect 605748 77930 605800 77936
rect 603724 60716 603776 60722
rect 603724 60658 603776 60664
rect 591304 57248 591356 57254
rect 591304 57190 591356 57196
rect 580264 55684 580316 55690
rect 580264 55626 580316 55632
rect 579068 53100 579120 53106
rect 579068 53042 579120 53048
rect 576122 44976 576178 44985
rect 576122 44911 576178 44920
rect 478786 44704 478842 44713
rect 478786 44639 478842 44648
rect 605852 43625 605880 100014
rect 607370 99770 607398 100028
rect 607324 99742 607398 99770
rect 607692 100014 608028 100042
rect 607220 95532 607272 95538
rect 607220 95474 607272 95480
rect 605838 43616 605894 43625
rect 605838 43551 605894 43560
rect 607232 43489 607260 95474
rect 607324 45257 607352 99742
rect 607692 95538 607720 100014
rect 608658 99770 608686 100028
rect 608612 99742 608686 99770
rect 608796 100014 609316 100042
rect 609960 100014 610020 100042
rect 607680 95532 607732 95538
rect 607680 95474 607732 95480
rect 607310 45248 607366 45257
rect 607310 45183 607366 45192
rect 608612 45121 608640 99742
rect 608598 45112 608654 45121
rect 608598 45047 608654 45056
rect 608796 44878 608824 100014
rect 608784 44872 608836 44878
rect 608784 44814 608836 44820
rect 607218 43480 607274 43489
rect 607218 43415 607274 43424
rect 473176 42528 473228 42534
rect 473176 42470 473228 42476
rect 518622 42392 518678 42401
rect 518678 42350 518834 42378
rect 518622 42327 518678 42336
rect 471610 42120 471666 42129
rect 471408 42078 471610 42106
rect 471610 42055 471666 42064
rect 514850 42120 514906 42129
rect 520370 42120 520426 42129
rect 514906 42078 515154 42106
rect 514850 42055 514906 42064
rect 521750 42120 521806 42129
rect 520426 42078 520674 42106
rect 520370 42055 520426 42064
rect 525982 42120 526038 42129
rect 521806 42078 521870 42106
rect 521750 42055 521806 42064
rect 529662 42120 529718 42129
rect 526038 42078 526194 42106
rect 529322 42078 529662 42106
rect 525982 42055 526038 42064
rect 529662 42055 529718 42064
rect 460570 41783 460626 41792
rect 609992 41449 610020 100014
rect 610176 100014 610604 100042
rect 610912 100014 611248 100042
rect 611372 100014 611892 100042
rect 612016 100014 612536 100042
rect 612752 100014 613180 100042
rect 613488 100014 613916 100042
rect 614560 100014 614896 100042
rect 615204 100014 615448 100042
rect 615848 100014 616184 100042
rect 616492 100014 616736 100042
rect 617136 100014 617472 100042
rect 617780 100014 618116 100042
rect 618424 100014 618760 100042
rect 619068 100014 619496 100042
rect 619712 100014 620048 100042
rect 620448 100014 620784 100042
rect 621092 100014 621428 100042
rect 621736 100014 622072 100042
rect 622380 100014 622716 100042
rect 623024 100014 623544 100042
rect 623668 100014 623728 100042
rect 624312 100014 624648 100042
rect 624956 100014 625108 100042
rect 625600 100014 625936 100042
rect 626244 100014 626396 100042
rect 610072 96960 610124 96966
rect 610072 96902 610124 96908
rect 610084 45529 610112 96902
rect 610070 45520 610126 45529
rect 610070 45455 610126 45464
rect 610176 45393 610204 100014
rect 610912 96966 610940 100014
rect 610900 96960 610952 96966
rect 610900 96902 610952 96908
rect 610162 45384 610218 45393
rect 610162 45319 610218 45328
rect 611372 41585 611400 100014
rect 612016 84194 612044 100014
rect 611464 84166 612044 84194
rect 611464 46481 611492 84166
rect 611450 46472 611506 46481
rect 611450 46407 611506 46416
rect 612752 46209 612780 100014
rect 613488 84194 613516 100014
rect 614868 97510 614896 100014
rect 614856 97504 614908 97510
rect 614856 97446 614908 97452
rect 612844 84166 613516 84194
rect 612844 46345 612872 84166
rect 615420 75206 615448 100014
rect 616156 96966 616184 100014
rect 616144 96960 616196 96966
rect 616144 96902 616196 96908
rect 616708 89690 616736 100014
rect 617444 96966 617472 100014
rect 616788 96960 616840 96966
rect 616788 96902 616840 96908
rect 617432 96960 617484 96966
rect 617432 96902 617484 96908
rect 616696 89684 616748 89690
rect 616696 89626 616748 89632
rect 616800 88330 616828 96902
rect 616788 88324 616840 88330
rect 616788 88266 616840 88272
rect 618088 84182 618116 100014
rect 618168 96960 618220 96966
rect 618168 96902 618220 96908
rect 618076 84176 618128 84182
rect 618076 84118 618128 84124
rect 618180 84114 618208 96902
rect 618732 96898 618760 100014
rect 618720 96892 618772 96898
rect 618720 96834 618772 96840
rect 619468 86290 619496 100014
rect 620020 96898 620048 100014
rect 620756 97442 620784 100014
rect 620744 97436 620796 97442
rect 620744 97378 620796 97384
rect 621400 97238 621428 100014
rect 621664 97504 621716 97510
rect 621664 97446 621716 97452
rect 621388 97232 621440 97238
rect 621388 97174 621440 97180
rect 619548 96892 619600 96898
rect 619548 96834 619600 96840
rect 620008 96892 620060 96898
rect 620008 96834 620060 96840
rect 620928 96892 620980 96898
rect 620928 96834 620980 96840
rect 619456 86284 619508 86290
rect 619456 86226 619508 86232
rect 619560 85542 619588 96834
rect 620940 88262 620968 96834
rect 620928 88256 620980 88262
rect 620928 88198 620980 88204
rect 619548 85536 619600 85542
rect 619548 85478 619600 85484
rect 618168 84108 618220 84114
rect 618168 84050 618220 84056
rect 615408 75200 615460 75206
rect 615408 75142 615460 75148
rect 618904 59900 618956 59906
rect 618904 59842 618956 59848
rect 618916 53854 618944 59842
rect 621676 58682 621704 97446
rect 622044 97306 622072 100014
rect 622032 97300 622084 97306
rect 622032 97242 622084 97248
rect 622688 96966 622716 100014
rect 623516 97050 623544 100014
rect 623700 97170 623728 100014
rect 624620 97918 624648 100014
rect 625080 97986 625108 100014
rect 625068 97980 625120 97986
rect 625068 97922 625120 97928
rect 624608 97912 624660 97918
rect 624608 97854 624660 97860
rect 625804 97912 625856 97918
rect 625804 97854 625856 97860
rect 623688 97164 623740 97170
rect 623688 97106 623740 97112
rect 624424 97164 624476 97170
rect 624424 97106 624476 97112
rect 623516 97022 623728 97050
rect 622676 96960 622728 96966
rect 622676 96902 622728 96908
rect 623596 96960 623648 96966
rect 623596 96902 623648 96908
rect 623608 76634 623636 96902
rect 623596 76628 623648 76634
rect 623596 76570 623648 76576
rect 623700 75274 623728 97022
rect 624436 76566 624464 97106
rect 625816 89729 625844 97854
rect 625908 96966 625936 100014
rect 625988 97980 626040 97986
rect 625988 97922 626040 97928
rect 625896 96960 625948 96966
rect 625896 96902 625948 96908
rect 626000 90681 626028 97922
rect 626368 92585 626396 100014
rect 626552 100014 626980 100042
rect 627624 100014 627868 100042
rect 628268 100014 628328 100042
rect 626448 96960 626500 96966
rect 626448 96902 626500 96908
rect 626354 92576 626410 92585
rect 626354 92511 626410 92520
rect 626460 91633 626488 96902
rect 626552 93537 626580 100014
rect 627840 94489 627868 100014
rect 628300 95985 628328 100014
rect 628760 100014 628912 100042
rect 629556 100014 629708 100042
rect 630200 100014 630628 100042
rect 630844 100014 631180 100042
rect 631488 100014 631824 100042
rect 632132 100014 632468 100042
rect 632776 100014 633112 100042
rect 633512 100014 633848 100042
rect 634156 100014 634492 100042
rect 634800 100014 635136 100042
rect 635444 100014 635780 100042
rect 636088 100014 636148 100042
rect 636732 100014 637068 100042
rect 637376 100014 637528 100042
rect 638020 100014 638356 100042
rect 638664 100014 638908 100042
rect 639308 100014 639644 100042
rect 639952 100014 640288 100042
rect 640688 100014 641024 100042
rect 641332 100014 641668 100042
rect 628286 95976 628342 95985
rect 628286 95911 628342 95920
rect 628760 95826 628788 100014
rect 628728 95798 628788 95826
rect 629680 95826 629708 100014
rect 630600 96642 630628 100014
rect 631152 97646 631180 100014
rect 631140 97640 631192 97646
rect 631140 97582 631192 97588
rect 631796 96762 631824 100014
rect 632440 97714 632468 100014
rect 633084 97918 633112 100014
rect 633072 97912 633124 97918
rect 633072 97854 633124 97860
rect 633820 97850 633848 100014
rect 634464 97986 634492 100014
rect 634452 97980 634504 97986
rect 634452 97922 634504 97928
rect 633808 97844 633860 97850
rect 633808 97786 633860 97792
rect 632428 97708 632480 97714
rect 632428 97650 632480 97656
rect 634084 97708 634136 97714
rect 634084 97650 634136 97656
rect 632152 97640 632204 97646
rect 632152 97582 632204 97588
rect 631784 96756 631836 96762
rect 631784 96698 631836 96704
rect 630600 96614 630720 96642
rect 630692 95826 630720 96614
rect 629680 95798 629832 95826
rect 630692 95798 631028 95826
rect 632164 95690 632192 97582
rect 632980 96756 633032 96762
rect 632980 96698 633032 96704
rect 632992 95826 633020 96698
rect 634096 95826 634124 97650
rect 635108 97578 635136 100014
rect 635280 97912 635332 97918
rect 635280 97854 635332 97860
rect 635096 97572 635148 97578
rect 635096 97514 635148 97520
rect 635292 95826 635320 97854
rect 635752 97714 635780 100014
rect 635740 97708 635792 97714
rect 635740 97650 635792 97656
rect 636120 96762 636148 100014
rect 636384 97844 636436 97850
rect 636384 97786 636436 97792
rect 636108 96756 636160 96762
rect 636108 96698 636160 96704
rect 636396 95826 636424 97786
rect 637040 97782 637068 100014
rect 637028 97776 637080 97782
rect 637028 97718 637080 97724
rect 637500 97646 637528 100014
rect 638328 97986 638356 100014
rect 637580 97980 637632 97986
rect 637580 97922 637632 97928
rect 638316 97980 638368 97986
rect 638316 97922 638368 97928
rect 637488 97640 637540 97646
rect 637488 97582 637540 97588
rect 637592 95826 637620 97922
rect 638880 96558 638908 100014
rect 639052 97572 639104 97578
rect 639052 97514 639104 97520
rect 638868 96552 638920 96558
rect 638868 96494 638920 96500
rect 632992 95798 633328 95826
rect 634096 95798 634432 95826
rect 635292 95798 635628 95826
rect 636396 95798 636732 95826
rect 637592 95798 637928 95826
rect 639064 95690 639092 97514
rect 639616 95946 639644 100014
rect 639880 97708 639932 97714
rect 639880 97650 639932 97656
rect 639604 95940 639656 95946
rect 639604 95882 639656 95888
rect 639892 95826 639920 97650
rect 640260 96626 640288 100014
rect 640996 96898 641024 100014
rect 640984 96892 641036 96898
rect 640984 96834 641036 96840
rect 640984 96756 641036 96762
rect 640984 96698 641036 96704
rect 640248 96620 640300 96626
rect 640248 96562 640300 96568
rect 640996 95826 641024 96698
rect 641640 95878 641668 100014
rect 641732 100014 641976 100042
rect 642284 100014 642620 100042
rect 643264 100014 643600 100042
rect 643908 100014 644428 100042
rect 644552 100014 644888 100042
rect 645196 100014 645716 100042
rect 645840 100014 646176 100042
rect 646484 100014 646820 100042
rect 647220 100014 647556 100042
rect 647864 100014 648200 100042
rect 648508 100014 648568 100042
rect 649152 100014 649488 100042
rect 649796 100014 649948 100042
rect 650440 100014 650776 100042
rect 651084 100014 651328 100042
rect 651728 100014 652064 100042
rect 652372 100014 652708 100042
rect 653016 100014 653352 100042
rect 653752 100014 653996 100042
rect 654396 100014 654732 100042
rect 655040 100014 655376 100042
rect 655684 100014 656020 100042
rect 656328 100014 656664 100042
rect 656972 100014 657308 100042
rect 641732 96665 641760 100014
rect 642180 97776 642232 97782
rect 642180 97718 642232 97724
rect 641718 96656 641774 96665
rect 641718 96591 641774 96600
rect 641628 95872 641680 95878
rect 639892 95798 640228 95826
rect 640996 95798 641332 95826
rect 641628 95814 641680 95820
rect 642192 95826 642220 97718
rect 642284 96529 642312 100014
rect 643572 97510 643600 100014
rect 643560 97504 643612 97510
rect 643560 97446 643612 97452
rect 643284 96892 643336 96898
rect 643284 96834 643336 96840
rect 643192 96620 643244 96626
rect 643192 96562 643244 96568
rect 643100 96552 643152 96558
rect 642270 96520 642326 96529
rect 643100 96494 643152 96500
rect 642270 96455 642326 96464
rect 642192 95798 642528 95826
rect 632132 95662 632192 95690
rect 639032 95662 639092 95690
rect 627826 94480 627882 94489
rect 627826 94415 627882 94424
rect 626538 93528 626594 93537
rect 626538 93463 626594 93472
rect 626446 91624 626502 91633
rect 626446 91559 626502 91568
rect 625986 90672 626042 90681
rect 625986 90607 626042 90616
rect 625802 89720 625858 89729
rect 625802 89655 625858 89664
rect 626448 89684 626500 89690
rect 626448 89626 626500 89632
rect 626460 88913 626488 89626
rect 643112 89593 643140 96494
rect 643098 89584 643154 89593
rect 643098 89519 643154 89528
rect 626446 88904 626502 88913
rect 626446 88839 626502 88848
rect 626448 88324 626500 88330
rect 626448 88266 626500 88272
rect 626356 88256 626408 88262
rect 626356 88198 626408 88204
rect 626368 87009 626396 88198
rect 626460 87961 626488 88266
rect 626446 87952 626502 87961
rect 626446 87887 626502 87896
rect 626354 87000 626410 87009
rect 626354 86935 626410 86944
rect 626448 86284 626500 86290
rect 626448 86226 626500 86232
rect 626460 86057 626488 86226
rect 626446 86048 626502 86057
rect 626446 85983 626502 85992
rect 626448 85536 626500 85542
rect 626448 85478 626500 85484
rect 626460 85105 626488 85478
rect 643204 85241 643232 96562
rect 643190 85232 643246 85241
rect 643190 85167 643246 85176
rect 626446 85096 626502 85105
rect 626446 85031 626502 85040
rect 625620 84176 625672 84182
rect 625618 84144 625620 84153
rect 625672 84144 625674 84153
rect 625618 84079 625674 84088
rect 626448 84108 626500 84114
rect 626448 84050 626500 84056
rect 626460 83201 626488 84050
rect 626446 83192 626502 83201
rect 626446 83127 626502 83136
rect 643296 82249 643324 96834
rect 644400 92478 644428 100014
rect 644664 97980 644716 97986
rect 644664 97922 644716 97928
rect 644572 97640 644624 97646
rect 644572 97582 644624 97588
rect 644480 95940 644532 95946
rect 644480 95882 644532 95888
rect 644388 92472 644440 92478
rect 644388 92414 644440 92420
rect 644492 87145 644520 95882
rect 644584 94625 644612 97582
rect 644570 94616 644626 94625
rect 644570 94551 644626 94560
rect 644676 92177 644704 97922
rect 644860 96966 644888 100014
rect 644848 96960 644900 96966
rect 644848 96902 644900 96908
rect 644662 92168 644718 92177
rect 644662 92103 644718 92112
rect 644478 87136 644534 87145
rect 644478 87071 644534 87080
rect 645688 86630 645716 100014
rect 646044 97436 646096 97442
rect 646044 97378 646096 97384
rect 645860 95872 645912 95878
rect 645860 95814 645912 95820
rect 645676 86624 645728 86630
rect 645676 86566 645728 86572
rect 626446 82240 626502 82249
rect 626446 82175 626502 82184
rect 643282 82240 643338 82249
rect 643282 82175 643338 82184
rect 626460 78198 626488 82175
rect 631520 80974 631856 81002
rect 638972 80974 639308 81002
rect 629206 80880 629262 80889
rect 629206 80815 629262 80824
rect 626448 78192 626500 78198
rect 626448 78134 626500 78140
rect 629220 78062 629248 80815
rect 631048 78124 631100 78130
rect 631048 78066 631100 78072
rect 629208 78056 629260 78062
rect 629208 77998 629260 78004
rect 628380 77648 628432 77654
rect 628380 77590 628432 77596
rect 628392 77382 628420 77590
rect 628380 77376 628432 77382
rect 628380 77318 628432 77324
rect 624424 76560 624476 76566
rect 624424 76502 624476 76508
rect 628392 75290 628420 77318
rect 631060 77314 631088 78066
rect 631520 77654 631548 80974
rect 638972 78130 639000 80974
rect 642456 78192 642508 78198
rect 642456 78134 642508 78140
rect 638960 78124 639012 78130
rect 638960 78066 639012 78072
rect 636752 77988 636804 77994
rect 636752 77930 636804 77936
rect 633898 77888 633954 77897
rect 633898 77823 633954 77832
rect 631508 77648 631560 77654
rect 631508 77590 631560 77596
rect 631048 77308 631100 77314
rect 631048 77250 631100 77256
rect 631060 75290 631088 77250
rect 633912 75290 633940 77823
rect 636764 75290 636792 77930
rect 639602 77752 639658 77761
rect 639602 77687 639658 77696
rect 639616 75290 639644 77687
rect 642468 75290 642496 78134
rect 645308 78056 645360 78062
rect 645308 77998 645360 78004
rect 645320 75290 645348 77998
rect 623688 75268 623740 75274
rect 628176 75262 628420 75290
rect 631028 75262 631088 75290
rect 633880 75276 633940 75290
rect 633866 75262 633940 75276
rect 636732 75262 636792 75290
rect 639584 75276 639644 75290
rect 639570 75262 639644 75276
rect 642436 75262 642496 75290
rect 645288 75262 645348 75290
rect 623688 75210 623740 75216
rect 623778 74760 623834 74769
rect 623778 74695 623834 74704
rect 633530 74760 633586 74769
rect 633866 74746 633894 75262
rect 639234 75168 639290 75177
rect 639570 75154 639598 75262
rect 639290 75140 639598 75154
rect 639290 75126 639584 75140
rect 639234 75103 639290 75112
rect 633586 74732 633894 74746
rect 633586 74718 633880 74732
rect 633530 74695 633586 74704
rect 623792 70446 623820 74695
rect 623044 70440 623096 70446
rect 623044 70382 623096 70388
rect 623780 70440 623832 70446
rect 623780 70382 623832 70388
rect 623056 59906 623084 70382
rect 645872 64874 645900 95814
rect 646056 66042 646084 97378
rect 646148 95946 646176 100014
rect 646504 96960 646556 96966
rect 646504 96902 646556 96908
rect 646136 95940 646188 95946
rect 646136 95882 646188 95888
rect 646516 93158 646544 96902
rect 646792 96082 646820 100014
rect 647528 97850 647556 100014
rect 647516 97844 647568 97850
rect 647516 97786 647568 97792
rect 648172 97374 648200 100014
rect 648160 97368 648212 97374
rect 648160 97310 648212 97316
rect 647424 97232 647476 97238
rect 647424 97174 647476 97180
rect 646780 96076 646832 96082
rect 646780 96018 646832 96024
rect 646504 93152 646556 93158
rect 646504 93094 646556 93100
rect 646320 76628 646372 76634
rect 646320 76570 646372 76576
rect 646136 75268 646188 75274
rect 646136 75210 646188 75216
rect 646148 71777 646176 75210
rect 646332 74526 646360 76570
rect 646964 76560 647016 76566
rect 646964 76502 647016 76508
rect 646872 75200 646924 75206
rect 646872 75142 646924 75148
rect 646320 74520 646372 74526
rect 646884 74497 646912 75142
rect 646320 74462 646372 74468
rect 646870 74488 646926 74497
rect 646870 74423 646926 74432
rect 646976 73001 647004 76502
rect 647240 74520 647292 74526
rect 647240 74462 647292 74468
rect 646962 72992 647018 73001
rect 646962 72927 647018 72936
rect 646134 71768 646190 71777
rect 646134 71703 646190 71712
rect 647252 70009 647280 74462
rect 647238 70000 647294 70009
rect 647238 69935 647294 69944
rect 647436 67017 647464 97174
rect 648540 86562 648568 100014
rect 649460 97442 649488 100014
rect 649448 97436 649500 97442
rect 649448 97378 649500 97384
rect 648804 97300 648856 97306
rect 648804 97242 648856 97248
rect 648528 86556 648580 86562
rect 648528 86498 648580 86504
rect 648816 68513 648844 97242
rect 649920 86834 649948 100014
rect 650748 96966 650776 100014
rect 650736 96960 650788 96966
rect 650736 96902 650788 96908
rect 651196 96960 651248 96966
rect 651196 96902 651248 96908
rect 649908 86828 649960 86834
rect 649908 86770 649960 86776
rect 651208 86766 651236 96902
rect 651300 86902 651328 100014
rect 652036 97306 652064 100014
rect 652024 97300 652076 97306
rect 652024 97242 652076 97248
rect 651288 86896 651340 86902
rect 651288 86838 651340 86844
rect 651196 86760 651248 86766
rect 651196 86702 651248 86708
rect 652680 86698 652708 100014
rect 653324 96014 653352 100014
rect 653312 96008 653364 96014
rect 653312 95950 653364 95956
rect 652668 86692 652720 86698
rect 652668 86634 652720 86640
rect 653968 86494 653996 100014
rect 654704 97238 654732 100014
rect 654784 97844 654836 97850
rect 654784 97786 654836 97792
rect 654692 97232 654744 97238
rect 654692 97174 654744 97180
rect 654796 92585 654824 97786
rect 655348 93401 655376 100014
rect 655428 96960 655480 96966
rect 655428 96902 655480 96908
rect 655334 93392 655390 93401
rect 655334 93327 655390 93336
rect 654876 93152 654928 93158
rect 654876 93094 654928 93100
rect 654782 92576 654838 92585
rect 654782 92511 654838 92520
rect 654324 92472 654376 92478
rect 654324 92414 654376 92420
rect 654336 91497 654364 92414
rect 654322 91488 654378 91497
rect 654322 91423 654378 91432
rect 654888 90681 654916 93094
rect 654874 90672 654930 90681
rect 654874 90607 654930 90616
rect 655440 89865 655468 96902
rect 655992 96830 656020 100014
rect 655980 96824 656032 96830
rect 655980 96766 656032 96772
rect 656636 96218 656664 100014
rect 656808 96620 656860 96626
rect 656808 96562 656860 96568
rect 656624 96212 656676 96218
rect 656624 96154 656676 96160
rect 655426 89856 655482 89865
rect 655426 89791 655482 89800
rect 656820 88874 656848 96562
rect 657280 95266 657308 100014
rect 657372 100014 657616 100042
rect 658260 100014 658320 100042
rect 658904 100014 659240 100042
rect 657268 95260 657320 95266
rect 657268 95202 657320 95208
rect 657372 94761 657400 100014
rect 657728 97164 657780 97170
rect 657728 97106 657780 97112
rect 657740 95132 657768 97106
rect 658292 96626 658320 100014
rect 658832 97436 658884 97442
rect 658832 97378 658884 97384
rect 658372 97232 658424 97238
rect 658372 97174 658424 97180
rect 658280 96620 658332 96626
rect 658280 96562 658332 96568
rect 658384 95146 658412 97174
rect 658306 95118 658412 95146
rect 658844 95132 658872 97378
rect 659212 97238 659240 100014
rect 659304 100014 659548 100042
rect 660284 100014 660620 100042
rect 659200 97232 659252 97238
rect 659200 97174 659252 97180
rect 659304 96966 659332 100014
rect 660396 97504 660448 97510
rect 660396 97446 660448 97452
rect 660120 97368 660172 97374
rect 660120 97310 660172 97316
rect 659292 96960 659344 96966
rect 659292 96902 659344 96908
rect 659568 96824 659620 96830
rect 659568 96766 659620 96772
rect 659580 95132 659608 96766
rect 660132 95132 660160 97310
rect 660408 95146 660436 97446
rect 660592 96898 660620 100014
rect 660684 100014 660928 100042
rect 661572 100014 661908 100042
rect 662216 100014 662368 100042
rect 662860 100014 663104 100042
rect 660684 97170 660712 100014
rect 660672 97164 660724 97170
rect 660672 97106 660724 97112
rect 660580 96892 660632 96898
rect 660580 96834 660632 96840
rect 661408 96892 661460 96898
rect 661408 96834 661460 96840
rect 660408 95118 660698 95146
rect 661420 95132 661448 96834
rect 661880 96762 661908 100014
rect 661960 97300 662012 97306
rect 661960 97242 662012 97248
rect 661868 96756 661920 96762
rect 661868 96698 661920 96704
rect 661972 95132 662000 97242
rect 662340 97170 662368 100014
rect 663076 97986 663104 100014
rect 663168 100014 663504 100042
rect 663064 97980 663116 97986
rect 663064 97922 663116 97928
rect 662512 97232 662564 97238
rect 662512 97174 662564 97180
rect 662328 97164 662380 97170
rect 662328 97106 662380 97112
rect 662524 95132 662552 97174
rect 663064 96756 663116 96762
rect 663064 96698 663116 96704
rect 663076 95132 663104 96698
rect 657358 94752 657414 94761
rect 657358 94687 657414 94696
rect 658108 88874 658306 88890
rect 656808 88868 656860 88874
rect 656808 88810 656860 88816
rect 658096 88868 658306 88874
rect 658148 88862 658306 88868
rect 661986 88874 662368 88890
rect 661986 88868 662380 88874
rect 661986 88862 662328 88868
rect 658096 88810 658148 88816
rect 662328 88810 662380 88816
rect 659488 88330 659594 88346
rect 663168 88330 663196 100014
rect 665364 97980 665416 97986
rect 665364 97922 665416 97928
rect 663984 97164 664036 97170
rect 663984 97106 664036 97112
rect 663892 96212 663944 96218
rect 663892 96154 663944 96160
rect 663800 96076 663852 96082
rect 663800 96018 663852 96024
rect 663812 92585 663840 96018
rect 663798 92576 663854 92585
rect 663798 92511 663854 92520
rect 663904 90681 663932 96154
rect 663890 90672 663946 90681
rect 663890 90607 663946 90616
rect 663996 88874 664024 97106
rect 665272 96008 665324 96014
rect 665272 95950 665324 95956
rect 665180 95940 665232 95946
rect 665180 95882 665232 95888
rect 664076 95260 664128 95266
rect 664076 95202 664128 95208
rect 664088 89049 664116 95202
rect 665192 91769 665220 95882
rect 665178 91760 665234 91769
rect 665178 91695 665234 91704
rect 665284 89865 665312 95950
rect 665376 93401 665404 97922
rect 665362 93392 665418 93401
rect 665362 93327 665418 93336
rect 665270 89856 665326 89865
rect 665270 89791 665326 89800
rect 664074 89040 664130 89049
rect 664074 88975 664130 88984
rect 663984 88868 664036 88874
rect 663984 88810 664036 88816
rect 659476 88324 659594 88330
rect 659528 88318 659594 88324
rect 663156 88324 663208 88330
rect 659476 88266 659528 88272
rect 663156 88266 663208 88272
rect 657188 86902 657216 88196
rect 657176 86896 657228 86902
rect 657176 86838 657228 86844
rect 657740 86766 657768 88196
rect 657728 86760 657780 86766
rect 657728 86702 657780 86708
rect 658844 86494 658872 88196
rect 660132 86630 660160 88196
rect 660684 86834 660712 88196
rect 660672 86828 660724 86834
rect 660672 86770 660724 86776
rect 660120 86624 660172 86630
rect 660120 86566 660172 86572
rect 661420 86562 661448 88196
rect 662524 86698 662552 88196
rect 662512 86692 662564 86698
rect 662512 86634 662564 86640
rect 661408 86556 661460 86562
rect 661408 86498 661460 86504
rect 653956 86488 654008 86494
rect 653956 86430 654008 86436
rect 658832 86488 658884 86494
rect 658832 86430 658884 86436
rect 648802 68504 648858 68513
rect 648802 68439 648858 68448
rect 647422 67008 647478 67017
rect 647422 66943 647478 66952
rect 646134 66056 646190 66065
rect 646056 66014 646134 66042
rect 646134 65991 646190 66000
rect 645872 64846 646176 64874
rect 646148 64433 646176 64846
rect 646134 64424 646190 64433
rect 646134 64359 646190 64368
rect 623044 59900 623096 59906
rect 623044 59842 623096 59848
rect 621664 58676 621716 58682
rect 621664 58618 621716 58624
rect 662420 58676 662472 58682
rect 662420 58618 662472 58624
rect 616328 53848 616380 53854
rect 616328 53790 616380 53796
rect 618904 53848 618956 53854
rect 618904 53790 618956 53796
rect 616340 52426 616368 53790
rect 616328 52420 616380 52426
rect 616328 52362 616380 52368
rect 661130 47560 661186 47569
rect 661130 47495 661186 47504
rect 648104 47126 649670 47188
rect 648104 46658 648157 47126
rect 649617 46658 649670 47126
rect 648104 46590 649670 46658
rect 612830 46336 612886 46345
rect 612830 46271 612886 46280
rect 612738 46200 612794 46209
rect 612738 46135 612794 46144
rect 661144 44849 661172 47495
rect 662432 47433 662460 58618
rect 669976 49094 670004 961862
rect 672736 938738 672764 975666
rect 675772 966521 675800 966723
rect 675758 966512 675814 966521
rect 675758 966447 675814 966456
rect 675758 966240 675814 966249
rect 675758 966175 675814 966184
rect 675772 966076 675800 966175
rect 675772 965025 675800 965435
rect 675758 965016 675814 965025
rect 675758 964951 675814 964960
rect 675772 963393 675800 963595
rect 675758 963384 675814 963393
rect 675758 963319 675814 963328
rect 675680 962849 675708 963016
rect 675666 962840 675722 962849
rect 675666 962775 675722 962784
rect 674840 961920 674892 961926
rect 675496 961897 675524 962404
rect 675482 961888 675538 961897
rect 674892 961868 675142 961874
rect 674840 961862 675142 961868
rect 674852 961846 675142 961862
rect 675482 961823 675538 961832
rect 675404 961382 675432 961755
rect 675024 961376 675076 961382
rect 675024 961318 675076 961324
rect 675392 961376 675444 961382
rect 675392 961318 675444 961324
rect 674748 958248 674800 958254
rect 674748 958190 674800 958196
rect 673368 957024 673420 957030
rect 673368 956966 673420 956972
rect 673184 956140 673236 956146
rect 673184 956082 673236 956088
rect 672724 938732 672776 938738
rect 672724 938674 672776 938680
rect 672356 935808 672408 935814
rect 672356 935750 672408 935756
rect 671344 927444 671396 927450
rect 671344 927386 671396 927392
rect 670056 921868 670108 921874
rect 670056 921810 670108 921816
rect 670068 760850 670096 921810
rect 670608 788044 670660 788050
rect 670608 787986 670660 787992
rect 670056 760844 670108 760850
rect 670056 760786 670108 760792
rect 670056 749420 670108 749426
rect 670056 749362 670108 749368
rect 670068 178838 670096 749362
rect 670620 711278 670648 787986
rect 670608 711272 670660 711278
rect 670608 711214 670660 711220
rect 670148 703860 670200 703866
rect 670148 703802 670200 703808
rect 670056 178832 670108 178838
rect 670056 178774 670108 178780
rect 670160 173670 670188 703802
rect 670608 686112 670660 686118
rect 670608 686054 670660 686060
rect 670620 621178 670648 686054
rect 670608 621172 670660 621178
rect 670608 621114 670660 621120
rect 670240 392012 670292 392018
rect 670240 391954 670292 391960
rect 670148 173664 670200 173670
rect 670148 173606 670200 173612
rect 670252 143342 670280 391954
rect 671356 184210 671384 927386
rect 671436 869440 671488 869446
rect 671436 869382 671488 869388
rect 671448 716174 671476 869382
rect 672172 773628 672224 773634
rect 672172 773570 672224 773576
rect 671988 743232 672040 743238
rect 671988 743174 672040 743180
rect 671436 716168 671488 716174
rect 671436 716110 671488 716116
rect 671436 709368 671488 709374
rect 671436 709310 671488 709316
rect 671448 579970 671476 709310
rect 671896 698216 671948 698222
rect 671896 698158 671948 698164
rect 671908 621314 671936 698158
rect 672000 665378 672028 743174
rect 672184 710054 672212 773570
rect 672368 759121 672396 935750
rect 672816 935740 672868 935746
rect 672816 935682 672868 935688
rect 672724 803208 672776 803214
rect 672724 803150 672776 803156
rect 672632 786752 672684 786758
rect 672632 786694 672684 786700
rect 672540 780768 672592 780774
rect 672540 780710 672592 780716
rect 672448 777368 672500 777374
rect 672448 777310 672500 777316
rect 672354 759112 672410 759121
rect 672264 759076 672316 759082
rect 672354 759047 672410 759056
rect 672264 759018 672316 759024
rect 672276 714542 672304 759018
rect 672356 742552 672408 742558
rect 672356 742494 672408 742500
rect 672264 714536 672316 714542
rect 672264 714478 672316 714484
rect 672264 714060 672316 714066
rect 672264 714002 672316 714008
rect 672172 710048 672224 710054
rect 672172 709990 672224 709996
rect 672276 669730 672304 714002
rect 672264 669724 672316 669730
rect 672264 669666 672316 669672
rect 672264 666596 672316 666602
rect 672264 666538 672316 666544
rect 671988 665372 672040 665378
rect 671988 665314 672040 665320
rect 671988 652792 672040 652798
rect 671988 652734 672040 652740
rect 671896 621308 671948 621314
rect 671896 621250 671948 621256
rect 671436 579964 671488 579970
rect 671436 579906 671488 579912
rect 672000 575618 672028 652734
rect 672276 622742 672304 666538
rect 672368 664018 672396 742494
rect 672460 708422 672488 777310
rect 672552 710462 672580 780710
rect 672644 712094 672672 786694
rect 672632 712088 672684 712094
rect 672632 712030 672684 712036
rect 672540 710456 672592 710462
rect 672540 710398 672592 710404
rect 672448 708416 672500 708422
rect 672448 708358 672500 708364
rect 672632 690464 672684 690470
rect 672632 690406 672684 690412
rect 672540 684276 672592 684282
rect 672540 684218 672592 684224
rect 672356 664012 672408 664018
rect 672356 663954 672408 663960
rect 672356 623892 672408 623898
rect 672356 623834 672408 623840
rect 672264 622736 672316 622742
rect 672264 622678 672316 622684
rect 672264 622464 672316 622470
rect 672264 622406 672316 622412
rect 672276 577046 672304 622406
rect 672368 578270 672396 623834
rect 672448 623824 672500 623830
rect 672448 623766 672500 623772
rect 672460 580106 672488 623766
rect 672552 619818 672580 684218
rect 672644 619954 672672 690406
rect 672736 670954 672764 803150
rect 672828 758441 672856 935682
rect 673196 931666 673224 956082
rect 673184 931660 673236 931666
rect 673184 931602 673236 931608
rect 673380 930306 673408 956966
rect 674196 948116 674248 948122
rect 674196 948058 674248 948064
rect 674208 939214 674236 948058
rect 674196 939208 674248 939214
rect 674196 939150 674248 939156
rect 674656 938324 674708 938330
rect 674656 938266 674708 938272
rect 673828 937508 673880 937514
rect 673828 937450 673880 937456
rect 673368 930300 673420 930306
rect 673368 930242 673420 930248
rect 673184 872704 673236 872710
rect 673184 872646 673236 872652
rect 673000 869712 673052 869718
rect 673000 869654 673052 869660
rect 672908 862844 672960 862850
rect 672908 862786 672960 862792
rect 672814 758432 672870 758441
rect 672814 758367 672870 758376
rect 672920 755002 672948 862786
rect 672908 754996 672960 755002
rect 672908 754938 672960 754944
rect 673012 752282 673040 869654
rect 673092 869644 673144 869650
rect 673092 869586 673144 869592
rect 673000 752276 673052 752282
rect 673000 752218 673052 752224
rect 673104 750922 673132 869586
rect 673196 753642 673224 872646
rect 673276 782944 673328 782950
rect 673276 782886 673328 782892
rect 673184 753636 673236 753642
rect 673184 753578 673236 753584
rect 673092 750916 673144 750922
rect 673092 750858 673144 750864
rect 672816 749488 672868 749494
rect 672816 749430 672868 749436
rect 672724 670948 672776 670954
rect 672724 670890 672776 670896
rect 672724 667956 672776 667962
rect 672724 667898 672776 667904
rect 672736 622606 672764 667898
rect 672828 625530 672856 749430
rect 673184 739152 673236 739158
rect 673184 739094 673236 739100
rect 673092 735004 673144 735010
rect 673092 734946 673144 734952
rect 672908 714876 672960 714882
rect 672908 714818 672960 714824
rect 672920 669594 672948 714818
rect 673000 688696 673052 688702
rect 673000 688638 673052 688644
rect 672908 669588 672960 669594
rect 672908 669530 672960 669536
rect 672908 645584 672960 645590
rect 672908 645526 672960 645532
rect 672816 625524 672868 625530
rect 672816 625466 672868 625472
rect 672724 622600 672776 622606
rect 672724 622542 672776 622548
rect 672632 619948 672684 619954
rect 672632 619890 672684 619896
rect 672540 619812 672592 619818
rect 672540 619754 672592 619760
rect 672724 614168 672776 614174
rect 672724 614110 672776 614116
rect 672632 595332 672684 595338
rect 672632 595274 672684 595280
rect 672448 580100 672500 580106
rect 672448 580042 672500 580048
rect 672356 578264 672408 578270
rect 672356 578206 672408 578212
rect 672264 577040 672316 577046
rect 672264 576982 672316 576988
rect 672540 576972 672592 576978
rect 672540 576914 672592 576920
rect 672448 576904 672500 576910
rect 672448 576846 672500 576852
rect 671988 575612 672040 575618
rect 671988 575554 672040 575560
rect 671988 561944 672040 561950
rect 671988 561886 672040 561892
rect 672000 484430 672028 561886
rect 672460 532914 672488 576846
rect 672448 532908 672500 532914
rect 672448 532850 672500 532856
rect 672552 531350 672580 576914
rect 672540 531344 672592 531350
rect 672540 531286 672592 531292
rect 672644 530058 672672 595274
rect 672632 530052 672684 530058
rect 672632 529994 672684 530000
rect 671988 484424 672040 484430
rect 671988 484366 672040 484372
rect 671528 456816 671580 456822
rect 671528 456758 671580 456764
rect 671436 390584 671488 390590
rect 671436 390526 671488 390532
rect 671448 223174 671476 390526
rect 671540 313546 671568 456758
rect 671620 324352 671672 324358
rect 671620 324294 671672 324300
rect 671528 313540 671580 313546
rect 671528 313482 671580 313488
rect 671528 284368 671580 284374
rect 671528 284310 671580 284316
rect 671436 223168 671488 223174
rect 671436 223110 671488 223116
rect 671436 211200 671488 211206
rect 671436 211142 671488 211148
rect 671344 184204 671396 184210
rect 671344 184146 671396 184152
rect 671344 167068 671396 167074
rect 671344 167010 671396 167016
rect 670240 143336 670292 143342
rect 670240 143278 670292 143284
rect 670148 121508 670200 121514
rect 670148 121450 670200 121456
rect 670056 120760 670108 120766
rect 670056 120702 670108 120708
rect 670068 110362 670096 120702
rect 670160 111314 670188 121450
rect 671356 114374 671384 167010
rect 671448 123894 671476 211142
rect 671540 132802 671568 284310
rect 671632 176866 671660 324294
rect 672632 221876 672684 221882
rect 672632 221818 672684 221824
rect 672540 221060 672592 221066
rect 672540 221002 672592 221008
rect 671620 176860 671672 176866
rect 671620 176802 671672 176808
rect 672552 176526 672580 221002
rect 672644 177002 672672 221818
rect 672632 176996 672684 177002
rect 672632 176938 672684 176944
rect 672540 176520 672592 176526
rect 672540 176462 672592 176468
rect 672736 164014 672764 614110
rect 672816 593428 672868 593434
rect 672816 593370 672868 593376
rect 672828 528698 672856 593370
rect 672920 574258 672948 645526
rect 673012 615534 673040 688638
rect 673104 661162 673132 734946
rect 673196 663814 673224 739094
rect 673288 707606 673316 782886
rect 673644 780020 673696 780026
rect 673644 779962 673696 779968
rect 673368 759144 673420 759150
rect 673368 759086 673420 759092
rect 673380 715358 673408 759086
rect 673368 715352 673420 715358
rect 673368 715294 673420 715300
rect 673460 713244 673512 713250
rect 673460 713186 673512 713192
rect 673276 707600 673328 707606
rect 673276 707542 673328 707548
rect 673276 692980 673328 692986
rect 673276 692922 673328 692928
rect 673184 663808 673236 663814
rect 673184 663750 673236 663756
rect 673092 661156 673144 661162
rect 673092 661098 673144 661104
rect 673184 647760 673236 647766
rect 673184 647702 673236 647708
rect 673092 643408 673144 643414
rect 673092 643350 673144 643356
rect 673000 615528 673052 615534
rect 673000 615470 673052 615476
rect 672908 574252 672960 574258
rect 672908 574194 672960 574200
rect 673104 569974 673132 643350
rect 673196 571538 673224 647702
rect 673288 616894 673316 692922
rect 673368 687336 673420 687342
rect 673368 687278 673420 687284
rect 673380 617098 673408 687278
rect 673472 668710 673500 713186
rect 673552 712428 673604 712434
rect 673552 712370 673604 712376
rect 673460 668704 673512 668710
rect 673460 668646 673512 668652
rect 673564 667894 673592 712370
rect 673656 707198 673684 779962
rect 673840 759558 673868 937450
rect 674472 873588 674524 873594
rect 674472 873530 674524 873536
rect 674288 869848 674340 869854
rect 674288 869790 674340 869796
rect 674196 787364 674248 787370
rect 674196 787306 674248 787312
rect 674012 784304 674064 784310
rect 674012 784246 674064 784252
rect 673920 778660 673972 778666
rect 673920 778602 673972 778608
rect 673828 759552 673880 759558
rect 673828 759494 673880 759500
rect 673736 738268 673788 738274
rect 673736 738210 673788 738216
rect 673644 707192 673696 707198
rect 673644 707134 673696 707140
rect 673552 667888 673604 667894
rect 673552 667830 673604 667836
rect 673748 662386 673776 738210
rect 673828 728680 673880 728686
rect 673828 728622 673880 728628
rect 673840 665038 673868 728622
rect 673932 706790 673960 778602
rect 674024 709238 674052 784246
rect 674208 709646 674236 787306
rect 674300 755614 674328 869790
rect 674380 868556 674432 868562
rect 674380 868498 674432 868504
rect 674288 755608 674340 755614
rect 674288 755550 674340 755556
rect 674392 753166 674420 868498
rect 674484 754390 674512 873530
rect 674564 872228 674616 872234
rect 674564 872170 674616 872176
rect 674472 754384 674524 754390
rect 674472 754326 674524 754332
rect 674380 753160 674432 753166
rect 674380 753102 674432 753108
rect 674576 752758 674604 872170
rect 674668 760374 674696 938266
rect 674760 930782 674788 958190
rect 675036 957953 675064 961318
rect 675772 959177 675800 959276
rect 675758 959168 675814 959177
rect 675758 959103 675814 959112
rect 675404 958254 675432 958732
rect 675392 958248 675444 958254
rect 675392 958190 675444 958196
rect 675022 957944 675078 957953
rect 675022 957879 675078 957888
rect 675024 957840 675076 957846
rect 675772 957817 675800 958052
rect 675024 957782 675076 957788
rect 675758 957808 675814 957817
rect 675036 955534 675064 957782
rect 675758 957743 675814 957752
rect 675404 957030 675432 957440
rect 675392 957024 675444 957030
rect 675392 956966 675444 956972
rect 675496 956146 675524 956216
rect 675484 956140 675536 956146
rect 675484 956082 675536 956088
rect 675024 955528 675076 955534
rect 675024 955470 675076 955476
rect 675484 955528 675536 955534
rect 675484 955470 675536 955476
rect 675496 955060 675524 955470
rect 675404 954009 675432 954380
rect 675390 954000 675446 954009
rect 675390 953935 675446 953944
rect 675772 952066 675800 952544
rect 675760 952060 675812 952066
rect 675760 952002 675812 952008
rect 675760 951788 675812 951794
rect 675760 951730 675812 951736
rect 675772 949482 675800 951730
rect 679806 949784 679862 949793
rect 679806 949719 679862 949728
rect 679622 949648 679678 949657
rect 679622 949583 679678 949592
rect 676862 949512 676918 949521
rect 675760 949476 675812 949482
rect 676862 949447 676918 949456
rect 678244 949476 678296 949482
rect 675760 949418 675812 949424
rect 676034 939992 676090 940001
rect 676034 939927 676090 939936
rect 676048 939826 676076 939927
rect 676036 939820 676088 939826
rect 676036 939762 676088 939768
rect 676218 939312 676274 939321
rect 676218 939247 676274 939256
rect 676036 939208 676088 939214
rect 676034 939176 676036 939185
rect 676088 939176 676090 939185
rect 676034 939111 676090 939120
rect 676034 938768 676090 938777
rect 676232 938738 676260 939247
rect 676034 938703 676090 938712
rect 676220 938732 676272 938738
rect 676048 938602 676076 938703
rect 676220 938674 676272 938680
rect 676036 938596 676088 938602
rect 676036 938538 676088 938544
rect 676034 938360 676090 938369
rect 676034 938295 676036 938304
rect 676088 938295 676090 938304
rect 676036 938266 676088 938272
rect 676218 937680 676274 937689
rect 676218 937615 676274 937624
rect 676034 937544 676090 937553
rect 676034 937479 676036 937488
rect 676088 937479 676090 937488
rect 676036 937450 676088 937456
rect 676232 937378 676260 937615
rect 676220 937372 676272 937378
rect 676220 937314 676272 937320
rect 676218 937272 676274 937281
rect 676218 937207 676220 937216
rect 676272 937207 676274 937216
rect 676220 937178 676272 937184
rect 676126 936456 676182 936465
rect 676126 936391 676182 936400
rect 676034 935912 676090 935921
rect 676034 935847 676090 935856
rect 676048 935814 676076 935847
rect 676036 935808 676088 935814
rect 676036 935750 676088 935756
rect 676140 935746 676168 936391
rect 676218 936048 676274 936057
rect 676218 935983 676274 935992
rect 676128 935740 676180 935746
rect 676128 935682 676180 935688
rect 676232 935678 676260 935983
rect 676220 935672 676272 935678
rect 676220 935614 676272 935620
rect 676876 935241 676904 949447
rect 678244 949418 678296 949424
rect 676862 935232 676918 935241
rect 676862 935167 676918 935176
rect 678256 933609 678284 949418
rect 678242 933600 678298 933609
rect 678242 933535 678298 933544
rect 679636 932385 679664 949583
rect 679820 932793 679848 949719
rect 703694 940508 703722 940644
rect 704154 940508 704182 940644
rect 704614 940508 704642 940644
rect 705074 940508 705102 940644
rect 705534 940508 705562 940644
rect 705994 940508 706022 940644
rect 706454 940508 706482 940644
rect 706914 940508 706942 940644
rect 707374 940508 707402 940644
rect 707834 940508 707862 940644
rect 708294 940508 708322 940644
rect 708754 940508 708782 940644
rect 709214 940508 709242 940644
rect 679806 932784 679862 932793
rect 679806 932719 679862 932728
rect 679622 932376 679678 932385
rect 679622 932311 679678 932320
rect 676034 931832 676090 931841
rect 676034 931767 676090 931776
rect 676048 931666 676076 931767
rect 676036 931660 676088 931666
rect 676036 931602 676088 931608
rect 674748 930776 674800 930782
rect 676220 930776 676272 930782
rect 674748 930718 674800 930724
rect 676218 930744 676220 930753
rect 676272 930744 676274 930753
rect 676218 930679 676274 930688
rect 676218 930336 676274 930345
rect 676218 930271 676220 930280
rect 676272 930271 676274 930280
rect 676220 930242 676272 930248
rect 683118 929520 683174 929529
rect 683118 929455 683174 929464
rect 683132 928713 683160 929455
rect 683118 928704 683174 928713
rect 683118 928639 683174 928648
rect 683132 927450 683160 928639
rect 683120 927444 683172 927450
rect 683120 927386 683172 927392
rect 675404 877305 675432 877540
rect 675390 877296 675446 877305
rect 675390 877231 675446 877240
rect 675772 876625 675800 876860
rect 675758 876616 675814 876625
rect 675758 876551 675814 876560
rect 675772 875945 675800 876248
rect 675758 875936 675814 875945
rect 675758 875871 675814 875880
rect 675772 874041 675800 874412
rect 675758 874032 675814 874041
rect 675758 873967 675814 873976
rect 675404 873594 675432 873868
rect 675392 873588 675444 873594
rect 675392 873530 675444 873536
rect 675404 872710 675432 873188
rect 675392 872704 675444 872710
rect 675392 872646 675444 872652
rect 675404 872234 675432 872576
rect 675392 872228 675444 872234
rect 675392 872170 675444 872176
rect 675404 869854 675432 870060
rect 675392 869848 675444 869854
rect 675392 869790 675444 869796
rect 675392 869712 675444 869718
rect 675392 869654 675444 869660
rect 674932 869644 674984 869650
rect 674932 869586 674984 869592
rect 674944 868766 674972 869586
rect 675404 869516 675432 869654
rect 674932 868760 674984 868766
rect 674932 868702 674984 868708
rect 675392 868760 675444 868766
rect 675392 868702 675444 868708
rect 674932 868624 674984 868630
rect 674932 868566 674984 868572
rect 674944 866250 674972 868566
rect 675404 868224 675432 868702
rect 675496 868562 675524 868875
rect 675484 868556 675536 868562
rect 675484 868498 675536 868504
rect 675772 866833 675800 867035
rect 675758 866824 675814 866833
rect 675758 866759 675814 866768
rect 674932 866244 674984 866250
rect 674932 866186 674984 866192
rect 675392 866244 675444 866250
rect 675392 866186 675444 866192
rect 675404 865844 675432 866186
rect 675772 864793 675800 865195
rect 675758 864784 675814 864793
rect 675758 864719 675814 864728
rect 675496 862850 675524 863328
rect 675484 862844 675536 862850
rect 675484 862786 675536 862792
rect 675404 788050 675432 788324
rect 675392 788044 675444 788050
rect 675392 787986 675444 787992
rect 675404 787370 675432 787679
rect 675392 787364 675444 787370
rect 675392 787306 675444 787312
rect 675404 786758 675432 787032
rect 675392 786752 675444 786758
rect 675392 786694 675444 786700
rect 675496 784825 675524 785196
rect 675482 784816 675538 784825
rect 675482 784751 675538 784760
rect 675404 784310 675432 784652
rect 675392 784304 675444 784310
rect 675392 784246 675444 784252
rect 675758 784136 675814 784145
rect 675758 784071 675814 784080
rect 675772 783972 675800 784071
rect 675496 782950 675524 783360
rect 675484 782944 675536 782950
rect 675484 782886 675536 782892
rect 675496 780774 675524 780844
rect 675484 780768 675536 780774
rect 675484 780710 675536 780716
rect 675496 780026 675524 780300
rect 675484 780020 675536 780026
rect 675484 779962 675536 779968
rect 675390 779920 675446 779929
rect 675390 779855 675446 779864
rect 675404 779686 675432 779855
rect 674748 779000 674800 779006
rect 674748 778942 674800 778948
rect 674760 777102 674788 778942
rect 675496 778666 675524 779008
rect 675484 778660 675536 778666
rect 675484 778602 675536 778608
rect 675404 777374 675432 777852
rect 675392 777368 675444 777374
rect 675392 777310 675444 777316
rect 674748 777096 674800 777102
rect 674748 777038 674800 777044
rect 675392 777096 675444 777102
rect 675392 777038 675444 777044
rect 675404 776628 675432 777038
rect 675404 775713 675432 776016
rect 675390 775704 675446 775713
rect 675390 775639 675446 775648
rect 675496 773634 675524 774180
rect 675484 773628 675536 773634
rect 675484 773570 675536 773576
rect 675758 773392 675814 773401
rect 675758 773327 675814 773336
rect 674656 760368 674708 760374
rect 674656 760310 674708 760316
rect 674656 758260 674708 758266
rect 674656 758202 674708 758208
rect 674564 752752 674616 752758
rect 674564 752694 674616 752700
rect 674288 735684 674340 735690
rect 674288 735626 674340 735632
rect 674196 709640 674248 709646
rect 674196 709582 674248 709588
rect 674012 709232 674064 709238
rect 674012 709174 674064 709180
rect 673920 706784 673972 706790
rect 673920 706726 673972 706732
rect 673920 690056 673972 690062
rect 673920 689998 673972 690004
rect 673828 665032 673880 665038
rect 673828 664974 673880 664980
rect 673736 662380 673788 662386
rect 673736 662322 673788 662328
rect 673644 622260 673696 622266
rect 673644 622202 673696 622208
rect 673368 617092 673420 617098
rect 673368 617034 673420 617040
rect 673276 616888 673328 616894
rect 673276 616830 673328 616836
rect 673368 607640 673420 607646
rect 673368 607582 673420 607588
rect 673276 603084 673328 603090
rect 673276 603026 673328 603032
rect 673184 571532 673236 571538
rect 673184 571474 673236 571480
rect 673092 569968 673144 569974
rect 673092 569910 673144 569916
rect 673092 560244 673144 560250
rect 673092 560186 673144 560192
rect 673000 554804 673052 554810
rect 673000 554746 673052 554752
rect 672908 553512 672960 553518
rect 672908 553454 672960 553460
rect 672816 528692 672868 528698
rect 672816 528634 672868 528640
rect 672920 481778 672948 553454
rect 673012 481914 673040 554746
rect 673104 484634 673132 560186
rect 673184 557592 673236 557598
rect 673184 557534 673236 557540
rect 673092 484628 673144 484634
rect 673092 484570 673144 484576
rect 673196 483138 673224 557534
rect 673288 525978 673316 603026
rect 673380 528834 673408 607582
rect 673656 577454 673684 622202
rect 673932 617030 673960 689998
rect 674196 668908 674248 668914
rect 674196 668850 674248 668856
rect 674012 639124 674064 639130
rect 674012 639066 674064 639072
rect 673920 617024 673972 617030
rect 673920 616966 673972 616972
rect 673828 603492 673880 603498
rect 673828 603434 673880 603440
rect 673736 579284 673788 579290
rect 673736 579226 673788 579232
rect 673644 577448 673696 577454
rect 673644 577390 673696 577396
rect 673748 534954 673776 579226
rect 673736 534948 673788 534954
rect 673736 534890 673788 534896
rect 673368 528828 673420 528834
rect 673368 528770 673420 528776
rect 673840 528426 673868 603434
rect 673920 578604 673972 578610
rect 673920 578546 673972 578552
rect 673932 534138 673960 578546
rect 674024 574598 674052 639066
rect 674208 624374 674236 668850
rect 674300 665310 674328 735626
rect 674564 734392 674616 734398
rect 674564 734334 674616 734340
rect 674472 733644 674524 733650
rect 674472 733586 674524 733592
rect 674484 731414 674512 733586
rect 674576 732086 674604 734334
rect 674564 732080 674616 732086
rect 674564 732022 674616 732028
rect 674484 731386 674604 731414
rect 674472 730516 674524 730522
rect 674472 730458 674524 730464
rect 674380 689376 674432 689382
rect 674380 689318 674432 689324
rect 674288 665304 674340 665310
rect 674288 665246 674340 665252
rect 674288 644836 674340 644842
rect 674288 644778 674340 644784
rect 674196 624368 674248 624374
rect 674196 624310 674248 624316
rect 674196 598460 674248 598466
rect 674196 598402 674248 598408
rect 674012 574592 674064 574598
rect 674012 574534 674064 574540
rect 673920 534132 673972 534138
rect 673920 534074 673972 534080
rect 673828 528420 673880 528426
rect 673828 528362 673880 528368
rect 674208 526386 674236 598402
rect 674300 571742 674328 644778
rect 674392 617846 674420 689318
rect 674484 666534 674512 730458
rect 674472 666528 674524 666534
rect 674472 666470 674524 666476
rect 674576 661638 674604 731386
rect 674668 713726 674696 758202
rect 674746 757480 674802 757489
rect 674746 757415 674802 757424
rect 674656 713720 674708 713726
rect 674656 713662 674708 713668
rect 674760 712881 674788 757415
rect 675772 756265 675800 773327
rect 679622 772712 679678 772721
rect 679622 772647 679678 772656
rect 676126 761288 676182 761297
rect 676126 761223 676182 761232
rect 676034 760744 676090 760753
rect 676140 760714 676168 761223
rect 676218 760880 676274 760889
rect 676218 760815 676220 760824
rect 676272 760815 676274 760824
rect 676220 760786 676272 760792
rect 676034 760679 676090 760688
rect 676128 760708 676180 760714
rect 676048 760578 676076 760679
rect 676128 760650 676180 760656
rect 676036 760572 676088 760578
rect 676036 760514 676088 760520
rect 676036 760368 676088 760374
rect 676034 760336 676036 760345
rect 676088 760336 676090 760345
rect 676034 760271 676090 760280
rect 676218 759656 676274 759665
rect 676218 759591 676274 759600
rect 676036 759552 676088 759558
rect 676034 759520 676036 759529
rect 676088 759520 676090 759529
rect 676034 759455 676090 759464
rect 676232 759150 676260 759591
rect 676220 759144 676272 759150
rect 676034 759112 676090 759121
rect 676220 759086 676272 759092
rect 676034 759047 676036 759056
rect 676088 759047 676090 759056
rect 676036 759018 676088 759024
rect 676034 758296 676090 758305
rect 676034 758231 676036 758240
rect 676088 758231 676090 758240
rect 676036 758202 676088 758208
rect 679636 756809 679664 772647
rect 703694 762076 703722 762212
rect 704154 762076 704182 762212
rect 704614 762076 704642 762212
rect 705074 762076 705102 762212
rect 705534 762076 705562 762212
rect 705994 762076 706022 762212
rect 706454 762076 706482 762212
rect 706914 762076 706942 762212
rect 707374 762076 707402 762212
rect 707834 762076 707862 762212
rect 708294 762076 708322 762212
rect 708754 762076 708782 762212
rect 709214 762076 709242 762212
rect 679622 756800 679678 756809
rect 679622 756735 679678 756744
rect 675758 756256 675814 756265
rect 675758 756191 675814 756200
rect 676220 755608 676272 755614
rect 676218 755576 676220 755585
rect 676272 755576 676274 755585
rect 676218 755511 676274 755520
rect 676034 755032 676090 755041
rect 676034 754967 676036 754976
rect 676088 754967 676090 754976
rect 676036 754938 676088 754944
rect 676220 754384 676272 754390
rect 676218 754352 676220 754361
rect 676272 754352 676274 754361
rect 676218 754287 676274 754296
rect 676034 753808 676090 753817
rect 676034 753743 676090 753752
rect 676048 753642 676076 753743
rect 676036 753636 676088 753642
rect 676036 753578 676088 753584
rect 676220 753160 676272 753166
rect 676218 753128 676220 753137
rect 676272 753128 676274 753137
rect 676218 753063 676274 753072
rect 676220 752752 676272 752758
rect 676218 752720 676220 752729
rect 676272 752720 676274 752729
rect 676218 752655 676274 752664
rect 676218 752312 676274 752321
rect 676218 752247 676220 752256
rect 676272 752247 676274 752256
rect 676220 752218 676272 752224
rect 676218 751496 676274 751505
rect 676218 751431 676274 751440
rect 676232 750922 676260 751431
rect 683118 751088 683174 751097
rect 683118 751023 683174 751032
rect 676220 750916 676272 750922
rect 676220 750858 676272 750864
rect 683132 750281 683160 751023
rect 683118 750272 683174 750281
rect 683118 750207 683174 750216
rect 683132 749426 683160 750207
rect 683120 749420 683172 749426
rect 683120 749362 683172 749368
rect 675404 743238 675432 743308
rect 675392 743232 675444 743238
rect 675392 743174 675444 743180
rect 675404 742558 675432 742696
rect 675392 742552 675444 742558
rect 675392 742494 675444 742500
rect 675496 741713 675524 742016
rect 675482 741704 675538 741713
rect 675482 741639 675538 741648
rect 675772 739945 675800 740180
rect 675758 739936 675814 739945
rect 675758 739871 675814 739880
rect 675404 739158 675432 739636
rect 675666 739256 675722 739265
rect 675666 739191 675722 739200
rect 675392 739152 675444 739158
rect 675392 739094 675444 739100
rect 675680 739024 675708 739191
rect 675404 738274 675432 738344
rect 675392 738268 675444 738274
rect 675392 738210 675444 738216
rect 675404 735690 675432 735896
rect 675392 735684 675444 735690
rect 675392 735626 675444 735632
rect 675404 735010 675432 735319
rect 675392 735004 675444 735010
rect 675392 734946 675444 734952
rect 675772 734369 675800 734672
rect 675758 734360 675814 734369
rect 675758 734295 675814 734304
rect 675404 733650 675432 734031
rect 675392 733644 675444 733650
rect 675392 733586 675444 733592
rect 675758 733000 675814 733009
rect 675758 732935 675814 732944
rect 675772 732836 675800 732935
rect 675392 732080 675444 732086
rect 675392 732022 675444 732028
rect 675404 731612 675432 732022
rect 675404 730522 675432 731000
rect 675392 730516 675444 730522
rect 675392 730458 675444 730464
rect 675496 728686 675524 729164
rect 675484 728680 675536 728686
rect 675484 728622 675536 728628
rect 678242 727288 678298 727297
rect 678242 727223 678298 727232
rect 676034 716544 676090 716553
rect 676034 716479 676090 716488
rect 676048 716310 676076 716479
rect 676036 716304 676088 716310
rect 676036 716246 676088 716252
rect 676036 716168 676088 716174
rect 676034 716136 676036 716145
rect 676088 716136 676090 716145
rect 676034 716071 676090 716080
rect 676034 715728 676090 715737
rect 676034 715663 676090 715672
rect 675944 715352 675996 715358
rect 675942 715320 675944 715329
rect 675996 715320 675998 715329
rect 675942 715255 675998 715264
rect 676048 715018 676076 715663
rect 676036 715012 676088 715018
rect 676036 714954 676088 714960
rect 676034 714912 676090 714921
rect 676034 714847 676036 714856
rect 676088 714847 676090 714856
rect 676036 714818 676088 714824
rect 676036 714536 676088 714542
rect 676034 714504 676036 714513
rect 676088 714504 676090 714513
rect 676034 714439 676090 714448
rect 676034 714096 676090 714105
rect 676034 714031 676036 714040
rect 676088 714031 676090 714040
rect 676036 714002 676088 714008
rect 676036 713720 676088 713726
rect 676034 713688 676036 713697
rect 676088 713688 676090 713697
rect 676034 713623 676090 713632
rect 677322 713488 677378 713497
rect 677322 713423 677378 713432
rect 676034 713280 676090 713289
rect 676034 713215 676036 713224
rect 676088 713215 676090 713224
rect 676036 713186 676088 713192
rect 674746 712872 674802 712881
rect 674746 712807 674802 712816
rect 676034 712464 676090 712473
rect 676034 712399 676036 712408
rect 676088 712399 676090 712408
rect 676036 712370 676088 712376
rect 676036 712088 676088 712094
rect 676034 712056 676036 712065
rect 676088 712056 676090 712065
rect 676034 711991 676090 712000
rect 676036 711272 676088 711278
rect 676034 711240 676036 711249
rect 676088 711240 676090 711249
rect 676034 711175 676090 711184
rect 675942 711104 675998 711113
rect 675942 711039 675998 711048
rect 675956 704449 675984 711039
rect 676036 710456 676088 710462
rect 676034 710424 676036 710433
rect 676088 710424 676090 710433
rect 676034 710359 676090 710368
rect 676036 710048 676088 710054
rect 676034 710016 676036 710025
rect 676088 710016 676090 710025
rect 676034 709951 676090 709960
rect 676036 709640 676088 709646
rect 676034 709608 676036 709617
rect 676088 709608 676090 709617
rect 676034 709543 676090 709552
rect 676036 709232 676088 709238
rect 676034 709200 676036 709209
rect 676088 709200 676090 709209
rect 676034 709135 676090 709144
rect 676036 708416 676088 708422
rect 676034 708384 676036 708393
rect 676088 708384 676090 708393
rect 676034 708319 676090 708328
rect 677336 708286 677364 713423
rect 678256 711657 678284 727223
rect 703694 717196 703722 717264
rect 704154 717196 704182 717264
rect 704614 717196 704642 717264
rect 705074 717196 705102 717264
rect 705534 717196 705562 717264
rect 705994 717196 706022 717264
rect 706454 717196 706482 717264
rect 706914 717196 706942 717264
rect 707374 717196 707402 717264
rect 707834 717196 707862 717264
rect 708294 717196 708322 717264
rect 708754 717196 708782 717264
rect 709214 717196 709242 717264
rect 678242 711648 678298 711657
rect 678242 711583 678298 711592
rect 676036 708280 676088 708286
rect 676036 708222 676088 708228
rect 677324 708280 677376 708286
rect 677324 708222 677376 708228
rect 676048 707985 676076 708222
rect 676034 707976 676090 707985
rect 676034 707911 676090 707920
rect 676036 707600 676088 707606
rect 676034 707568 676036 707577
rect 676088 707568 676090 707577
rect 676034 707503 676090 707512
rect 676036 707192 676088 707198
rect 676034 707160 676036 707169
rect 676088 707160 676090 707169
rect 676034 707095 676090 707104
rect 676036 706784 676088 706790
rect 676034 706752 676036 706761
rect 676088 706752 676090 706761
rect 676034 706687 676090 706696
rect 676034 706344 676090 706353
rect 676034 706279 676090 706288
rect 676048 705129 676076 706279
rect 676034 705120 676090 705129
rect 676034 705055 676090 705064
rect 675942 704440 675998 704449
rect 675942 704375 675998 704384
rect 676048 703866 676076 705055
rect 676036 703860 676088 703866
rect 676036 703802 676088 703808
rect 675404 698222 675432 698323
rect 675392 698216 675444 698222
rect 675392 698158 675444 698164
rect 675404 697377 675432 697680
rect 675390 697368 675446 697377
rect 675390 697303 675446 697312
rect 675680 696969 675708 697035
rect 675666 696960 675722 696969
rect 675666 696895 675722 696904
rect 675772 695065 675800 695195
rect 675758 695056 675814 695065
rect 675758 694991 675814 695000
rect 675496 694210 675524 694620
rect 675758 694240 675814 694249
rect 674656 694204 674708 694210
rect 674656 694146 674708 694152
rect 675484 694204 675536 694210
rect 675758 694175 675814 694184
rect 675484 694146 675536 694152
rect 674564 661632 674616 661638
rect 674564 661574 674616 661580
rect 674564 649868 674616 649874
rect 674564 649810 674616 649816
rect 674472 643748 674524 643754
rect 674472 643690 674524 643696
rect 674484 641918 674512 643690
rect 674472 641912 674524 641918
rect 674472 641854 674524 641860
rect 674380 617840 674432 617846
rect 674380 617782 674432 617788
rect 674472 604784 674524 604790
rect 674472 604726 674524 604732
rect 674380 599820 674432 599826
rect 674380 599762 674432 599768
rect 674288 571736 674340 571742
rect 674288 571678 674340 571684
rect 674288 555280 674340 555286
rect 674288 555222 674340 555228
rect 674196 526380 674248 526386
rect 674196 526322 674248 526328
rect 673276 525972 673328 525978
rect 673276 525914 673328 525920
rect 674300 486062 674328 555222
rect 674392 526794 674420 599762
rect 674484 530466 674512 604726
rect 674576 575414 674604 649810
rect 674668 619206 674696 694146
rect 675772 694008 675800 694175
rect 675496 692986 675524 693328
rect 675484 692980 675536 692986
rect 675484 692922 675536 692928
rect 675404 690470 675432 690880
rect 675392 690464 675444 690470
rect 675392 690406 675444 690412
rect 675404 690062 675432 690336
rect 675392 690056 675444 690062
rect 675392 689998 675444 690004
rect 675496 689382 675524 689656
rect 675484 689376 675536 689382
rect 675484 689318 675536 689324
rect 674748 689308 674800 689314
rect 674748 689250 674800 689256
rect 674760 687070 674788 689250
rect 675404 688702 675432 689044
rect 675392 688696 675444 688702
rect 675392 688638 675444 688644
rect 675404 687342 675432 687820
rect 675392 687336 675444 687342
rect 675392 687278 675444 687284
rect 674748 687064 674800 687070
rect 674748 687006 674800 687012
rect 675484 687064 675536 687070
rect 675484 687006 675536 687012
rect 675496 686664 675524 687006
rect 675392 686112 675444 686118
rect 675392 686054 675444 686060
rect 675404 685984 675432 686054
rect 675392 684276 675444 684282
rect 675392 684218 675444 684224
rect 675404 684148 675432 684218
rect 678242 679008 678298 679017
rect 678242 678943 678298 678952
rect 676218 671120 676274 671129
rect 676218 671055 676274 671064
rect 676034 670984 676090 670993
rect 676232 670954 676260 671055
rect 676034 670919 676090 670928
rect 676220 670948 676272 670954
rect 676048 670818 676076 670919
rect 676220 670890 676272 670896
rect 676036 670812 676088 670818
rect 676036 670754 676088 670760
rect 676310 670304 676366 670313
rect 676310 670239 676366 670248
rect 676126 669896 676182 669905
rect 676126 669831 676182 669840
rect 674746 669760 674802 669769
rect 674746 669695 674802 669704
rect 674760 625161 674788 669695
rect 676140 669594 676168 669831
rect 676220 669724 676272 669730
rect 676220 669666 676272 669672
rect 676128 669588 676180 669594
rect 676128 669530 676180 669536
rect 676232 669497 676260 669666
rect 676218 669488 676274 669497
rect 676324 669458 676352 670239
rect 676218 669423 676274 669432
rect 676312 669452 676364 669458
rect 676312 669394 676364 669400
rect 676034 668944 676090 668953
rect 676034 668879 676036 668888
rect 676088 668879 676090 668888
rect 676036 668850 676088 668856
rect 676220 668704 676272 668710
rect 676218 668672 676220 668681
rect 676272 668672 676274 668681
rect 676218 668607 676274 668616
rect 676034 668128 676090 668137
rect 676034 668063 676090 668072
rect 676048 667962 676076 668063
rect 676036 667956 676088 667962
rect 676036 667898 676088 667904
rect 676220 667888 676272 667894
rect 676218 667856 676220 667865
rect 676272 667856 676274 667865
rect 676218 667791 676274 667800
rect 678256 667049 678284 678943
rect 703694 671908 703722 672044
rect 704154 671908 704182 672044
rect 704614 671908 704642 672044
rect 705074 671908 705102 672044
rect 705534 671908 705562 672044
rect 705994 671908 706022 672044
rect 706454 671908 706482 672044
rect 706914 671908 706942 672044
rect 707374 671908 707402 672044
rect 707834 671908 707862 672044
rect 708294 671908 708322 672044
rect 708754 671908 708782 672044
rect 709214 671908 709242 672044
rect 676218 667040 676274 667049
rect 676218 666975 676274 666984
rect 678242 667040 678298 667049
rect 678242 666975 678298 666984
rect 676232 666602 676260 666975
rect 676220 666596 676272 666602
rect 676220 666538 676272 666544
rect 676036 666528 676088 666534
rect 676034 666496 676036 666505
rect 676088 666496 676090 666505
rect 676034 666431 676090 666440
rect 676218 665816 676274 665825
rect 676218 665751 676274 665760
rect 676232 665378 676260 665751
rect 676220 665372 676272 665378
rect 676220 665314 676272 665320
rect 676036 665304 676088 665310
rect 676034 665272 676036 665281
rect 676088 665272 676090 665281
rect 676034 665207 676090 665216
rect 676220 665032 676272 665038
rect 676218 665000 676220 665009
rect 676272 665000 676274 665009
rect 676218 664935 676274 664944
rect 676218 664184 676274 664193
rect 676218 664119 676274 664128
rect 676232 664018 676260 664119
rect 676220 664012 676272 664018
rect 676220 663954 676272 663960
rect 676220 663808 676272 663814
rect 676218 663776 676220 663785
rect 676272 663776 676274 663785
rect 676218 663711 676274 663720
rect 676034 662416 676090 662425
rect 676034 662351 676036 662360
rect 676088 662351 676090 662360
rect 676036 662322 676088 662328
rect 676218 661736 676274 661745
rect 676218 661671 676274 661680
rect 676036 661632 676088 661638
rect 676034 661600 676036 661609
rect 676088 661600 676090 661609
rect 676034 661535 676090 661544
rect 676232 661162 676260 661671
rect 676220 661156 676272 661162
rect 676220 661098 676272 661104
rect 683118 660920 683174 660929
rect 683118 660855 683174 660864
rect 683132 660113 683160 660855
rect 683118 660104 683174 660113
rect 683118 660039 683174 660048
rect 675404 652798 675432 653140
rect 675392 652792 675444 652798
rect 675392 652734 675444 652740
rect 675496 652225 675524 652460
rect 675482 652216 675538 652225
rect 675482 652151 675538 652160
rect 675772 651545 675800 651848
rect 675758 651536 675814 651545
rect 675758 651471 675814 651480
rect 675404 649874 675432 650012
rect 675392 649868 675444 649874
rect 675392 649810 675444 649816
rect 675404 649233 675432 649468
rect 675390 649224 675446 649233
rect 675390 649159 675446 649168
rect 675772 648689 675800 648788
rect 675758 648680 675814 648689
rect 675758 648615 675814 648624
rect 675496 647766 675524 648176
rect 675484 647760 675536 647766
rect 675484 647702 675536 647708
rect 675404 645590 675432 645660
rect 675392 645584 675444 645590
rect 675392 645526 675444 645532
rect 675404 644842 675432 645116
rect 675392 644836 675444 644842
rect 675392 644778 675444 644784
rect 675758 644736 675814 644745
rect 675758 644671 675814 644680
rect 675772 644475 675800 644671
rect 675404 643414 675432 643824
rect 675392 643408 675444 643414
rect 675392 643350 675444 643356
rect 675666 643104 675722 643113
rect 675666 643039 675722 643048
rect 675680 642635 675708 643039
rect 675392 641912 675444 641918
rect 675392 641854 675444 641860
rect 675404 641444 675432 641854
rect 675496 640393 675524 640795
rect 675482 640384 675538 640393
rect 675482 640319 675538 640328
rect 675392 639124 675444 639130
rect 675392 639066 675444 639072
rect 675404 638928 675432 639066
rect 675666 638208 675722 638217
rect 675666 638143 675722 638152
rect 674746 625152 674802 625161
rect 674746 625087 674802 625096
rect 674656 619200 674708 619206
rect 674656 619142 674708 619148
rect 675680 610706 675708 638143
rect 678242 633448 678298 633457
rect 678242 633383 678298 633392
rect 676126 626104 676182 626113
rect 676126 626039 676182 626048
rect 676140 625530 676168 626039
rect 676218 625696 676274 625705
rect 676218 625631 676274 625640
rect 676128 625524 676180 625530
rect 676128 625466 676180 625472
rect 676232 625394 676260 625631
rect 676220 625388 676272 625394
rect 676220 625330 676272 625336
rect 676218 625288 676274 625297
rect 676218 625223 676274 625232
rect 676232 625190 676260 625223
rect 676220 625184 676272 625190
rect 676220 625126 676272 625132
rect 676218 624472 676274 624481
rect 676218 624407 676274 624416
rect 676036 624368 676088 624374
rect 676034 624336 676036 624345
rect 676088 624336 676090 624345
rect 676034 624271 676090 624280
rect 676034 623928 676090 623937
rect 676034 623863 676036 623872
rect 676088 623863 676090 623872
rect 676036 623834 676088 623840
rect 676232 623830 676260 624407
rect 676220 623824 676272 623830
rect 676220 623766 676272 623772
rect 676126 623248 676182 623257
rect 676126 623183 676182 623192
rect 676036 622736 676088 622742
rect 676034 622704 676036 622713
rect 676088 622704 676090 622713
rect 676034 622639 676090 622648
rect 676140 622606 676168 623183
rect 676218 622840 676274 622849
rect 676218 622775 676274 622784
rect 676128 622600 676180 622606
rect 676128 622542 676180 622548
rect 676232 622470 676260 622775
rect 676220 622464 676272 622470
rect 676220 622406 676272 622412
rect 676034 622296 676090 622305
rect 676034 622231 676036 622240
rect 676088 622231 676090 622240
rect 676036 622202 676088 622208
rect 678256 622033 678284 633383
rect 703694 626892 703722 627028
rect 704154 626892 704182 627028
rect 704614 626892 704642 627028
rect 705074 626892 705102 627028
rect 705534 626892 705562 627028
rect 705994 626892 706022 627028
rect 706454 626892 706482 627028
rect 706914 626892 706942 627028
rect 707374 626892 707402 627028
rect 707834 626892 707862 627028
rect 708294 626892 708322 627028
rect 708754 626892 708782 627028
rect 709214 626892 709242 627028
rect 678242 622024 678298 622033
rect 678242 621959 678298 621968
rect 676034 621480 676090 621489
rect 676034 621415 676090 621424
rect 676048 621178 676076 621415
rect 676220 621308 676272 621314
rect 676220 621250 676272 621256
rect 676232 621217 676260 621250
rect 676218 621208 676274 621217
rect 676036 621172 676088 621178
rect 676218 621143 676274 621152
rect 676036 621114 676088 621120
rect 676218 619984 676274 619993
rect 676218 619919 676220 619928
rect 676272 619919 676274 619928
rect 676220 619890 676272 619896
rect 676034 619848 676090 619857
rect 676034 619783 676036 619792
rect 676088 619783 676090 619792
rect 676036 619754 676088 619760
rect 676220 619200 676272 619206
rect 676218 619168 676220 619177
rect 676272 619168 676274 619177
rect 676218 619103 676274 619112
rect 676126 617944 676182 617953
rect 676126 617879 676182 617888
rect 676036 617840 676088 617846
rect 676034 617808 676036 617817
rect 676088 617808 676090 617817
rect 676034 617743 676090 617752
rect 676140 617098 676168 617879
rect 676218 617128 676274 617137
rect 676128 617092 676180 617098
rect 676218 617063 676274 617072
rect 676128 617034 676180 617040
rect 676036 617024 676088 617030
rect 676034 616992 676036 617001
rect 676088 616992 676090 617001
rect 676034 616927 676090 616936
rect 676232 616894 676260 617063
rect 676220 616888 676272 616894
rect 676220 616830 676272 616836
rect 676218 616312 676274 616321
rect 676218 616247 676274 616256
rect 676232 615534 676260 616247
rect 683118 615904 683174 615913
rect 683118 615839 683174 615848
rect 676220 615528 676272 615534
rect 676220 615470 676272 615476
rect 683132 615097 683160 615839
rect 683118 615088 683174 615097
rect 683118 615023 683174 615032
rect 683132 614174 683160 615023
rect 683120 614168 683172 614174
rect 683120 614110 683172 614116
rect 675208 610700 675260 610706
rect 675208 610642 675260 610648
rect 675668 610700 675720 610706
rect 675668 610642 675720 610648
rect 674656 604376 674708 604382
rect 674656 604318 674708 604324
rect 674564 575408 674616 575414
rect 674564 575350 674616 575356
rect 674564 554192 674616 554198
rect 674564 554134 674616 554140
rect 674472 530460 674524 530466
rect 674472 530402 674524 530408
rect 674380 526788 674432 526794
rect 674380 526730 674432 526736
rect 674288 486056 674340 486062
rect 674288 485998 674340 486004
rect 674576 483614 674604 554134
rect 674668 528902 674696 604318
rect 675220 600953 675248 610642
rect 675496 607889 675524 608124
rect 675482 607880 675538 607889
rect 675482 607815 675538 607824
rect 675392 607640 675444 607646
rect 675392 607582 675444 607588
rect 675404 607479 675432 607582
rect 675404 606529 675432 606832
rect 675390 606520 675446 606529
rect 675390 606455 675446 606464
rect 675404 604790 675432 604996
rect 675392 604784 675444 604790
rect 675392 604726 675444 604732
rect 675404 604382 675432 604452
rect 675392 604376 675444 604382
rect 675392 604318 675444 604324
rect 675496 603498 675524 603772
rect 675484 603492 675536 603498
rect 675484 603434 675536 603440
rect 675404 603090 675432 603160
rect 675392 603084 675444 603090
rect 675392 603026 675444 603032
rect 675206 600944 675262 600953
rect 675206 600879 675262 600888
rect 675588 600273 675616 600644
rect 675574 600264 675630 600273
rect 675574 600199 675630 600208
rect 675496 599826 675524 600100
rect 675484 599820 675536 599826
rect 675484 599762 675536 599768
rect 674748 599208 674800 599214
rect 674748 599150 674800 599156
rect 674760 596902 674788 599150
rect 675772 599049 675800 599488
rect 675758 599040 675814 599049
rect 675758 598975 675814 598984
rect 675496 598466 675524 598808
rect 675484 598460 675536 598466
rect 675484 598402 675536 598408
rect 675758 597816 675814 597825
rect 675758 597751 675814 597760
rect 675772 597652 675800 597751
rect 674748 596896 674800 596902
rect 674748 596838 674800 596844
rect 675392 596896 675444 596902
rect 675392 596838 675444 596844
rect 675404 596428 675432 596838
rect 675404 595338 675432 595816
rect 675392 595332 675444 595338
rect 675392 595274 675444 595280
rect 675496 593434 675524 593980
rect 675484 593428 675536 593434
rect 675484 593370 675536 593376
rect 675482 593192 675538 593201
rect 675482 593127 675538 593136
rect 675666 593192 675722 593201
rect 675666 593127 675722 593136
rect 675496 568585 675524 593127
rect 675680 576201 675708 593127
rect 678242 589248 678298 589257
rect 678242 589183 678298 589192
rect 676034 581088 676090 581097
rect 676034 581023 676036 581032
rect 676088 581023 676090 581032
rect 676036 580994 676088 581000
rect 676126 580544 676182 580553
rect 676126 580479 676182 580488
rect 676034 580272 676090 580281
rect 676034 580207 676090 580216
rect 676048 579834 676076 580207
rect 676140 579970 676168 580479
rect 676218 580136 676274 580145
rect 676218 580071 676220 580080
rect 676272 580071 676274 580080
rect 676220 580042 676272 580048
rect 676128 579964 676180 579970
rect 676128 579906 676180 579912
rect 676036 579828 676088 579834
rect 676036 579770 676088 579776
rect 676218 579320 676274 579329
rect 676218 579255 676220 579264
rect 676272 579255 676274 579264
rect 676220 579226 676272 579232
rect 676218 578912 676274 578921
rect 676218 578847 676274 578856
rect 676034 578640 676090 578649
rect 676034 578575 676036 578584
rect 676088 578575 676090 578584
rect 676036 578546 676088 578552
rect 676232 578270 676260 578847
rect 676220 578264 676272 578270
rect 676220 578206 676272 578212
rect 676218 578096 676274 578105
rect 676218 578031 676274 578040
rect 676126 577688 676182 577697
rect 676126 577623 676182 577632
rect 676036 577448 676088 577454
rect 676034 577416 676036 577425
rect 676088 577416 676090 577425
rect 676034 577351 676090 577360
rect 676034 577008 676090 577017
rect 676034 576943 676036 576952
rect 676088 576943 676090 576952
rect 676036 576914 676088 576920
rect 676140 576910 676168 577623
rect 676232 577046 676260 578031
rect 676220 577040 676272 577046
rect 676220 576982 676272 576988
rect 676128 576904 676180 576910
rect 678256 576881 678284 589183
rect 703694 581740 703722 581876
rect 704154 581740 704182 581876
rect 704614 581740 704642 581876
rect 705074 581740 705102 581876
rect 705534 581740 705562 581876
rect 705994 581740 706022 581876
rect 706454 581740 706482 581876
rect 706914 581740 706942 581876
rect 707374 581740 707402 581876
rect 707834 581740 707862 581876
rect 708294 581740 708322 581876
rect 708754 581740 708782 581876
rect 709214 581740 709242 581876
rect 676128 576846 676180 576852
rect 678242 576872 678298 576881
rect 678242 576807 678298 576816
rect 675666 576192 675722 576201
rect 675666 576127 675722 576136
rect 676218 575648 676274 575657
rect 676218 575583 676220 575592
rect 676272 575583 676274 575592
rect 676220 575554 676272 575560
rect 676036 575408 676088 575414
rect 676034 575376 676036 575385
rect 676088 575376 676090 575385
rect 676034 575311 676090 575320
rect 676218 574832 676274 574841
rect 676218 574767 676274 574776
rect 676036 574592 676088 574598
rect 676034 574560 676036 574569
rect 676088 574560 676090 574569
rect 676034 574495 676090 574504
rect 676232 574258 676260 574767
rect 676220 574252 676272 574258
rect 676220 574194 676272 574200
rect 676218 571976 676274 571985
rect 676218 571911 676274 571920
rect 676036 571736 676088 571742
rect 676034 571704 676036 571713
rect 676088 571704 676090 571713
rect 676034 571639 676090 571648
rect 676232 571538 676260 571911
rect 676220 571532 676272 571538
rect 676220 571474 676272 571480
rect 676218 571160 676274 571169
rect 676218 571095 676274 571104
rect 676232 569974 676260 571095
rect 683118 570752 683174 570761
rect 683118 570687 683174 570696
rect 676220 569968 676272 569974
rect 683132 569945 683160 570687
rect 676220 569910 676272 569916
rect 683118 569936 683174 569945
rect 683118 569871 683174 569880
rect 683132 568614 683160 569871
rect 683120 568608 683172 568614
rect 675482 568576 675538 568585
rect 683120 568550 683172 568556
rect 675482 568511 675538 568520
rect 675772 562737 675800 562904
rect 675758 562728 675814 562737
rect 675758 562663 675814 562672
rect 675404 561950 675432 562292
rect 675392 561944 675444 561950
rect 675392 561886 675444 561892
rect 675772 561241 675800 561612
rect 675758 561232 675814 561241
rect 675758 561167 675814 561176
rect 675208 560244 675260 560250
rect 675208 560186 675260 560192
rect 675220 559706 675248 560186
rect 675208 559700 675260 559706
rect 675208 559642 675260 559648
rect 675392 559700 675444 559706
rect 675392 559642 675444 559648
rect 675404 559232 675432 559642
rect 675496 559609 675524 559776
rect 675482 559600 675538 559609
rect 675482 559535 675538 559544
rect 675772 558385 675800 558620
rect 675758 558376 675814 558385
rect 675758 558311 675814 558320
rect 675496 557598 675524 557940
rect 675484 557592 675536 557598
rect 675484 557534 675536 557540
rect 675404 555286 675432 555492
rect 675392 555280 675444 555286
rect 675392 555222 675444 555228
rect 675312 554905 675418 554933
rect 675312 554810 675340 554905
rect 675300 554804 675352 554810
rect 675300 554746 675352 554752
rect 675312 554254 675418 554282
rect 675312 554198 675340 554254
rect 675300 554192 675352 554198
rect 675300 554134 675352 554140
rect 675300 554056 675352 554062
rect 675300 553998 675352 554004
rect 675312 551253 675340 553998
rect 675404 553518 675432 553656
rect 675392 553512 675444 553518
rect 675392 553454 675444 553460
rect 675772 551993 675800 552432
rect 675758 551984 675814 551993
rect 675758 551919 675814 551928
rect 675312 551225 675418 551253
rect 675312 550582 675418 550610
rect 675312 549234 675340 550582
rect 674932 549228 674984 549234
rect 674932 549170 674984 549176
rect 675300 549228 675352 549234
rect 675300 549170 675352 549176
rect 674748 548344 674800 548350
rect 674748 548286 674800 548292
rect 674656 528896 674708 528902
rect 674656 528838 674708 528844
rect 674760 485625 674788 548286
rect 674944 488374 674972 549170
rect 675312 548746 675418 548774
rect 675312 548350 675340 548746
rect 675300 548344 675352 548350
rect 675300 548286 675352 548292
rect 681002 546544 681058 546553
rect 681002 546479 681058 546488
rect 678242 543824 678298 543833
rect 678242 543759 678298 543768
rect 676218 535936 676274 535945
rect 676218 535871 676274 535880
rect 676232 535770 676260 535871
rect 676220 535764 676272 535770
rect 676034 535732 676090 535741
rect 676220 535706 676272 535712
rect 676034 535667 676090 535676
rect 676048 535634 676076 535667
rect 676036 535628 676088 535634
rect 676036 535570 676088 535576
rect 676218 535120 676274 535129
rect 676218 535055 676274 535064
rect 676036 534948 676088 534954
rect 676034 534916 676036 534925
rect 676088 534916 676090 534925
rect 676034 534851 676090 534860
rect 676232 534274 676260 535055
rect 676220 534268 676272 534274
rect 676220 534210 676272 534216
rect 676036 534132 676088 534138
rect 676034 534100 676036 534109
rect 676088 534100 676090 534109
rect 676034 534035 676090 534044
rect 676218 533080 676274 533089
rect 676218 533015 676274 533024
rect 676232 532914 676260 533015
rect 676220 532908 676272 532914
rect 676220 532850 676272 532856
rect 677322 532672 677378 532681
rect 677322 532607 677378 532616
rect 676218 532264 676274 532273
rect 676218 532199 676274 532208
rect 676232 531350 676260 532199
rect 676220 531344 676272 531350
rect 676220 531286 676272 531292
rect 676218 531040 676274 531049
rect 676218 530975 676274 530984
rect 676036 530460 676088 530466
rect 676034 530428 676036 530437
rect 676088 530428 676090 530437
rect 676034 530363 676090 530372
rect 676232 530058 676260 530975
rect 676220 530052 676272 530058
rect 676220 529994 676272 530000
rect 676126 529408 676182 529417
rect 676126 529343 676182 529352
rect 676036 528896 676088 528902
rect 676036 528838 676088 528844
rect 676048 528805 676076 528838
rect 676034 528796 676090 528805
rect 676034 528731 676090 528740
rect 676140 528698 676168 529343
rect 676218 529000 676274 529009
rect 676218 528935 676274 528944
rect 676232 528834 676260 528935
rect 676220 528828 676272 528834
rect 676220 528770 676272 528776
rect 676128 528692 676180 528698
rect 676128 528634 676180 528640
rect 676036 528420 676088 528426
rect 676034 528388 676036 528397
rect 676088 528388 676090 528397
rect 676034 528323 676090 528332
rect 676218 526960 676274 526969
rect 676218 526895 676274 526904
rect 676036 526788 676088 526794
rect 676034 526756 676036 526765
rect 676088 526756 676090 526765
rect 676034 526691 676090 526700
rect 676036 526380 676088 526386
rect 676034 526348 676036 526357
rect 676088 526348 676090 526357
rect 676034 526283 676090 526292
rect 676232 525978 676260 526895
rect 676220 525972 676272 525978
rect 676220 525914 676272 525920
rect 676128 521008 676180 521014
rect 676128 520950 676180 520956
rect 676036 520940 676088 520946
rect 676036 520882 676088 520888
rect 676048 499574 676076 520882
rect 675864 499546 676076 499574
rect 675864 490113 675892 499546
rect 675942 492144 675998 492153
rect 675942 492079 675998 492088
rect 675956 491706 675984 492079
rect 676034 491736 676090 491745
rect 675944 491700 675996 491706
rect 676034 491671 676090 491680
rect 675944 491642 675996 491648
rect 676048 491570 676076 491671
rect 676036 491564 676088 491570
rect 676036 491506 676088 491512
rect 676036 491428 676088 491434
rect 676036 491370 676088 491376
rect 676048 491337 676076 491370
rect 676034 491328 676090 491337
rect 676034 491263 676090 491272
rect 676034 490920 676090 490929
rect 676140 490906 676168 520950
rect 676090 490878 676168 490906
rect 676034 490855 676090 490864
rect 676034 490512 676090 490521
rect 676034 490447 676090 490456
rect 675850 490104 675906 490113
rect 675850 490039 675906 490048
rect 675944 489320 675996 489326
rect 675942 489288 675944 489297
rect 675996 489288 675998 489297
rect 675942 489223 675998 489232
rect 675942 488880 675998 488889
rect 675942 488815 675998 488824
rect 675956 488646 675984 488815
rect 675944 488640 675996 488646
rect 675944 488582 675996 488588
rect 675944 488504 675996 488510
rect 675942 488472 675944 488481
rect 675996 488472 675998 488481
rect 675942 488407 675998 488416
rect 674932 488368 674984 488374
rect 674932 488310 674984 488316
rect 675944 488368 675996 488374
rect 675944 488310 675996 488316
rect 675850 488064 675906 488073
rect 675850 487999 675852 488008
rect 675904 487999 675906 488008
rect 675852 487970 675904 487976
rect 675956 487257 675984 488310
rect 675942 487248 675998 487257
rect 675942 487183 675998 487192
rect 675944 486056 675996 486062
rect 675942 486024 675944 486033
rect 675996 486024 675998 486033
rect 675942 485959 675998 485968
rect 674746 485616 674802 485625
rect 674746 485551 674802 485560
rect 675850 485208 675906 485217
rect 675850 485143 675906 485152
rect 675864 484430 675892 485143
rect 675942 484800 675998 484809
rect 675942 484735 675998 484744
rect 675956 484634 675984 484735
rect 675944 484628 675996 484634
rect 675944 484570 675996 484576
rect 675852 484424 675904 484430
rect 675852 484366 675904 484372
rect 674564 483608 674616 483614
rect 675944 483608 675996 483614
rect 674564 483550 674616 483556
rect 675942 483576 675944 483585
rect 675996 483576 675998 483585
rect 675942 483511 675998 483520
rect 675942 483168 675998 483177
rect 673184 483132 673236 483138
rect 675942 483103 675944 483112
rect 673184 483074 673236 483080
rect 675996 483103 675998 483112
rect 675944 483074 675996 483080
rect 675850 482760 675906 482769
rect 675850 482695 675906 482704
rect 675864 481914 675892 482695
rect 675942 482352 675998 482361
rect 675942 482287 675998 482296
rect 673000 481908 673052 481914
rect 673000 481850 673052 481856
rect 675852 481908 675904 481914
rect 675852 481850 675904 481856
rect 675956 481778 675984 482287
rect 672908 481772 672960 481778
rect 672908 481714 672960 481720
rect 675944 481772 675996 481778
rect 675944 481714 675996 481720
rect 674196 480276 674248 480282
rect 674196 480218 674248 480224
rect 673184 401668 673236 401674
rect 673184 401610 673236 401616
rect 673092 393372 673144 393378
rect 673092 393314 673144 393320
rect 673104 376786 673132 393314
rect 673092 376780 673144 376786
rect 673092 376722 673144 376728
rect 673196 357542 673224 401610
rect 673368 400308 673420 400314
rect 673368 400250 673420 400256
rect 673276 400240 673328 400246
rect 673276 400182 673328 400188
rect 673184 357536 673236 357542
rect 673184 357478 673236 357484
rect 673288 356726 673316 400182
rect 673276 356720 673328 356726
rect 673276 356662 673328 356668
rect 673380 355910 673408 400250
rect 673368 355904 673420 355910
rect 673368 355846 673420 355852
rect 672908 355428 672960 355434
rect 672908 355370 672960 355376
rect 672816 346452 672868 346458
rect 672816 346394 672868 346400
rect 672724 164008 672776 164014
rect 672724 163950 672776 163956
rect 672828 138242 672856 346394
rect 672920 310690 672948 355370
rect 673276 354612 673328 354618
rect 673276 354554 673328 354560
rect 673184 349308 673236 349314
rect 673184 349250 673236 349256
rect 673092 348900 673144 348906
rect 673092 348842 673144 348848
rect 673000 338156 673052 338162
rect 673000 338098 673052 338104
rect 672908 310684 672960 310690
rect 672908 310626 672960 310632
rect 672908 310548 672960 310554
rect 672908 310490 672960 310496
rect 672816 138236 672868 138242
rect 672816 138178 672868 138184
rect 672920 132938 672948 310490
rect 673012 178226 673040 338098
rect 673104 331634 673132 348842
rect 673196 332654 673224 349250
rect 673184 332648 673236 332654
rect 673184 332590 673236 332596
rect 673092 331628 673144 331634
rect 673092 331570 673144 331576
rect 673288 325694 673316 354554
rect 673368 350940 673420 350946
rect 673368 350882 673420 350888
rect 673380 336598 673408 350882
rect 674104 350600 674156 350606
rect 674104 350542 674156 350548
rect 673368 336592 673420 336598
rect 673368 336534 673420 336540
rect 673288 325666 673408 325694
rect 673276 309460 673328 309466
rect 673276 309402 673328 309408
rect 673184 303748 673236 303754
rect 673184 303690 673236 303696
rect 673092 303680 673144 303686
rect 673092 303622 673144 303628
rect 673104 287978 673132 303622
rect 673092 287972 673144 287978
rect 673092 287914 673144 287920
rect 673196 286618 673224 303690
rect 673184 286612 673236 286618
rect 673184 286554 673236 286560
rect 673288 265130 673316 309402
rect 673380 309398 673408 325666
rect 673368 309392 673420 309398
rect 673368 309334 673420 309340
rect 673368 309256 673420 309262
rect 673368 309198 673420 309204
rect 673380 265266 673408 309198
rect 673368 265260 673420 265266
rect 673368 265202 673420 265208
rect 673276 265124 673328 265130
rect 673276 265066 673328 265072
rect 673368 264988 673420 264994
rect 673368 264930 673420 264936
rect 673276 263628 673328 263634
rect 673276 263570 673328 263576
rect 673184 258120 673236 258126
rect 673184 258062 673236 258068
rect 673092 256760 673144 256766
rect 673092 256702 673144 256708
rect 673000 178220 673052 178226
rect 673000 178162 673052 178168
rect 673000 167884 673052 167890
rect 673000 167826 673052 167832
rect 672908 132932 672960 132938
rect 672908 132874 672960 132880
rect 671528 132796 671580 132802
rect 671528 132738 671580 132744
rect 672724 129940 672776 129946
rect 672724 129882 672776 129888
rect 671436 123888 671488 123894
rect 671436 123830 671488 123836
rect 671344 114368 671396 114374
rect 671344 114310 671396 114316
rect 670148 111308 670200 111314
rect 670148 111250 670200 111256
rect 670056 110356 670108 110362
rect 670056 110298 670108 110304
rect 672736 106146 672764 129882
rect 673012 117298 673040 167826
rect 673104 128178 673132 256702
rect 673196 241262 673224 258062
rect 673184 241256 673236 241262
rect 673184 241198 673236 241204
rect 673288 219910 673316 263570
rect 673380 220726 673408 264930
rect 673918 251696 673974 251705
rect 673918 251631 673974 251640
rect 673644 249892 673696 249898
rect 673644 249834 673696 249840
rect 673656 242894 673684 249834
rect 673734 249792 673790 249801
rect 673734 249727 673790 249736
rect 673748 244274 673776 249727
rect 673826 249656 673882 249665
rect 673826 249591 673882 249600
rect 673840 246129 673868 249591
rect 673932 246265 673960 251631
rect 674012 251524 674064 251530
rect 674012 251466 674064 251472
rect 674024 246566 674052 251466
rect 674012 246560 674064 246566
rect 674012 246502 674064 246508
rect 673918 246256 673974 246265
rect 673918 246191 673974 246200
rect 673826 246120 673882 246129
rect 673826 246055 673882 246064
rect 673748 244246 673960 244274
rect 673932 243642 673960 244246
rect 673920 243636 673972 243642
rect 673920 243578 673972 243584
rect 673644 242888 673696 242894
rect 673644 242830 673696 242836
rect 673368 220720 673420 220726
rect 673368 220662 673420 220668
rect 673276 219904 673328 219910
rect 673276 219846 673328 219852
rect 673184 214124 673236 214130
rect 673184 214066 673236 214072
rect 673196 197470 673224 214066
rect 673184 197464 673236 197470
rect 673184 197406 673236 197412
rect 674116 178090 674144 350542
rect 674104 178084 674156 178090
rect 674104 178026 674156 178032
rect 674012 176792 674064 176798
rect 674012 176734 674064 176740
rect 673368 174412 673420 174418
rect 673368 174354 673420 174360
rect 673184 169516 673236 169522
rect 673184 169458 673236 169464
rect 673196 155514 673224 169458
rect 673276 168700 673328 168706
rect 673276 168642 673328 168648
rect 673184 155508 673236 155514
rect 673184 155450 673236 155456
rect 673288 151434 673316 168642
rect 673276 151428 673328 151434
rect 673276 151370 673328 151376
rect 673380 128586 673408 174354
rect 674024 132326 674052 176734
rect 674104 168292 674156 168298
rect 674104 168234 674156 168240
rect 674012 132320 674064 132326
rect 674012 132262 674064 132268
rect 673368 128580 673420 128586
rect 673368 128522 673420 128528
rect 673092 128172 673144 128178
rect 673092 128114 673144 128120
rect 673368 123004 673420 123010
rect 673368 122946 673420 122952
rect 673000 117292 673052 117298
rect 673000 117234 673052 117240
rect 673380 106350 673408 122946
rect 674116 117842 674144 168234
rect 674208 148578 674236 480218
rect 676048 402665 676076 490447
rect 677336 489326 677364 532607
rect 678256 531865 678284 543759
rect 677506 531856 677562 531865
rect 677506 531791 677562 531800
rect 678242 531856 678298 531865
rect 678242 531791 678298 531800
rect 677414 489928 677470 489937
rect 677414 489863 677470 489872
rect 677324 489320 677376 489326
rect 677324 489262 677376 489268
rect 676128 488640 676180 488646
rect 676128 488582 676180 488588
rect 676034 402656 676090 402665
rect 676034 402591 676090 402600
rect 676140 401962 676168 488582
rect 677232 488028 677284 488034
rect 677232 487970 677284 487976
rect 676218 403744 676274 403753
rect 676218 403679 676274 403688
rect 676232 403442 676260 403679
rect 676220 403436 676272 403442
rect 676220 403378 676272 403384
rect 676218 403336 676274 403345
rect 676218 403271 676220 403280
rect 676272 403271 676274 403280
rect 676402 403336 676458 403345
rect 676402 403271 676458 403280
rect 676220 403242 676272 403248
rect 676416 403170 676444 403271
rect 676404 403164 676456 403170
rect 676404 403106 676456 403112
rect 676218 402112 676274 402121
rect 676218 402047 676274 402056
rect 676048 401934 676168 401962
rect 676048 401033 676076 401934
rect 676232 401674 676260 402047
rect 676220 401668 676272 401674
rect 676220 401610 676272 401616
rect 676126 401296 676182 401305
rect 676126 401231 676182 401240
rect 676034 401024 676090 401033
rect 676034 400959 676090 400968
rect 676140 400246 676168 401231
rect 677244 400489 677272 487970
rect 677428 470594 677456 489863
rect 677520 488510 677548 531791
rect 681016 531049 681044 546479
rect 703694 536724 703722 536860
rect 704154 536724 704182 536860
rect 704614 536724 704642 536860
rect 705074 536724 705102 536860
rect 705534 536724 705562 536860
rect 705994 536724 706022 536860
rect 706454 536724 706482 536860
rect 706914 536724 706942 536860
rect 707374 536724 707402 536860
rect 707834 536724 707862 536860
rect 708294 536724 708322 536860
rect 708754 536724 708782 536860
rect 709214 536724 709242 536860
rect 683302 534304 683358 534313
rect 683302 534239 683358 534248
rect 681002 531040 681058 531049
rect 681002 530975 681058 530984
rect 683118 525736 683174 525745
rect 683118 525671 683174 525680
rect 683132 524929 683160 525671
rect 683118 524920 683174 524929
rect 683118 524855 683174 524864
rect 683132 524482 683160 524855
rect 683120 524476 683172 524482
rect 683120 524418 683172 524424
rect 683316 521014 683344 534239
rect 683670 533488 683726 533497
rect 683670 533423 683726 533432
rect 683304 521008 683356 521014
rect 683304 520950 683356 520956
rect 683684 520946 683712 533423
rect 683672 520940 683724 520946
rect 683672 520882 683724 520888
rect 679622 503704 679678 503713
rect 679622 503639 679678 503648
rect 677508 488504 677560 488510
rect 677508 488446 677560 488452
rect 679636 486849 679664 503639
rect 679806 503568 679862 503577
rect 679806 503503 679862 503512
rect 679622 486840 679678 486849
rect 679622 486775 679678 486784
rect 679820 486441 679848 503503
rect 703694 492796 703722 492864
rect 704154 492796 704182 492864
rect 704614 492796 704642 492864
rect 705074 492796 705102 492864
rect 705534 492796 705562 492864
rect 705994 492796 706022 492864
rect 706454 492796 706482 492864
rect 706914 492796 706942 492864
rect 707374 492796 707402 492864
rect 707834 492796 707862 492864
rect 708294 492796 708322 492864
rect 708754 492796 708782 492864
rect 709214 492796 709242 492864
rect 679806 486432 679862 486441
rect 679806 486367 679862 486376
rect 678978 480720 679034 480729
rect 678978 480655 679034 480664
rect 678992 480282 679020 480655
rect 678980 480276 679032 480282
rect 678980 480218 679032 480224
rect 677336 470566 677456 470594
rect 677336 402121 677364 470566
rect 703694 404532 703722 404668
rect 704154 404532 704182 404668
rect 704614 404532 704642 404668
rect 705074 404532 705102 404668
rect 705534 404532 705562 404668
rect 705994 404532 706022 404668
rect 706454 404532 706482 404668
rect 706914 404532 706942 404668
rect 707374 404532 707402 404668
rect 707834 404532 707862 404668
rect 708294 404532 708322 404668
rect 708754 404532 708782 404668
rect 709214 404532 709242 404668
rect 677322 402112 677378 402121
rect 677322 402047 677378 402056
rect 676218 400480 676274 400489
rect 676218 400415 676274 400424
rect 677230 400480 677286 400489
rect 677230 400415 677286 400424
rect 676232 400314 676260 400415
rect 676220 400308 676272 400314
rect 676220 400250 676272 400256
rect 676128 400240 676180 400246
rect 676128 400182 676180 400188
rect 676218 399664 676274 399673
rect 674748 399628 674800 399634
rect 676218 399599 676220 399608
rect 674748 399570 674800 399576
rect 676272 399599 676274 399608
rect 676220 399570 676272 399576
rect 674656 394052 674708 394058
rect 674656 393994 674708 394000
rect 674668 376718 674696 393994
rect 674656 376712 674708 376718
rect 674656 376654 674708 376660
rect 674380 364404 674432 364410
rect 674380 364346 674432 364352
rect 674288 302252 674340 302258
rect 674288 302194 674340 302200
rect 674196 148572 674248 148578
rect 674196 148514 674248 148520
rect 674300 133006 674328 302194
rect 674392 222766 674420 364346
rect 674656 357060 674708 357066
rect 674656 357002 674708 357008
rect 674472 356244 674524 356250
rect 674472 356186 674524 356192
rect 674484 311710 674512 356186
rect 674564 350600 674616 350606
rect 674564 350542 674616 350548
rect 674576 330614 674604 350542
rect 674564 330608 674616 330614
rect 674564 330550 674616 330556
rect 674668 312526 674696 357002
rect 674760 355065 674788 399570
rect 676034 398576 676090 398585
rect 676034 398511 676090 398520
rect 676048 398274 676076 398511
rect 675024 398268 675076 398274
rect 675024 398210 675076 398216
rect 676036 398268 676088 398274
rect 676036 398210 676088 398216
rect 674932 397520 674984 397526
rect 674932 397462 674984 397468
rect 674944 383110 674972 397462
rect 675036 386170 675064 398210
rect 676034 398168 676090 398177
rect 676034 398103 676090 398112
rect 676048 397526 676076 398103
rect 676862 397624 676918 397633
rect 676862 397559 676918 397568
rect 676036 397520 676088 397526
rect 676036 397462 676088 397468
rect 676494 394768 676550 394777
rect 676494 394703 676550 394712
rect 676218 394360 676274 394369
rect 676218 394295 676274 394304
rect 676034 394088 676090 394097
rect 676034 394023 676036 394032
rect 676088 394023 676090 394032
rect 676036 393994 676088 394000
rect 676232 393378 676260 394295
rect 676220 393372 676272 393378
rect 676220 393314 676272 393320
rect 675208 387796 675260 387802
rect 675208 387738 675260 387744
rect 675116 387728 675168 387734
rect 675116 387670 675168 387676
rect 675024 386164 675076 386170
rect 675024 386106 675076 386112
rect 675024 386028 675076 386034
rect 675024 385970 675076 385976
rect 675036 383926 675064 385970
rect 675024 383920 675076 383926
rect 675024 383862 675076 383868
rect 674932 383104 674984 383110
rect 674932 383046 674984 383052
rect 675128 381138 675156 387670
rect 675220 385830 675248 387738
rect 676508 387734 676536 394703
rect 676876 388521 676904 397559
rect 676954 396808 677010 396817
rect 676954 396743 677010 396752
rect 676862 388512 676918 388521
rect 676862 388447 676918 388456
rect 676968 387802 676996 396743
rect 679622 396400 679678 396409
rect 679622 396335 679678 396344
rect 678242 395992 678298 396001
rect 678242 395927 678298 395936
rect 676956 387796 677008 387802
rect 676956 387738 677008 387744
rect 676496 387728 676548 387734
rect 676496 387670 676548 387676
rect 678256 387666 678284 395927
rect 679636 388249 679664 396335
rect 683118 393544 683174 393553
rect 683118 393479 683174 393488
rect 683132 392329 683160 393479
rect 683118 392320 683174 392329
rect 683118 392255 683174 392264
rect 683132 392018 683160 392255
rect 683120 392012 683172 392018
rect 683120 391954 683172 391960
rect 679622 388240 679678 388249
rect 679622 388175 679678 388184
rect 675300 387660 675352 387666
rect 675300 387602 675352 387608
rect 678244 387660 678296 387666
rect 678244 387602 678296 387608
rect 675312 386034 675340 387602
rect 675392 386164 675444 386170
rect 675392 386106 675444 386112
rect 675300 386028 675352 386034
rect 675300 385970 675352 385976
rect 675208 385824 675260 385830
rect 675208 385766 675260 385772
rect 675404 385696 675432 386106
rect 675392 385620 675444 385626
rect 675392 385562 675444 385568
rect 675404 385084 675432 385562
rect 675758 384976 675814 384985
rect 675758 384911 675814 384920
rect 675772 384435 675800 384911
rect 675300 383920 675352 383926
rect 675300 383862 675352 383868
rect 675312 381426 675340 383862
rect 675392 383104 675444 383110
rect 675392 383046 675444 383052
rect 675404 382568 675432 383046
rect 675390 382256 675446 382265
rect 675390 382191 675446 382200
rect 675404 382024 675432 382191
rect 675312 381398 675418 381426
rect 675116 381132 675168 381138
rect 675116 381074 675168 381080
rect 675392 381132 675444 381138
rect 675392 381074 675444 381080
rect 675404 380732 675432 381074
rect 675482 378720 675538 378729
rect 675482 378655 675538 378664
rect 675496 378284 675524 378655
rect 675404 377210 675432 377740
rect 675758 377360 675814 377369
rect 675758 377295 675814 377304
rect 675312 377182 675432 377210
rect 675312 376786 675340 377182
rect 675772 377060 675800 377295
rect 675300 376780 675352 376786
rect 675300 376722 675352 376728
rect 675484 376712 675536 376718
rect 675484 376654 675536 376660
rect 675496 376448 675524 376654
rect 675772 375057 675800 375224
rect 675758 375048 675814 375057
rect 675758 374983 675814 374992
rect 675758 373688 675814 373697
rect 675758 373623 675814 373632
rect 675772 373388 675800 373623
rect 675758 372056 675814 372065
rect 675758 371991 675814 372000
rect 675772 371552 675800 371991
rect 703694 359380 703722 359516
rect 704154 359380 704182 359516
rect 704614 359380 704642 359516
rect 705074 359380 705102 359516
rect 705534 359380 705562 359516
rect 705994 359380 706022 359516
rect 706454 359380 706482 359516
rect 706914 359380 706942 359516
rect 707374 359380 707402 359516
rect 707834 359380 707862 359516
rect 708294 359380 708322 359516
rect 708754 359380 708782 359516
rect 709214 359380 709242 359516
rect 675850 358728 675906 358737
rect 675850 358663 675906 358672
rect 675864 357610 675892 358663
rect 675942 358320 675998 358329
rect 675942 358255 675998 358264
rect 675956 357882 675984 358255
rect 676034 357912 676090 357921
rect 675944 357876 675996 357882
rect 676034 357847 676090 357856
rect 675944 357818 675996 357824
rect 676048 357746 676076 357847
rect 676036 357740 676088 357746
rect 676036 357682 676088 357688
rect 675852 357604 675904 357610
rect 675852 357546 675904 357552
rect 676036 357536 676088 357542
rect 676034 357504 676036 357513
rect 676088 357504 676090 357513
rect 676034 357439 676090 357448
rect 676034 357096 676090 357105
rect 676034 357031 676036 357040
rect 676088 357031 676090 357040
rect 676036 357002 676088 357008
rect 676036 356720 676088 356726
rect 676034 356688 676036 356697
rect 676088 356688 676090 356697
rect 676034 356623 676090 356632
rect 676034 356280 676090 356289
rect 676034 356215 676036 356224
rect 676088 356215 676090 356224
rect 676036 356186 676088 356192
rect 676036 355904 676088 355910
rect 676034 355872 676036 355881
rect 676088 355872 676090 355881
rect 676034 355807 676090 355816
rect 676034 355464 676090 355473
rect 676034 355399 676036 355408
rect 676088 355399 676090 355408
rect 676036 355370 676088 355376
rect 674746 355056 674802 355065
rect 674746 354991 674802 355000
rect 676034 354648 676090 354657
rect 676034 354583 676036 354592
rect 676088 354583 676090 354592
rect 676036 354554 676088 354560
rect 679622 352608 679678 352617
rect 679622 352543 679678 352552
rect 676034 351384 676090 351393
rect 676034 351319 676090 351328
rect 676048 351082 676076 351319
rect 676036 351076 676088 351082
rect 676036 351018 676088 351024
rect 676772 351076 676824 351082
rect 676772 351018 676824 351024
rect 676034 350976 676090 350985
rect 676034 350911 676036 350920
rect 676088 350911 676090 350920
rect 676036 350882 676088 350888
rect 676036 350600 676088 350606
rect 676034 350568 676036 350577
rect 676088 350568 676090 350577
rect 676034 350503 676090 350512
rect 676034 350160 676090 350169
rect 676090 350118 676168 350146
rect 676034 350095 676090 350104
rect 675942 349752 675998 349761
rect 675942 349687 675998 349696
rect 675956 346633 675984 349687
rect 676034 349344 676090 349353
rect 676034 349279 676036 349288
rect 676088 349279 676090 349288
rect 676036 349250 676088 349256
rect 676034 348936 676090 348945
rect 676034 348871 676036 348880
rect 676088 348871 676090 348880
rect 676036 348842 676088 348848
rect 676034 348528 676090 348537
rect 676034 348463 676090 348472
rect 676048 347313 676076 348463
rect 676034 347304 676090 347313
rect 676034 347239 676090 347248
rect 675942 346624 675998 346633
rect 675942 346559 675998 346568
rect 676048 346458 676076 347239
rect 676140 346497 676168 350118
rect 676784 346497 676812 351018
rect 676126 346488 676182 346497
rect 676036 346452 676088 346458
rect 676126 346423 676182 346432
rect 676770 346488 676826 346497
rect 676770 346423 676826 346432
rect 676036 346394 676088 346400
rect 679636 342417 679664 352543
rect 679806 351792 679862 351801
rect 679806 351727 679862 351736
rect 679622 342408 679678 342417
rect 679622 342343 679678 342352
rect 679820 342281 679848 351727
rect 675298 342272 675354 342281
rect 675298 342207 675354 342216
rect 679806 342272 679862 342281
rect 679806 342207 679862 342216
rect 675312 339878 675340 342207
rect 675666 340776 675722 340785
rect 675666 340711 675722 340720
rect 675680 340544 675708 340711
rect 675312 339850 675418 339878
rect 675758 339416 675814 339425
rect 675758 339351 675814 339360
rect 675772 339252 675800 339351
rect 675482 337920 675538 337929
rect 675482 337855 675538 337864
rect 675496 337416 675524 337855
rect 675404 336734 675432 336843
rect 674840 336728 674892 336734
rect 674840 336670 674892 336676
rect 675392 336728 675444 336734
rect 675392 336670 675444 336676
rect 674852 335345 674880 336670
rect 675392 336592 675444 336598
rect 675392 336534 675444 336540
rect 675404 336192 675432 336534
rect 675758 335880 675814 335889
rect 675758 335815 675814 335824
rect 675772 335580 675800 335815
rect 674838 335336 674894 335345
rect 674838 335271 674894 335280
rect 675758 333568 675814 333577
rect 675758 333503 675814 333512
rect 675772 333064 675800 333503
rect 675392 332648 675444 332654
rect 675392 332590 675444 332596
rect 675404 332520 675432 332590
rect 675758 332208 675814 332217
rect 675758 332143 675814 332152
rect 675772 331875 675800 332143
rect 675392 331628 675444 331634
rect 675392 331570 675444 331576
rect 675404 331228 675432 331570
rect 675392 330608 675444 330614
rect 675392 330550 675444 330556
rect 675404 330035 675432 330550
rect 675496 327690 675524 328168
rect 675116 327684 675168 327690
rect 675116 327626 675168 327632
rect 675484 327684 675536 327690
rect 675484 327626 675536 327632
rect 675128 325689 675156 327626
rect 675772 325854 675800 326332
rect 675760 325848 675812 325854
rect 675760 325790 675812 325796
rect 675114 325680 675170 325689
rect 675114 325615 675170 325624
rect 675760 325644 675812 325650
rect 675760 325586 675812 325592
rect 675772 325553 675800 325586
rect 675758 325544 675814 325553
rect 675758 325479 675814 325488
rect 703694 314364 703722 314500
rect 704154 314364 704182 314500
rect 704614 314364 704642 314500
rect 705074 314364 705102 314500
rect 705534 314364 705562 314500
rect 705994 314364 706022 314500
rect 706454 314364 706482 314500
rect 706914 314364 706942 314500
rect 707374 314364 707402 314500
rect 707834 314364 707862 314500
rect 708294 314364 708322 314500
rect 708754 314364 708782 314500
rect 709214 314364 709242 314500
rect 676218 313576 676274 313585
rect 676218 313511 676220 313520
rect 676272 313511 676274 313520
rect 676220 313482 676272 313488
rect 676036 313404 676088 313410
rect 676036 313346 676088 313352
rect 676048 313313 676076 313346
rect 676034 313304 676090 313313
rect 676034 313239 676090 313248
rect 676218 312760 676274 312769
rect 676218 312695 676274 312704
rect 674656 312520 674708 312526
rect 676036 312520 676088 312526
rect 674656 312462 674708 312468
rect 676034 312488 676036 312497
rect 676088 312488 676090 312497
rect 676034 312423 676090 312432
rect 676232 312050 676260 312695
rect 676220 312044 676272 312050
rect 676220 311986 676272 311992
rect 676218 311944 676274 311953
rect 674748 311908 674800 311914
rect 676218 311879 676220 311888
rect 674748 311850 674800 311856
rect 676272 311879 676274 311888
rect 676220 311850 676272 311856
rect 674472 311704 674524 311710
rect 674472 311646 674524 311652
rect 674656 311092 674708 311098
rect 674656 311034 674708 311040
rect 674564 304564 674616 304570
rect 674564 304506 674616 304512
rect 674576 291106 674604 304506
rect 674564 291100 674616 291106
rect 674564 291042 674616 291048
rect 674668 266694 674696 311034
rect 674760 267481 674788 311850
rect 676036 311704 676088 311710
rect 676034 311672 676036 311681
rect 676088 311672 676090 311681
rect 676034 311607 676090 311616
rect 676218 311128 676274 311137
rect 676218 311063 676220 311072
rect 676272 311063 676274 311072
rect 676220 311034 676272 311040
rect 676218 310720 676274 310729
rect 676218 310655 676220 310664
rect 676272 310655 676274 310664
rect 676220 310626 676272 310632
rect 676310 310312 676366 310321
rect 676310 310247 676366 310256
rect 676126 309904 676182 309913
rect 676126 309839 676182 309848
rect 676140 309398 676168 309839
rect 676218 309496 676274 309505
rect 676218 309431 676220 309440
rect 676272 309431 676274 309440
rect 676220 309402 676272 309408
rect 676128 309392 676180 309398
rect 676128 309334 676180 309340
rect 676324 309262 676352 310247
rect 676312 309256 676364 309262
rect 676312 309198 676364 309204
rect 681002 309088 681058 309097
rect 681002 309023 681058 309032
rect 679714 308272 679770 308281
rect 679714 308207 679770 308216
rect 679622 307864 679678 307873
rect 679622 307799 679678 307808
rect 676862 306640 676918 306649
rect 676862 306575 676918 306584
rect 676310 306232 676366 306241
rect 676310 306167 676366 306176
rect 676218 304600 676274 304609
rect 676218 304535 676220 304544
rect 676272 304535 676274 304544
rect 676220 304506 676272 304512
rect 676126 304192 676182 304201
rect 676126 304127 676182 304136
rect 676140 303686 676168 304127
rect 676218 303784 676274 303793
rect 676218 303719 676220 303728
rect 676272 303719 676274 303728
rect 676220 303690 676272 303696
rect 676128 303680 676180 303686
rect 676128 303622 676180 303628
rect 675116 298172 675168 298178
rect 675116 298114 675168 298120
rect 675128 294098 675156 298114
rect 675760 298104 675812 298110
rect 675760 298046 675812 298052
rect 675208 298036 675260 298042
rect 675208 297978 675260 297984
rect 675220 295254 675248 297978
rect 675772 296206 675800 298046
rect 676324 297401 676352 306167
rect 676402 305824 676458 305833
rect 676402 305759 676458 305768
rect 676416 298178 676444 305759
rect 676404 298172 676456 298178
rect 676404 298114 676456 298120
rect 676876 298042 676904 306575
rect 677598 305416 677654 305425
rect 677598 305351 677654 305360
rect 676864 298036 676916 298042
rect 676864 297978 676916 297984
rect 677612 297537 677640 305351
rect 679636 297809 679664 307799
rect 679728 298110 679756 308207
rect 681016 299441 681044 309023
rect 683118 303376 683174 303385
rect 683118 303311 683174 303320
rect 683132 302569 683160 303311
rect 683118 302560 683174 302569
rect 683118 302495 683174 302504
rect 683132 302258 683160 302495
rect 683120 302252 683172 302258
rect 683120 302194 683172 302200
rect 681002 299432 681058 299441
rect 681002 299367 681058 299376
rect 679716 298104 679768 298110
rect 679716 298046 679768 298052
rect 679622 297800 679678 297809
rect 679622 297735 679678 297744
rect 677598 297528 677654 297537
rect 677598 297463 677654 297472
rect 676310 297392 676366 297401
rect 676310 297327 676366 297336
rect 675760 296200 675812 296206
rect 675760 296142 675812 296148
rect 675760 295996 675812 296002
rect 675760 295938 675812 295944
rect 675772 295528 675800 295938
rect 675208 295248 675260 295254
rect 675208 295190 675260 295196
rect 675392 295248 675444 295254
rect 675392 295190 675444 295196
rect 675404 294879 675432 295190
rect 675758 294808 675814 294817
rect 675758 294743 675814 294752
rect 675772 294236 675800 294743
rect 675116 294092 675168 294098
rect 675116 294034 675168 294040
rect 675024 294024 675076 294030
rect 675024 293966 675076 293972
rect 675036 291786 675064 293966
rect 675666 292632 675722 292641
rect 675666 292567 675722 292576
rect 675680 292400 675708 292567
rect 675482 292088 675538 292097
rect 675482 292023 675538 292032
rect 675496 291856 675524 292023
rect 675024 291780 675076 291786
rect 675024 291722 675076 291728
rect 675392 291780 675444 291786
rect 675392 291722 675444 291728
rect 675404 291176 675432 291722
rect 675392 291100 675444 291106
rect 675392 291042 675444 291048
rect 675404 290564 675432 291042
rect 675758 288416 675814 288425
rect 675758 288351 675814 288360
rect 675772 288048 675800 288351
rect 675392 287972 675444 287978
rect 675392 287914 675444 287920
rect 675404 287504 675432 287914
rect 675758 287328 675814 287337
rect 675758 287263 675814 287272
rect 675772 286892 675800 287263
rect 675392 286612 675444 286618
rect 675392 286554 675444 286560
rect 675404 286212 675432 286554
rect 675482 285560 675538 285569
rect 675482 285495 675538 285504
rect 675496 285056 675524 285495
rect 675758 283656 675814 283665
rect 675758 283591 675814 283600
rect 675772 283220 675800 283591
rect 675758 281480 675814 281489
rect 675758 281415 675814 281424
rect 675772 281355 675800 281415
rect 703694 269348 703722 269484
rect 704154 269348 704182 269484
rect 704614 269348 704642 269484
rect 705074 269348 705102 269484
rect 705534 269348 705562 269484
rect 705994 269348 706022 269484
rect 706454 269348 706482 269484
rect 706914 269348 706942 269484
rect 707374 269348 707402 269484
rect 707834 269348 707862 269484
rect 708294 269348 708322 269484
rect 708754 269348 708782 269484
rect 709214 269348 709242 269484
rect 676218 268560 676274 268569
rect 676218 268495 676274 268504
rect 676126 268152 676182 268161
rect 676232 268122 676260 268495
rect 676126 268087 676182 268096
rect 676220 268116 676272 268122
rect 676140 267782 676168 268087
rect 676220 268058 676272 268064
rect 676220 267980 676272 267986
rect 676220 267922 676272 267928
rect 676128 267776 676180 267782
rect 676232 267753 676260 267922
rect 676128 267718 676180 267724
rect 676218 267744 676274 267753
rect 676218 267679 676274 267688
rect 674746 267472 674802 267481
rect 674746 267407 674802 267416
rect 676218 266928 676274 266937
rect 674748 266892 674800 266898
rect 676218 266863 676220 266872
rect 674748 266834 674800 266840
rect 676272 266863 676274 266872
rect 676220 266834 676272 266840
rect 674656 266688 674708 266694
rect 674656 266630 674708 266636
rect 674656 266076 674708 266082
rect 674656 266018 674708 266024
rect 674564 259140 674616 259146
rect 674564 259082 674616 259088
rect 674472 250028 674524 250034
rect 674472 249970 674524 249976
rect 674484 247314 674512 249970
rect 674576 249898 674604 259082
rect 674564 249892 674616 249898
rect 674564 249834 674616 249840
rect 674564 249756 674616 249762
rect 674564 249698 674616 249704
rect 674472 247308 674524 247314
rect 674472 247250 674524 247256
rect 674576 247110 674604 249698
rect 674564 247104 674616 247110
rect 674564 247046 674616 247052
rect 674380 222760 674432 222766
rect 674380 222702 674432 222708
rect 674668 221542 674696 266018
rect 674760 222329 674788 266834
rect 676036 266688 676088 266694
rect 676034 266656 676036 266665
rect 676088 266656 676090 266665
rect 676034 266591 676090 266600
rect 676218 266112 676274 266121
rect 676218 266047 676220 266056
rect 676272 266047 676274 266056
rect 676220 266018 676272 266024
rect 676218 265704 676274 265713
rect 676218 265639 676274 265648
rect 676126 265296 676182 265305
rect 676232 265266 676260 265639
rect 676126 265231 676182 265240
rect 676220 265260 676272 265266
rect 676036 265124 676088 265130
rect 676036 265066 676088 265072
rect 676048 265033 676076 265066
rect 676034 265024 676090 265033
rect 676140 264994 676168 265231
rect 676220 265202 676272 265208
rect 676034 264959 676090 264968
rect 676128 264988 676180 264994
rect 676128 264930 676180 264936
rect 676218 264480 676274 264489
rect 676218 264415 676274 264424
rect 676232 263634 676260 264415
rect 676220 263628 676272 263634
rect 676220 263570 676272 263576
rect 678242 263256 678298 263265
rect 678242 263191 678298 263200
rect 676862 261216 676918 261225
rect 676862 261151 676918 261160
rect 676402 259992 676458 260001
rect 676402 259927 676458 259936
rect 676218 259176 676274 259185
rect 676218 259111 676220 259120
rect 676272 259111 676274 259120
rect 676220 259082 676272 259088
rect 676218 258768 676274 258777
rect 676218 258703 676274 258712
rect 676232 258126 676260 258703
rect 676220 258120 676272 258126
rect 676220 258062 676272 258068
rect 675760 252612 675812 252618
rect 675760 252554 675812 252560
rect 675208 251660 675260 251666
rect 675208 251602 675260 251608
rect 675024 251592 675076 251598
rect 675024 251534 675076 251540
rect 675036 249762 675064 251534
rect 675220 250034 675248 251602
rect 675772 251258 675800 252554
rect 676416 251705 676444 259927
rect 676494 259584 676550 259593
rect 676494 259519 676550 259528
rect 676402 251696 676458 251705
rect 676508 251666 676536 259519
rect 676402 251631 676458 251640
rect 676496 251660 676548 251666
rect 676496 251602 676548 251608
rect 676876 251598 676904 261151
rect 676954 260808 677010 260817
rect 676954 260743 677010 260752
rect 676968 251598 676996 260743
rect 678256 252618 678284 263191
rect 678334 262440 678390 262449
rect 678334 262375 678390 262384
rect 678348 252657 678376 262375
rect 683118 258360 683174 258369
rect 683118 258295 683174 258304
rect 683132 257553 683160 258295
rect 683118 257544 683174 257553
rect 683118 257479 683174 257488
rect 683132 256766 683160 257479
rect 683120 256760 683172 256766
rect 683120 256702 683172 256708
rect 678334 252648 678390 252657
rect 678244 252612 678296 252618
rect 678334 252583 678390 252592
rect 678244 252554 678296 252560
rect 676864 251592 676916 251598
rect 676864 251534 676916 251540
rect 676956 251592 677008 251598
rect 676956 251534 677008 251540
rect 675760 251252 675812 251258
rect 675760 251194 675812 251200
rect 675760 250980 675812 250986
rect 675760 250922 675812 250928
rect 675772 250512 675800 250922
rect 675758 250336 675814 250345
rect 675758 250271 675814 250280
rect 675208 250028 675260 250034
rect 675208 249970 675260 249976
rect 675772 249900 675800 250271
rect 675758 249792 675814 249801
rect 675024 249756 675076 249762
rect 675758 249727 675814 249736
rect 675024 249698 675076 249704
rect 675022 249656 675078 249665
rect 675022 249591 675078 249600
rect 675036 247926 675064 249591
rect 675206 249520 675262 249529
rect 675206 249455 675262 249464
rect 675220 248538 675248 249455
rect 675772 249220 675800 249727
rect 675208 248532 675260 248538
rect 675208 248474 675260 248480
rect 675208 248328 675260 248334
rect 675208 248270 675260 248276
rect 675024 247920 675076 247926
rect 675024 247862 675076 247868
rect 675116 247308 675168 247314
rect 675116 247250 675168 247256
rect 675128 246090 675156 247250
rect 675220 246265 675248 248270
rect 675484 247920 675536 247926
rect 675484 247862 675536 247868
rect 675496 247384 675524 247862
rect 675392 247104 675444 247110
rect 675392 247046 675444 247052
rect 675404 246840 675432 247046
rect 675392 246560 675444 246566
rect 675392 246502 675444 246508
rect 675206 246256 675262 246265
rect 675206 246191 675262 246200
rect 675404 246199 675432 246502
rect 675116 246084 675168 246090
rect 675116 246026 675168 246032
rect 675392 246084 675444 246090
rect 675392 246026 675444 246032
rect 675404 245548 675432 246026
rect 675300 243636 675352 243642
rect 675300 243578 675352 243584
rect 675312 243085 675340 243578
rect 675312 243057 675418 243085
rect 675300 242888 675352 242894
rect 675300 242830 675352 242836
rect 675312 242533 675340 242830
rect 675312 242505 675418 242533
rect 675298 241904 675354 241913
rect 675354 241862 675418 241890
rect 675298 241839 675354 241848
rect 675300 241256 675352 241262
rect 675352 241217 675418 241245
rect 675300 241198 675352 241204
rect 675390 240272 675446 240281
rect 675390 240207 675446 240216
rect 675404 240040 675432 240207
rect 675758 238504 675814 238513
rect 675758 238439 675814 238448
rect 675772 238204 675800 238439
rect 675758 236872 675814 236881
rect 675758 236807 675814 236816
rect 675772 236368 675800 236807
rect 703694 224196 703722 224264
rect 704154 224196 704182 224264
rect 704614 224196 704642 224264
rect 705074 224196 705102 224264
rect 705534 224196 705562 224264
rect 705994 224196 706022 224264
rect 706454 224196 706482 224264
rect 706914 224196 706942 224264
rect 707374 224196 707402 224264
rect 707834 224196 707862 224264
rect 708294 224196 708322 224264
rect 708754 224196 708782 224264
rect 709214 224196 709242 224264
rect 676034 223544 676090 223553
rect 676034 223479 676090 223488
rect 675944 223168 675996 223174
rect 675942 223136 675944 223145
rect 675996 223136 675998 223145
rect 675942 223071 675998 223080
rect 675944 222760 675996 222766
rect 675942 222728 675944 222737
rect 675996 222728 675998 222737
rect 675942 222663 675998 222672
rect 674746 222320 674802 222329
rect 674746 222255 674802 222264
rect 676048 222222 676076 223479
rect 676036 222216 676088 222222
rect 676036 222158 676088 222164
rect 676034 221912 676090 221921
rect 676034 221847 676036 221856
rect 676088 221847 676090 221856
rect 676036 221818 676088 221824
rect 674656 221536 674708 221542
rect 676036 221536 676088 221542
rect 674656 221478 674708 221484
rect 676034 221504 676036 221513
rect 676088 221504 676090 221513
rect 676034 221439 676090 221448
rect 676034 221096 676090 221105
rect 676034 221031 676036 221040
rect 676088 221031 676090 221040
rect 676036 221002 676088 221008
rect 676036 220720 676088 220726
rect 676034 220688 676036 220697
rect 676088 220688 676090 220697
rect 676034 220623 676090 220632
rect 676034 220280 676090 220289
rect 674656 220244 674708 220250
rect 676034 220215 676036 220224
rect 674656 220186 674708 220192
rect 676088 220215 676090 220224
rect 676036 220186 676088 220192
rect 674380 216164 674432 216170
rect 674380 216106 674432 216112
rect 674392 201890 674420 216106
rect 674472 215756 674524 215762
rect 674472 215698 674524 215704
rect 674380 201884 674432 201890
rect 674380 201826 674432 201832
rect 674484 201482 674512 215698
rect 674564 213716 674616 213722
rect 674564 213658 674616 213664
rect 674472 201476 674524 201482
rect 674472 201418 674524 201424
rect 674576 196586 674604 213658
rect 674564 196580 674616 196586
rect 674564 196522 674616 196528
rect 674564 176044 674616 176050
rect 674564 175986 674616 175992
rect 674576 175386 674604 175986
rect 674668 175710 674696 220186
rect 676036 219904 676088 219910
rect 676034 219872 676036 219881
rect 676088 219872 676090 219881
rect 676034 219807 676090 219816
rect 674746 219464 674802 219473
rect 674746 219399 674802 219408
rect 674656 175704 674708 175710
rect 674656 175646 674708 175652
rect 674576 175358 674696 175386
rect 674564 175228 674616 175234
rect 674564 175170 674616 175176
rect 674472 170332 674524 170338
rect 674472 170274 674524 170280
rect 674380 169108 674432 169114
rect 674380 169050 674432 169056
rect 674392 152590 674420 169050
rect 674380 152584 674432 152590
rect 674380 152526 674432 152532
rect 674484 150414 674512 170274
rect 674472 150408 674524 150414
rect 674472 150350 674524 150356
rect 674288 133000 674340 133006
rect 674288 132942 674340 132948
rect 674576 130558 674604 175170
rect 674668 131374 674696 175358
rect 674760 174865 674788 219399
rect 676034 219056 676090 219065
rect 676090 219014 676352 219042
rect 676034 218991 676090 219000
rect 676034 216608 676090 216617
rect 676090 216566 676260 216594
rect 676034 216543 676090 216552
rect 676034 216200 676090 216209
rect 676034 216135 676036 216144
rect 676088 216135 676090 216144
rect 676036 216106 676088 216112
rect 676232 215966 676260 216566
rect 676220 215960 676272 215966
rect 676220 215902 676272 215908
rect 676034 215792 676090 215801
rect 676034 215727 676036 215736
rect 676088 215727 676090 215736
rect 676036 215698 676088 215704
rect 675942 215384 675998 215393
rect 675942 215319 675998 215328
rect 675850 214976 675906 214985
rect 675850 214911 675906 214920
rect 675864 211313 675892 214911
rect 675956 211449 675984 215319
rect 676034 214160 676090 214169
rect 676034 214095 676036 214104
rect 676088 214095 676090 214104
rect 676036 214066 676088 214072
rect 676034 214024 676090 214033
rect 676324 214010 676352 219014
rect 679622 217424 679678 217433
rect 679622 217359 679678 217368
rect 676864 215960 676916 215966
rect 676864 215902 676916 215908
rect 676090 213982 676352 214010
rect 676034 213959 676090 213968
rect 676034 213752 676090 213761
rect 676034 213687 676036 213696
rect 676088 213687 676090 213696
rect 676036 213658 676088 213664
rect 676034 213344 676090 213353
rect 676034 213279 676090 213288
rect 676048 212129 676076 213279
rect 676034 212120 676090 212129
rect 676034 212055 676090 212064
rect 675942 211440 675998 211449
rect 675942 211375 675998 211384
rect 675850 211304 675906 211313
rect 675850 211239 675906 211248
rect 676048 211206 676076 212055
rect 676036 211200 676088 211206
rect 676036 211142 676088 211148
rect 676876 208321 676904 215902
rect 676862 208312 676918 208321
rect 676862 208247 676918 208256
rect 679636 207233 679664 217359
rect 679622 207224 679678 207233
rect 679622 207159 679678 207168
rect 675390 205592 675446 205601
rect 675390 205527 675446 205536
rect 675404 205323 675432 205527
rect 675758 205048 675814 205057
rect 675758 204983 675814 204992
rect 675772 204680 675800 204983
rect 675758 204232 675814 204241
rect 675758 204167 675814 204176
rect 675772 204035 675800 204167
rect 675114 202872 675170 202881
rect 675114 202807 675170 202816
rect 674838 201376 674894 201385
rect 674838 201311 674894 201320
rect 674852 197062 674880 201311
rect 675128 200734 675156 202807
rect 675758 202736 675814 202745
rect 675758 202671 675814 202680
rect 675772 202195 675800 202671
rect 675392 201884 675444 201890
rect 675392 201826 675444 201832
rect 675404 201620 675432 201826
rect 675392 201476 675444 201482
rect 675392 201418 675444 201424
rect 675404 201008 675432 201418
rect 675116 200728 675168 200734
rect 675116 200670 675168 200676
rect 675392 200728 675444 200734
rect 675392 200670 675444 200676
rect 675404 200328 675432 200670
rect 675482 198384 675538 198393
rect 675482 198319 675538 198328
rect 675496 197880 675524 198319
rect 675484 197464 675536 197470
rect 675484 197406 675536 197412
rect 675496 197336 675524 197406
rect 674840 197056 674892 197062
rect 674840 196998 674892 197004
rect 675392 197056 675444 197062
rect 675392 196998 675444 197004
rect 675404 196656 675432 196998
rect 675392 196580 675444 196586
rect 675392 196522 675444 196528
rect 675404 196044 675432 196522
rect 675758 195392 675814 195401
rect 675758 195327 675814 195336
rect 675772 194820 675800 195327
rect 675404 192506 675432 192984
rect 674840 192500 674892 192506
rect 674840 192442 674892 192448
rect 675392 192500 675444 192506
rect 675392 192442 675444 192448
rect 674852 190233 674880 192442
rect 675772 190670 675800 191148
rect 675760 190664 675812 190670
rect 675760 190606 675812 190612
rect 675760 190392 675812 190398
rect 675758 190360 675760 190369
rect 675812 190360 675814 190369
rect 675758 190295 675814 190304
rect 674838 190224 674894 190233
rect 674838 190159 674894 190168
rect 703694 179180 703722 179316
rect 704154 179180 704182 179316
rect 704614 179180 704642 179316
rect 705074 179180 705102 179316
rect 705534 179180 705562 179316
rect 705994 179180 706022 179316
rect 706454 179180 706482 179316
rect 706914 179180 706942 179316
rect 707374 179180 707402 179316
rect 707834 179180 707862 179316
rect 708294 179180 708322 179316
rect 708754 179180 708782 179316
rect 709214 179180 709242 179316
rect 676034 178528 676090 178537
rect 676034 178463 676090 178472
rect 676048 178226 676076 178463
rect 676036 178220 676088 178226
rect 676036 178162 676088 178168
rect 676034 178120 676090 178129
rect 676034 178055 676036 178064
rect 676088 178055 676090 178064
rect 676036 178026 676088 178032
rect 675942 177712 675998 177721
rect 675942 177647 675998 177656
rect 675956 176866 675984 177647
rect 676034 177304 676090 177313
rect 676034 177239 676090 177248
rect 676048 177002 676076 177239
rect 676036 176996 676088 177002
rect 676036 176938 676088 176944
rect 676034 176896 676090 176905
rect 675944 176860 675996 176866
rect 676034 176831 676090 176840
rect 675944 176802 675996 176808
rect 676048 176798 676076 176831
rect 676036 176792 676088 176798
rect 676036 176734 676088 176740
rect 676036 176520 676088 176526
rect 676034 176488 676036 176497
rect 676088 176488 676090 176497
rect 676034 176423 676090 176432
rect 676034 176080 676090 176089
rect 676034 176015 676036 176024
rect 676088 176015 676090 176024
rect 676036 175986 676088 175992
rect 676036 175704 676088 175710
rect 676034 175672 676036 175681
rect 676088 175672 676090 175681
rect 676034 175607 676090 175616
rect 676034 175264 676090 175273
rect 676034 175199 676036 175208
rect 676088 175199 676090 175208
rect 676036 175170 676088 175176
rect 674746 174856 674802 174865
rect 674746 174791 674802 174800
rect 676034 174448 676090 174457
rect 676034 174383 676036 174392
rect 676088 174383 676090 174392
rect 676036 174354 676088 174360
rect 678242 174040 678298 174049
rect 678242 173975 678298 173984
rect 676034 173224 676090 173233
rect 676034 173159 676090 173168
rect 676048 172582 676076 173159
rect 674840 172576 674892 172582
rect 674840 172518 674892 172524
rect 676036 172576 676088 172582
rect 676036 172518 676088 172524
rect 674852 160818 674880 172518
rect 676862 171592 676918 171601
rect 676862 171527 676918 171536
rect 676034 170776 676090 170785
rect 676090 170734 676260 170762
rect 676034 170711 676090 170720
rect 676034 170368 676090 170377
rect 676034 170303 676036 170312
rect 676088 170303 676090 170312
rect 676036 170274 676088 170280
rect 676034 169552 676090 169561
rect 676034 169487 676036 169496
rect 676088 169487 676090 169496
rect 676036 169458 676088 169464
rect 676034 169144 676090 169153
rect 676034 169079 676036 169088
rect 676088 169079 676090 169088
rect 676036 169050 676088 169056
rect 676034 168736 676090 168745
rect 676034 168671 676036 168680
rect 676088 168671 676090 168680
rect 676036 168642 676088 168648
rect 676034 168328 676090 168337
rect 676034 168263 676036 168272
rect 676088 168263 676090 168272
rect 676036 168234 676088 168240
rect 676034 167920 676090 167929
rect 676034 167855 676036 167864
rect 676088 167855 676090 167864
rect 676036 167826 676088 167832
rect 676034 167104 676090 167113
rect 676034 167039 676036 167048
rect 676088 167039 676090 167048
rect 676036 167010 676088 167016
rect 676232 162761 676260 170734
rect 676586 169960 676642 169969
rect 676586 169895 676642 169904
rect 676600 166433 676628 169895
rect 676876 166433 676904 171527
rect 676586 166424 676642 166433
rect 676586 166359 676642 166368
rect 676862 166424 676918 166433
rect 676862 166359 676918 166368
rect 676218 162752 676274 162761
rect 676218 162687 676274 162696
rect 678256 162625 678284 173975
rect 681002 172408 681058 172417
rect 681002 172343 681058 172352
rect 678426 171184 678482 171193
rect 678426 171119 678482 171128
rect 678242 162616 678298 162625
rect 678242 162551 678298 162560
rect 678440 162489 678468 171119
rect 678426 162480 678482 162489
rect 678426 162415 678482 162424
rect 681016 162353 681044 172343
rect 681002 162344 681058 162353
rect 681002 162279 681058 162288
rect 674840 160812 674892 160818
rect 674840 160754 674892 160760
rect 675484 160812 675536 160818
rect 675484 160754 675536 160760
rect 675496 160344 675524 160754
rect 675758 160032 675814 160041
rect 675758 159967 675814 159976
rect 675772 159664 675800 159967
rect 675758 159488 675814 159497
rect 675758 159423 675814 159432
rect 675772 159052 675800 159423
rect 675758 157448 675814 157457
rect 675758 157383 675814 157392
rect 675772 157216 675800 157383
rect 675666 157040 675722 157049
rect 675666 156975 675722 156984
rect 675680 156643 675708 156975
rect 675574 156496 675630 156505
rect 675574 156431 675630 156440
rect 675588 155992 675616 156431
rect 675484 155508 675536 155514
rect 675484 155450 675536 155456
rect 675496 155380 675524 155450
rect 675390 153096 675446 153105
rect 675390 153031 675446 153040
rect 675404 152864 675432 153031
rect 675392 152584 675444 152590
rect 675392 152526 675444 152532
rect 675404 152320 675432 152526
rect 675772 151609 675800 151675
rect 675758 151600 675814 151609
rect 675758 151535 675814 151544
rect 675392 151428 675444 151434
rect 675392 151370 675444 151376
rect 675404 151028 675432 151370
rect 675392 150408 675444 150414
rect 675392 150350 675444 150356
rect 675404 149835 675432 150350
rect 675758 148472 675814 148481
rect 675758 148407 675814 148416
rect 675772 147968 675800 148407
rect 675758 146296 675814 146305
rect 675758 146231 675814 146240
rect 675772 146132 675800 146231
rect 703694 133892 703722 134028
rect 704154 133892 704182 134028
rect 704614 133892 704642 134028
rect 705074 133892 705102 134028
rect 705534 133892 705562 134028
rect 705994 133892 706022 134028
rect 706454 133892 706482 134028
rect 706914 133892 706942 134028
rect 707374 133892 707402 134028
rect 707834 133892 707862 134028
rect 708294 133892 708322 134028
rect 708754 133892 708782 134028
rect 709214 133892 709242 134028
rect 676126 133104 676182 133113
rect 676126 133039 676182 133048
rect 676034 132968 676090 132977
rect 676034 132903 676036 132912
rect 676088 132903 676090 132912
rect 676036 132874 676088 132880
rect 676140 132666 676168 133039
rect 676220 132796 676272 132802
rect 676220 132738 676272 132744
rect 676232 132705 676260 132738
rect 676218 132696 676274 132705
rect 676128 132660 676180 132666
rect 676218 132631 676274 132640
rect 676128 132602 676180 132608
rect 676220 132320 676272 132326
rect 676218 132288 676220 132297
rect 676272 132288 676274 132297
rect 676218 132223 676274 132232
rect 676218 131472 676274 131481
rect 676218 131407 676274 131416
rect 674656 131368 674708 131374
rect 676036 131368 676088 131374
rect 674656 131310 674708 131316
rect 676034 131336 676036 131345
rect 676088 131336 676090 131345
rect 676034 131271 676090 131280
rect 676232 131170 676260 131407
rect 676220 131164 676272 131170
rect 676220 131106 676272 131112
rect 676218 130656 676274 130665
rect 676218 130591 676274 130600
rect 674564 130552 674616 130558
rect 676036 130552 676088 130558
rect 674564 130494 674616 130500
rect 676034 130520 676036 130529
rect 676088 130520 676090 130529
rect 676034 130455 676090 130464
rect 676232 129946 676260 130591
rect 676220 129940 676272 129946
rect 676220 129882 676272 129888
rect 676218 129840 676274 129849
rect 676218 129775 676220 129784
rect 676272 129775 676274 129784
rect 676220 129746 676272 129752
rect 676126 129432 676182 129441
rect 676126 129367 676182 129376
rect 676140 128586 676168 129367
rect 676218 129024 676274 129033
rect 676218 128959 676274 128968
rect 676128 128580 676180 128586
rect 676128 128522 676180 128528
rect 676232 128382 676260 128959
rect 676220 128376 676272 128382
rect 676220 128318 676272 128324
rect 683670 128208 683726 128217
rect 683670 128143 683726 128152
rect 676034 128072 676090 128081
rect 676034 128007 676090 128016
rect 676048 127022 676076 128007
rect 683118 127392 683174 127401
rect 683118 127327 683174 127336
rect 675116 127016 675168 127022
rect 675116 126958 675168 126964
rect 676036 127016 676088 127022
rect 676036 126958 676088 126964
rect 676862 126984 676918 126993
rect 674746 123584 674802 123593
rect 674746 123519 674802 123528
rect 674104 117836 674156 117842
rect 674104 117778 674156 117784
rect 674656 116272 674708 116278
rect 674656 116214 674708 116220
rect 674668 114646 674696 116214
rect 674656 114640 674708 114646
rect 674656 114582 674708 114588
rect 673368 106344 673420 106350
rect 673368 106286 673420 106292
rect 674760 106282 674788 123519
rect 675128 115598 675156 126958
rect 676862 126919 676918 126928
rect 676402 125352 676458 125361
rect 676402 125287 676458 125296
rect 676218 123720 676274 123729
rect 676218 123655 676274 123664
rect 676232 123010 676260 123655
rect 676220 123004 676272 123010
rect 676220 122946 676272 122952
rect 676218 122904 676274 122913
rect 676218 122839 676220 122848
rect 676272 122839 676274 122848
rect 676220 122810 676272 122816
rect 676126 122496 676182 122505
rect 676126 122431 676182 122440
rect 676140 121514 676168 122431
rect 676218 121680 676274 121689
rect 676218 121615 676274 121624
rect 676128 121508 676180 121514
rect 676128 121450 676180 121456
rect 676232 120766 676260 121615
rect 676220 120760 676272 120766
rect 676220 120702 676272 120708
rect 676416 117337 676444 125287
rect 676876 118017 676904 126919
rect 679622 125760 679678 125769
rect 679622 125695 679678 125704
rect 678242 125352 678298 125361
rect 678242 125287 678298 125296
rect 677598 124128 677654 124137
rect 677598 124063 677654 124072
rect 676862 118008 676918 118017
rect 676862 117943 676918 117952
rect 676402 117328 676458 117337
rect 676402 117263 676458 117272
rect 675208 116612 675260 116618
rect 675208 116554 675260 116560
rect 675116 115592 675168 115598
rect 675116 115534 675168 115540
rect 675116 115456 675168 115462
rect 675116 115398 675168 115404
rect 675128 114730 675156 115398
rect 675220 114850 675248 116554
rect 677612 116278 677640 124063
rect 677600 116272 677652 116278
rect 677600 116214 677652 116220
rect 678256 116210 678284 125287
rect 679636 117201 679664 125695
rect 683132 124953 683160 127327
rect 683302 126168 683358 126177
rect 683302 126103 683358 126112
rect 683118 124944 683174 124953
rect 683118 124879 683174 124888
rect 679622 117192 679678 117201
rect 679622 117127 679678 117136
rect 683316 116618 683344 126103
rect 683684 121689 683712 128143
rect 683670 121680 683726 121689
rect 683670 121615 683726 121624
rect 683304 116612 683356 116618
rect 683304 116554 683356 116560
rect 678244 116204 678296 116210
rect 678244 116146 678296 116152
rect 675392 115592 675444 115598
rect 675392 115534 675444 115540
rect 675404 115124 675432 115534
rect 675208 114844 675260 114850
rect 675208 114786 675260 114792
rect 675392 114844 675444 114850
rect 675392 114786 675444 114792
rect 675128 114702 675248 114730
rect 675116 114640 675168 114646
rect 675116 114582 675168 114588
rect 675128 110702 675156 114582
rect 675220 111178 675248 114702
rect 675404 114479 675432 114786
rect 675758 114200 675814 114209
rect 675758 114135 675814 114144
rect 675772 113832 675800 114135
rect 675758 112568 675814 112577
rect 675758 112503 675814 112512
rect 675772 111996 675800 112503
rect 675482 111752 675538 111761
rect 675482 111687 675538 111696
rect 675496 111452 675524 111687
rect 675208 111172 675260 111178
rect 675208 111114 675260 111120
rect 675392 111172 675444 111178
rect 675392 111114 675444 111120
rect 675404 110772 675432 111114
rect 675116 110696 675168 110702
rect 675116 110638 675168 110644
rect 675392 110696 675444 110702
rect 675392 110638 675444 110644
rect 675404 110160 675432 110638
rect 675114 109032 675170 109041
rect 675114 108967 675170 108976
rect 675128 107030 675156 108967
rect 675758 108216 675814 108225
rect 675758 108151 675814 108160
rect 675772 107644 675800 108151
rect 675116 107024 675168 107030
rect 675116 106966 675168 106972
rect 675392 107024 675444 107030
rect 675392 106966 675444 106972
rect 675404 106488 675432 106966
rect 675496 106622 675524 107100
rect 675484 106616 675536 106622
rect 675484 106558 675536 106564
rect 674748 106276 674800 106282
rect 674748 106218 674800 106224
rect 675392 106276 675444 106282
rect 675392 106218 675444 106224
rect 672724 106140 672776 106146
rect 672724 106082 672776 106088
rect 675404 105808 675432 106218
rect 675482 104816 675538 104825
rect 675482 104751 675538 104760
rect 675496 104652 675524 104751
rect 675758 103184 675814 103193
rect 675758 103119 675814 103128
rect 675772 102816 675800 103119
rect 675758 101416 675814 101425
rect 675758 101351 675814 101360
rect 675772 100980 675800 101351
rect 664444 49088 664496 49094
rect 664444 49030 664496 49036
rect 669964 49088 670016 49094
rect 669964 49030 670016 49036
rect 664456 48521 664484 49030
rect 664442 48512 664498 48521
rect 664442 48447 664498 48456
rect 662418 47424 662474 47433
rect 662418 47359 662474 47368
rect 661130 44840 661186 44849
rect 661130 44775 661186 44784
rect 611358 41576 611414 41585
rect 611358 41511 611414 41520
rect 609978 41440 610034 41449
rect 609978 41375 610034 41384
rect 141698 40352 141754 40361
rect 141698 40287 141754 40296
rect 141712 39984 141740 40287
<< via2 >>
rect 154578 1007140 154634 1007176
rect 154578 1007120 154580 1007140
rect 154580 1007120 154632 1007140
rect 154632 1007120 154634 1007140
rect 80978 995696 81034 995752
rect 82358 995696 82414 995752
rect 92478 995696 92534 995752
rect 41786 968768 41842 968824
rect 41786 967272 41842 967328
rect 41786 965096 41842 965152
rect 41786 963464 41842 963520
rect 41786 962104 41842 962160
rect 42062 958432 42118 958488
rect 41786 957752 41842 957808
rect 31022 952856 31078 952912
rect 27618 943744 27674 943800
rect 36726 952312 36782 952368
rect 36542 952176 36598 952232
rect 35806 943064 35862 943120
rect 35714 942656 35770 942712
rect 32402 938168 32458 938224
rect 31022 937352 31078 937408
rect 41970 943744 42026 943800
rect 41786 941840 41842 941896
rect 37922 936536 37978 936592
rect 36726 936128 36782 936184
rect 36542 935312 36598 935368
rect 39946 933272 40002 933328
rect 41234 817944 41290 818000
rect 41326 817264 41382 817320
rect 41786 941024 41842 941080
rect 41694 939256 41750 939312
rect 41694 932204 41750 932240
rect 41694 932184 41696 932204
rect 41696 932184 41748 932204
rect 41748 932184 41750 932204
rect 41878 940208 41934 940264
rect 42154 938984 42210 939040
rect 41970 938576 42026 938632
rect 42982 935720 43038 935776
rect 44822 940616 44878 940672
rect 46202 942248 46258 942304
rect 47582 941432 47638 941488
rect 84658 995560 84714 995616
rect 85210 995560 85266 995616
rect 86038 995560 86094 995616
rect 88890 995424 88946 995480
rect 87510 995152 87566 995208
rect 93122 995832 93178 995888
rect 94778 997192 94834 997248
rect 94502 996920 94558 996976
rect 93306 995560 93362 995616
rect 103150 1006460 103206 1006496
rect 103150 1006440 103152 1006460
rect 103152 1006440 103204 1006460
rect 103204 1006440 103206 1006460
rect 103610 1006476 103612 1006496
rect 103612 1006476 103664 1006496
rect 103664 1006476 103666 1006496
rect 103610 1006440 103666 1006476
rect 98274 1006068 98276 1006088
rect 98276 1006068 98328 1006088
rect 98328 1006068 98330 1006088
rect 98274 1006032 98330 1006068
rect 99102 1006068 99104 1006088
rect 99104 1006068 99156 1006088
rect 99156 1006068 99158 1006088
rect 99102 1006032 99158 1006068
rect 99470 1002124 99472 1002144
rect 99472 1002124 99524 1002144
rect 99524 1002124 99526 1002144
rect 99470 1002088 99526 1002124
rect 99930 1001972 99986 1002008
rect 99930 1001952 99932 1001972
rect 99932 1001952 99984 1001972
rect 99984 1001952 99986 1001972
rect 100666 1006324 100722 1006360
rect 100666 1006304 100668 1006324
rect 100668 1006304 100720 1006324
rect 100720 1006304 100722 1006324
rect 104346 1006340 104348 1006360
rect 104348 1006340 104400 1006360
rect 104400 1006340 104402 1006360
rect 104346 1006304 104402 1006340
rect 108854 1006324 108910 1006360
rect 108854 1006304 108856 1006324
rect 108856 1006304 108908 1006324
rect 108908 1006304 108910 1006324
rect 101954 1006204 101956 1006224
rect 101956 1006204 102008 1006224
rect 102008 1006204 102010 1006224
rect 101954 1006168 102010 1006204
rect 100298 1002244 100354 1002280
rect 100298 1002224 100300 1002244
rect 100300 1002224 100352 1002244
rect 100352 1002224 100354 1002244
rect 101494 1002108 101550 1002144
rect 101494 1002088 101496 1002108
rect 101496 1002088 101548 1002108
rect 101548 1002088 101550 1002108
rect 101126 1001988 101128 1002008
rect 101128 1001988 101180 1002008
rect 101180 1001988 101182 1002008
rect 101126 1001952 101182 1001988
rect 102322 1001972 102378 1002008
rect 102322 1001952 102324 1001972
rect 102324 1001952 102376 1001972
rect 102376 1001952 102378 1001972
rect 98642 995152 98698 995208
rect 80150 995016 80206 995072
rect 95882 995016 95938 995072
rect 104806 1006188 104862 1006224
rect 104806 1006168 104808 1006188
rect 104808 1006168 104860 1006188
rect 104860 1006168 104862 1006188
rect 108486 1006204 108488 1006224
rect 108488 1006204 108540 1006224
rect 108540 1006204 108542 1006224
rect 108486 1006168 108542 1006204
rect 103150 1004692 103206 1004728
rect 103150 1004672 103152 1004692
rect 103152 1004672 103204 1004692
rect 103204 1004672 103206 1004692
rect 106830 1002380 106886 1002416
rect 106830 1002360 106832 1002380
rect 106832 1002360 106884 1002380
rect 106884 1002360 106886 1002380
rect 106002 1002244 106058 1002280
rect 108486 1002260 108488 1002280
rect 108488 1002260 108540 1002280
rect 108540 1002260 108542 1002280
rect 106002 1002224 106004 1002244
rect 106004 1002224 106056 1002244
rect 106056 1002224 106058 1002244
rect 105634 1002108 105690 1002144
rect 105634 1002088 105636 1002108
rect 105636 1002088 105688 1002108
rect 105688 1002088 105690 1002108
rect 104346 1001988 104348 1002008
rect 104348 1001988 104400 1002008
rect 104400 1001988 104402 1002008
rect 104346 1001952 104402 1001988
rect 108486 1002224 108542 1002260
rect 107658 1002124 107660 1002144
rect 107660 1002124 107712 1002144
rect 107712 1002124 107714 1002144
rect 107658 1002088 107714 1002124
rect 106462 1001972 106518 1002008
rect 107198 1001988 107200 1002008
rect 107200 1001988 107252 1002008
rect 107252 1001988 107254 1002008
rect 106462 1001952 106464 1001972
rect 106464 1001952 106516 1001972
rect 106516 1001952 106518 1001972
rect 107198 1001952 107254 1001988
rect 108026 1001972 108082 1002008
rect 108026 1001952 108028 1001972
rect 108028 1001952 108080 1001972
rect 108080 1001952 108082 1001972
rect 111798 1001952 111854 1002008
rect 109866 997192 109922 997248
rect 112994 997192 113050 997248
rect 116122 997228 116124 997248
rect 116124 997228 116176 997248
rect 116176 997228 116178 997248
rect 116122 997192 116178 997228
rect 116122 997092 116124 997112
rect 116124 997092 116176 997112
rect 116176 997092 116178 997112
rect 116122 997056 116178 997092
rect 122102 990936 122158 990992
rect 129370 995696 129426 995752
rect 133142 995696 133198 995752
rect 143998 1000592 144054 1000648
rect 143814 997192 143870 997248
rect 136546 995560 136602 995616
rect 130014 995424 130070 995480
rect 132130 995288 132186 995344
rect 131578 995152 131634 995208
rect 144826 995696 144882 995752
rect 145654 997056 145710 997112
rect 203890 1007004 203946 1007040
rect 203890 1006984 203892 1007004
rect 203892 1006984 203944 1007004
rect 203944 1006984 203946 1007004
rect 308954 1007004 309010 1007040
rect 308954 1006984 308956 1007004
rect 308956 1006984 309008 1007004
rect 309008 1006984 309010 1007004
rect 154118 1006460 154174 1006496
rect 154118 1006440 154120 1006460
rect 154120 1006440 154172 1006460
rect 154172 1006440 154174 1006460
rect 149702 1006068 149704 1006088
rect 149704 1006068 149756 1006088
rect 149756 1006068 149758 1006088
rect 149702 1006032 149758 1006068
rect 150438 1006068 150440 1006088
rect 150440 1006068 150492 1006088
rect 150492 1006068 150494 1006088
rect 150438 1006032 150494 1006068
rect 156142 1006188 156198 1006224
rect 156142 1006168 156144 1006188
rect 156144 1006168 156196 1006188
rect 156196 1006168 156198 1006188
rect 151726 1006032 151782 1006088
rect 157430 1006068 157432 1006088
rect 157432 1006068 157484 1006088
rect 157484 1006068 157486 1006088
rect 157430 1006032 157486 1006068
rect 159086 1006068 159088 1006088
rect 159088 1006068 159140 1006088
rect 159140 1006068 159142 1006088
rect 159086 1006032 159142 1006068
rect 160650 1006052 160706 1006088
rect 160650 1006032 160652 1006052
rect 160652 1006032 160704 1006052
rect 160704 1006032 160706 1006052
rect 152554 1005388 152556 1005408
rect 152556 1005388 152608 1005408
rect 152608 1005388 152610 1005408
rect 152554 1005352 152610 1005388
rect 152922 1004964 152978 1005000
rect 152922 1004944 152924 1004964
rect 152924 1004944 152976 1004964
rect 152976 1004944 152978 1004964
rect 146942 996104 146998 996160
rect 148506 1000592 148562 1000648
rect 153750 1004828 153806 1004864
rect 153750 1004808 153752 1004828
rect 153752 1004808 153804 1004828
rect 153804 1004808 153806 1004828
rect 150898 1001972 150954 1002008
rect 150898 1001952 150900 1001972
rect 150900 1001952 150952 1001972
rect 150952 1001952 150954 1001972
rect 152094 1004708 152096 1004728
rect 152096 1004708 152148 1004728
rect 152148 1004708 152150 1004728
rect 152094 1004672 152150 1004708
rect 153290 1004692 153346 1004728
rect 153290 1004672 153292 1004692
rect 153292 1004672 153344 1004692
rect 153344 1004672 153346 1004692
rect 151082 995832 151138 995888
rect 148322 995560 148378 995616
rect 145562 995424 145618 995480
rect 151726 1001988 151728 1002008
rect 151728 1001988 151780 1002008
rect 151780 1001988 151782 1002008
rect 151726 1001952 151782 1001988
rect 151266 995288 151322 995344
rect 136270 995016 136326 995072
rect 140134 995016 140190 995072
rect 160650 1004964 160706 1005000
rect 160650 1004944 160652 1004964
rect 160652 1004944 160704 1004964
rect 160704 1004944 160706 1004964
rect 159454 1004828 159510 1004864
rect 159454 1004808 159456 1004828
rect 159456 1004808 159508 1004828
rect 159508 1004808 159510 1004828
rect 159822 1004692 159878 1004728
rect 159822 1004672 159824 1004692
rect 159824 1004672 159876 1004692
rect 159876 1004672 159878 1004692
rect 160282 1004708 160284 1004728
rect 160284 1004708 160336 1004728
rect 160336 1004708 160338 1004728
rect 160282 1004672 160338 1004708
rect 155774 1002108 155830 1002144
rect 155774 1002088 155776 1002108
rect 155776 1002088 155828 1002108
rect 155828 1002088 155830 1002108
rect 157430 1002108 157486 1002144
rect 157430 1002088 157432 1002108
rect 157432 1002088 157484 1002108
rect 157484 1002088 157486 1002108
rect 158258 1002124 158260 1002144
rect 158260 1002124 158312 1002144
rect 158312 1002124 158314 1002144
rect 158258 1002088 158314 1002124
rect 155774 1001952 155830 1002008
rect 156970 1001972 157026 1002008
rect 156970 1001952 156972 1001972
rect 156972 1001952 157024 1001972
rect 157024 1001952 157026 1001972
rect 158626 1001988 158628 1002008
rect 158628 1001988 158680 1002008
rect 158680 1001988 158682 1002008
rect 158626 1001952 158682 1001988
rect 162122 997328 162178 997384
rect 161110 997056 161166 997112
rect 164422 997328 164478 997384
rect 164422 997092 164424 997112
rect 164424 997092 164476 997112
rect 164476 997092 164478 997112
rect 164422 997056 164478 997092
rect 167550 997228 167552 997248
rect 167552 997228 167604 997248
rect 167604 997228 167606 997248
rect 167550 997192 167606 997228
rect 167550 997092 167552 997112
rect 167552 997092 167604 997112
rect 167604 997092 167606 997112
rect 167550 997056 167606 997092
rect 165986 995036 166042 995072
rect 165986 995016 165988 995036
rect 165988 995016 166040 995036
rect 166040 995016 166042 995036
rect 167550 995036 167606 995072
rect 167550 995016 167552 995036
rect 167552 995016 167604 995036
rect 167604 995016 167606 995036
rect 195058 1001816 195114 1001872
rect 195242 1001816 195298 1001872
rect 261022 1006868 261078 1006904
rect 261022 1006848 261024 1006868
rect 261024 1006848 261076 1006868
rect 261076 1006848 261078 1006868
rect 203522 1006596 203578 1006632
rect 203522 1006576 203524 1006596
rect 203524 1006576 203576 1006596
rect 203576 1006576 203578 1006596
rect 184662 995696 184718 995752
rect 188158 995696 188214 995752
rect 188802 995560 188858 995616
rect 195242 997192 195298 997248
rect 195242 995560 195298 995616
rect 181120 995152 181176 995208
rect 184478 995424 184534 995480
rect 187284 995288 187340 995344
rect 195058 995424 195114 995480
rect 204718 1006324 204774 1006360
rect 204718 1006304 204720 1006324
rect 204720 1006304 204772 1006324
rect 204772 1006304 204774 1006324
rect 258170 1006324 258226 1006360
rect 258170 1006304 258172 1006324
rect 258172 1006304 258224 1006324
rect 258224 1006304 258226 1006324
rect 205546 1006188 205602 1006224
rect 205546 1006168 205548 1006188
rect 205548 1006168 205600 1006188
rect 205600 1006168 205602 1006188
rect 201038 1006052 201094 1006088
rect 201038 1006032 201040 1006052
rect 201040 1006032 201092 1006052
rect 201092 1006032 201094 1006052
rect 201866 1006052 201922 1006088
rect 201866 1006032 201868 1006052
rect 201868 1006032 201920 1006052
rect 201920 1006032 201922 1006052
rect 204350 1006068 204352 1006088
rect 204352 1006068 204404 1006088
rect 204404 1006068 204406 1006088
rect 204350 1006032 204406 1006068
rect 208766 1006052 208822 1006088
rect 208766 1006032 208768 1006052
rect 208768 1006032 208820 1006052
rect 208820 1006032 208822 1006052
rect 209594 1006068 209596 1006088
rect 209596 1006068 209648 1006088
rect 209648 1006068 209650 1006088
rect 209594 1006032 209650 1006068
rect 215206 1006032 215262 1006088
rect 202326 1004692 202382 1004728
rect 202326 1004672 202328 1004692
rect 202328 1004672 202380 1004692
rect 202380 1004672 202382 1004692
rect 200210 997092 200212 997112
rect 200212 997092 200264 997112
rect 200264 997092 200266 997112
rect 200210 997056 200266 997092
rect 197358 996240 197414 996296
rect 200762 995696 200818 995752
rect 202694 1001988 202696 1002008
rect 202696 1001988 202748 1002008
rect 202748 1001988 202750 1002008
rect 202694 1001952 202750 1001988
rect 203062 1001972 203118 1002008
rect 203062 1001952 203064 1001972
rect 203064 1001952 203116 1001972
rect 203116 1001952 203118 1001972
rect 208398 1004844 208400 1004864
rect 208400 1004844 208452 1004864
rect 208452 1004844 208454 1004864
rect 208398 1004808 208454 1004844
rect 208766 1004708 208768 1004728
rect 208768 1004708 208820 1004728
rect 208820 1004708 208822 1004728
rect 208766 1004672 208822 1004708
rect 207202 1002532 207204 1002552
rect 207204 1002532 207256 1002552
rect 207256 1002532 207258 1002552
rect 207202 1002496 207258 1002532
rect 205178 1002108 205234 1002144
rect 205178 1002088 205180 1002108
rect 205180 1002088 205232 1002108
rect 205232 1002088 205234 1002108
rect 206742 1002108 206798 1002144
rect 206742 1002088 206744 1002108
rect 206744 1002088 206796 1002108
rect 206796 1002088 206798 1002108
rect 205914 1001972 205970 1002008
rect 205914 1001952 205916 1001972
rect 205916 1001952 205968 1001972
rect 205968 1001952 205970 1001972
rect 206742 1001952 206798 1002008
rect 207570 1001952 207626 1002008
rect 203522 995288 203578 995344
rect 202418 995152 202474 995208
rect 186502 995016 186558 995072
rect 191746 995016 191802 995072
rect 210422 1002244 210478 1002280
rect 210422 1002224 210424 1002244
rect 210424 1002224 210476 1002244
rect 210476 1002224 210478 1002244
rect 210054 1002124 210056 1002144
rect 210056 1002124 210108 1002144
rect 210108 1002124 210110 1002144
rect 210054 1002088 210110 1002124
rect 211250 1002108 211306 1002144
rect 211250 1002088 211252 1002108
rect 211252 1002088 211304 1002108
rect 211304 1002088 211306 1002108
rect 210882 1001952 210938 1002008
rect 211710 1001988 211712 1002008
rect 211712 1001988 211764 1002008
rect 211764 1001988 211766 1002008
rect 211710 1001952 211766 1001988
rect 212078 1001972 212134 1002008
rect 212078 1001952 212080 1001972
rect 212080 1001952 212132 1001972
rect 212132 1001952 212134 1001972
rect 213366 997328 213422 997384
rect 215758 997348 215814 997384
rect 215758 997328 215760 997348
rect 215760 997328 215812 997348
rect 215812 997328 215814 997348
rect 218886 997192 218942 997248
rect 217414 995052 217416 995072
rect 217416 995052 217468 995072
rect 217468 995052 217470 995072
rect 217414 995016 217470 995052
rect 218886 995052 218888 995072
rect 218888 995052 218940 995072
rect 218940 995052 218942 995072
rect 218886 995016 218942 995052
rect 252466 1006204 252468 1006224
rect 252468 1006204 252520 1006224
rect 252520 1006204 252522 1006224
rect 252466 1006168 252522 1006204
rect 253294 1006204 253296 1006224
rect 253296 1006204 253348 1006224
rect 253348 1006204 253350 1006224
rect 253294 1006168 253350 1006204
rect 246578 997192 246634 997248
rect 235262 995696 235318 995752
rect 243818 995696 243874 995752
rect 232226 995560 232282 995616
rect 242070 995560 242126 995616
rect 234618 995152 234674 995208
rect 236550 995424 236606 995480
rect 238712 995288 238768 995344
rect 247038 995424 247094 995480
rect 247682 996376 247738 996432
rect 249062 995560 249118 995616
rect 253662 1002652 253718 1002688
rect 253662 1002632 253664 1002652
rect 253664 1002632 253716 1002652
rect 253716 1002632 253718 1002652
rect 250442 996104 250498 996160
rect 250350 995968 250406 996024
rect 251362 995288 251418 995344
rect 254122 1001972 254178 1002008
rect 254122 1001952 254124 1001972
rect 254124 1001952 254176 1001972
rect 254176 1001952 254178 1001972
rect 254490 1001988 254492 1002008
rect 254492 1001988 254544 1002008
rect 254544 1001988 254546 1002008
rect 254490 1001952 254546 1001988
rect 256514 1006188 256570 1006224
rect 256514 1006168 256516 1006188
rect 256516 1006168 256568 1006188
rect 256568 1006168 256570 1006188
rect 255318 1006052 255374 1006088
rect 258538 1006068 258540 1006088
rect 258540 1006068 258592 1006088
rect 258592 1006068 258594 1006088
rect 255318 1006032 255320 1006052
rect 255320 1006032 255372 1006052
rect 255372 1006032 255374 1006052
rect 258538 1006032 258594 1006068
rect 258998 1006052 259054 1006088
rect 258998 1006032 259000 1006052
rect 259000 1006032 259052 1006052
rect 259052 1006032 259054 1006052
rect 262678 1006052 262734 1006088
rect 262678 1006032 262680 1006052
rect 262680 1006032 262732 1006052
rect 262732 1006032 262734 1006052
rect 263046 1006068 263048 1006088
rect 263048 1006068 263100 1006088
rect 263100 1006068 263102 1006088
rect 263046 1006032 263102 1006068
rect 254950 1002532 254952 1002552
rect 254952 1002532 255004 1002552
rect 255004 1002532 255006 1002552
rect 254950 1002496 255006 1002532
rect 255686 1002108 255742 1002144
rect 255686 1002088 255688 1002108
rect 255688 1002088 255740 1002108
rect 255740 1002088 255742 1002108
rect 256146 1002124 256148 1002144
rect 256148 1002124 256200 1002144
rect 256200 1002124 256202 1002144
rect 256146 1002088 256202 1002124
rect 256974 1001988 256976 1002008
rect 256976 1001988 257028 1002008
rect 257028 1001988 257030 1002008
rect 256974 1001952 257030 1001988
rect 245658 995016 245714 995072
rect 260194 1002244 260250 1002280
rect 260194 1002224 260196 1002244
rect 260196 1002224 260248 1002244
rect 260248 1002224 260250 1002244
rect 261482 1002108 261538 1002144
rect 261482 1002088 261484 1002108
rect 261484 1002088 261536 1002108
rect 261536 1002088 261538 1002108
rect 261850 1002124 261852 1002144
rect 261852 1002124 261904 1002144
rect 261904 1002124 261906 1002144
rect 261850 1002088 261906 1002124
rect 257802 1001972 257858 1002008
rect 257802 1001952 257804 1001972
rect 257804 1001952 257856 1001972
rect 257856 1001952 257858 1001972
rect 259826 1001972 259882 1002008
rect 259826 1001952 259828 1001972
rect 259828 1001952 259880 1001972
rect 259880 1001952 259882 1001972
rect 260654 1001988 260656 1002008
rect 260656 1001988 260708 1002008
rect 260708 1001988 260710 1002008
rect 260654 1001952 260710 1001988
rect 261850 1001952 261906 1002008
rect 263506 1001972 263562 1002008
rect 263506 1001952 263508 1001972
rect 263508 1001952 263560 1001972
rect 263560 1001952 263562 1001972
rect 267002 1001952 267058 1002008
rect 270314 997228 270316 997248
rect 270316 997228 270368 997248
rect 270368 997228 270370 997248
rect 270314 997192 270370 997228
rect 287978 995696 288034 995752
rect 291750 995696 291806 995752
rect 293590 995696 293646 995752
rect 298098 997736 298154 997792
rect 298374 997192 298430 997248
rect 291106 995560 291162 995616
rect 283470 995152 283526 995208
rect 292394 995424 292450 995480
rect 295338 995424 295394 995480
rect 290278 995288 290334 995344
rect 298742 996240 298798 996296
rect 298926 995560 298982 995616
rect 300122 995832 300178 995888
rect 299018 995424 299074 995480
rect 426346 1006884 426348 1006904
rect 426348 1006884 426400 1006904
rect 426400 1006884 426402 1006904
rect 426346 1006848 426402 1006884
rect 427174 1006868 427230 1006904
rect 427174 1006848 427176 1006868
rect 427176 1006848 427228 1006868
rect 427228 1006848 427230 1006868
rect 425150 1006748 425152 1006768
rect 425152 1006748 425204 1006768
rect 425204 1006748 425206 1006768
rect 425150 1006712 425206 1006748
rect 427542 1006732 427598 1006768
rect 427542 1006712 427544 1006732
rect 427544 1006712 427596 1006732
rect 427596 1006712 427598 1006732
rect 428002 1006612 428004 1006632
rect 428004 1006612 428056 1006632
rect 428056 1006612 428058 1006632
rect 428002 1006576 428058 1006612
rect 423494 1006476 423496 1006496
rect 423496 1006476 423548 1006496
rect 423548 1006476 423550 1006496
rect 423494 1006440 423550 1006476
rect 428370 1006440 428426 1006496
rect 308126 1006324 308182 1006360
rect 308126 1006304 308128 1006324
rect 308128 1006304 308180 1006324
rect 308180 1006304 308182 1006324
rect 310150 1006340 310152 1006360
rect 310152 1006340 310204 1006360
rect 310204 1006340 310206 1006360
rect 310150 1006304 310206 1006340
rect 423862 1006324 423918 1006360
rect 423862 1006304 423864 1006324
rect 423864 1006304 423916 1006324
rect 423916 1006304 423918 1006324
rect 425978 1006340 425980 1006360
rect 425980 1006340 426032 1006360
rect 426032 1006340 426034 1006360
rect 425978 1006304 426034 1006340
rect 306102 1006188 306158 1006224
rect 306102 1006168 306104 1006188
rect 306104 1006168 306156 1006188
rect 306156 1006168 306158 1006188
rect 357346 1006204 357348 1006224
rect 357348 1006204 357400 1006224
rect 357400 1006204 357402 1006224
rect 357346 1006168 357402 1006204
rect 361394 1006188 361450 1006224
rect 361394 1006168 361396 1006188
rect 361396 1006168 361448 1006188
rect 361448 1006168 361450 1006188
rect 304078 1006052 304134 1006088
rect 304078 1006032 304080 1006052
rect 304080 1006032 304132 1006052
rect 304132 1006032 304134 1006052
rect 304906 1006052 304962 1006088
rect 304906 1006032 304908 1006052
rect 304908 1006032 304960 1006052
rect 304960 1006032 304962 1006052
rect 305642 1006068 305644 1006088
rect 305644 1006068 305696 1006088
rect 305696 1006068 305698 1006088
rect 305642 1006032 305698 1006068
rect 306470 1006052 306526 1006088
rect 306470 1006032 306472 1006052
rect 306472 1006032 306524 1006052
rect 306524 1006032 306526 1006052
rect 310610 1006052 310666 1006088
rect 310610 1006032 310612 1006052
rect 310612 1006032 310664 1006052
rect 310664 1006032 310666 1006052
rect 314658 1006052 314714 1006088
rect 314658 1006032 314660 1006052
rect 314660 1006032 314712 1006052
rect 314712 1006032 314714 1006052
rect 354494 1006052 354550 1006088
rect 354494 1006032 354496 1006052
rect 354496 1006032 354548 1006052
rect 354548 1006032 354550 1006052
rect 355230 1006032 355286 1006088
rect 356058 1006052 356114 1006088
rect 356058 1006032 356060 1006052
rect 356060 1006032 356112 1006052
rect 356112 1006032 356114 1006052
rect 358542 1006068 358544 1006088
rect 358544 1006068 358596 1006088
rect 358596 1006068 358598 1006088
rect 358542 1006032 358598 1006068
rect 303250 997772 303252 997792
rect 303252 997772 303304 997792
rect 303304 997772 303306 997792
rect 303250 997736 303306 997772
rect 302882 997056 302938 997112
rect 300306 995288 300362 995344
rect 298282 995152 298338 995208
rect 285954 995016 286010 995072
rect 304262 995696 304318 995752
rect 306930 1004828 306986 1004864
rect 306930 1004808 306932 1004828
rect 306932 1004808 306984 1004828
rect 306984 1004808 306986 1004828
rect 305274 1001972 305330 1002008
rect 305274 1001952 305276 1001972
rect 305276 1001952 305328 1001972
rect 305328 1001952 305330 1001972
rect 307298 1004844 307300 1004864
rect 307300 1004844 307352 1004864
rect 307352 1004844 307354 1004864
rect 307298 1004808 307354 1004844
rect 307758 1004692 307814 1004728
rect 307758 1004672 307760 1004692
rect 307760 1004672 307812 1004692
rect 307812 1004672 307814 1004692
rect 308586 1004708 308588 1004728
rect 308588 1004708 308640 1004728
rect 308640 1004708 308642 1004728
rect 308586 1004672 308642 1004708
rect 310150 1001972 310206 1002008
rect 310150 1001952 310152 1001972
rect 310152 1001952 310204 1001972
rect 310204 1001952 310206 1001972
rect 311438 1001988 311440 1002008
rect 311440 1001988 311492 1002008
rect 311492 1001988 311494 1002008
rect 311438 1001952 311494 1001988
rect 312174 997908 312176 997928
rect 312176 997908 312228 997928
rect 312228 997908 312230 997928
rect 312174 997872 312230 997908
rect 313002 997772 313004 997792
rect 313004 997772 313056 997792
rect 313056 997772 313058 997792
rect 313002 997736 313058 997772
rect 313830 997892 313886 997928
rect 313830 997872 313832 997892
rect 313832 997872 313884 997892
rect 313884 997872 313886 997892
rect 315118 997772 315120 997792
rect 315120 997772 315172 997792
rect 315172 997772 315174 997792
rect 315118 997736 315174 997772
rect 318062 997736 318118 997792
rect 360566 1005372 360622 1005408
rect 360566 1005352 360568 1005372
rect 360568 1005352 360620 1005372
rect 360620 1005352 360622 1005372
rect 356518 1005252 356520 1005272
rect 356520 1005252 356572 1005272
rect 356572 1005252 356574 1005272
rect 356518 1005216 356574 1005252
rect 356518 1004572 356520 1004592
rect 356520 1004572 356572 1004592
rect 356572 1004572 356574 1004592
rect 356518 1004536 356574 1004572
rect 358082 1003892 358084 1003912
rect 358084 1003892 358136 1003912
rect 358136 1003892 358138 1003912
rect 358082 1003856 358138 1003892
rect 357346 1001952 357402 1002008
rect 358542 1001972 358598 1002008
rect 358910 1001988 358912 1002008
rect 358912 1001988 358964 1002008
rect 358964 1001988 358966 1002008
rect 358542 1001952 358544 1001972
rect 358544 1001952 358596 1001972
rect 358596 1001952 358598 1001972
rect 358910 1001952 358966 1001988
rect 359370 1001972 359426 1002008
rect 359370 1001952 359372 1001972
rect 359372 1001952 359424 1001972
rect 359424 1001952 359426 1001972
rect 360198 1001972 360254 1002008
rect 360198 1001952 360200 1001972
rect 360200 1001952 360252 1001972
rect 360252 1001952 360254 1001972
rect 361762 1004828 361818 1004864
rect 361762 1004808 361764 1004828
rect 361764 1004808 361816 1004828
rect 361816 1004808 361818 1004828
rect 363418 1004844 363420 1004864
rect 363420 1004844 363472 1004864
rect 363472 1004844 363474 1004864
rect 363418 1004808 363474 1004844
rect 362590 1004692 362646 1004728
rect 362590 1004672 362592 1004692
rect 362592 1004672 362644 1004692
rect 362644 1004672 362646 1004692
rect 364246 1004708 364248 1004728
rect 364248 1004708 364300 1004728
rect 364300 1004708 364302 1004728
rect 364246 1004672 364302 1004708
rect 361026 1001988 361028 1002008
rect 361028 1001988 361080 1002008
rect 361080 1001988 361082 1002008
rect 361026 1001952 361082 1001988
rect 360198 995288 360254 995344
rect 365074 1001988 365076 1002008
rect 365076 1001988 365128 1002008
rect 365128 1001988 365130 1002008
rect 365074 1001952 365130 1001988
rect 365442 1001972 365498 1002008
rect 365442 1001952 365444 1001972
rect 365444 1001952 365496 1001972
rect 365496 1001952 365498 1001972
rect 369122 1001952 369178 1002008
rect 366546 997328 366602 997384
rect 363602 995424 363658 995480
rect 362222 995152 362278 995208
rect 369214 997348 369270 997384
rect 369214 997328 369216 997348
rect 369216 997328 369268 997348
rect 369268 997328 369270 997348
rect 369214 995460 369216 995480
rect 369216 995460 369268 995480
rect 369268 995460 369270 995480
rect 369214 995424 369270 995460
rect 372342 998316 372344 998336
rect 372344 998316 372396 998336
rect 372396 998316 372398 998336
rect 372342 998280 372398 998316
rect 372342 997192 372398 997248
rect 372342 996956 372344 996976
rect 372344 996956 372396 996976
rect 372396 996956 372398 996976
rect 372342 996920 372398 996956
rect 372342 996240 372398 996296
rect 424690 1006188 424746 1006224
rect 424690 1006168 424692 1006188
rect 424692 1006168 424744 1006188
rect 424744 1006168 424746 1006188
rect 430026 1006204 430028 1006224
rect 430028 1006204 430080 1006224
rect 430080 1006204 430082 1006224
rect 430026 1006168 430082 1006204
rect 422666 1006052 422722 1006088
rect 422666 1006032 422668 1006052
rect 422668 1006032 422720 1006052
rect 422720 1006032 422722 1006052
rect 425518 1006068 425520 1006088
rect 425520 1006068 425572 1006088
rect 425572 1006068 425574 1006088
rect 425518 1006032 425574 1006068
rect 377402 996104 377458 996160
rect 374642 995832 374698 995888
rect 428830 1005388 428832 1005408
rect 428832 1005388 428884 1005408
rect 428884 1005388 428886 1005408
rect 428830 1005352 428886 1005388
rect 432878 1005372 432934 1005408
rect 432878 1005352 432880 1005372
rect 432880 1005352 432932 1005372
rect 432932 1005352 432934 1005372
rect 432510 1005252 432512 1005272
rect 432512 1005252 432564 1005272
rect 432564 1005252 432566 1005272
rect 432510 1005216 432566 1005252
rect 421470 1001972 421526 1002008
rect 421470 1001952 421472 1001972
rect 421472 1001952 421524 1001972
rect 421524 1001952 421526 1001972
rect 424322 1001972 424378 1002008
rect 424322 1001952 424324 1001972
rect 424324 1001952 424376 1001972
rect 424376 1001952 424378 1001972
rect 426346 1001952 426402 1002008
rect 383474 998280 383530 998336
rect 378322 995696 378378 995752
rect 383566 997736 383622 997792
rect 399942 997192 399998 997248
rect 400034 996920 400090 996976
rect 388626 995696 388682 995752
rect 389362 995696 389418 995752
rect 392398 995696 392454 995752
rect 393410 995696 393466 995752
rect 372434 995560 372490 995616
rect 391938 995560 391994 995616
rect 372342 995460 372344 995480
rect 372344 995460 372396 995480
rect 372396 995460 372398 995480
rect 372342 995424 372398 995460
rect 370778 995324 370780 995344
rect 370780 995324 370832 995344
rect 370832 995324 370834 995344
rect 370778 995288 370834 995324
rect 372342 995324 372344 995344
rect 372344 995324 372396 995344
rect 372396 995324 372398 995344
rect 372342 995288 372398 995324
rect 370778 995188 370780 995208
rect 370780 995188 370832 995208
rect 370832 995188 370834 995208
rect 370778 995152 370834 995188
rect 372342 995188 372344 995208
rect 372344 995188 372396 995208
rect 372396 995188 372398 995208
rect 372342 995152 372398 995188
rect 387798 995152 387854 995208
rect 396722 995424 396778 995480
rect 395158 995288 395214 995344
rect 388074 995016 388130 995072
rect 430854 998164 430910 998200
rect 430854 998144 430856 998164
rect 430856 998144 430908 998164
rect 430908 998144 430910 998164
rect 429658 998044 429660 998064
rect 429660 998044 429712 998064
rect 429712 998044 429714 998064
rect 429658 998008 429714 998044
rect 430854 998028 430910 998064
rect 430854 998008 430856 998028
rect 430856 998008 430908 998028
rect 430908 998008 430910 998028
rect 431682 998028 431738 998064
rect 431682 998008 431684 998028
rect 431684 998008 431736 998028
rect 431736 998008 431738 998028
rect 429198 997892 429254 997928
rect 429198 997872 429200 997892
rect 429200 997872 429252 997892
rect 429252 997872 429254 997892
rect 430394 997908 430396 997928
rect 430396 997908 430448 997928
rect 430448 997908 430450 997928
rect 430394 997872 430450 997908
rect 432050 997892 432106 997928
rect 432050 997872 432052 997892
rect 432052 997872 432104 997892
rect 432104 997872 432106 997892
rect 435362 997736 435418 997792
rect 433982 997328 434038 997384
rect 436558 997328 436614 997384
rect 439686 997228 439688 997248
rect 439688 997228 439740 997248
rect 439740 997228 439742 997248
rect 439686 997192 439742 997228
rect 439686 995324 439688 995344
rect 439688 995324 439740 995344
rect 439740 995324 439742 995344
rect 439686 995288 439742 995324
rect 443642 998280 443698 998336
rect 440882 995152 440938 995208
rect 448610 996240 448666 996296
rect 454682 996104 454738 996160
rect 451922 995424 451978 995480
rect 446310 995016 446366 995072
rect 508686 1006460 508742 1006496
rect 508686 1006440 508688 1006460
rect 508688 1006440 508740 1006460
rect 508740 1006440 508742 1006460
rect 501326 1006324 501382 1006360
rect 501326 1006304 501328 1006324
rect 501328 1006304 501380 1006324
rect 501380 1006304 501382 1006324
rect 505834 1006204 505836 1006224
rect 505836 1006204 505888 1006224
rect 505888 1006204 505890 1006224
rect 505834 1006168 505890 1006204
rect 499670 1006068 499672 1006088
rect 499672 1006068 499724 1006088
rect 499724 1006068 499726 1006088
rect 499670 1006032 499726 1006068
rect 504546 1006068 504548 1006088
rect 504548 1006068 504600 1006088
rect 504600 1006068 504602 1006088
rect 504546 1006032 504602 1006068
rect 505374 1006052 505430 1006088
rect 505374 1006032 505376 1006052
rect 505376 1006032 505428 1006052
rect 505428 1006032 505430 1006052
rect 509882 1005372 509938 1005408
rect 509882 1005352 509884 1005372
rect 509884 1005352 509936 1005372
rect 509936 1005352 509938 1005372
rect 502890 1005252 502892 1005272
rect 502892 1005252 502944 1005272
rect 502944 1005252 502946 1005272
rect 502890 1005216 502946 1005252
rect 501694 1004828 501750 1004864
rect 501694 1004808 501696 1004828
rect 501696 1004808 501748 1004828
rect 501748 1004808 501750 1004828
rect 469862 995560 469918 995616
rect 472714 998280 472770 998336
rect 488906 997192 488962 997248
rect 481546 995696 481602 995752
rect 482650 995696 482706 995752
rect 485594 995696 485650 995752
rect 483754 995560 483810 995616
rect 476946 995424 477002 995480
rect 478602 995288 478658 995344
rect 481086 995152 481142 995208
rect 487802 995016 487858 995072
rect 498474 1001952 498530 1002008
rect 500498 1004708 500500 1004728
rect 500500 1004708 500552 1004728
rect 500552 1004708 500554 1004728
rect 500498 1004672 500554 1004708
rect 500498 1004572 500500 1004592
rect 500500 1004572 500552 1004592
rect 500552 1004572 500554 1004592
rect 500498 1004536 500554 1004572
rect 501326 1004556 501382 1004592
rect 501326 1004536 501328 1004556
rect 501328 1004536 501380 1004556
rect 501380 1004536 501382 1004556
rect 502522 1002108 502578 1002144
rect 502522 1002088 502524 1002108
rect 502524 1002088 502576 1002108
rect 502576 1002088 502578 1002108
rect 502890 1001972 502946 1002008
rect 502890 1001952 502892 1001972
rect 502892 1001952 502944 1001972
rect 502944 1001952 502946 1001972
rect 503350 1001988 503352 1002008
rect 503352 1001988 503404 1002008
rect 503404 1001988 503406 1002008
rect 503350 1001952 503406 1001988
rect 500958 995152 501014 995208
rect 505006 1001972 505062 1002008
rect 505006 1001952 505008 1001972
rect 505008 1001952 505060 1001972
rect 505060 1001952 505062 1001972
rect 507030 998044 507032 998064
rect 507032 998044 507084 998064
rect 507084 998044 507086 998064
rect 507030 998008 507086 998044
rect 508226 998028 508282 998064
rect 508226 998008 508228 998028
rect 508228 998008 508280 998028
rect 508280 998008 508282 998028
rect 506202 997892 506258 997928
rect 506202 997872 506204 997892
rect 506204 997872 506256 997892
rect 506256 997872 506258 997892
rect 507858 997908 507860 997928
rect 507860 997908 507912 997928
rect 507912 997908 507914 997928
rect 507858 997872 507914 997908
rect 509054 997892 509110 997928
rect 509054 997872 509056 997892
rect 509056 997872 509108 997892
rect 509108 997872 509110 997892
rect 506570 997736 506626 997792
rect 507398 997772 507400 997792
rect 507400 997772 507452 997792
rect 507452 997772 507454 997792
rect 507398 997736 507454 997772
rect 509514 997772 509516 997792
rect 509516 997772 509568 997792
rect 509568 997772 509570 997792
rect 509514 997736 509570 997772
rect 512642 997736 512698 997792
rect 511078 995832 511134 995888
rect 551926 1006340 551928 1006360
rect 551928 1006340 551980 1006360
rect 551980 1006340 551982 1006360
rect 551926 1006304 551982 1006340
rect 553950 1006324 554006 1006360
rect 553950 1006304 553952 1006324
rect 553952 1006304 554004 1006324
rect 554004 1006304 554006 1006324
rect 555974 1006204 555976 1006224
rect 555976 1006204 556028 1006224
rect 556028 1006204 556030 1006224
rect 555974 1006168 556030 1006204
rect 557170 1006188 557226 1006224
rect 557170 1006168 557172 1006188
rect 557172 1006168 557224 1006188
rect 557224 1006168 557226 1006188
rect 517978 998416 518034 998472
rect 516690 998300 516746 998336
rect 516690 998280 516692 998300
rect 516692 998280 516744 998300
rect 516744 998280 516746 998300
rect 516690 997228 516692 997248
rect 516692 997228 516744 997248
rect 516744 997228 516746 997248
rect 516690 997192 516746 997228
rect 550270 1006068 550272 1006088
rect 550272 1006068 550324 1006088
rect 550324 1006068 550326 1006088
rect 516690 995732 516692 995752
rect 516692 995732 516744 995752
rect 516744 995732 516746 995752
rect 516690 995696 516746 995732
rect 516690 995596 516692 995616
rect 516692 995596 516744 995616
rect 516744 995596 516746 995616
rect 516690 995560 516746 995596
rect 516690 995460 516692 995480
rect 516692 995460 516744 995480
rect 516744 995460 516746 995480
rect 516690 995424 516746 995460
rect 515218 995324 515220 995344
rect 515220 995324 515272 995344
rect 515272 995324 515274 995344
rect 515218 995288 515274 995324
rect 516690 995324 516692 995344
rect 516692 995324 516744 995344
rect 516744 995324 516746 995344
rect 516690 995288 516746 995324
rect 515218 995172 515274 995208
rect 515218 995152 515220 995172
rect 515220 995152 515272 995172
rect 515272 995152 515274 995172
rect 516690 995172 516746 995208
rect 516690 995152 516692 995172
rect 516692 995152 516744 995172
rect 516744 995152 516746 995172
rect 523958 998416 524014 998472
rect 524050 998280 524106 998336
rect 523958 996376 524014 996432
rect 540886 997192 540942 997248
rect 525338 995696 525394 995752
rect 526166 995696 526222 995752
rect 529018 995560 529074 995616
rect 532146 995288 532202 995344
rect 532606 995152 532662 995208
rect 538954 995424 539010 995480
rect 550270 1006032 550326 1006068
rect 551098 1006068 551100 1006088
rect 551100 1006068 551152 1006088
rect 551152 1006068 551154 1006088
rect 551098 1006032 551154 1006068
rect 553122 1006052 553178 1006088
rect 556802 1006068 556804 1006088
rect 556804 1006068 556856 1006088
rect 556856 1006068 556858 1006088
rect 553122 1006032 553124 1006052
rect 553124 1006032 553176 1006052
rect 553176 1006032 553178 1006052
rect 556802 1006032 556858 1006068
rect 556342 1004708 556344 1004728
rect 556344 1004708 556396 1004728
rect 556396 1004708 556398 1004728
rect 556342 1004672 556398 1004708
rect 552754 1002652 552810 1002688
rect 552754 1002632 552756 1002652
rect 552756 1002632 552808 1002652
rect 552808 1002632 552810 1002652
rect 552294 1002532 552296 1002552
rect 552296 1002532 552348 1002552
rect 552348 1002532 552350 1002552
rect 552294 1002496 552350 1002532
rect 554778 1002108 554834 1002144
rect 554778 1002088 554780 1002108
rect 554780 1002088 554832 1002108
rect 554832 1002088 554834 1002108
rect 553122 1001972 553178 1002008
rect 553122 1001952 553124 1001972
rect 553124 1001952 553176 1001972
rect 553176 1001952 553178 1001972
rect 553950 1001988 553952 1002008
rect 553952 1001988 554004 1002008
rect 554004 1001988 554006 1002008
rect 553950 1001952 554006 1001988
rect 554318 1001952 554374 1002008
rect 555146 1001952 555202 1002008
rect 557630 1004692 557686 1004728
rect 557630 1004672 557632 1004692
rect 557632 1004672 557684 1004692
rect 557684 1004672 557686 1004692
rect 559194 1002260 559196 1002280
rect 559196 1002260 559248 1002280
rect 559248 1002260 559250 1002280
rect 559194 1002224 559250 1002260
rect 558458 1002124 558460 1002144
rect 558460 1002124 558512 1002144
rect 558512 1002124 558514 1002144
rect 558458 1002088 558514 1002124
rect 557998 1001988 558000 1002008
rect 558000 1001988 558052 1002008
rect 558052 1001988 558054 1002008
rect 557998 1001952 558054 1001988
rect 558826 1001972 558882 1002008
rect 558826 1001952 558828 1001972
rect 558828 1001952 558880 1001972
rect 558880 1001952 558882 1001972
rect 559654 1002244 559710 1002280
rect 559654 1002224 559656 1002244
rect 559656 1002224 559708 1002244
rect 559708 1002224 559710 1002244
rect 560022 1002108 560078 1002144
rect 561310 1002124 561312 1002144
rect 561312 1002124 561364 1002144
rect 561364 1002124 561366 1002144
rect 560022 1002088 560024 1002108
rect 560024 1002088 560076 1002108
rect 560076 1002088 560078 1002108
rect 560482 1001972 560538 1002008
rect 560482 1001952 560484 1001972
rect 560484 1001952 560536 1001972
rect 560536 1001952 560538 1001972
rect 560850 1001988 560852 1002008
rect 560852 1001988 560904 1002008
rect 560904 1001988 560906 1002008
rect 560850 1001952 560906 1001988
rect 561310 1002088 561366 1002124
rect 561678 997328 561734 997384
rect 561678 996920 561734 996976
rect 564346 1006032 564402 1006088
rect 564990 997328 565046 997384
rect 564990 996940 565046 996976
rect 564990 996920 564992 996940
rect 564992 996920 565044 996940
rect 565044 996920 565046 996940
rect 568118 997228 568120 997248
rect 568120 997228 568172 997248
rect 568172 997228 568174 997248
rect 568118 997192 568174 997228
rect 568118 996784 568174 996840
rect 575202 997212 575258 997248
rect 575202 997192 575204 997212
rect 575204 997192 575256 997212
rect 575256 997192 575258 997212
rect 575478 996820 575480 996840
rect 575480 996820 575532 996840
rect 575532 996820 575534 996840
rect 575478 996784 575534 996820
rect 580906 997212 580962 997248
rect 580906 997192 580908 997212
rect 580908 997192 580960 997212
rect 580960 997192 580962 997212
rect 585138 997228 585140 997248
rect 585140 997228 585192 997248
rect 585192 997228 585194 997248
rect 585138 997192 585194 997228
rect 590934 997228 590936 997248
rect 590936 997228 590988 997248
rect 590988 997228 590990 997248
rect 590934 997192 590990 997228
rect 580722 996820 580724 996840
rect 580724 996820 580776 996840
rect 580776 996820 580778 996840
rect 580722 996784 580778 996820
rect 585506 996820 585508 996840
rect 585508 996820 585560 996840
rect 585560 996820 585562 996840
rect 585506 996784 585562 996820
rect 590566 996820 590568 996840
rect 590568 996820 590620 996840
rect 590620 996820 590622 996840
rect 590566 996784 590622 996820
rect 605930 996240 605986 996296
rect 623686 996648 623742 996704
rect 625894 996648 625950 996704
rect 633990 995696 634046 995752
rect 640798 995696 640854 995752
rect 635186 995560 635242 995616
rect 622398 995016 622454 995072
rect 629666 995016 629722 995072
rect 638958 994880 639014 994936
rect 640798 994880 640854 994936
rect 62118 975976 62174 976032
rect 62118 962920 62174 962976
rect 62118 949864 62174 949920
rect 55862 939800 55918 939856
rect 62118 936980 62120 937000
rect 62120 936980 62172 937000
rect 62172 936980 62174 937000
rect 62118 936944 62174 936980
rect 44178 934496 44234 934552
rect 42890 934088 42946 934144
rect 42798 933680 42854 933736
rect 41694 816584 41750 816640
rect 41878 815632 41934 815688
rect 41970 814816 42026 814872
rect 41786 814000 41842 814056
rect 40682 813184 40738 813240
rect 33782 812368 33838 812424
rect 33046 810328 33102 810384
rect 32402 809104 32458 809160
rect 33046 802440 33102 802496
rect 34426 810736 34482 810792
rect 35162 808696 35218 808752
rect 34426 802576 34482 802632
rect 39854 807288 39910 807328
rect 39854 807272 39856 807288
rect 39856 807272 39908 807288
rect 39908 807272 39910 807288
rect 42154 812776 42210 812832
rect 41786 811572 41842 811608
rect 41786 811552 41788 811572
rect 41788 811552 41840 811572
rect 41840 811552 41842 811572
rect 40682 801624 40738 801680
rect 33782 800944 33838 801000
rect 42062 809512 42118 809568
rect 41786 806248 41842 806304
rect 42338 811144 42394 811200
rect 42798 809920 42854 809976
rect 42430 796728 42486 796784
rect 42338 791968 42394 792024
rect 43442 806248 43498 806304
rect 42706 791832 42762 791888
rect 42706 788160 42762 788216
rect 42430 788024 42486 788080
rect 41786 786120 41842 786176
rect 35806 774288 35862 774344
rect 42798 771976 42854 772032
rect 33782 769392 33838 769448
rect 32402 768576 32458 768632
rect 31022 767760 31078 767816
rect 30378 764088 30434 764144
rect 30378 763272 30434 763328
rect 32494 766536 32550 766592
rect 40682 768984 40738 769040
rect 35162 767352 35218 767408
rect 35162 758240 35218 758296
rect 41510 762864 41566 762920
rect 40682 757696 40738 757752
rect 42706 756472 42762 756528
rect 41786 753072 41842 753128
rect 41786 751712 41842 751768
rect 41786 750352 41842 750408
rect 42706 749264 42762 749320
rect 42614 746544 42670 746600
rect 41786 742328 41842 742384
rect 31482 731060 31538 731096
rect 31482 731040 31484 731060
rect 31484 731040 31536 731060
rect 31536 731040 31538 731060
rect 31666 731040 31722 731096
rect 31574 730632 31630 730688
rect 31390 730224 31446 730280
rect 42890 767080 42946 767136
rect 42982 765856 43038 765912
rect 42798 729272 42854 729328
rect 42798 727232 42854 727288
rect 31022 726552 31078 726608
rect 40682 726144 40738 726200
rect 33782 725328 33838 725384
rect 34426 723288 34482 723344
rect 33782 715536 33838 715592
rect 31022 715400 31078 715456
rect 42154 725192 42210 725248
rect 40866 724512 40922 724568
rect 40774 723288 40830 723344
rect 42062 723968 42118 724024
rect 41510 720840 41566 720896
rect 41510 719652 41512 719672
rect 41512 719652 41564 719672
rect 41564 719652 41566 719672
rect 41510 719616 41566 719652
rect 40774 714040 40830 714096
rect 42062 713768 42118 713824
rect 42430 713224 42486 713280
rect 42522 712272 42578 712328
rect 42154 711728 42210 711784
rect 42522 710776 42578 710832
rect 41786 709824 41842 709880
rect 42522 708464 42578 708520
rect 42522 706560 42578 706616
rect 42246 704928 42302 704984
rect 42430 702888 42486 702944
rect 41786 699352 41842 699408
rect 35622 688336 35678 688392
rect 35806 687656 35862 687712
rect 35714 687248 35770 687304
rect 42890 724376 42946 724432
rect 42982 722336 43038 722392
rect 42798 684392 42854 684448
rect 42798 683984 42854 684040
rect 39302 683576 39358 683632
rect 32402 682760 32458 682816
rect 31022 681536 31078 681592
rect 30470 676864 30526 676866
rect 30470 676812 30472 676864
rect 30472 676812 30524 676864
rect 30524 676812 30526 676864
rect 30470 676810 30526 676812
rect 35162 680312 35218 680368
rect 32402 671336 32458 671392
rect 41694 683052 41750 683088
rect 41694 683032 41696 683052
rect 41696 683032 41748 683052
rect 41748 683032 41750 683052
rect 39302 670928 39358 670984
rect 41694 681828 41750 681864
rect 41694 681808 41696 681828
rect 41696 681808 41748 681828
rect 41748 681808 41750 681828
rect 41970 680720 42026 680776
rect 42062 670656 42118 670712
rect 42430 670112 42486 670168
rect 42706 669432 42762 669488
rect 42062 668480 42118 668536
rect 41786 665352 41842 665408
rect 41786 664536 41842 664592
rect 42062 663312 42118 663368
rect 42706 661272 42762 661328
rect 42154 660456 42210 660512
rect 42522 660320 42578 660376
rect 42338 658280 42394 658336
rect 35622 644680 35678 644736
rect 35806 644680 35862 644736
rect 42890 679088 42946 679144
rect 42982 678680 43038 678736
rect 42798 641416 42854 641472
rect 33782 639784 33838 639840
rect 32402 638152 32458 638208
rect 40682 639376 40738 639432
rect 35162 637744 35218 637800
rect 35162 629856 35218 629912
rect 40866 638968 40922 639024
rect 40682 629040 40738 629096
rect 42798 638560 42854 638616
rect 41050 637336 41106 637392
rect 41050 629176 41106 629232
rect 40866 628904 40922 628960
rect 42522 625096 42578 625152
rect 42522 623736 42578 623792
rect 42890 635704 42946 635760
rect 41786 621424 41842 621480
rect 43074 635296 43130 635352
rect 42246 618976 42302 619032
rect 42522 616800 42578 616856
rect 42246 615984 42302 616040
rect 41878 614080 41934 614136
rect 41786 612720 41842 612776
rect 35806 601840 35862 601896
rect 35806 601432 35862 601488
rect 35806 601024 35862 601080
rect 35714 600616 35770 600672
rect 42798 597624 42854 597680
rect 39302 596944 39358 597000
rect 33782 594904 33838 594960
rect 32402 593272 32458 593328
rect 40682 596536 40738 596592
rect 39302 585112 39358 585168
rect 40774 595720 40830 595776
rect 42062 593952 42118 594008
rect 41510 591232 41566 591288
rect 41510 590008 41566 590064
rect 41786 584160 41842 584216
rect 41970 584160 42026 584216
rect 42430 583616 42486 583672
rect 41970 582120 42026 582176
rect 41786 580216 41842 580272
rect 41786 578992 41842 579048
rect 41786 577496 41842 577552
rect 42706 576816 42762 576872
rect 42338 575864 42394 575920
rect 42338 573688 42394 573744
rect 41970 572736 42026 572792
rect 42706 571512 42762 571568
rect 42154 570424 42210 570480
rect 35622 558320 35678 558376
rect 35806 558320 35862 558376
rect 35714 557912 35770 557968
rect 42890 594360 42946 594416
rect 42982 592728 43038 592784
rect 42982 556824 43038 556880
rect 42890 556008 42946 556064
rect 42798 554784 42854 554840
rect 40866 553832 40922 553888
rect 40682 553424 40738 553480
rect 32402 552608 32458 552664
rect 31022 551792 31078 551848
rect 31666 548120 31722 548176
rect 35806 546896 35862 546952
rect 32402 542816 32458 542872
rect 40774 552200 40830 552256
rect 40958 553016 41014 553072
rect 40866 545128 40922 545184
rect 40958 542952 41014 543008
rect 40774 542272 40830 542328
rect 42614 535880 42670 535936
rect 41786 534520 41842 534576
rect 42614 533840 42670 533896
rect 42338 532616 42394 532672
rect 41786 530712 41842 530768
rect 42338 529488 42394 529544
rect 42614 529352 42670 529408
rect 41786 430480 41842 430536
rect 41786 430108 41788 430128
rect 41788 430108 41840 430128
rect 41840 430108 41842 430128
rect 41786 430072 41842 430108
rect 42982 551112 43038 551168
rect 43074 549888 43130 549944
rect 43350 430888 43406 430944
rect 42890 429664 42946 429720
rect 42798 428848 42854 428904
rect 43166 427624 43222 427680
rect 42890 426808 42946 426864
rect 41786 426400 41842 426456
rect 35162 425176 35218 425232
rect 32402 424360 32458 424416
rect 31022 422320 31078 422376
rect 40774 425012 40830 425068
rect 41326 425012 41382 425068
rect 42798 421912 42854 421968
rect 41786 419484 41842 419520
rect 41786 419464 41788 419484
rect 41788 419464 41840 419484
rect 41840 419464 41842 419484
rect 41326 417968 41382 418024
rect 35162 414568 35218 414624
rect 42154 411168 42210 411224
rect 41786 409400 41842 409456
rect 41786 406272 41842 406328
rect 41786 402464 41842 402520
rect 41970 401784 42026 401840
rect 41786 400016 41842 400072
rect 41786 399608 41842 399664
rect 41786 398792 41842 398848
rect 35622 387096 35678 387152
rect 35806 387504 35862 387560
rect 35806 387096 35862 387152
rect 35714 386688 35770 386744
rect 43074 421096 43130 421152
rect 43166 384784 43222 384840
rect 42890 383968 42946 384024
rect 42798 383560 42854 383616
rect 40866 382608 40922 382664
rect 37922 381384 37978 381440
rect 31022 380976 31078 381032
rect 33782 378120 33838 378176
rect 35806 377304 35862 377360
rect 33782 371864 33838 371920
rect 40682 379344 40738 379400
rect 37922 371320 37978 371376
rect 41510 376080 41566 376136
rect 41786 370232 41842 370288
rect 41878 366288 41934 366344
rect 41970 363704 42026 363760
rect 41786 362888 41842 362944
rect 41786 360032 41842 360088
rect 41786 358672 41842 358728
rect 41786 356904 41842 356960
rect 41786 355680 41842 355736
rect 35622 344256 35678 344312
rect 35806 344292 35808 344312
rect 35808 344292 35860 344312
rect 35860 344292 35862 344312
rect 35806 344256 35862 344292
rect 35714 343848 35770 343904
rect 42890 380296 42946 380352
rect 42982 378664 43038 378720
rect 43074 377848 43130 377904
rect 42798 340856 42854 340912
rect 42798 340448 42854 340504
rect 40866 339360 40922 339416
rect 40682 338136 40738 338192
rect 30378 334056 30434 334112
rect 30378 333260 30434 333296
rect 30378 333240 30380 333260
rect 30380 333240 30432 333260
rect 30432 333240 30434 333260
rect 40866 334056 40922 334112
rect 40682 328344 40738 328400
rect 41786 324808 41842 324864
rect 41786 321136 41842 321192
rect 41970 319912 42026 319968
rect 41786 317328 41842 317384
rect 41786 315832 41842 315888
rect 41786 315424 41842 315480
rect 41878 313792 41934 313848
rect 41786 313112 41842 313168
rect 41786 312296 41842 312352
rect 42062 301280 42118 301336
rect 41970 300872 42026 300928
rect 43074 338000 43130 338056
rect 42982 336368 43038 336424
rect 42890 334736 42946 334792
rect 43074 298832 43130 298888
rect 42798 297608 42854 297664
rect 33782 296384 33838 296440
rect 42430 294752 42486 294808
rect 33782 284824 33838 284880
rect 42982 293120 43038 293176
rect 42890 291896 42946 291952
rect 41786 281424 41842 281480
rect 42706 278704 42762 278760
rect 41786 277344 41842 277400
rect 41786 276664 41842 276720
rect 41786 272312 41842 272368
rect 41970 270408 42026 270464
rect 41786 269728 41842 269784
rect 41786 269048 41842 269104
rect 35806 258304 35862 258360
rect 31666 257896 31722 257952
rect 31666 257488 31722 257544
rect 31574 257080 31630 257136
rect 42890 256400 42946 256456
rect 31022 251776 31078 251832
rect 42706 251504 42762 251560
rect 39946 250552 40002 250608
rect 35806 246472 35862 246528
rect 31022 243480 31078 243536
rect 42798 245792 42854 245848
rect 40038 244568 40094 244624
rect 40038 244160 40094 244216
rect 40498 243480 40554 243536
rect 39946 241576 40002 241632
rect 40498 240896 40554 240952
rect 42706 245656 42762 245712
rect 42706 238856 42762 238912
rect 41878 238448 41934 238504
rect 42798 238040 42854 238096
rect 42706 237904 42762 237960
rect 41786 236680 41842 236736
rect 41786 234776 41842 234832
rect 41786 233280 41842 233336
rect 41786 230424 41842 230480
rect 42154 229880 42210 229936
rect 41786 228928 41842 228984
rect 42062 227296 42118 227352
rect 41786 226072 41842 226128
rect 35622 214648 35678 214704
rect 35806 214648 35862 214704
rect 35714 214240 35770 214296
rect 31206 210160 31262 210216
rect 31022 209752 31078 209808
rect 31022 199416 31078 199472
rect 39302 208528 39358 208584
rect 35806 203224 35862 203280
rect 31206 199280 31262 199336
rect 44270 815224 44326 815280
rect 44178 813592 44234 813648
rect 43626 773608 43682 773664
rect 44362 808288 44418 808344
rect 44730 772792 44786 772848
rect 44270 772384 44326 772440
rect 44178 770752 44234 770808
rect 44638 770344 44694 770400
rect 44362 769936 44418 769992
rect 44454 768304 44510 768360
rect 44546 765448 44602 765504
rect 44178 728864 44234 728920
rect 44638 727640 44694 727696
rect 44546 722744 44602 722800
rect 44362 721928 44418 721984
rect 44270 686432 44326 686488
rect 44178 686024 44234 686080
rect 44178 685616 44234 685672
rect 44362 681128 44418 681184
rect 44454 679904 44510 679960
rect 44270 643728 44326 643784
rect 44362 643184 44418 643240
rect 44178 643048 44234 643104
rect 44178 642232 44234 642288
rect 44086 599800 44142 599856
rect 44270 640736 44326 640792
rect 44178 599664 44234 599720
rect 44454 636928 44510 636984
rect 44546 599256 44602 599312
rect 44270 598032 44326 598088
rect 44362 595584 44418 595640
rect 44454 593136 44510 593192
rect 44178 557232 44234 557288
rect 44546 556416 44602 556472
rect 44178 555192 44234 555248
rect 44638 554376 44694 554432
rect 44362 551520 44418 551576
rect 44546 550296 44602 550352
rect 44454 548664 44510 548720
rect 44362 429256 44418 429312
rect 44270 428440 44326 428496
rect 44178 428032 44234 428088
rect 44638 427216 44694 427272
rect 44362 423136 44418 423192
rect 44454 421504 44510 421560
rect 44270 386008 44326 386064
rect 44178 385600 44234 385656
rect 44178 384376 44234 384432
rect 44638 385192 44694 385248
rect 44454 380704 44510 380760
rect 44546 379072 44602 379128
rect 44270 343304 44326 343360
rect 44362 342896 44418 342952
rect 44270 342080 44326 342136
rect 44178 341672 44234 341728
rect 43626 300464 43682 300520
rect 43074 255992 43130 256048
rect 43074 255584 43130 255640
rect 42982 250280 43038 250336
rect 42890 213696 42946 213752
rect 43166 241576 43222 241632
rect 44638 342488 44694 342544
rect 44362 341264 44418 341320
rect 44270 300056 44326 300112
rect 44178 299240 44234 299296
rect 44454 336776 44510 336832
rect 44546 335144 44602 335200
rect 44730 299648 44786 299704
rect 44362 298424 44418 298480
rect 44270 298016 44326 298072
rect 44178 291488 44234 291544
rect 43994 291080 44050 291136
rect 43810 290672 43866 290728
rect 44638 297200 44694 297256
rect 44454 293528 44510 293584
rect 44546 292304 44602 292360
rect 44270 255176 44326 255232
rect 44546 254768 44602 254824
rect 44270 253952 44326 254008
rect 43074 212880 43130 212936
rect 42798 212472 42854 212528
rect 41786 211656 41842 211712
rect 44362 251096 44418 251152
rect 44454 248648 44510 248704
rect 45006 289856 45062 289912
rect 44638 254360 44694 254416
rect 44546 248240 44602 248296
rect 62118 923752 62174 923808
rect 62118 910696 62174 910752
rect 50342 773880 50398 773936
rect 62118 897776 62174 897832
rect 62118 884720 62174 884776
rect 62118 871664 62174 871720
rect 62118 858608 62174 858664
rect 62118 845552 62174 845608
rect 62118 832496 62174 832552
rect 62118 819440 62174 819496
rect 54482 816856 54538 816912
rect 62118 806520 62174 806576
rect 62118 793600 62174 793656
rect 62118 780408 62174 780464
rect 62118 767372 62174 767408
rect 62118 767352 62120 767372
rect 62120 767352 62172 767372
rect 62172 767352 62174 767372
rect 62118 754296 62174 754352
rect 62118 741240 62174 741296
rect 62118 728184 62174 728240
rect 62118 715264 62174 715320
rect 62762 702208 62818 702264
rect 62118 689152 62174 689208
rect 62118 676096 62174 676152
rect 62118 663040 62174 663096
rect 62118 650020 62120 650040
rect 62120 650020 62172 650040
rect 62172 650020 62174 650040
rect 53102 633392 53158 633448
rect 46570 213288 46626 213344
rect 44638 212064 44694 212120
rect 44270 211248 44326 211304
rect 41326 210976 41382 211032
rect 42798 209208 42854 209264
rect 40866 204856 40922 204912
rect 40682 204448 40738 204504
rect 39302 197648 39358 197704
rect 41878 197104 41934 197160
rect 41786 195200 41842 195256
rect 41786 190168 41842 190224
rect 41786 187312 41842 187368
rect 44178 207984 44234 208040
rect 42890 207576 42946 207632
rect 42982 206352 43038 206408
rect 43074 205536 43130 205592
rect 41786 184048 41842 184104
rect 44454 206760 44510 206816
rect 44270 205944 44326 206000
rect 44362 205128 44418 205184
rect 41786 182960 41842 183016
rect 62118 649984 62174 650020
rect 62762 643456 62818 643512
rect 62118 637064 62174 637120
rect 62118 624008 62174 624064
rect 62118 610952 62174 611008
rect 62118 597896 62174 597952
rect 62118 584840 62174 584896
rect 62118 571784 62174 571840
rect 62118 558728 62174 558784
rect 53102 218320 53158 218376
rect 55034 222808 55090 222864
rect 62762 545808 62818 545864
rect 62118 532772 62174 532808
rect 62118 532752 62120 532772
rect 62120 532752 62172 532772
rect 62172 532752 62174 532772
rect 62118 519696 62174 519752
rect 62118 506640 62174 506696
rect 62118 493584 62174 493640
rect 62118 480528 62174 480584
rect 62118 467472 62174 467528
rect 62118 454552 62174 454608
rect 62118 441496 62174 441552
rect 62118 428440 62174 428496
rect 62118 415420 62120 415440
rect 62120 415420 62172 415440
rect 62172 415420 62174 415440
rect 62118 415384 62174 415420
rect 62118 402328 62174 402384
rect 62118 389272 62174 389328
rect 62118 376216 62174 376272
rect 62118 363296 62174 363352
rect 62118 350240 62174 350296
rect 62118 337184 62174 337240
rect 62118 324128 62174 324184
rect 62118 311072 62174 311128
rect 62118 298172 62174 298208
rect 62118 298152 62120 298172
rect 62120 298152 62172 298172
rect 62172 298152 62174 298172
rect 62118 285096 62174 285152
rect 350262 270136 350318 270192
rect 350354 268912 350410 268968
rect 357990 267416 358046 267472
rect 365994 267280 366050 267336
rect 368386 275440 368442 275496
rect 368202 268776 368258 268832
rect 371146 275304 371202 275360
rect 373906 275168 373962 275224
rect 379242 271360 379298 271416
rect 380714 267008 380770 267064
rect 382094 271224 382150 271280
rect 383290 271088 383346 271144
rect 383382 270000 383438 270056
rect 386234 273808 386290 273864
rect 388258 269864 388314 269920
rect 388442 267008 388498 267064
rect 389638 265920 389694 265976
rect 391386 266328 391442 266384
rect 392582 266328 392638 266384
rect 392306 265784 392362 265840
rect 397642 267688 397698 267744
rect 398470 268640 398526 268696
rect 401598 269728 401654 269784
rect 402518 268504 402574 268560
rect 404266 272720 404322 272776
rect 403438 267552 403494 267608
rect 405186 268368 405242 268424
rect 406934 272584 406990 272640
rect 406566 265648 406622 265704
rect 407394 266328 407450 266384
rect 408314 272448 408370 272504
rect 409234 265512 409290 265568
rect 411074 273944 411130 274000
rect 410430 266328 410486 266384
rect 411902 267688 411958 267744
rect 411442 267144 411498 267200
rect 411902 267008 411958 267064
rect 419538 273944 419594 274000
rect 433338 268912 433394 268968
rect 469310 267552 469366 267608
rect 484398 270136 484454 270192
rect 493322 267416 493378 267472
rect 518990 267280 519046 267336
rect 530490 275440 530546 275496
rect 537574 275304 537630 275360
rect 532698 268776 532754 268832
rect 544658 275168 544714 275224
rect 561218 271360 561274 271416
rect 568302 271224 568358 271280
rect 571798 271088 571854 271144
rect 572718 270000 572774 270056
rect 580078 273808 580134 273864
rect 585138 269864 585194 269920
rect 589278 265920 589334 265976
rect 596178 265784 596234 265840
rect 396998 264152 397054 264208
rect 401230 264172 401286 264208
rect 612738 268640 612794 268696
rect 401230 264152 401232 264172
rect 401232 264152 401284 264172
rect 401284 264152 401286 264172
rect 618258 269728 618314 269784
rect 623778 268504 623834 268560
rect 628562 272720 628618 272776
rect 630678 268368 630734 268424
rect 635646 272584 635702 272640
rect 639234 272448 639290 272504
rect 633438 265648 633494 265704
rect 647238 267144 647294 267200
rect 640522 265512 640578 265568
rect 415306 262268 415362 262304
rect 415306 262248 415308 262268
rect 415308 262248 415360 262268
rect 415360 262248 415362 262268
rect 414202 259120 414258 259176
rect 189078 258576 189134 258632
rect 415306 255856 415362 255912
rect 414386 252728 414442 252784
rect 414202 249464 414258 249520
rect 85026 247288 85082 247344
rect 84842 247152 84898 247208
rect 66902 229880 66958 229936
rect 58622 229744 58678 229800
rect 56874 221448 56930 221504
rect 59266 226888 59322 226944
rect 58714 222944 58770 223000
rect 62762 227024 62818 227080
rect 62026 224168 62082 224224
rect 190366 247968 190422 248024
rect 69478 224304 69534 224360
rect 66994 221584 67050 221640
rect 67546 220088 67602 220144
rect 70214 221720 70270 221776
rect 72974 227160 73030 227216
rect 72054 224440 72110 224496
rect 73710 221856 73766 221912
rect 74446 220224 74502 220280
rect 78494 224576 78550 224632
rect 90546 228384 90602 228440
rect 86866 228248 86922 228304
rect 89534 225528 89590 225584
rect 93030 225664 93086 225720
rect 92294 223080 92350 223136
rect 99010 223216 99066 223272
rect 189078 237396 189080 237416
rect 189080 237396 189132 237416
rect 189132 237396 189134 237416
rect 189078 237360 189134 237396
rect 415306 246336 415362 246392
rect 414386 243072 414442 243128
rect 414294 239944 414350 240000
rect 414202 233552 414258 233608
rect 414938 236680 414994 236736
rect 192390 222808 192446 222864
rect 194046 222944 194102 223000
rect 193402 221448 193458 221504
rect 194782 229744 194838 229800
rect 196162 229880 196218 229936
rect 195794 226888 195850 226944
rect 195426 224168 195482 224224
rect 196622 230288 196678 230344
rect 197266 227024 197322 227080
rect 197726 221584 197782 221640
rect 196622 220088 196678 220144
rect 199014 230288 199070 230344
rect 199750 224440 199806 224496
rect 200118 224304 200174 224360
rect 199106 221720 199162 221776
rect 201498 227160 201554 227216
rect 200578 221856 200634 221912
rect 202602 224576 202658 224632
rect 201590 220224 201646 220280
rect 206558 228248 206614 228304
rect 207938 228384 207994 228440
rect 208030 223080 208086 223136
rect 208674 225528 208730 225584
rect 210054 225664 210110 225720
rect 211158 223216 211214 223272
rect 375838 230016 375894 230072
rect 376942 230288 376998 230344
rect 377310 230152 377366 230208
rect 378690 229880 378746 229936
rect 377678 224576 377734 224632
rect 376206 223352 376262 223408
rect 379058 223216 379114 223272
rect 380162 229744 380218 229800
rect 380530 227296 380586 227352
rect 381910 224440 381966 224496
rect 383014 227160 383070 227216
rect 382186 220360 382242 220416
rect 381910 220224 381966 220280
rect 384026 224304 384082 224360
rect 384854 220088 384910 220144
rect 387246 228656 387302 228712
rect 388350 227024 388406 227080
rect 389178 220496 389234 220552
rect 389362 223080 389418 223136
rect 390834 225936 390890 225992
rect 390466 222944 390522 223000
rect 394054 225800 394110 225856
rect 392858 221720 392914 221776
rect 396446 225664 396502 225720
rect 397182 221584 397238 221640
rect 399390 228520 399446 228576
rect 400494 225528 400550 225584
rect 402610 228384 402666 228440
rect 400954 221856 401010 221912
rect 405002 221448 405058 221504
rect 407946 226888 408002 226944
rect 409602 224168 409658 224224
rect 411166 228248 411222 228304
rect 410982 222808 411038 222864
rect 428646 230288 428702 230344
rect 478142 230152 478198 230208
rect 486422 230016 486478 230072
rect 493322 229880 493378 229936
rect 496082 229744 496138 229800
rect 487802 223352 487858 223408
rect 490194 224576 490250 224632
rect 489090 216824 489146 216880
rect 494058 223216 494114 223272
rect 495622 220496 495678 220552
rect 496910 227296 496966 227352
rect 502522 227160 502578 227216
rect 499578 224440 499634 224496
rect 498658 220360 498714 220416
rect 499670 220224 499726 220280
rect 505374 224304 505430 224360
rect 507214 220088 507270 220144
rect 507214 219408 507270 219464
rect 513378 228656 513434 228712
rect 515494 227024 515550 227080
rect 521658 225936 521714 225992
rect 518162 223080 518218 223136
rect 520462 222944 520518 223000
rect 495990 216688 496046 216744
rect 525890 221720 525946 221776
rect 528926 225800 528982 225856
rect 528098 221856 528154 221912
rect 534078 225664 534134 225720
rect 536010 221584 536066 221640
rect 541530 228520 541586 228576
rect 544014 225528 544070 225584
rect 549258 228384 549314 228440
rect 546682 221448 546738 221504
rect 561678 226888 561734 226944
rect 556710 224168 556766 224224
rect 564438 228248 564494 228304
rect 569314 222808 569370 222864
rect 578882 216144 578938 216200
rect 578422 211656 578478 211712
rect 578514 210160 578570 210216
rect 579066 214648 579122 214704
rect 578974 213152 579030 213208
rect 579526 208664 579582 208720
rect 578790 207168 578846 207224
rect 579434 205672 579490 205728
rect 578882 204176 578938 204232
rect 579250 202680 579306 202736
rect 578238 201184 578294 201240
rect 578422 199688 578478 199744
rect 579066 198192 579122 198248
rect 579526 196696 579582 196752
rect 579526 195236 579528 195256
rect 579528 195236 579580 195256
rect 579580 195236 579582 195256
rect 579526 195200 579582 195236
rect 579526 193568 579582 193624
rect 579526 192072 579582 192128
rect 579250 190576 579306 190632
rect 578238 189080 578294 189136
rect 579250 187584 579306 187640
rect 578790 184592 578846 184648
rect 578238 177112 578294 177168
rect 578330 175616 578386 175672
rect 579066 181600 579122 181656
rect 578974 180104 579030 180160
rect 578422 174120 578478 174176
rect 579526 186088 579582 186144
rect 579342 183096 579398 183152
rect 579250 178608 579306 178664
rect 578790 172624 578846 172680
rect 578698 171128 578754 171184
rect 578698 166504 578754 166560
rect 578238 164328 578294 164384
rect 579250 168000 579306 168056
rect 579158 162016 579214 162072
rect 579434 169496 579490 169552
rect 579526 163512 579582 163568
rect 579342 160520 579398 160576
rect 579066 159024 579122 159080
rect 578974 157528 579030 157584
rect 578882 156032 578938 156088
rect 578514 154536 578570 154592
rect 578514 148552 578570 148608
rect 578514 146920 578570 146976
rect 578606 143928 578662 143984
rect 579250 153076 579252 153096
rect 579252 153076 579304 153096
rect 579304 153076 579306 153096
rect 579250 153040 579306 153076
rect 579526 151544 579582 151600
rect 579434 150048 579490 150104
rect 603078 209480 603134 209536
rect 603170 208528 603226 208584
rect 603078 207440 603134 207496
rect 603078 206488 603134 206544
rect 603078 205400 603134 205456
rect 603170 204448 603226 204504
rect 603078 203360 603134 203416
rect 603078 202408 603134 202464
rect 603078 201356 603080 201376
rect 603080 201356 603132 201376
rect 603132 201356 603134 201376
rect 603078 201320 603134 201356
rect 603170 200368 603226 200424
rect 603078 199280 603134 199336
rect 603078 198328 603134 198384
rect 603078 197240 603134 197296
rect 603170 196288 603226 196344
rect 603078 195236 603080 195256
rect 603080 195236 603132 195256
rect 603132 195236 603134 195256
rect 603078 195200 603134 195236
rect 603078 194248 603134 194304
rect 603078 193160 603134 193216
rect 603078 192208 603134 192264
rect 603078 191120 603134 191176
rect 603170 190168 603226 190224
rect 603078 189116 603080 189136
rect 603080 189116 603132 189136
rect 603132 189116 603134 189136
rect 603078 189080 603134 189116
rect 603078 188128 603134 188184
rect 603078 187040 603134 187096
rect 603170 186088 603226 186144
rect 603078 185020 603134 185056
rect 603078 185000 603080 185020
rect 603080 185000 603132 185020
rect 603132 185000 603134 185020
rect 603078 184048 603134 184104
rect 603078 182960 603134 183016
rect 603170 182008 603226 182064
rect 603078 180920 603134 180976
rect 603078 179968 603134 180024
rect 603078 178880 603134 178936
rect 603170 177928 603226 177984
rect 603078 176840 603134 176896
rect 603078 175888 603134 175944
rect 603078 174800 603134 174856
rect 603722 173848 603778 173904
rect 603078 172760 603134 172816
rect 603078 171808 603134 171864
rect 603170 170720 603226 170776
rect 603078 169804 603080 169824
rect 603080 169804 603132 169824
rect 603132 169804 603134 169824
rect 603078 169768 603134 169804
rect 603078 168680 603134 168736
rect 603078 167728 603134 167784
rect 603078 166640 603134 166696
rect 603078 164600 603134 164656
rect 603814 165688 603870 165744
rect 603078 163648 603134 163704
rect 603078 162560 603134 162616
rect 603722 161608 603778 161664
rect 603078 160520 603134 160576
rect 603078 159568 603134 159624
rect 603170 158480 603226 158536
rect 603078 157528 603134 157584
rect 579526 145424 579582 145480
rect 579526 142432 579582 142488
rect 579342 140936 579398 140992
rect 579250 139440 579306 139496
rect 579526 137964 579582 138000
rect 579526 137944 579528 137964
rect 579528 137944 579580 137964
rect 579580 137944 579582 137964
rect 579526 136484 579528 136504
rect 579528 136484 579580 136504
rect 579580 136484 579582 136504
rect 579526 136448 579582 136484
rect 579158 134952 579214 135008
rect 579066 133456 579122 133512
rect 578974 131960 579030 132016
rect 579250 130464 579306 130520
rect 578882 128968 578938 129024
rect 578882 127472 578938 127528
rect 579066 125976 579122 126032
rect 578422 124480 578478 124536
rect 579250 122848 579306 122904
rect 579526 121388 579528 121408
rect 579528 121388 579580 121408
rect 579580 121388 579582 121408
rect 579526 121352 579582 121388
rect 579250 119856 579306 119912
rect 578606 118396 578608 118416
rect 578608 118396 578660 118416
rect 578660 118396 578662 118416
rect 578606 118360 578662 118396
rect 578422 112376 578478 112432
rect 578698 110880 578754 110936
rect 578514 103436 578516 103456
rect 578516 103436 578568 103456
rect 578568 103436 578570 103456
rect 578514 103400 578570 103436
rect 578330 101904 578386 101960
rect 578698 100272 578754 100328
rect 578606 95784 578662 95840
rect 578698 94288 578754 94344
rect 578514 80824 578570 80880
rect 189078 51720 189134 51776
rect 281446 50496 281502 50552
rect 216126 50360 216182 50416
rect 85118 50224 85174 50280
rect 543002 50224 543058 50280
rect 412454 46552 412510 46608
rect 473174 46280 473230 46336
rect 470138 46144 470194 46200
rect 419722 45464 419778 45520
rect 415398 45328 415454 45384
rect 241518 44956 241520 44976
rect 241520 44956 241572 44976
rect 241572 44956 241574 44976
rect 241518 44920 241574 44956
rect 246118 44956 246120 44976
rect 246120 44956 246172 44976
rect 246172 44956 246174 44976
rect 246118 44920 246174 44956
rect 251086 44940 251142 44976
rect 251086 44920 251088 44940
rect 251088 44920 251140 44940
rect 251140 44920 251142 44940
rect 255870 44940 255926 44976
rect 255870 44920 255872 44940
rect 255872 44920 255924 44940
rect 255924 44920 255926 44940
rect 241518 44820 241520 44840
rect 241520 44820 241572 44840
rect 241572 44820 241574 44840
rect 241518 44784 241574 44820
rect 246118 44820 246120 44840
rect 246120 44820 246172 44840
rect 246172 44820 246174 44840
rect 246118 44784 246174 44820
rect 251086 44804 251142 44840
rect 251086 44784 251088 44804
rect 251088 44784 251140 44804
rect 251140 44784 251142 44804
rect 255870 44804 255926 44840
rect 255870 44784 255872 44804
rect 255872 44784 255924 44804
rect 255924 44784 255926 44804
rect 142342 44240 142398 44296
rect 361762 43560 361818 43616
rect 307298 43424 307354 43480
rect 187514 42064 187570 42120
rect 194322 42064 194378 42120
rect 310104 42336 310160 42392
rect 365074 42064 365130 42120
rect 416686 41792 416742 41848
rect 460570 41792 460626 41848
rect 579526 116864 579582 116920
rect 579526 115368 579582 115424
rect 579250 113872 579306 113928
rect 579434 109384 579490 109440
rect 579250 107888 579306 107944
rect 579526 106392 579582 106448
rect 579526 104896 579582 104952
rect 579526 98776 579582 98832
rect 579526 97280 579582 97336
rect 579526 92792 579582 92848
rect 579526 91296 579582 91352
rect 579526 89800 579582 89856
rect 579526 88304 579582 88360
rect 579526 86808 579582 86864
rect 579526 85312 579582 85368
rect 579526 83816 579582 83872
rect 579158 82320 579214 82376
rect 579066 79328 579122 79384
rect 579526 77832 579582 77888
rect 578974 76200 579030 76256
rect 578882 73208 578938 73264
rect 578330 68720 578386 68776
rect 578698 61240 578754 61296
rect 578974 59744 579030 59800
rect 578882 58248 578938 58304
rect 578238 55256 578294 55312
rect 578882 56752 578938 56808
rect 578330 53760 578386 53816
rect 579526 74704 579582 74760
rect 579526 71732 579582 71768
rect 579526 71712 579528 71732
rect 579528 71712 579580 71732
rect 579580 71712 579582 71732
rect 579526 70216 579582 70272
rect 579526 67224 579582 67280
rect 579250 65764 579252 65784
rect 579252 65764 579304 65784
rect 579304 65764 579306 65784
rect 579250 65728 579306 65764
rect 579526 64268 579528 64288
rect 579528 64268 579580 64288
rect 579580 64268 579582 64288
rect 579526 64232 579582 64268
rect 579526 62736 579582 62792
rect 603078 156440 603134 156496
rect 603078 155488 603134 155544
rect 603170 154400 603226 154456
rect 603078 153448 603134 153504
rect 603078 152360 603134 152416
rect 603078 151408 603134 151464
rect 603170 150320 603226 150376
rect 603078 149368 603134 149424
rect 603078 148280 603134 148336
rect 603078 147328 603134 147384
rect 603170 146240 603226 146296
rect 603906 145288 603962 145344
rect 603078 144200 603134 144256
rect 603722 143248 603778 143304
rect 603078 142180 603134 142216
rect 603078 142160 603080 142180
rect 603080 142160 603132 142180
rect 603132 142160 603134 142180
rect 603078 141208 603134 141264
rect 603078 140120 603134 140176
rect 603170 139168 603226 139224
rect 603078 138080 603134 138136
rect 603078 137128 603134 137184
rect 603078 136040 603134 136096
rect 603170 135088 603226 135144
rect 603078 134000 603134 134056
rect 603078 133048 603134 133104
rect 603078 131960 603134 132016
rect 603078 131008 603134 131064
rect 603078 128968 603134 129024
rect 603078 127880 603134 127936
rect 603170 126928 603226 126984
rect 603078 125840 603134 125896
rect 603078 124888 603134 124944
rect 602434 123800 602490 123856
rect 602342 118768 602398 118824
rect 603078 122868 603134 122904
rect 603078 122848 603080 122868
rect 603080 122848 603132 122868
rect 603132 122848 603134 122868
rect 603078 121760 603134 121816
rect 603078 120808 603134 120864
rect 603078 119720 603134 119776
rect 603078 117680 603134 117736
rect 603814 129920 603870 129976
rect 603446 116728 603502 116784
rect 603078 115640 603134 115696
rect 603170 114688 603226 114744
rect 603078 113600 603134 113656
rect 603078 112648 603134 112704
rect 603078 111560 603134 111616
rect 603814 110608 603870 110664
rect 603078 109520 603134 109576
rect 603078 108568 603134 108624
rect 603078 107480 603134 107536
rect 603170 106528 603226 106584
rect 603078 105440 603134 105496
rect 603722 104488 603778 104544
rect 603170 103400 603226 103456
rect 603078 102448 603134 102504
rect 603078 101360 603134 101416
rect 603078 100408 603134 100464
rect 610346 216824 610402 216880
rect 622490 216688 622546 216744
rect 623962 219408 624018 219464
rect 648618 267008 648674 267064
rect 647330 230424 647386 230480
rect 648526 213016 648582 213072
rect 651654 975840 651710 975896
rect 652022 962512 652078 962568
rect 651562 949320 651618 949376
rect 651562 936128 651618 936184
rect 651562 922664 651618 922720
rect 651562 909492 651618 909528
rect 651562 909472 651564 909492
rect 651564 909472 651616 909492
rect 651616 909472 651618 909492
rect 651562 896144 651618 896200
rect 652022 882816 652078 882872
rect 651562 869624 651618 869680
rect 651562 856296 651618 856352
rect 651562 842968 651618 843024
rect 651562 829776 651618 829832
rect 651562 816448 651618 816504
rect 651562 803256 651618 803312
rect 651654 789928 651710 789984
rect 651562 776600 651618 776656
rect 651562 763272 651618 763328
rect 651562 750080 651618 750136
rect 651562 736752 651618 736808
rect 652022 723424 652078 723480
rect 651562 710232 651618 710288
rect 652022 696904 652078 696960
rect 651838 683576 651894 683632
rect 651562 670384 651618 670440
rect 651562 657056 651618 657112
rect 651562 643728 651618 643784
rect 651562 630536 651618 630592
rect 651562 603880 651618 603936
rect 651562 590708 651618 590744
rect 651562 590688 651564 590708
rect 651564 590688 651616 590708
rect 651616 590688 651618 590708
rect 652390 617208 652446 617264
rect 651562 577360 651618 577416
rect 652114 564032 652170 564088
rect 651562 550840 651618 550896
rect 651562 537512 651618 537568
rect 651562 524184 651618 524240
rect 651562 510992 651618 511048
rect 651562 497664 651618 497720
rect 651562 484472 651618 484528
rect 651654 471144 651710 471200
rect 651562 457816 651618 457872
rect 651562 444488 651618 444544
rect 651562 431296 651618 431352
rect 651562 417968 651618 418024
rect 652022 404640 652078 404696
rect 651562 391448 651618 391504
rect 651562 378156 651564 378176
rect 651564 378156 651616 378176
rect 651616 378156 651618 378176
rect 651562 378120 651618 378156
rect 652022 364792 652078 364848
rect 651562 351600 651618 351656
rect 651654 338272 651710 338328
rect 651562 324944 651618 325000
rect 652390 311752 652446 311808
rect 652022 298424 652078 298480
rect 651562 285232 651618 285288
rect 654138 218456 654194 218512
rect 666926 209208 666982 209264
rect 666834 204176 666890 204232
rect 666834 200776 666890 200832
rect 666742 199008 666798 199064
rect 666650 193976 666706 194032
rect 666650 190576 666706 190632
rect 666558 188944 666614 189000
rect 666558 185544 666614 185600
rect 666558 163512 666614 163568
rect 666558 161472 666614 161528
rect 666558 153312 666614 153368
rect 666558 151816 666614 151872
rect 666558 151544 666614 151600
rect 666558 149912 666614 149968
rect 666558 142024 666614 142080
rect 666558 139712 666614 139768
rect 667938 209208 667994 209264
rect 667938 205808 667994 205864
rect 667938 199008 667994 199064
rect 667938 195608 667994 195664
rect 668030 183776 668086 183832
rect 668030 180376 668086 180432
rect 667938 178780 667940 178800
rect 667940 178780 667992 178800
rect 667992 178780 667994 178800
rect 667938 178744 667994 178780
rect 667938 175344 667994 175400
rect 667938 173612 667940 173632
rect 667940 173612 667992 173632
rect 667992 173612 667994 173632
rect 667938 173576 667994 173612
rect 667938 171128 667994 171184
rect 667938 168544 667994 168600
rect 667938 165144 667994 165200
rect 667938 158344 667994 158400
rect 667938 154944 667994 155000
rect 667938 143112 667994 143168
rect 668030 138080 668086 138136
rect 668030 134680 668086 134736
rect 666558 132368 666614 132424
rect 666558 129512 666614 129568
rect 668030 127880 668086 127936
rect 668030 124480 668086 124536
rect 667938 122848 667994 122904
rect 666558 122712 666614 122768
rect 666558 119448 666614 119504
rect 667938 110880 667994 110936
rect 667938 109248 667994 109304
rect 668306 183776 668362 183832
rect 668398 163512 668454 163568
rect 668582 158344 668638 158400
rect 668674 153312 668730 153368
rect 668306 148144 668362 148200
rect 668306 144880 668362 144936
rect 668582 132948 668584 132968
rect 668584 132948 668636 132968
rect 668636 132948 668638 132968
rect 668582 132912 668638 132948
rect 668490 116048 668546 116104
rect 668490 114316 668492 114336
rect 668492 114316 668544 114336
rect 668544 114316 668546 114336
rect 668490 114280 668546 114316
rect 668122 107480 668178 107536
rect 668674 104080 668730 104136
rect 669226 117680 669282 117736
rect 668858 112648 668914 112704
rect 669226 105848 669282 105904
rect 668766 102448 668822 102504
rect 668582 100816 668638 100872
rect 576122 44920 576178 44976
rect 478786 44648 478842 44704
rect 605838 43560 605894 43616
rect 607310 45192 607366 45248
rect 608598 45056 608654 45112
rect 607218 43424 607274 43480
rect 518622 42336 518678 42392
rect 471610 42064 471666 42120
rect 514850 42064 514906 42120
rect 520370 42064 520426 42120
rect 521750 42064 521806 42120
rect 525982 42064 526038 42120
rect 529662 42064 529718 42120
rect 610070 45464 610126 45520
rect 610162 45328 610218 45384
rect 611450 46416 611506 46472
rect 626354 92520 626410 92576
rect 628286 95920 628342 95976
rect 641718 96600 641774 96656
rect 642270 96464 642326 96520
rect 627826 94424 627882 94480
rect 626538 93472 626594 93528
rect 626446 91568 626502 91624
rect 625986 90616 626042 90672
rect 625802 89664 625858 89720
rect 643098 89528 643154 89584
rect 626446 88848 626502 88904
rect 626446 87896 626502 87952
rect 626354 86944 626410 87000
rect 626446 85992 626502 86048
rect 643190 85176 643246 85232
rect 626446 85040 626502 85096
rect 625618 84124 625620 84144
rect 625620 84124 625672 84144
rect 625672 84124 625674 84144
rect 625618 84088 625674 84124
rect 626446 83136 626502 83192
rect 644570 94560 644626 94616
rect 644662 92112 644718 92168
rect 644478 87080 644534 87136
rect 626446 82184 626502 82240
rect 643282 82184 643338 82240
rect 629206 80824 629262 80880
rect 633898 77832 633954 77888
rect 639602 77696 639658 77752
rect 623778 74704 623834 74760
rect 633530 74704 633586 74760
rect 639234 75112 639290 75168
rect 646870 74432 646926 74488
rect 646962 72936 647018 72992
rect 646134 71712 646190 71768
rect 647238 69944 647294 70000
rect 655334 93336 655390 93392
rect 654782 92520 654838 92576
rect 654322 91432 654378 91488
rect 654874 90616 654930 90672
rect 655426 89800 655482 89856
rect 657358 94696 657414 94752
rect 663798 92520 663854 92576
rect 663890 90616 663946 90672
rect 665178 91704 665234 91760
rect 665362 93336 665418 93392
rect 665270 89800 665326 89856
rect 664074 88984 664130 89040
rect 648802 68448 648858 68504
rect 647422 66952 647478 67008
rect 646134 66000 646190 66056
rect 646134 64368 646190 64424
rect 661130 47504 661186 47560
rect 648159 46664 649615 47120
rect 612830 46280 612886 46336
rect 612738 46144 612794 46200
rect 675758 966456 675814 966512
rect 675758 966184 675814 966240
rect 675758 964960 675814 965016
rect 675758 963328 675814 963384
rect 675666 962784 675722 962840
rect 675482 961832 675538 961888
rect 672354 759056 672410 759112
rect 672814 758376 672870 758432
rect 675758 959112 675814 959168
rect 675022 957888 675078 957944
rect 675758 957752 675814 957808
rect 675390 953944 675446 954000
rect 679806 949728 679862 949784
rect 679622 949592 679678 949648
rect 676862 949456 676918 949512
rect 676034 939936 676090 939992
rect 676218 939256 676274 939312
rect 676034 939156 676036 939176
rect 676036 939156 676088 939176
rect 676088 939156 676090 939176
rect 676034 939120 676090 939156
rect 676034 938712 676090 938768
rect 676034 938324 676090 938360
rect 676034 938304 676036 938324
rect 676036 938304 676088 938324
rect 676088 938304 676090 938324
rect 676218 937624 676274 937680
rect 676034 937508 676090 937544
rect 676034 937488 676036 937508
rect 676036 937488 676088 937508
rect 676088 937488 676090 937508
rect 676218 937236 676274 937272
rect 676218 937216 676220 937236
rect 676220 937216 676272 937236
rect 676272 937216 676274 937236
rect 676126 936400 676182 936456
rect 676034 935856 676090 935912
rect 676218 935992 676274 936048
rect 676862 935176 676918 935232
rect 678242 933544 678298 933600
rect 679806 932728 679862 932784
rect 679622 932320 679678 932376
rect 676034 931776 676090 931832
rect 676218 930724 676220 930744
rect 676220 930724 676272 930744
rect 676272 930724 676274 930744
rect 676218 930688 676274 930724
rect 676218 930300 676274 930336
rect 676218 930280 676220 930300
rect 676220 930280 676272 930300
rect 676272 930280 676274 930300
rect 683118 929464 683174 929520
rect 683118 928648 683174 928704
rect 675390 877240 675446 877296
rect 675758 876560 675814 876616
rect 675758 875880 675814 875936
rect 675758 873976 675814 874032
rect 675758 866768 675814 866824
rect 675758 864728 675814 864784
rect 675482 784760 675538 784816
rect 675758 784080 675814 784136
rect 675390 779864 675446 779920
rect 675390 775648 675446 775704
rect 675758 773336 675814 773392
rect 674746 757424 674802 757480
rect 679622 772656 679678 772712
rect 676126 761232 676182 761288
rect 676034 760688 676090 760744
rect 676218 760844 676274 760880
rect 676218 760824 676220 760844
rect 676220 760824 676272 760844
rect 676272 760824 676274 760844
rect 676034 760316 676036 760336
rect 676036 760316 676088 760336
rect 676088 760316 676090 760336
rect 676034 760280 676090 760316
rect 676218 759600 676274 759656
rect 676034 759500 676036 759520
rect 676036 759500 676088 759520
rect 676088 759500 676090 759520
rect 676034 759464 676090 759500
rect 676034 759076 676090 759112
rect 676034 759056 676036 759076
rect 676036 759056 676088 759076
rect 676088 759056 676090 759076
rect 676034 758260 676090 758296
rect 676034 758240 676036 758260
rect 676036 758240 676088 758260
rect 676088 758240 676090 758260
rect 679622 756744 679678 756800
rect 675758 756200 675814 756256
rect 676218 755556 676220 755576
rect 676220 755556 676272 755576
rect 676272 755556 676274 755576
rect 676218 755520 676274 755556
rect 676034 754996 676090 755032
rect 676034 754976 676036 754996
rect 676036 754976 676088 754996
rect 676088 754976 676090 754996
rect 676218 754332 676220 754352
rect 676220 754332 676272 754352
rect 676272 754332 676274 754352
rect 676218 754296 676274 754332
rect 676034 753752 676090 753808
rect 676218 753108 676220 753128
rect 676220 753108 676272 753128
rect 676272 753108 676274 753128
rect 676218 753072 676274 753108
rect 676218 752700 676220 752720
rect 676220 752700 676272 752720
rect 676272 752700 676274 752720
rect 676218 752664 676274 752700
rect 676218 752276 676274 752312
rect 676218 752256 676220 752276
rect 676220 752256 676272 752276
rect 676272 752256 676274 752276
rect 676218 751440 676274 751496
rect 683118 751032 683174 751088
rect 683118 750216 683174 750272
rect 675482 741648 675538 741704
rect 675758 739880 675814 739936
rect 675666 739200 675722 739256
rect 675758 734304 675814 734360
rect 675758 732944 675814 733000
rect 678242 727232 678298 727288
rect 676034 716488 676090 716544
rect 676034 716116 676036 716136
rect 676036 716116 676088 716136
rect 676088 716116 676090 716136
rect 676034 716080 676090 716116
rect 676034 715672 676090 715728
rect 675942 715300 675944 715320
rect 675944 715300 675996 715320
rect 675996 715300 675998 715320
rect 675942 715264 675998 715300
rect 676034 714876 676090 714912
rect 676034 714856 676036 714876
rect 676036 714856 676088 714876
rect 676088 714856 676090 714876
rect 676034 714484 676036 714504
rect 676036 714484 676088 714504
rect 676088 714484 676090 714504
rect 676034 714448 676090 714484
rect 676034 714060 676090 714096
rect 676034 714040 676036 714060
rect 676036 714040 676088 714060
rect 676088 714040 676090 714060
rect 676034 713668 676036 713688
rect 676036 713668 676088 713688
rect 676088 713668 676090 713688
rect 676034 713632 676090 713668
rect 677322 713432 677378 713488
rect 676034 713244 676090 713280
rect 676034 713224 676036 713244
rect 676036 713224 676088 713244
rect 676088 713224 676090 713244
rect 674746 712816 674802 712872
rect 676034 712428 676090 712464
rect 676034 712408 676036 712428
rect 676036 712408 676088 712428
rect 676088 712408 676090 712428
rect 676034 712036 676036 712056
rect 676036 712036 676088 712056
rect 676088 712036 676090 712056
rect 676034 712000 676090 712036
rect 676034 711220 676036 711240
rect 676036 711220 676088 711240
rect 676088 711220 676090 711240
rect 676034 711184 676090 711220
rect 675942 711048 675998 711104
rect 676034 710404 676036 710424
rect 676036 710404 676088 710424
rect 676088 710404 676090 710424
rect 676034 710368 676090 710404
rect 676034 709996 676036 710016
rect 676036 709996 676088 710016
rect 676088 709996 676090 710016
rect 676034 709960 676090 709996
rect 676034 709588 676036 709608
rect 676036 709588 676088 709608
rect 676088 709588 676090 709608
rect 676034 709552 676090 709588
rect 676034 709180 676036 709200
rect 676036 709180 676088 709200
rect 676088 709180 676090 709200
rect 676034 709144 676090 709180
rect 676034 708364 676036 708384
rect 676036 708364 676088 708384
rect 676088 708364 676090 708384
rect 676034 708328 676090 708364
rect 678242 711592 678298 711648
rect 676034 707920 676090 707976
rect 676034 707548 676036 707568
rect 676036 707548 676088 707568
rect 676088 707548 676090 707568
rect 676034 707512 676090 707548
rect 676034 707140 676036 707160
rect 676036 707140 676088 707160
rect 676088 707140 676090 707160
rect 676034 707104 676090 707140
rect 676034 706732 676036 706752
rect 676036 706732 676088 706752
rect 676088 706732 676090 706752
rect 676034 706696 676090 706732
rect 676034 706288 676090 706344
rect 676034 705064 676090 705120
rect 675942 704384 675998 704440
rect 675390 697312 675446 697368
rect 675666 696904 675722 696960
rect 675758 695000 675814 695056
rect 675758 694184 675814 694240
rect 678242 678952 678298 679008
rect 676218 671064 676274 671120
rect 676034 670928 676090 670984
rect 676310 670248 676366 670304
rect 676126 669840 676182 669896
rect 674746 669704 674802 669760
rect 676218 669432 676274 669488
rect 676034 668908 676090 668944
rect 676034 668888 676036 668908
rect 676036 668888 676088 668908
rect 676088 668888 676090 668908
rect 676218 668652 676220 668672
rect 676220 668652 676272 668672
rect 676272 668652 676274 668672
rect 676218 668616 676274 668652
rect 676034 668072 676090 668128
rect 676218 667836 676220 667856
rect 676220 667836 676272 667856
rect 676272 667836 676274 667856
rect 676218 667800 676274 667836
rect 676218 666984 676274 667040
rect 678242 666984 678298 667040
rect 676034 666476 676036 666496
rect 676036 666476 676088 666496
rect 676088 666476 676090 666496
rect 676034 666440 676090 666476
rect 676218 665760 676274 665816
rect 676034 665252 676036 665272
rect 676036 665252 676088 665272
rect 676088 665252 676090 665272
rect 676034 665216 676090 665252
rect 676218 664980 676220 665000
rect 676220 664980 676272 665000
rect 676272 664980 676274 665000
rect 676218 664944 676274 664980
rect 676218 664128 676274 664184
rect 676218 663756 676220 663776
rect 676220 663756 676272 663776
rect 676272 663756 676274 663776
rect 676218 663720 676274 663756
rect 676034 662380 676090 662416
rect 676034 662360 676036 662380
rect 676036 662360 676088 662380
rect 676088 662360 676090 662380
rect 676218 661680 676274 661736
rect 676034 661580 676036 661600
rect 676036 661580 676088 661600
rect 676088 661580 676090 661600
rect 676034 661544 676090 661580
rect 683118 660864 683174 660920
rect 683118 660048 683174 660104
rect 675482 652160 675538 652216
rect 675758 651480 675814 651536
rect 675390 649168 675446 649224
rect 675758 648624 675814 648680
rect 675758 644680 675814 644736
rect 675666 643048 675722 643104
rect 675482 640328 675538 640384
rect 675666 638152 675722 638208
rect 674746 625096 674802 625152
rect 678242 633392 678298 633448
rect 676126 626048 676182 626104
rect 676218 625640 676274 625696
rect 676218 625232 676274 625288
rect 676218 624416 676274 624472
rect 676034 624316 676036 624336
rect 676036 624316 676088 624336
rect 676088 624316 676090 624336
rect 676034 624280 676090 624316
rect 676034 623892 676090 623928
rect 676034 623872 676036 623892
rect 676036 623872 676088 623892
rect 676088 623872 676090 623892
rect 676126 623192 676182 623248
rect 676034 622684 676036 622704
rect 676036 622684 676088 622704
rect 676088 622684 676090 622704
rect 676034 622648 676090 622684
rect 676218 622784 676274 622840
rect 676034 622260 676090 622296
rect 676034 622240 676036 622260
rect 676036 622240 676088 622260
rect 676088 622240 676090 622260
rect 678242 621968 678298 622024
rect 676034 621424 676090 621480
rect 676218 621152 676274 621208
rect 676218 619948 676274 619984
rect 676218 619928 676220 619948
rect 676220 619928 676272 619948
rect 676272 619928 676274 619948
rect 676034 619812 676090 619848
rect 676034 619792 676036 619812
rect 676036 619792 676088 619812
rect 676088 619792 676090 619812
rect 676218 619148 676220 619168
rect 676220 619148 676272 619168
rect 676272 619148 676274 619168
rect 676218 619112 676274 619148
rect 676126 617888 676182 617944
rect 676034 617788 676036 617808
rect 676036 617788 676088 617808
rect 676088 617788 676090 617808
rect 676034 617752 676090 617788
rect 676218 617072 676274 617128
rect 676034 616972 676036 616992
rect 676036 616972 676088 616992
rect 676088 616972 676090 616992
rect 676034 616936 676090 616972
rect 676218 616256 676274 616312
rect 683118 615848 683174 615904
rect 683118 615032 683174 615088
rect 675482 607824 675538 607880
rect 675390 606464 675446 606520
rect 675206 600888 675262 600944
rect 675574 600208 675630 600264
rect 675758 598984 675814 599040
rect 675758 597760 675814 597816
rect 675482 593136 675538 593192
rect 675666 593136 675722 593192
rect 678242 589192 678298 589248
rect 676034 581052 676090 581088
rect 676034 581032 676036 581052
rect 676036 581032 676088 581052
rect 676088 581032 676090 581052
rect 676126 580488 676182 580544
rect 676034 580216 676090 580272
rect 676218 580100 676274 580136
rect 676218 580080 676220 580100
rect 676220 580080 676272 580100
rect 676272 580080 676274 580100
rect 676218 579284 676274 579320
rect 676218 579264 676220 579284
rect 676220 579264 676272 579284
rect 676272 579264 676274 579284
rect 676218 578856 676274 578912
rect 676034 578604 676090 578640
rect 676034 578584 676036 578604
rect 676036 578584 676088 578604
rect 676088 578584 676090 578604
rect 676218 578040 676274 578096
rect 676126 577632 676182 577688
rect 676034 577396 676036 577416
rect 676036 577396 676088 577416
rect 676088 577396 676090 577416
rect 676034 577360 676090 577396
rect 676034 576972 676090 577008
rect 676034 576952 676036 576972
rect 676036 576952 676088 576972
rect 676088 576952 676090 576972
rect 678242 576816 678298 576872
rect 675666 576136 675722 576192
rect 676218 575612 676274 575648
rect 676218 575592 676220 575612
rect 676220 575592 676272 575612
rect 676272 575592 676274 575612
rect 676034 575356 676036 575376
rect 676036 575356 676088 575376
rect 676088 575356 676090 575376
rect 676034 575320 676090 575356
rect 676218 574776 676274 574832
rect 676034 574540 676036 574560
rect 676036 574540 676088 574560
rect 676088 574540 676090 574560
rect 676034 574504 676090 574540
rect 676218 571920 676274 571976
rect 676034 571684 676036 571704
rect 676036 571684 676088 571704
rect 676088 571684 676090 571704
rect 676034 571648 676090 571684
rect 676218 571104 676274 571160
rect 683118 570696 683174 570752
rect 683118 569880 683174 569936
rect 675482 568520 675538 568576
rect 675758 562672 675814 562728
rect 675758 561176 675814 561232
rect 675482 559544 675538 559600
rect 675758 558320 675814 558376
rect 675758 551928 675814 551984
rect 681002 546488 681058 546544
rect 678242 543768 678298 543824
rect 676218 535880 676274 535936
rect 676034 535676 676090 535732
rect 676218 535064 676274 535120
rect 676034 534896 676036 534916
rect 676036 534896 676088 534916
rect 676088 534896 676090 534916
rect 676034 534860 676090 534896
rect 676034 534080 676036 534100
rect 676036 534080 676088 534100
rect 676088 534080 676090 534100
rect 676034 534044 676090 534080
rect 676218 533024 676274 533080
rect 677322 532616 677378 532672
rect 676218 532208 676274 532264
rect 676218 530984 676274 531040
rect 676034 530408 676036 530428
rect 676036 530408 676088 530428
rect 676088 530408 676090 530428
rect 676034 530372 676090 530408
rect 676126 529352 676182 529408
rect 676034 528740 676090 528796
rect 676218 528944 676274 529000
rect 676034 528368 676036 528388
rect 676036 528368 676088 528388
rect 676088 528368 676090 528388
rect 676034 528332 676090 528368
rect 676218 526904 676274 526960
rect 676034 526736 676036 526756
rect 676036 526736 676088 526756
rect 676088 526736 676090 526756
rect 676034 526700 676090 526736
rect 676034 526328 676036 526348
rect 676036 526328 676088 526348
rect 676088 526328 676090 526348
rect 676034 526292 676090 526328
rect 675942 492088 675998 492144
rect 676034 491680 676090 491736
rect 676034 491272 676090 491328
rect 676034 490864 676090 490920
rect 676034 490456 676090 490512
rect 675850 490048 675906 490104
rect 675942 489268 675944 489288
rect 675944 489268 675996 489288
rect 675996 489268 675998 489288
rect 675942 489232 675998 489268
rect 675942 488824 675998 488880
rect 675942 488452 675944 488472
rect 675944 488452 675996 488472
rect 675996 488452 675998 488472
rect 675942 488416 675998 488452
rect 675850 488028 675906 488064
rect 675850 488008 675852 488028
rect 675852 488008 675904 488028
rect 675904 488008 675906 488028
rect 675942 487192 675998 487248
rect 675942 486004 675944 486024
rect 675944 486004 675996 486024
rect 675996 486004 675998 486024
rect 675942 485968 675998 486004
rect 674746 485560 674802 485616
rect 675850 485152 675906 485208
rect 675942 484744 675998 484800
rect 675942 483556 675944 483576
rect 675944 483556 675996 483576
rect 675996 483556 675998 483576
rect 675942 483520 675998 483556
rect 675942 483132 675998 483168
rect 675942 483112 675944 483132
rect 675944 483112 675996 483132
rect 675996 483112 675998 483132
rect 675850 482704 675906 482760
rect 675942 482296 675998 482352
rect 673918 251640 673974 251696
rect 673734 249736 673790 249792
rect 673826 249600 673882 249656
rect 673918 246200 673974 246256
rect 673826 246064 673882 246120
rect 677506 531800 677562 531856
rect 678242 531800 678298 531856
rect 677414 489872 677470 489928
rect 676034 402600 676090 402656
rect 676218 403688 676274 403744
rect 676218 403300 676274 403336
rect 676218 403280 676220 403300
rect 676220 403280 676272 403300
rect 676272 403280 676274 403300
rect 676402 403280 676458 403336
rect 676218 402056 676274 402112
rect 676126 401240 676182 401296
rect 676034 400968 676090 401024
rect 683302 534248 683358 534304
rect 681002 530984 681058 531040
rect 683118 525680 683174 525736
rect 683118 524864 683174 524920
rect 683670 533432 683726 533488
rect 679622 503648 679678 503704
rect 679806 503512 679862 503568
rect 679622 486784 679678 486840
rect 679806 486376 679862 486432
rect 678978 480664 679034 480720
rect 677322 402056 677378 402112
rect 676218 400424 676274 400480
rect 677230 400424 677286 400480
rect 676218 399628 676274 399664
rect 676218 399608 676220 399628
rect 676220 399608 676272 399628
rect 676272 399608 676274 399628
rect 676034 398520 676090 398576
rect 676034 398112 676090 398168
rect 676862 397568 676918 397624
rect 676494 394712 676550 394768
rect 676218 394304 676274 394360
rect 676034 394052 676090 394088
rect 676034 394032 676036 394052
rect 676036 394032 676088 394052
rect 676088 394032 676090 394052
rect 676954 396752 677010 396808
rect 676862 388456 676918 388512
rect 679622 396344 679678 396400
rect 678242 395936 678298 395992
rect 683118 393488 683174 393544
rect 683118 392264 683174 392320
rect 679622 388184 679678 388240
rect 675758 384920 675814 384976
rect 675390 382200 675446 382256
rect 675482 378664 675538 378720
rect 675758 377304 675814 377360
rect 675758 374992 675814 375048
rect 675758 373632 675814 373688
rect 675758 372000 675814 372056
rect 675850 358672 675906 358728
rect 675942 358264 675998 358320
rect 676034 357856 676090 357912
rect 676034 357484 676036 357504
rect 676036 357484 676088 357504
rect 676088 357484 676090 357504
rect 676034 357448 676090 357484
rect 676034 357060 676090 357096
rect 676034 357040 676036 357060
rect 676036 357040 676088 357060
rect 676088 357040 676090 357060
rect 676034 356668 676036 356688
rect 676036 356668 676088 356688
rect 676088 356668 676090 356688
rect 676034 356632 676090 356668
rect 676034 356244 676090 356280
rect 676034 356224 676036 356244
rect 676036 356224 676088 356244
rect 676088 356224 676090 356244
rect 676034 355852 676036 355872
rect 676036 355852 676088 355872
rect 676088 355852 676090 355872
rect 676034 355816 676090 355852
rect 676034 355428 676090 355464
rect 676034 355408 676036 355428
rect 676036 355408 676088 355428
rect 676088 355408 676090 355428
rect 674746 355000 674802 355056
rect 676034 354612 676090 354648
rect 676034 354592 676036 354612
rect 676036 354592 676088 354612
rect 676088 354592 676090 354612
rect 679622 352552 679678 352608
rect 676034 351328 676090 351384
rect 676034 350940 676090 350976
rect 676034 350920 676036 350940
rect 676036 350920 676088 350940
rect 676088 350920 676090 350940
rect 676034 350548 676036 350568
rect 676036 350548 676088 350568
rect 676088 350548 676090 350568
rect 676034 350512 676090 350548
rect 676034 350104 676090 350160
rect 675942 349696 675998 349752
rect 676034 349308 676090 349344
rect 676034 349288 676036 349308
rect 676036 349288 676088 349308
rect 676088 349288 676090 349308
rect 676034 348900 676090 348936
rect 676034 348880 676036 348900
rect 676036 348880 676088 348900
rect 676088 348880 676090 348900
rect 676034 348472 676090 348528
rect 676034 347248 676090 347304
rect 675942 346568 675998 346624
rect 676126 346432 676182 346488
rect 676770 346432 676826 346488
rect 679806 351736 679862 351792
rect 679622 342352 679678 342408
rect 675298 342216 675354 342272
rect 679806 342216 679862 342272
rect 675666 340720 675722 340776
rect 675758 339360 675814 339416
rect 675482 337864 675538 337920
rect 675758 335824 675814 335880
rect 674838 335280 674894 335336
rect 675758 333512 675814 333568
rect 675758 332152 675814 332208
rect 675114 325624 675170 325680
rect 675758 325488 675814 325544
rect 676218 313540 676274 313576
rect 676218 313520 676220 313540
rect 676220 313520 676272 313540
rect 676272 313520 676274 313540
rect 676034 313248 676090 313304
rect 676218 312704 676274 312760
rect 676034 312468 676036 312488
rect 676036 312468 676088 312488
rect 676088 312468 676090 312488
rect 676034 312432 676090 312468
rect 676218 311908 676274 311944
rect 676218 311888 676220 311908
rect 676220 311888 676272 311908
rect 676272 311888 676274 311908
rect 676034 311652 676036 311672
rect 676036 311652 676088 311672
rect 676088 311652 676090 311672
rect 676034 311616 676090 311652
rect 676218 311092 676274 311128
rect 676218 311072 676220 311092
rect 676220 311072 676272 311092
rect 676272 311072 676274 311092
rect 676218 310684 676274 310720
rect 676218 310664 676220 310684
rect 676220 310664 676272 310684
rect 676272 310664 676274 310684
rect 676310 310256 676366 310312
rect 676126 309848 676182 309904
rect 676218 309460 676274 309496
rect 676218 309440 676220 309460
rect 676220 309440 676272 309460
rect 676272 309440 676274 309460
rect 681002 309032 681058 309088
rect 679714 308216 679770 308272
rect 679622 307808 679678 307864
rect 676862 306584 676918 306640
rect 676310 306176 676366 306232
rect 676218 304564 676274 304600
rect 676218 304544 676220 304564
rect 676220 304544 676272 304564
rect 676272 304544 676274 304564
rect 676126 304136 676182 304192
rect 676218 303748 676274 303784
rect 676218 303728 676220 303748
rect 676220 303728 676272 303748
rect 676272 303728 676274 303748
rect 676402 305768 676458 305824
rect 677598 305360 677654 305416
rect 683118 303320 683174 303376
rect 683118 302504 683174 302560
rect 681002 299376 681058 299432
rect 679622 297744 679678 297800
rect 677598 297472 677654 297528
rect 676310 297336 676366 297392
rect 675758 294752 675814 294808
rect 675666 292576 675722 292632
rect 675482 292032 675538 292088
rect 675758 288360 675814 288416
rect 675758 287272 675814 287328
rect 675482 285504 675538 285560
rect 675758 283600 675814 283656
rect 675758 281424 675814 281480
rect 676218 268504 676274 268560
rect 676126 268096 676182 268152
rect 676218 267688 676274 267744
rect 674746 267416 674802 267472
rect 676218 266892 676274 266928
rect 676218 266872 676220 266892
rect 676220 266872 676272 266892
rect 676272 266872 676274 266892
rect 676034 266636 676036 266656
rect 676036 266636 676088 266656
rect 676088 266636 676090 266656
rect 676034 266600 676090 266636
rect 676218 266076 676274 266112
rect 676218 266056 676220 266076
rect 676220 266056 676272 266076
rect 676272 266056 676274 266076
rect 676218 265648 676274 265704
rect 676126 265240 676182 265296
rect 676034 264968 676090 265024
rect 676218 264424 676274 264480
rect 678242 263200 678298 263256
rect 676862 261160 676918 261216
rect 676402 259936 676458 259992
rect 676218 259140 676274 259176
rect 676218 259120 676220 259140
rect 676220 259120 676272 259140
rect 676272 259120 676274 259140
rect 676218 258712 676274 258768
rect 676494 259528 676550 259584
rect 676402 251640 676458 251696
rect 676954 260752 677010 260808
rect 678334 262384 678390 262440
rect 683118 258304 683174 258360
rect 683118 257488 683174 257544
rect 678334 252592 678390 252648
rect 675758 250280 675814 250336
rect 675758 249736 675814 249792
rect 675022 249600 675078 249656
rect 675206 249464 675262 249520
rect 675206 246200 675262 246256
rect 675298 241848 675354 241904
rect 675390 240216 675446 240272
rect 675758 238448 675814 238504
rect 675758 236816 675814 236872
rect 676034 223488 676090 223544
rect 675942 223116 675944 223136
rect 675944 223116 675996 223136
rect 675996 223116 675998 223136
rect 675942 223080 675998 223116
rect 675942 222708 675944 222728
rect 675944 222708 675996 222728
rect 675996 222708 675998 222728
rect 675942 222672 675998 222708
rect 674746 222264 674802 222320
rect 676034 221876 676090 221912
rect 676034 221856 676036 221876
rect 676036 221856 676088 221876
rect 676088 221856 676090 221876
rect 676034 221484 676036 221504
rect 676036 221484 676088 221504
rect 676088 221484 676090 221504
rect 676034 221448 676090 221484
rect 676034 221060 676090 221096
rect 676034 221040 676036 221060
rect 676036 221040 676088 221060
rect 676088 221040 676090 221060
rect 676034 220668 676036 220688
rect 676036 220668 676088 220688
rect 676088 220668 676090 220688
rect 676034 220632 676090 220668
rect 676034 220244 676090 220280
rect 676034 220224 676036 220244
rect 676036 220224 676088 220244
rect 676088 220224 676090 220244
rect 676034 219852 676036 219872
rect 676036 219852 676088 219872
rect 676088 219852 676090 219872
rect 676034 219816 676090 219852
rect 674746 219408 674802 219464
rect 676034 219000 676090 219056
rect 676034 216552 676090 216608
rect 676034 216164 676090 216200
rect 676034 216144 676036 216164
rect 676036 216144 676088 216164
rect 676088 216144 676090 216164
rect 676034 215756 676090 215792
rect 676034 215736 676036 215756
rect 676036 215736 676088 215756
rect 676088 215736 676090 215756
rect 675942 215328 675998 215384
rect 675850 214920 675906 214976
rect 676034 214124 676090 214160
rect 676034 214104 676036 214124
rect 676036 214104 676088 214124
rect 676088 214104 676090 214124
rect 676034 213968 676090 214024
rect 679622 217368 679678 217424
rect 676034 213716 676090 213752
rect 676034 213696 676036 213716
rect 676036 213696 676088 213716
rect 676088 213696 676090 213716
rect 676034 213288 676090 213344
rect 676034 212064 676090 212120
rect 675942 211384 675998 211440
rect 675850 211248 675906 211304
rect 676862 208256 676918 208312
rect 679622 207168 679678 207224
rect 675390 205536 675446 205592
rect 675758 204992 675814 205048
rect 675758 204176 675814 204232
rect 675114 202816 675170 202872
rect 674838 201320 674894 201376
rect 675758 202680 675814 202736
rect 675482 198328 675538 198384
rect 675758 195336 675814 195392
rect 675758 190340 675760 190360
rect 675760 190340 675812 190360
rect 675812 190340 675814 190360
rect 675758 190304 675814 190340
rect 674838 190168 674894 190224
rect 676034 178472 676090 178528
rect 676034 178084 676090 178120
rect 676034 178064 676036 178084
rect 676036 178064 676088 178084
rect 676088 178064 676090 178084
rect 675942 177656 675998 177712
rect 676034 177248 676090 177304
rect 676034 176840 676090 176896
rect 676034 176468 676036 176488
rect 676036 176468 676088 176488
rect 676088 176468 676090 176488
rect 676034 176432 676090 176468
rect 676034 176044 676090 176080
rect 676034 176024 676036 176044
rect 676036 176024 676088 176044
rect 676088 176024 676090 176044
rect 676034 175652 676036 175672
rect 676036 175652 676088 175672
rect 676088 175652 676090 175672
rect 676034 175616 676090 175652
rect 676034 175228 676090 175264
rect 676034 175208 676036 175228
rect 676036 175208 676088 175228
rect 676088 175208 676090 175228
rect 674746 174800 674802 174856
rect 676034 174412 676090 174448
rect 676034 174392 676036 174412
rect 676036 174392 676088 174412
rect 676088 174392 676090 174412
rect 678242 173984 678298 174040
rect 676034 173168 676090 173224
rect 676862 171536 676918 171592
rect 676034 170720 676090 170776
rect 676034 170332 676090 170368
rect 676034 170312 676036 170332
rect 676036 170312 676088 170332
rect 676088 170312 676090 170332
rect 676034 169516 676090 169552
rect 676034 169496 676036 169516
rect 676036 169496 676088 169516
rect 676088 169496 676090 169516
rect 676034 169108 676090 169144
rect 676034 169088 676036 169108
rect 676036 169088 676088 169108
rect 676088 169088 676090 169108
rect 676034 168700 676090 168736
rect 676034 168680 676036 168700
rect 676036 168680 676088 168700
rect 676088 168680 676090 168700
rect 676034 168292 676090 168328
rect 676034 168272 676036 168292
rect 676036 168272 676088 168292
rect 676088 168272 676090 168292
rect 676034 167884 676090 167920
rect 676034 167864 676036 167884
rect 676036 167864 676088 167884
rect 676088 167864 676090 167884
rect 676034 167068 676090 167104
rect 676034 167048 676036 167068
rect 676036 167048 676088 167068
rect 676088 167048 676090 167068
rect 676586 169904 676642 169960
rect 676586 166368 676642 166424
rect 676862 166368 676918 166424
rect 676218 162696 676274 162752
rect 681002 172352 681058 172408
rect 678426 171128 678482 171184
rect 678242 162560 678298 162616
rect 678426 162424 678482 162480
rect 681002 162288 681058 162344
rect 675758 159976 675814 160032
rect 675758 159432 675814 159488
rect 675758 157392 675814 157448
rect 675666 156984 675722 157040
rect 675574 156440 675630 156496
rect 675390 153040 675446 153096
rect 675758 151544 675814 151600
rect 675758 148416 675814 148472
rect 675758 146240 675814 146296
rect 676126 133048 676182 133104
rect 676034 132932 676090 132968
rect 676034 132912 676036 132932
rect 676036 132912 676088 132932
rect 676088 132912 676090 132932
rect 676218 132640 676274 132696
rect 676218 132268 676220 132288
rect 676220 132268 676272 132288
rect 676272 132268 676274 132288
rect 676218 132232 676274 132268
rect 676218 131416 676274 131472
rect 676034 131316 676036 131336
rect 676036 131316 676088 131336
rect 676088 131316 676090 131336
rect 676034 131280 676090 131316
rect 676218 130600 676274 130656
rect 676034 130500 676036 130520
rect 676036 130500 676088 130520
rect 676088 130500 676090 130520
rect 676034 130464 676090 130500
rect 676218 129804 676274 129840
rect 676218 129784 676220 129804
rect 676220 129784 676272 129804
rect 676272 129784 676274 129804
rect 676126 129376 676182 129432
rect 676218 128968 676274 129024
rect 683670 128152 683726 128208
rect 676034 128016 676090 128072
rect 683118 127336 683174 127392
rect 674746 123528 674802 123584
rect 676862 126928 676918 126984
rect 676402 125296 676458 125352
rect 676218 123664 676274 123720
rect 676218 122868 676274 122904
rect 676218 122848 676220 122868
rect 676220 122848 676272 122868
rect 676272 122848 676274 122868
rect 676126 122440 676182 122496
rect 676218 121624 676274 121680
rect 679622 125704 679678 125760
rect 678242 125296 678298 125352
rect 677598 124072 677654 124128
rect 676862 117952 676918 118008
rect 676402 117272 676458 117328
rect 683302 126112 683358 126168
rect 683118 124888 683174 124944
rect 679622 117136 679678 117192
rect 683670 121624 683726 121680
rect 675758 114144 675814 114200
rect 675758 112512 675814 112568
rect 675482 111696 675538 111752
rect 675114 108976 675170 109032
rect 675758 108160 675814 108216
rect 675482 104760 675538 104816
rect 675758 103128 675814 103184
rect 675758 101360 675814 101416
rect 664442 48456 664498 48512
rect 662418 47368 662474 47424
rect 661130 44784 661186 44840
rect 611358 41520 611414 41576
rect 609978 41384 610034 41440
rect 141698 40296 141754 40352
<< metal3 >>
rect 114782 1031568 115982 1031696
rect 114782 1030864 114809 1031568
rect 115953 1030864 115982 1031568
rect 113182 1030370 114382 1030482
rect 113182 1029666 113213 1030370
rect 114357 1029666 114382 1030370
rect 103145 1006498 103211 1006501
rect 103605 1006498 103671 1006501
rect 103145 1006496 103408 1006498
rect 103145 1006440 103150 1006496
rect 103206 1006440 103408 1006496
rect 103145 1006438 103408 1006440
rect 103605 1006496 103776 1006498
rect 103605 1006440 103610 1006496
rect 103666 1006440 103776 1006496
rect 103605 1006438 103776 1006440
rect 103145 1006435 103211 1006438
rect 103605 1006435 103671 1006438
rect 100661 1006362 100727 1006365
rect 104341 1006362 104407 1006365
rect 108849 1006362 108915 1006365
rect 100661 1006360 100924 1006362
rect 100661 1006304 100666 1006360
rect 100722 1006304 100924 1006360
rect 100661 1006302 100924 1006304
rect 104341 1006360 104604 1006362
rect 104341 1006304 104346 1006360
rect 104402 1006304 104604 1006360
rect 104341 1006302 104604 1006304
rect 108849 1006360 109112 1006362
rect 108849 1006304 108854 1006360
rect 108910 1006304 109112 1006360
rect 108849 1006302 109112 1006304
rect 100661 1006299 100727 1006302
rect 104341 1006299 104407 1006302
rect 108849 1006299 108915 1006302
rect 101949 1006226 102015 1006229
rect 104801 1006226 104867 1006229
rect 108481 1006226 108547 1006229
rect 101949 1006224 102212 1006226
rect 101949 1006168 101954 1006224
rect 102010 1006168 102212 1006224
rect 101949 1006166 102212 1006168
rect 104801 1006224 104972 1006226
rect 104801 1006168 104806 1006224
rect 104862 1006168 104972 1006224
rect 104801 1006166 104972 1006168
rect 108284 1006224 108547 1006226
rect 108284 1006168 108486 1006224
rect 108542 1006168 108547 1006224
rect 108284 1006166 108547 1006168
rect 101949 1006163 102015 1006166
rect 104801 1006163 104867 1006166
rect 108481 1006163 108547 1006166
rect 98269 1006090 98335 1006093
rect 99097 1006090 99163 1006093
rect 98072 1006088 98335 1006090
rect 98072 1006032 98274 1006088
rect 98330 1006032 98335 1006088
rect 98072 1006030 98335 1006032
rect 98532 1006030 98900 1006090
rect 99097 1006088 99268 1006090
rect 99097 1006032 99102 1006088
rect 99158 1006032 99268 1006088
rect 99097 1006030 99268 1006032
rect 98269 1006027 98335 1006030
rect 99097 1006027 99163 1006030
rect 103145 1004730 103211 1004733
rect 102948 1004728 103211 1004730
rect 102948 1004672 103150 1004728
rect 103206 1004672 103211 1004728
rect 102948 1004670 103211 1004672
rect 103145 1004667 103211 1004670
rect 106825 1002418 106891 1002421
rect 106628 1002416 106891 1002418
rect 106628 1002360 106830 1002416
rect 106886 1002360 106891 1002416
rect 106628 1002358 106891 1002360
rect 106825 1002355 106891 1002358
rect 100293 1002282 100359 1002285
rect 105997 1002282 106063 1002285
rect 100293 1002280 100556 1002282
rect 100293 1002224 100298 1002280
rect 100354 1002224 100556 1002280
rect 100293 1002222 100556 1002224
rect 105892 1002280 106063 1002282
rect 105892 1002224 106002 1002280
rect 106058 1002224 106063 1002280
rect 105892 1002222 106063 1002224
rect 100293 1002219 100359 1002222
rect 105997 1002219 106063 1002222
rect 108481 1002282 108547 1002285
rect 108481 1002280 108652 1002282
rect 108481 1002224 108486 1002280
rect 108542 1002224 108652 1002280
rect 108481 1002222 108652 1002224
rect 108481 1002219 108547 1002222
rect 99465 1002146 99531 1002149
rect 101489 1002146 101555 1002149
rect 105629 1002146 105695 1002149
rect 107653 1002146 107719 1002149
rect 99465 1002144 99728 1002146
rect 99465 1002088 99470 1002144
rect 99526 1002088 99728 1002144
rect 99465 1002086 99728 1002088
rect 101489 1002144 101752 1002146
rect 101489 1002088 101494 1002144
rect 101550 1002088 101752 1002144
rect 101489 1002086 101752 1002088
rect 105432 1002144 105695 1002146
rect 105432 1002088 105634 1002144
rect 105690 1002088 105695 1002144
rect 105432 1002086 105695 1002088
rect 107456 1002144 107719 1002146
rect 107456 1002088 107658 1002144
rect 107714 1002088 107719 1002144
rect 107456 1002086 107719 1002088
rect 99465 1002083 99531 1002086
rect 101489 1002083 101555 1002086
rect 105629 1002083 105695 1002086
rect 107653 1002083 107719 1002086
rect 99925 1002010 99991 1002013
rect 101121 1002010 101187 1002013
rect 102317 1002010 102383 1002013
rect 104341 1002010 104407 1002013
rect 106457 1002010 106523 1002013
rect 107193 1002010 107259 1002013
rect 108021 1002010 108087 1002013
rect 111793 1002010 111859 1002013
rect 99925 1002008 100096 1002010
rect 99925 1001952 99930 1002008
rect 99986 1001952 100096 1002008
rect 99925 1001950 100096 1001952
rect 101121 1002008 101292 1002010
rect 101121 1001952 101126 1002008
rect 101182 1001952 101292 1002008
rect 101121 1001950 101292 1001952
rect 102317 1002008 102580 1002010
rect 102317 1001952 102322 1002008
rect 102378 1001952 102580 1002008
rect 102317 1001950 102580 1001952
rect 104236 1002008 104407 1002010
rect 104236 1001952 104346 1002008
rect 104402 1001952 104407 1002008
rect 104236 1001950 104407 1001952
rect 106260 1002008 106523 1002010
rect 106260 1001952 106462 1002008
rect 106518 1001952 106523 1002008
rect 106260 1001950 106523 1001952
rect 107088 1002008 107259 1002010
rect 107088 1001952 107198 1002008
rect 107254 1001952 107259 1002008
rect 107088 1001950 107259 1001952
rect 107916 1002008 108087 1002010
rect 107916 1001952 108026 1002008
rect 108082 1001952 108087 1002008
rect 107916 1001950 108087 1001952
rect 109480 1002008 111859 1002010
rect 109480 1001952 111798 1002008
rect 111854 1001952 111859 1002008
rect 109480 1001950 111859 1001952
rect 99925 1001947 99991 1001950
rect 101121 1001947 101187 1001950
rect 102317 1001947 102383 1001950
rect 104341 1001947 104407 1001950
rect 106457 1001947 106523 1001950
rect 107193 1001947 107259 1001950
rect 108021 1001947 108087 1001950
rect 111793 1001947 111859 1001950
rect 85246 997188 85252 997252
rect 85316 997250 85322 997252
rect 94773 997250 94839 997253
rect 85316 997248 94839 997250
rect 85316 997192 94778 997248
rect 94834 997192 94839 997248
rect 85316 997190 94839 997192
rect 85316 997188 85322 997190
rect 94773 997187 94839 997190
rect 109861 997250 109927 997253
rect 112989 997250 113055 997253
rect 109861 997248 113055 997250
rect 109861 997192 109866 997248
rect 109922 997192 112994 997248
rect 113050 997192 113055 997248
rect 109861 997190 113055 997192
rect 109861 997187 109927 997190
rect 112989 997187 113055 997190
rect 84694 996916 84700 996980
rect 84764 996978 84770 996980
rect 94497 996978 94563 996981
rect 84764 996976 94563 996978
rect 84764 996920 94502 996976
rect 94558 996920 94563 996976
rect 84764 996918 94563 996920
rect 84764 996916 84770 996918
rect 94497 996915 94563 996918
rect 113182 996677 114382 1029666
rect 93117 995890 93183 995893
rect 82126 995888 93183 995890
rect 82126 995832 93122 995888
rect 93178 995832 93183 995888
rect 82126 995830 93183 995832
rect 80973 995754 81039 995757
rect 82126 995754 82186 995830
rect 93117 995827 93183 995830
rect 80973 995752 82186 995754
rect 80973 995696 80978 995752
rect 81034 995696 82186 995752
rect 80973 995694 82186 995696
rect 82353 995754 82419 995757
rect 92473 995754 92539 995757
rect 82353 995752 92539 995754
rect 82353 995696 82358 995752
rect 82414 995696 92478 995752
rect 92534 995696 92539 995752
rect 82353 995694 92539 995696
rect 80973 995691 81039 995694
rect 82353 995691 82419 995694
rect 92473 995691 92539 995694
rect 84653 995620 84719 995621
rect 85205 995620 85271 995621
rect 84653 995618 84700 995620
rect 84608 995616 84700 995618
rect 84608 995560 84658 995616
rect 84608 995558 84700 995560
rect 84653 995556 84700 995558
rect 84764 995556 84770 995620
rect 85205 995618 85252 995620
rect 85160 995616 85252 995618
rect 85160 995560 85210 995616
rect 85160 995558 85252 995560
rect 85205 995556 85252 995558
rect 85316 995556 85322 995620
rect 86033 995618 86099 995621
rect 93301 995618 93367 995621
rect 86033 995616 93367 995618
rect 86033 995560 86038 995616
rect 86094 995560 93306 995616
rect 93362 995560 93367 995616
rect 86033 995558 93367 995560
rect 84653 995555 84719 995556
rect 85205 995555 85271 995556
rect 86033 995555 86099 995558
rect 93301 995555 93367 995558
rect 113182 995573 113227 996677
rect 114331 995573 114382 996677
rect 113182 995502 114382 995573
rect 88885 995484 88951 995485
rect 88885 995482 88932 995484
rect 88840 995480 88932 995482
rect 88840 995424 88890 995480
rect 88840 995422 88932 995424
rect 88885 995420 88932 995422
rect 88996 995420 89002 995484
rect 88885 995419 88951 995420
rect 87505 995210 87571 995213
rect 98637 995210 98703 995213
rect 87505 995208 98703 995210
rect 87505 995152 87510 995208
rect 87566 995152 98642 995208
rect 98698 995152 98703 995208
rect 87505 995150 98703 995152
rect 87505 995147 87571 995150
rect 98637 995147 98703 995150
rect 114782 995083 115982 1030864
rect 166182 1031568 167382 1031696
rect 166182 1030864 166209 1031568
rect 167353 1030864 167382 1031568
rect 164582 1030370 165782 1030482
rect 164582 1029666 164613 1030370
rect 165757 1029666 165782 1030370
rect 154573 1007178 154639 1007181
rect 154573 1007176 154836 1007178
rect 154573 1007120 154578 1007176
rect 154634 1007120 154836 1007176
rect 154573 1007118 154836 1007120
rect 154573 1007115 154639 1007118
rect 154113 1006498 154179 1006501
rect 154113 1006496 154376 1006498
rect 154113 1006440 154118 1006496
rect 154174 1006440 154376 1006496
rect 154113 1006438 154376 1006440
rect 154113 1006435 154179 1006438
rect 156137 1006226 156203 1006229
rect 156137 1006224 156400 1006226
rect 156137 1006168 156142 1006224
rect 156198 1006168 156400 1006224
rect 156137 1006166 156400 1006168
rect 156137 1006163 156203 1006166
rect 149697 1006090 149763 1006093
rect 150433 1006090 150499 1006093
rect 151721 1006090 151787 1006093
rect 157425 1006090 157491 1006093
rect 159081 1006090 159147 1006093
rect 149500 1006088 149763 1006090
rect 149500 1006032 149702 1006088
rect 149758 1006032 149763 1006088
rect 149500 1006030 149763 1006032
rect 149868 1006030 150328 1006090
rect 150433 1006088 150696 1006090
rect 150433 1006032 150438 1006088
rect 150494 1006032 150696 1006088
rect 150433 1006030 150696 1006032
rect 151721 1006088 151892 1006090
rect 151721 1006032 151726 1006088
rect 151782 1006032 151892 1006088
rect 151721 1006030 151892 1006032
rect 157425 1006088 157596 1006090
rect 157425 1006032 157430 1006088
rect 157486 1006032 157596 1006088
rect 157425 1006030 157596 1006032
rect 158884 1006088 159147 1006090
rect 158884 1006032 159086 1006088
rect 159142 1006032 159147 1006088
rect 158884 1006030 159147 1006032
rect 149697 1006027 149763 1006030
rect 150433 1006027 150499 1006030
rect 151721 1006027 151787 1006030
rect 157425 1006027 157491 1006030
rect 159081 1006027 159147 1006030
rect 160645 1006090 160711 1006093
rect 160645 1006088 160908 1006090
rect 160645 1006032 160650 1006088
rect 160706 1006032 160908 1006088
rect 160645 1006030 160908 1006032
rect 160645 1006027 160711 1006030
rect 152549 1005410 152615 1005413
rect 152549 1005408 152720 1005410
rect 152549 1005352 152554 1005408
rect 152610 1005352 152720 1005408
rect 152549 1005350 152720 1005352
rect 152549 1005347 152615 1005350
rect 152917 1005002 152983 1005005
rect 160645 1005002 160711 1005005
rect 152917 1005000 153180 1005002
rect 152917 1004944 152922 1005000
rect 152978 1004944 153180 1005000
rect 152917 1004942 153180 1004944
rect 160540 1005000 160711 1005002
rect 160540 1004944 160650 1005000
rect 160706 1004944 160711 1005000
rect 160540 1004942 160711 1004944
rect 152917 1004939 152983 1004942
rect 160645 1004939 160711 1004942
rect 153745 1004866 153811 1004869
rect 159449 1004866 159515 1004869
rect 153745 1004864 153916 1004866
rect 153745 1004808 153750 1004864
rect 153806 1004808 153916 1004864
rect 153745 1004806 153916 1004808
rect 159252 1004864 159515 1004866
rect 159252 1004808 159454 1004864
rect 159510 1004808 159515 1004864
rect 159252 1004806 159515 1004808
rect 153745 1004803 153811 1004806
rect 159449 1004803 159515 1004806
rect 152089 1004730 152155 1004733
rect 153285 1004730 153351 1004733
rect 159817 1004730 159883 1004733
rect 160277 1004730 160343 1004733
rect 152089 1004728 152352 1004730
rect 152089 1004672 152094 1004728
rect 152150 1004672 152352 1004728
rect 152089 1004670 152352 1004672
rect 153285 1004728 153548 1004730
rect 153285 1004672 153290 1004728
rect 153346 1004672 153548 1004728
rect 153285 1004670 153548 1004672
rect 159712 1004728 159883 1004730
rect 159712 1004672 159822 1004728
rect 159878 1004672 159883 1004728
rect 159712 1004670 159883 1004672
rect 160080 1004728 160343 1004730
rect 160080 1004672 160282 1004728
rect 160338 1004672 160343 1004728
rect 160080 1004670 160343 1004672
rect 152089 1004667 152155 1004670
rect 153285 1004667 153351 1004670
rect 159817 1004667 159883 1004670
rect 160277 1004667 160343 1004670
rect 155769 1002146 155835 1002149
rect 157425 1002146 157491 1002149
rect 158253 1002146 158319 1002149
rect 155572 1002144 155835 1002146
rect 155572 1002088 155774 1002144
rect 155830 1002088 155835 1002144
rect 155572 1002086 155835 1002088
rect 157228 1002144 157491 1002146
rect 157228 1002088 157430 1002144
rect 157486 1002088 157491 1002144
rect 157228 1002086 157491 1002088
rect 158056 1002144 158319 1002146
rect 158056 1002088 158258 1002144
rect 158314 1002088 158319 1002144
rect 158056 1002086 158319 1002088
rect 155769 1002083 155835 1002086
rect 157425 1002083 157491 1002086
rect 158253 1002083 158319 1002086
rect 150893 1002010 150959 1002013
rect 151721 1002010 151787 1002013
rect 150893 1002008 151156 1002010
rect 150893 1001952 150898 1002008
rect 150954 1001952 151156 1002008
rect 150893 1001950 151156 1001952
rect 151524 1002008 151787 1002010
rect 151524 1001952 151726 1002008
rect 151782 1001952 151787 1002008
rect 151524 1001950 151787 1001952
rect 150893 1001947 150959 1001950
rect 151721 1001947 151787 1001950
rect 155769 1002010 155835 1002013
rect 156965 1002010 157031 1002013
rect 158621 1002010 158687 1002013
rect 155769 1002008 156032 1002010
rect 155769 1001952 155774 1002008
rect 155830 1001952 156032 1002008
rect 155769 1001950 156032 1001952
rect 156860 1002008 157031 1002010
rect 156860 1001952 156970 1002008
rect 157026 1001952 157031 1002008
rect 156860 1001950 157031 1001952
rect 158516 1002008 158687 1002010
rect 158516 1001952 158626 1002008
rect 158682 1001952 158687 1002008
rect 158516 1001950 158687 1001952
rect 155769 1001947 155835 1001950
rect 156965 1001947 157031 1001950
rect 158621 1001947 158687 1001950
rect 143993 1000650 144059 1000653
rect 148501 1000650 148567 1000653
rect 143993 1000648 148567 1000650
rect 143993 1000592 143998 1000648
rect 144054 1000592 148506 1000648
rect 148562 1000592 148567 1000648
rect 143993 1000590 148567 1000592
rect 143993 1000587 144059 1000590
rect 148501 1000587 148567 1000590
rect 162117 997386 162183 997389
rect 164417 997386 164483 997389
rect 162117 997384 164483 997386
rect 162117 997328 162122 997384
rect 162178 997328 164422 997384
rect 164478 997328 164483 997384
rect 162117 997326 164483 997328
rect 162117 997323 162183 997326
rect 164417 997323 164483 997326
rect 116117 997250 116183 997253
rect 143809 997250 143875 997253
rect 116117 997248 143875 997250
rect 116117 997192 116122 997248
rect 116178 997192 143814 997248
rect 143870 997192 143875 997248
rect 116117 997190 143875 997192
rect 116117 997187 116183 997190
rect 143809 997187 143875 997190
rect 116117 997114 116183 997117
rect 145649 997114 145715 997117
rect 116117 997112 145715 997114
rect 116117 997056 116122 997112
rect 116178 997056 145654 997112
rect 145710 997056 145715 997112
rect 116117 997054 145715 997056
rect 116117 997051 116183 997054
rect 145649 997051 145715 997054
rect 161105 997114 161171 997117
rect 164417 997114 164483 997117
rect 161105 997112 164483 997114
rect 161105 997056 161110 997112
rect 161166 997056 164422 997112
rect 164478 997056 164483 997112
rect 161105 997054 164483 997056
rect 161105 997051 161171 997054
rect 164417 997051 164483 997054
rect 164582 996677 165782 1029666
rect 136766 996100 136772 996164
rect 136836 996162 136842 996164
rect 146937 996162 147003 996165
rect 136836 996160 147003 996162
rect 136836 996104 146942 996160
rect 146998 996104 147003 996160
rect 136836 996102 147003 996104
rect 136836 996100 136842 996102
rect 146937 996099 147003 996102
rect 151077 995890 151143 995893
rect 132450 995888 151143 995890
rect 132450 995832 151082 995888
rect 151138 995832 151143 995888
rect 132450 995830 151143 995832
rect 129365 995754 129431 995757
rect 132450 995754 132510 995830
rect 151077 995827 151143 995830
rect 129365 995752 132510 995754
rect 129365 995696 129370 995752
rect 129426 995696 132510 995752
rect 129365 995694 132510 995696
rect 133137 995754 133203 995757
rect 144821 995754 144887 995757
rect 133137 995752 144887 995754
rect 133137 995696 133142 995752
rect 133198 995696 144826 995752
rect 144882 995696 144887 995752
rect 133137 995694 144887 995696
rect 129365 995691 129431 995694
rect 133137 995691 133203 995694
rect 144821 995691 144887 995694
rect 136541 995618 136607 995621
rect 148317 995618 148383 995621
rect 136541 995616 148383 995618
rect 136541 995560 136546 995616
rect 136602 995560 148322 995616
rect 148378 995560 148383 995616
rect 136541 995558 148383 995560
rect 136541 995555 136607 995558
rect 148317 995555 148383 995558
rect 130009 995482 130075 995485
rect 145557 995482 145623 995485
rect 130009 995480 145623 995482
rect 130009 995424 130014 995480
rect 130070 995424 145562 995480
rect 145618 995424 145623 995480
rect 130009 995422 145623 995424
rect 130009 995419 130075 995422
rect 145557 995419 145623 995422
rect 132125 995346 132191 995349
rect 151261 995346 151327 995349
rect 132125 995344 151327 995346
rect 132125 995288 132130 995344
rect 132186 995288 151266 995344
rect 151322 995288 151327 995344
rect 132125 995286 151327 995288
rect 132125 995283 132191 995286
rect 151261 995283 151327 995286
rect 131573 995210 131639 995213
rect 155174 995210 155234 996132
rect 164582 995573 164627 996677
rect 165731 995573 165782 996677
rect 164582 995502 165782 995573
rect 131573 995208 155234 995210
rect 131573 995152 131578 995208
rect 131634 995152 155234 995208
rect 131573 995150 155234 995152
rect 131573 995147 131639 995150
rect 80145 995074 80211 995077
rect 95877 995074 95943 995077
rect 80145 995072 95943 995074
rect 80145 995016 80150 995072
rect 80206 995016 95882 995072
rect 95938 995016 95943 995072
rect 80145 995014 95943 995016
rect 80145 995011 80211 995014
rect 95877 995011 95943 995014
rect 114782 993979 114845 995083
rect 115949 993979 115982 995083
rect 166182 995083 167382 1030864
rect 217582 1031568 218782 1031696
rect 217582 1030864 217609 1031568
rect 218753 1030864 218782 1031568
rect 215982 1030370 217182 1030482
rect 215982 1029666 216013 1030370
rect 217157 1029666 217182 1030370
rect 203885 1007042 203951 1007045
rect 203885 1007040 204148 1007042
rect 203885 1006984 203890 1007040
rect 203946 1006984 204148 1007040
rect 203885 1006982 204148 1006984
rect 203885 1006979 203951 1006982
rect 203517 1006634 203583 1006637
rect 203517 1006632 203780 1006634
rect 203517 1006576 203522 1006632
rect 203578 1006576 203780 1006632
rect 203517 1006574 203780 1006576
rect 203517 1006571 203583 1006574
rect 204713 1006362 204779 1006365
rect 204713 1006360 204976 1006362
rect 204713 1006304 204718 1006360
rect 204774 1006304 204976 1006360
rect 204713 1006302 204976 1006304
rect 204713 1006299 204779 1006302
rect 205541 1006226 205607 1006229
rect 205541 1006224 205804 1006226
rect 205541 1006168 205546 1006224
rect 205602 1006168 205804 1006224
rect 205541 1006166 205804 1006168
rect 205541 1006163 205607 1006166
rect 201033 1006090 201099 1006093
rect 201861 1006090 201927 1006093
rect 204345 1006090 204411 1006093
rect 208761 1006090 208827 1006093
rect 209589 1006090 209655 1006093
rect 215201 1006090 215267 1006093
rect 200836 1006088 201099 1006090
rect 200836 1006032 201038 1006088
rect 201094 1006032 201099 1006088
rect 200836 1006030 201099 1006032
rect 201296 1006030 201756 1006090
rect 201861 1006088 202124 1006090
rect 201861 1006032 201866 1006088
rect 201922 1006032 202124 1006088
rect 201861 1006030 202124 1006032
rect 204345 1006088 204516 1006090
rect 204345 1006032 204350 1006088
rect 204406 1006032 204516 1006088
rect 204345 1006030 204516 1006032
rect 208761 1006088 209024 1006090
rect 208761 1006032 208766 1006088
rect 208822 1006032 209024 1006088
rect 208761 1006030 209024 1006032
rect 209484 1006088 209655 1006090
rect 209484 1006032 209594 1006088
rect 209650 1006032 209655 1006088
rect 209484 1006030 209655 1006032
rect 212336 1006088 215267 1006090
rect 212336 1006032 215206 1006088
rect 215262 1006032 215267 1006088
rect 212336 1006030 215267 1006032
rect 201033 1006027 201099 1006030
rect 201861 1006027 201927 1006030
rect 204345 1006027 204411 1006030
rect 208761 1006027 208827 1006030
rect 209589 1006027 209655 1006030
rect 215201 1006027 215267 1006030
rect 208393 1004866 208459 1004869
rect 208196 1004864 208459 1004866
rect 208196 1004808 208398 1004864
rect 208454 1004808 208459 1004864
rect 208196 1004806 208459 1004808
rect 208393 1004803 208459 1004806
rect 202321 1004730 202387 1004733
rect 208761 1004730 208827 1004733
rect 202321 1004728 202492 1004730
rect 202321 1004672 202326 1004728
rect 202382 1004672 202492 1004728
rect 202321 1004670 202492 1004672
rect 208656 1004728 208827 1004730
rect 208656 1004672 208766 1004728
rect 208822 1004672 208827 1004728
rect 208656 1004670 208827 1004672
rect 202321 1004667 202387 1004670
rect 208761 1004667 208827 1004670
rect 207197 1002554 207263 1002557
rect 207197 1002552 207460 1002554
rect 207197 1002496 207202 1002552
rect 207258 1002496 207460 1002552
rect 207197 1002494 207460 1002496
rect 207197 1002491 207263 1002494
rect 210417 1002282 210483 1002285
rect 210220 1002280 210483 1002282
rect 210220 1002224 210422 1002280
rect 210478 1002224 210483 1002280
rect 210220 1002222 210483 1002224
rect 210417 1002219 210483 1002222
rect 205173 1002146 205239 1002149
rect 206737 1002146 206803 1002149
rect 210049 1002146 210115 1002149
rect 211245 1002146 211311 1002149
rect 205173 1002144 205344 1002146
rect 205173 1002088 205178 1002144
rect 205234 1002088 205344 1002144
rect 205173 1002086 205344 1002088
rect 206540 1002144 206803 1002146
rect 206540 1002088 206742 1002144
rect 206798 1002088 206803 1002144
rect 206540 1002086 206803 1002088
rect 209852 1002144 210115 1002146
rect 209852 1002088 210054 1002144
rect 210110 1002088 210115 1002144
rect 209852 1002086 210115 1002088
rect 211140 1002144 211311 1002146
rect 211140 1002088 211250 1002144
rect 211306 1002088 211311 1002144
rect 211140 1002086 211311 1002088
rect 205173 1002083 205239 1002086
rect 206737 1002083 206803 1002086
rect 210049 1002083 210115 1002086
rect 211245 1002083 211311 1002086
rect 202689 1002010 202755 1002013
rect 203057 1002010 203123 1002013
rect 205909 1002010 205975 1002013
rect 206737 1002010 206803 1002013
rect 207565 1002010 207631 1002013
rect 210877 1002010 210943 1002013
rect 211705 1002010 211771 1002013
rect 212073 1002010 212139 1002013
rect 202689 1002008 202952 1002010
rect 202689 1001952 202694 1002008
rect 202750 1001952 202952 1002008
rect 202689 1001950 202952 1001952
rect 203057 1002008 203320 1002010
rect 203057 1001952 203062 1002008
rect 203118 1001952 203320 1002008
rect 203057 1001950 203320 1001952
rect 205909 1002008 206172 1002010
rect 205909 1001952 205914 1002008
rect 205970 1001952 206172 1002008
rect 205909 1001950 206172 1001952
rect 206737 1002008 207000 1002010
rect 206737 1001952 206742 1002008
rect 206798 1001952 207000 1002008
rect 206737 1001950 207000 1001952
rect 207565 1002008 207828 1002010
rect 207565 1001952 207570 1002008
rect 207626 1001952 207828 1002008
rect 207565 1001950 207828 1001952
rect 210680 1002008 210943 1002010
rect 210680 1001952 210882 1002008
rect 210938 1001952 210943 1002008
rect 210680 1001950 210943 1001952
rect 211508 1002008 211771 1002010
rect 211508 1001952 211710 1002008
rect 211766 1001952 211771 1002008
rect 211508 1001950 211771 1001952
rect 211876 1002008 212139 1002010
rect 211876 1001952 212078 1002008
rect 212134 1001952 212139 1002008
rect 211876 1001950 212139 1001952
rect 202689 1001947 202755 1001950
rect 203057 1001947 203123 1001950
rect 205909 1001947 205975 1001950
rect 206737 1001947 206803 1001950
rect 207565 1001947 207631 1001950
rect 210877 1001947 210943 1001950
rect 211705 1001947 211771 1001950
rect 212073 1001947 212139 1001950
rect 195053 1001874 195119 1001877
rect 195237 1001874 195303 1001877
rect 195053 1001872 195303 1001874
rect 195053 1001816 195058 1001872
rect 195114 1001816 195242 1001872
rect 195298 1001816 195303 1001872
rect 195053 1001814 195303 1001816
rect 195053 1001811 195119 1001814
rect 195237 1001811 195303 1001814
rect 213361 997386 213427 997389
rect 215753 997386 215819 997389
rect 213361 997384 215819 997386
rect 213361 997328 213366 997384
rect 213422 997328 215758 997384
rect 215814 997328 215819 997384
rect 213361 997326 215819 997328
rect 213361 997323 213427 997326
rect 215753 997323 215819 997326
rect 167545 997250 167611 997253
rect 195237 997250 195303 997253
rect 167545 997248 195303 997250
rect 167545 997192 167550 997248
rect 167606 997192 195242 997248
rect 195298 997192 195303 997248
rect 167545 997190 195303 997192
rect 167545 997187 167611 997190
rect 195237 997187 195303 997190
rect 167545 997114 167611 997117
rect 200205 997114 200271 997117
rect 167545 997112 200271 997114
rect 167545 997056 167550 997112
rect 167606 997056 200210 997112
rect 200266 997056 200271 997112
rect 167545 997054 200271 997056
rect 167545 997051 167611 997054
rect 200205 997051 200271 997054
rect 215982 996677 217182 1029666
rect 184614 996374 186330 996434
rect 184614 995757 184674 996374
rect 186270 996298 186330 996374
rect 197353 996298 197419 996301
rect 186270 996296 197419 996298
rect 186270 996240 197358 996296
rect 197414 996240 197419 996296
rect 186270 996238 197419 996240
rect 197353 996235 197419 996238
rect 184614 995752 184723 995757
rect 184614 995696 184662 995752
rect 184718 995696 184723 995752
rect 184614 995694 184723 995696
rect 184657 995691 184723 995694
rect 188153 995754 188219 995757
rect 200757 995754 200823 995757
rect 188153 995752 200823 995754
rect 188153 995696 188158 995752
rect 188214 995696 200762 995752
rect 200818 995696 200823 995752
rect 188153 995694 200823 995696
rect 188153 995691 188219 995694
rect 200757 995691 200823 995694
rect 188797 995618 188863 995621
rect 195237 995618 195303 995621
rect 188797 995616 195303 995618
rect 188797 995560 188802 995616
rect 188858 995560 195242 995616
rect 195298 995560 195303 995616
rect 188797 995558 195303 995560
rect 188797 995555 188863 995558
rect 195237 995555 195303 995558
rect 215982 995573 216027 996677
rect 217131 995573 217182 996677
rect 215982 995502 217182 995573
rect 184473 995482 184539 995485
rect 195053 995482 195119 995485
rect 184473 995480 195119 995482
rect 184473 995424 184478 995480
rect 184534 995424 195058 995480
rect 195114 995424 195119 995480
rect 184473 995422 195119 995424
rect 184473 995419 184539 995422
rect 195053 995419 195119 995422
rect 187279 995346 187345 995349
rect 203517 995346 203583 995349
rect 187279 995344 203583 995346
rect 187279 995288 187284 995344
rect 187340 995288 203522 995344
rect 203578 995288 203583 995344
rect 187279 995286 203583 995288
rect 187279 995283 187345 995286
rect 203517 995283 203583 995286
rect 181115 995210 181181 995213
rect 202413 995210 202479 995213
rect 181115 995208 202479 995210
rect 181115 995152 181120 995208
rect 181176 995152 202418 995208
rect 202474 995152 202479 995208
rect 181115 995150 202479 995152
rect 181115 995147 181181 995150
rect 202413 995147 202479 995150
rect 136265 995074 136331 995077
rect 136766 995074 136772 995076
rect 136265 995072 136772 995074
rect 136265 995016 136270 995072
rect 136326 995016 136772 995072
rect 136265 995014 136772 995016
rect 136265 995011 136331 995014
rect 136766 995012 136772 995014
rect 136836 995012 136842 995076
rect 140129 995074 140195 995077
rect 165981 995074 166047 995077
rect 140129 995072 166047 995074
rect 140129 995016 140134 995072
rect 140190 995016 165986 995072
rect 166042 995016 166047 995072
rect 140129 995014 166047 995016
rect 140129 995011 140195 995014
rect 165981 995011 166047 995014
rect 114782 993858 115982 993979
rect 166182 993979 166245 995083
rect 167349 993979 167382 995083
rect 217582 995083 218782 1030864
rect 268982 1031568 270182 1031696
rect 268982 1030864 269009 1031568
rect 270153 1030864 270182 1031568
rect 267382 1030370 268582 1030482
rect 267382 1029666 267413 1030370
rect 268557 1029666 268582 1030370
rect 261017 1006906 261083 1006909
rect 260820 1006904 261083 1006906
rect 260820 1006848 261022 1006904
rect 261078 1006848 261083 1006904
rect 260820 1006846 261083 1006848
rect 261017 1006843 261083 1006846
rect 258165 1006362 258231 1006365
rect 258165 1006360 258428 1006362
rect 258165 1006304 258170 1006360
rect 258226 1006304 258428 1006360
rect 258165 1006302 258428 1006304
rect 258165 1006299 258231 1006302
rect 252461 1006226 252527 1006229
rect 252264 1006224 252527 1006226
rect 252264 1006168 252466 1006224
rect 252522 1006168 252527 1006224
rect 252264 1006166 252527 1006168
rect 252461 1006163 252527 1006166
rect 253289 1006226 253355 1006229
rect 256509 1006226 256575 1006229
rect 253289 1006224 253460 1006226
rect 253289 1006168 253294 1006224
rect 253350 1006168 253460 1006224
rect 253289 1006166 253460 1006168
rect 256509 1006224 256772 1006226
rect 256509 1006168 256514 1006224
rect 256570 1006168 256772 1006224
rect 256509 1006166 256772 1006168
rect 253289 1006163 253355 1006166
rect 256509 1006163 256575 1006166
rect 255313 1006090 255379 1006093
rect 258533 1006090 258599 1006093
rect 258993 1006090 259059 1006093
rect 262673 1006090 262739 1006093
rect 263041 1006090 263107 1006093
rect 252724 1006030 253092 1006090
rect 255313 1006088 255576 1006090
rect 255313 1006032 255318 1006088
rect 255374 1006032 255576 1006088
rect 255313 1006030 255576 1006032
rect 258533 1006088 258796 1006090
rect 258533 1006032 258538 1006088
rect 258594 1006032 258796 1006088
rect 258533 1006030 258796 1006032
rect 258993 1006088 259164 1006090
rect 258993 1006032 258998 1006088
rect 259054 1006032 259164 1006088
rect 258993 1006030 259164 1006032
rect 262476 1006088 262739 1006090
rect 262476 1006032 262678 1006088
rect 262734 1006032 262739 1006088
rect 262476 1006030 262739 1006032
rect 262844 1006088 263107 1006090
rect 262844 1006032 263046 1006088
rect 263102 1006032 263107 1006088
rect 262844 1006030 263107 1006032
rect 255313 1006027 255379 1006030
rect 258533 1006027 258599 1006030
rect 258993 1006027 259059 1006030
rect 262673 1006027 262739 1006030
rect 263041 1006027 263107 1006030
rect 253657 1002690 253723 1002693
rect 253657 1002688 253920 1002690
rect 253657 1002632 253662 1002688
rect 253718 1002632 253920 1002688
rect 253657 1002630 253920 1002632
rect 253657 1002627 253723 1002630
rect 254945 1002554 255011 1002557
rect 254945 1002552 255116 1002554
rect 254945 1002496 254950 1002552
rect 255006 1002496 255116 1002552
rect 254945 1002494 255116 1002496
rect 254945 1002491 255011 1002494
rect 260189 1002282 260255 1002285
rect 260084 1002280 260255 1002282
rect 260084 1002224 260194 1002280
rect 260250 1002224 260255 1002280
rect 260084 1002222 260255 1002224
rect 260189 1002219 260255 1002222
rect 255681 1002146 255747 1002149
rect 256141 1002146 256207 1002149
rect 261477 1002146 261543 1002149
rect 261845 1002146 261911 1002149
rect 255681 1002144 255944 1002146
rect 255681 1002088 255686 1002144
rect 255742 1002088 255944 1002144
rect 255681 1002086 255944 1002088
rect 256141 1002144 256404 1002146
rect 256141 1002088 256146 1002144
rect 256202 1002088 256404 1002144
rect 256141 1002086 256404 1002088
rect 261280 1002144 261543 1002146
rect 261280 1002088 261482 1002144
rect 261538 1002088 261543 1002144
rect 261280 1002086 261543 1002088
rect 261648 1002144 261911 1002146
rect 261648 1002088 261850 1002144
rect 261906 1002088 261911 1002144
rect 261648 1002086 261911 1002088
rect 255681 1002083 255747 1002086
rect 256141 1002083 256207 1002086
rect 261477 1002083 261543 1002086
rect 261845 1002083 261911 1002086
rect 254117 1002010 254183 1002013
rect 254485 1002010 254551 1002013
rect 256969 1002010 257035 1002013
rect 257797 1002010 257863 1002013
rect 259821 1002010 259887 1002013
rect 260649 1002010 260715 1002013
rect 254117 1002008 254380 1002010
rect 254117 1001952 254122 1002008
rect 254178 1001952 254380 1002008
rect 254117 1001950 254380 1001952
rect 254485 1002008 254748 1002010
rect 254485 1001952 254490 1002008
rect 254546 1001952 254748 1002008
rect 254485 1001950 254748 1001952
rect 256969 1002008 257140 1002010
rect 256969 1001952 256974 1002008
rect 257030 1001952 257140 1002008
rect 256969 1001950 257140 1001952
rect 257600 1002008 257863 1002010
rect 257600 1001952 257802 1002008
rect 257858 1001952 257863 1002008
rect 257600 1001950 257863 1001952
rect 259624 1002008 259887 1002010
rect 259624 1001952 259826 1002008
rect 259882 1001952 259887 1002008
rect 259624 1001950 259887 1001952
rect 260452 1002008 260715 1002010
rect 260452 1001952 260654 1002008
rect 260710 1001952 260715 1002008
rect 260452 1001950 260715 1001952
rect 254117 1001947 254183 1001950
rect 254485 1001947 254551 1001950
rect 256969 1001947 257035 1001950
rect 257797 1001947 257863 1001950
rect 259821 1001947 259887 1001950
rect 260649 1001947 260715 1001950
rect 261845 1002010 261911 1002013
rect 263501 1002010 263567 1002013
rect 266997 1002010 267063 1002013
rect 261845 1002008 262108 1002010
rect 261845 1001952 261850 1002008
rect 261906 1001952 262108 1002008
rect 261845 1001950 262108 1001952
rect 263304 1002008 263567 1002010
rect 263304 1001952 263506 1002008
rect 263562 1001952 263567 1002008
rect 263304 1001950 263567 1001952
rect 263764 1002008 267063 1002010
rect 263764 1001952 267002 1002008
rect 267058 1001952 267063 1002008
rect 263764 1001950 267063 1001952
rect 261845 1001947 261911 1001950
rect 263501 1001947 263567 1001950
rect 266997 1001947 267063 1001950
rect 218881 997250 218947 997253
rect 246573 997250 246639 997253
rect 218881 997248 246639 997250
rect 218881 997192 218886 997248
rect 218942 997192 246578 997248
rect 246634 997192 246639 997248
rect 218881 997190 246639 997192
rect 218881 997187 218947 997190
rect 246573 997187 246639 997190
rect 267382 996677 268582 1029666
rect 243854 996372 243860 996436
rect 243924 996434 243930 996436
rect 247677 996434 247743 996437
rect 243924 996432 247743 996434
rect 243924 996376 247682 996432
rect 247738 996376 247743 996432
rect 243924 996374 247743 996376
rect 243924 996372 243930 996374
rect 247677 996371 247743 996374
rect 250437 996162 250503 996165
rect 236870 996160 250503 996162
rect 236870 996104 250442 996160
rect 250498 996104 250503 996160
rect 236870 996102 250503 996104
rect 235257 995754 235323 995757
rect 236870 995754 236930 996102
rect 250437 996099 250503 996102
rect 250345 996026 250411 996029
rect 235257 995752 236930 995754
rect 235257 995696 235262 995752
rect 235318 995696 236930 995752
rect 235257 995694 236930 995696
rect 238710 996024 250411 996026
rect 238710 995968 250350 996024
rect 250406 995968 250411 996024
rect 238710 995966 250411 995968
rect 235257 995691 235323 995694
rect 232221 995618 232287 995621
rect 238710 995618 238770 995966
rect 250345 995963 250411 995966
rect 243813 995756 243879 995757
rect 243813 995754 243860 995756
rect 243768 995752 243860 995754
rect 243768 995696 243818 995752
rect 243768 995694 243860 995696
rect 243813 995692 243860 995694
rect 243924 995692 243930 995756
rect 243813 995691 243879 995692
rect 232221 995616 238770 995618
rect 232221 995560 232226 995616
rect 232282 995560 238770 995616
rect 232221 995558 238770 995560
rect 242065 995618 242131 995621
rect 249057 995618 249123 995621
rect 242065 995616 249123 995618
rect 242065 995560 242070 995616
rect 242126 995560 249062 995616
rect 249118 995560 249123 995616
rect 242065 995558 249123 995560
rect 232221 995555 232287 995558
rect 242065 995555 242131 995558
rect 249057 995555 249123 995558
rect 236545 995482 236611 995485
rect 247033 995482 247099 995485
rect 236545 995480 247099 995482
rect 236545 995424 236550 995480
rect 236606 995424 247038 995480
rect 247094 995424 247099 995480
rect 236545 995422 247099 995424
rect 236545 995419 236611 995422
rect 247033 995419 247099 995422
rect 238707 995346 238773 995349
rect 251357 995346 251423 995349
rect 238707 995344 251423 995346
rect 238707 995288 238712 995344
rect 238768 995288 251362 995344
rect 251418 995288 251423 995344
rect 238707 995286 251423 995288
rect 238707 995283 238773 995286
rect 251357 995283 251423 995286
rect 234613 995210 234679 995213
rect 257938 995210 257998 996132
rect 267382 995573 267427 996677
rect 268531 995573 268582 996677
rect 267382 995502 268582 995573
rect 234613 995208 257998 995210
rect 234613 995152 234618 995208
rect 234674 995152 257998 995208
rect 234613 995150 257998 995152
rect 234613 995147 234679 995150
rect 167545 995074 167611 995077
rect 186497 995074 186563 995077
rect 167545 995072 186563 995074
rect 167545 995016 167550 995072
rect 167606 995016 186502 995072
rect 186558 995016 186563 995072
rect 167545 995014 186563 995016
rect 167545 995011 167611 995014
rect 186497 995011 186563 995014
rect 191741 995074 191807 995077
rect 217409 995074 217475 995077
rect 191741 995072 217475 995074
rect 191741 995016 191746 995072
rect 191802 995016 217414 995072
rect 217470 995016 217475 995072
rect 191741 995014 217475 995016
rect 191741 995011 191807 995014
rect 217409 995011 217475 995014
rect 166182 993858 167382 993979
rect 217582 993979 217645 995083
rect 218749 993979 218782 995083
rect 268982 995083 270182 1030864
rect 320582 1031568 321782 1031696
rect 320582 1030864 320609 1031568
rect 321753 1030864 321782 1031568
rect 318982 1030370 320182 1030482
rect 318982 1029666 319013 1030370
rect 320157 1029666 320182 1030370
rect 308949 1007042 309015 1007045
rect 308949 1007040 309212 1007042
rect 308949 1006984 308954 1007040
rect 309010 1006984 309212 1007040
rect 308949 1006982 309212 1006984
rect 308949 1006979 309015 1006982
rect 308121 1006362 308187 1006365
rect 310145 1006362 310211 1006365
rect 308121 1006360 308384 1006362
rect 308121 1006304 308126 1006360
rect 308182 1006304 308384 1006360
rect 308121 1006302 308384 1006304
rect 310145 1006360 310408 1006362
rect 310145 1006304 310150 1006360
rect 310206 1006304 310408 1006360
rect 310145 1006302 310408 1006304
rect 308121 1006299 308187 1006302
rect 310145 1006299 310211 1006302
rect 306097 1006226 306163 1006229
rect 306097 1006224 306360 1006226
rect 306097 1006168 306102 1006224
rect 306158 1006168 306360 1006224
rect 306097 1006166 306360 1006168
rect 306097 1006163 306163 1006166
rect 304073 1006090 304139 1006093
rect 304901 1006090 304967 1006093
rect 305637 1006090 305703 1006093
rect 306465 1006090 306531 1006093
rect 310605 1006090 310671 1006093
rect 314653 1006090 314719 1006093
rect 303876 1006088 304139 1006090
rect 303876 1006032 304078 1006088
rect 304134 1006032 304139 1006088
rect 303876 1006030 304139 1006032
rect 304244 1006030 304704 1006090
rect 304901 1006088 305164 1006090
rect 304901 1006032 304906 1006088
rect 304962 1006032 305164 1006088
rect 304901 1006030 305164 1006032
rect 305637 1006088 305900 1006090
rect 305637 1006032 305642 1006088
rect 305698 1006032 305900 1006088
rect 305637 1006030 305900 1006032
rect 306465 1006088 306728 1006090
rect 306465 1006032 306470 1006088
rect 306526 1006032 306728 1006088
rect 306465 1006030 306728 1006032
rect 310605 1006088 310868 1006090
rect 310605 1006032 310610 1006088
rect 310666 1006032 310868 1006088
rect 310605 1006030 310868 1006032
rect 314548 1006088 314719 1006090
rect 314548 1006032 314658 1006088
rect 314714 1006032 314719 1006088
rect 314548 1006030 314719 1006032
rect 304073 1006027 304139 1006030
rect 304901 1006027 304967 1006030
rect 305637 1006027 305703 1006030
rect 306465 1006027 306531 1006030
rect 310605 1006027 310671 1006030
rect 314653 1006027 314719 1006030
rect 306925 1004866 306991 1004869
rect 307293 1004866 307359 1004869
rect 306925 1004864 307188 1004866
rect 306925 1004808 306930 1004864
rect 306986 1004808 307188 1004864
rect 306925 1004806 307188 1004808
rect 307293 1004864 307556 1004866
rect 307293 1004808 307298 1004864
rect 307354 1004808 307556 1004864
rect 307293 1004806 307556 1004808
rect 306925 1004803 306991 1004806
rect 307293 1004803 307359 1004806
rect 307753 1004730 307819 1004733
rect 308581 1004730 308647 1004733
rect 307753 1004728 307924 1004730
rect 307753 1004672 307758 1004728
rect 307814 1004672 307924 1004728
rect 307753 1004670 307924 1004672
rect 308581 1004728 308752 1004730
rect 308581 1004672 308586 1004728
rect 308642 1004672 308752 1004728
rect 308581 1004670 308752 1004672
rect 307753 1004667 307819 1004670
rect 308581 1004667 308647 1004670
rect 305269 1002010 305335 1002013
rect 310145 1002010 310211 1002013
rect 311433 1002010 311499 1002013
rect 305269 1002008 305532 1002010
rect 305269 1001952 305274 1002008
rect 305330 1001952 305532 1002008
rect 305269 1001950 305532 1001952
rect 309948 1002008 310211 1002010
rect 309948 1001952 310150 1002008
rect 310206 1001952 310211 1002008
rect 309948 1001950 310211 1001952
rect 311236 1002008 311499 1002010
rect 311236 1001952 311438 1002008
rect 311494 1001952 311499 1002008
rect 311236 1001950 311499 1001952
rect 305269 1001947 305335 1001950
rect 310145 1001947 310211 1001950
rect 311433 1001947 311499 1001950
rect 312169 997930 312235 997933
rect 313825 997930 313891 997933
rect 312064 997928 312235 997930
rect 312064 997872 312174 997928
rect 312230 997872 312235 997928
rect 312064 997870 312235 997872
rect 313628 997928 313891 997930
rect 313628 997872 313830 997928
rect 313886 997872 313891 997928
rect 313628 997870 313891 997872
rect 312169 997867 312235 997870
rect 313825 997867 313891 997870
rect 298093 997794 298159 997797
rect 303245 997794 303311 997797
rect 312997 997794 313063 997797
rect 315113 997794 315179 997797
rect 318057 997794 318123 997797
rect 298093 997792 303311 997794
rect 298093 997736 298098 997792
rect 298154 997736 303250 997792
rect 303306 997736 303311 997792
rect 298093 997734 303311 997736
rect 312892 997792 313063 997794
rect 312892 997736 313002 997792
rect 313058 997736 313063 997792
rect 312892 997734 313063 997736
rect 314916 997792 315179 997794
rect 314916 997736 315118 997792
rect 315174 997736 315179 997792
rect 314916 997734 315179 997736
rect 315284 997792 318123 997794
rect 315284 997736 318062 997792
rect 318118 997736 318123 997792
rect 315284 997734 318123 997736
rect 298093 997731 298159 997734
rect 303245 997731 303311 997734
rect 312997 997731 313063 997734
rect 315113 997731 315179 997734
rect 318057 997731 318123 997734
rect 270309 997250 270375 997253
rect 298369 997250 298435 997253
rect 270309 997248 298435 997250
rect 270309 997192 270314 997248
rect 270370 997192 298374 997248
rect 298430 997192 298435 997248
rect 270309 997190 298435 997192
rect 270309 997187 270375 997190
rect 298369 997187 298435 997190
rect 292430 997052 292436 997116
rect 292500 997114 292506 997116
rect 302877 997114 302943 997117
rect 292500 997112 302943 997114
rect 292500 997056 302882 997112
rect 302938 997056 302943 997112
rect 292500 997054 302943 997056
rect 292500 997052 292506 997054
rect 302877 997051 302943 997054
rect 318982 996677 320182 1029666
rect 288022 996374 291210 996434
rect 288022 995757 288082 996374
rect 291150 996298 291210 996374
rect 298737 996298 298803 996301
rect 291150 996296 298803 996298
rect 291150 996240 298742 996296
rect 298798 996240 298803 996296
rect 291150 996238 298803 996240
rect 298737 996235 298803 996238
rect 300117 995890 300183 995893
rect 293358 995888 300183 995890
rect 293358 995832 300122 995888
rect 300178 995832 300183 995888
rect 293358 995830 300183 995832
rect 287973 995752 288082 995757
rect 287973 995696 287978 995752
rect 288034 995696 288082 995752
rect 287973 995694 288082 995696
rect 291745 995754 291811 995757
rect 293358 995754 293418 995830
rect 300117 995827 300183 995830
rect 291745 995752 293418 995754
rect 291745 995696 291750 995752
rect 291806 995696 293418 995752
rect 291745 995694 293418 995696
rect 293585 995754 293651 995757
rect 304257 995754 304323 995757
rect 293585 995752 304323 995754
rect 293585 995696 293590 995752
rect 293646 995696 304262 995752
rect 304318 995696 304323 995752
rect 293585 995694 304323 995696
rect 287973 995691 288039 995694
rect 291745 995691 291811 995694
rect 293585 995691 293651 995694
rect 304257 995691 304323 995694
rect 291101 995618 291167 995621
rect 298921 995618 298987 995621
rect 291101 995616 298987 995618
rect 291101 995560 291106 995616
rect 291162 995560 298926 995616
rect 298982 995560 298987 995616
rect 291101 995558 298987 995560
rect 291101 995555 291167 995558
rect 298921 995555 298987 995558
rect 292389 995484 292455 995485
rect 292389 995482 292436 995484
rect 292344 995480 292436 995482
rect 292344 995424 292394 995480
rect 292344 995422 292436 995424
rect 292389 995420 292436 995422
rect 292500 995420 292506 995484
rect 295333 995482 295399 995485
rect 299013 995482 299079 995485
rect 295333 995480 299079 995482
rect 295333 995424 295338 995480
rect 295394 995424 299018 995480
rect 299074 995424 299079 995480
rect 295333 995422 299079 995424
rect 292389 995419 292455 995420
rect 295333 995419 295399 995422
rect 299013 995419 299079 995422
rect 290273 995346 290339 995349
rect 300301 995346 300367 995349
rect 290273 995344 300367 995346
rect 290273 995288 290278 995344
rect 290334 995288 300306 995344
rect 300362 995288 300367 995344
rect 290273 995286 300367 995288
rect 290273 995283 290339 995286
rect 300301 995283 300367 995286
rect 283465 995210 283531 995213
rect 298277 995210 298343 995213
rect 283465 995208 298343 995210
rect 283465 995152 283470 995208
rect 283526 995152 298282 995208
rect 298338 995152 298343 995208
rect 283465 995150 298343 995152
rect 283465 995147 283531 995150
rect 298277 995147 298343 995150
rect 218881 995074 218947 995077
rect 245653 995074 245719 995077
rect 218881 995072 245719 995074
rect 218881 995016 218886 995072
rect 218942 995016 245658 995072
rect 245714 995016 245719 995072
rect 218881 995014 245719 995016
rect 218881 995011 218947 995014
rect 245653 995011 245719 995014
rect 217582 993858 218782 993979
rect 268982 993979 269045 995083
rect 270149 993979 270182 995083
rect 285949 995074 286015 995077
rect 309550 995074 309610 996132
rect 318982 995573 319027 996677
rect 320131 995573 320182 996677
rect 318982 995502 320182 995573
rect 285949 995072 309610 995074
rect 285949 995016 285954 995072
rect 286010 995016 309610 995072
rect 285949 995014 309610 995016
rect 320582 995083 321782 1030864
rect 370982 1031568 372182 1031696
rect 370982 1030864 371009 1031568
rect 372153 1030864 372182 1031568
rect 369382 1030370 370582 1030482
rect 369382 1029666 369413 1030370
rect 370557 1029666 370582 1030370
rect 357341 1006226 357407 1006229
rect 361389 1006226 361455 1006229
rect 357144 1006224 357407 1006226
rect 357144 1006168 357346 1006224
rect 357402 1006168 357407 1006224
rect 357144 1006166 357407 1006168
rect 361192 1006224 361455 1006226
rect 361192 1006168 361394 1006224
rect 361450 1006168 361455 1006224
rect 361192 1006166 361455 1006168
rect 357341 1006163 357407 1006166
rect 361389 1006163 361455 1006166
rect 354489 1006090 354555 1006093
rect 355225 1006090 355291 1006093
rect 356053 1006090 356119 1006093
rect 358537 1006090 358603 1006093
rect 354292 1006088 354555 1006090
rect 354292 1006032 354494 1006088
rect 354550 1006032 354555 1006088
rect 354292 1006030 354555 1006032
rect 354660 1006030 355120 1006090
rect 355225 1006088 355488 1006090
rect 355225 1006032 355230 1006088
rect 355286 1006032 355488 1006088
rect 355225 1006030 355488 1006032
rect 355948 1006088 356119 1006090
rect 355948 1006032 356058 1006088
rect 356114 1006032 356119 1006088
rect 355948 1006030 356119 1006032
rect 358340 1006088 358603 1006090
rect 358340 1006032 358542 1006088
rect 358598 1006032 358603 1006088
rect 358340 1006030 358603 1006032
rect 354489 1006027 354555 1006030
rect 355225 1006027 355291 1006030
rect 356053 1006027 356119 1006030
rect 358537 1006027 358603 1006030
rect 360561 1005410 360627 1005413
rect 360364 1005408 360627 1005410
rect 360364 1005352 360566 1005408
rect 360622 1005352 360627 1005408
rect 360364 1005350 360627 1005352
rect 360561 1005347 360627 1005350
rect 356513 1005274 356579 1005277
rect 356316 1005272 356579 1005274
rect 356316 1005216 356518 1005272
rect 356574 1005216 356579 1005272
rect 356316 1005214 356579 1005216
rect 356513 1005211 356579 1005214
rect 361757 1004866 361823 1004869
rect 363413 1004866 363479 1004869
rect 361652 1004864 361823 1004866
rect 361652 1004808 361762 1004864
rect 361818 1004808 361823 1004864
rect 361652 1004806 361823 1004808
rect 363308 1004864 363479 1004866
rect 363308 1004808 363418 1004864
rect 363474 1004808 363479 1004864
rect 363308 1004806 363479 1004808
rect 361757 1004803 361823 1004806
rect 363413 1004803 363479 1004806
rect 362585 1004730 362651 1004733
rect 364241 1004730 364307 1004733
rect 362388 1004728 362651 1004730
rect 362388 1004672 362590 1004728
rect 362646 1004672 362651 1004728
rect 362388 1004670 362651 1004672
rect 364044 1004728 364307 1004730
rect 364044 1004672 364246 1004728
rect 364302 1004672 364307 1004728
rect 364044 1004670 364307 1004672
rect 362585 1004667 362651 1004670
rect 364241 1004667 364307 1004670
rect 356513 1004594 356579 1004597
rect 356513 1004592 356684 1004594
rect 356513 1004536 356518 1004592
rect 356574 1004536 356684 1004592
rect 356513 1004534 356684 1004536
rect 356513 1004531 356579 1004534
rect 358077 1003914 358143 1003917
rect 357972 1003912 358143 1003914
rect 357972 1003856 358082 1003912
rect 358138 1003856 358143 1003912
rect 357972 1003854 358143 1003856
rect 358077 1003851 358143 1003854
rect 357341 1002010 357407 1002013
rect 358537 1002010 358603 1002013
rect 358905 1002010 358971 1002013
rect 359365 1002010 359431 1002013
rect 360193 1002010 360259 1002013
rect 361021 1002010 361087 1002013
rect 365069 1002010 365135 1002013
rect 365437 1002010 365503 1002013
rect 369117 1002010 369183 1002013
rect 357341 1002008 357604 1002010
rect 357341 1001952 357346 1002008
rect 357402 1001952 357604 1002008
rect 357341 1001950 357604 1001952
rect 358537 1002008 358800 1002010
rect 358537 1001952 358542 1002008
rect 358598 1001952 358800 1002008
rect 358537 1001950 358800 1001952
rect 358905 1002008 359168 1002010
rect 358905 1001952 358910 1002008
rect 358966 1001952 359168 1002008
rect 358905 1001950 359168 1001952
rect 359365 1002008 359628 1002010
rect 359365 1001952 359370 1002008
rect 359426 1001952 359628 1002008
rect 359365 1001950 359628 1001952
rect 359996 1002008 360259 1002010
rect 359996 1001952 360198 1002008
rect 360254 1001952 360259 1002008
rect 359996 1001950 360259 1001952
rect 360824 1002008 361087 1002010
rect 360824 1001952 361026 1002008
rect 361082 1001952 361087 1002008
rect 360824 1001950 361087 1001952
rect 364872 1002008 365135 1002010
rect 364872 1001952 365074 1002008
rect 365130 1001952 365135 1002008
rect 364872 1001950 365135 1001952
rect 365332 1002008 365503 1002010
rect 365332 1001952 365442 1002008
rect 365498 1001952 365503 1002008
rect 365332 1001950 365503 1001952
rect 365700 1002008 369183 1002010
rect 365700 1001952 369122 1002008
rect 369178 1001952 369183 1002008
rect 365700 1001950 369183 1001952
rect 357341 1001947 357407 1001950
rect 358537 1001947 358603 1001950
rect 358905 1001947 358971 1001950
rect 359365 1001947 359431 1001950
rect 360193 1001947 360259 1001950
rect 361021 1001947 361087 1001950
rect 365069 1001947 365135 1001950
rect 365437 1001947 365503 1001950
rect 369117 1001947 369183 1001950
rect 366541 997386 366607 997389
rect 369209 997386 369275 997389
rect 366541 997384 369275 997386
rect 366541 997328 366546 997384
rect 366602 997328 369214 997384
rect 369270 997328 369275 997384
rect 366541 997326 369275 997328
rect 366541 997323 366607 997326
rect 369209 997323 369275 997326
rect 369382 996677 370582 1029666
rect 369382 995573 369427 996677
rect 370531 995573 370582 996677
rect 369382 995502 370582 995573
rect 363597 995482 363663 995485
rect 369209 995482 369275 995485
rect 363597 995480 369275 995482
rect 363597 995424 363602 995480
rect 363658 995424 369214 995480
rect 369270 995424 369275 995480
rect 363597 995422 369275 995424
rect 363597 995419 363663 995422
rect 369209 995419 369275 995422
rect 360193 995346 360259 995349
rect 370773 995346 370839 995349
rect 360193 995344 370839 995346
rect 360193 995288 360198 995344
rect 360254 995288 370778 995344
rect 370834 995288 370839 995344
rect 360193 995286 370839 995288
rect 360193 995283 360259 995286
rect 370773 995283 370839 995286
rect 362217 995210 362283 995213
rect 370773 995210 370839 995213
rect 362217 995208 370839 995210
rect 362217 995152 362222 995208
rect 362278 995152 370778 995208
rect 370834 995152 370839 995208
rect 362217 995150 370839 995152
rect 362217 995147 362283 995150
rect 370773 995147 370839 995150
rect 285949 995011 286015 995014
rect 268982 993858 270182 993979
rect 320582 993979 320645 995083
rect 321749 993979 321782 995083
rect 320582 993858 321782 993979
rect 370982 995083 372182 1030864
rect 438382 1031568 439582 1031696
rect 438382 1030864 438409 1031568
rect 439553 1030864 439582 1031568
rect 436782 1030370 437982 1030482
rect 436782 1029666 436813 1030370
rect 437957 1029666 437982 1030370
rect 426341 1006906 426407 1006909
rect 427169 1006906 427235 1006909
rect 426144 1006904 426407 1006906
rect 426144 1006848 426346 1006904
rect 426402 1006848 426407 1006904
rect 426144 1006846 426407 1006848
rect 426972 1006904 427235 1006906
rect 426972 1006848 427174 1006904
rect 427230 1006848 427235 1006904
rect 426972 1006846 427235 1006848
rect 426341 1006843 426407 1006846
rect 427169 1006843 427235 1006846
rect 425145 1006770 425211 1006773
rect 427537 1006770 427603 1006773
rect 424948 1006768 425211 1006770
rect 424948 1006712 425150 1006768
rect 425206 1006712 425211 1006768
rect 424948 1006710 425211 1006712
rect 427340 1006768 427603 1006770
rect 427340 1006712 427542 1006768
rect 427598 1006712 427603 1006768
rect 427340 1006710 427603 1006712
rect 425145 1006707 425211 1006710
rect 427537 1006707 427603 1006710
rect 427997 1006634 428063 1006637
rect 427800 1006632 428063 1006634
rect 427800 1006576 428002 1006632
rect 428058 1006576 428063 1006632
rect 427800 1006574 428063 1006576
rect 427997 1006571 428063 1006574
rect 423489 1006498 423555 1006501
rect 428365 1006498 428431 1006501
rect 423292 1006496 423555 1006498
rect 423292 1006440 423494 1006496
rect 423550 1006440 423555 1006496
rect 423292 1006438 423555 1006440
rect 428260 1006496 428431 1006498
rect 428260 1006440 428370 1006496
rect 428426 1006440 428431 1006496
rect 428260 1006438 428431 1006440
rect 423489 1006435 423555 1006438
rect 428365 1006435 428431 1006438
rect 423857 1006362 423923 1006365
rect 425973 1006362 426039 1006365
rect 423752 1006360 423923 1006362
rect 423752 1006304 423862 1006360
rect 423918 1006304 423923 1006360
rect 423752 1006302 423923 1006304
rect 425776 1006360 426039 1006362
rect 425776 1006304 425978 1006360
rect 426034 1006304 426039 1006360
rect 425776 1006302 426039 1006304
rect 423857 1006299 423923 1006302
rect 425973 1006299 426039 1006302
rect 424685 1006226 424751 1006229
rect 430021 1006226 430087 1006229
rect 424580 1006224 424751 1006226
rect 424580 1006168 424690 1006224
rect 424746 1006168 424751 1006224
rect 424580 1006166 424751 1006168
rect 429824 1006224 430087 1006226
rect 429824 1006168 430026 1006224
rect 430082 1006168 430087 1006224
rect 429824 1006166 430087 1006168
rect 424685 1006163 424751 1006166
rect 430021 1006163 430087 1006166
rect 422661 1006090 422727 1006093
rect 425513 1006090 425579 1006093
rect 422096 1006030 422556 1006090
rect 422661 1006088 422924 1006090
rect 422661 1006032 422666 1006088
rect 422722 1006032 422924 1006088
rect 422661 1006030 422924 1006032
rect 425316 1006088 425579 1006090
rect 425316 1006032 425518 1006088
rect 425574 1006032 425579 1006088
rect 425316 1006030 425579 1006032
rect 422661 1006027 422727 1006030
rect 425513 1006027 425579 1006030
rect 428825 1005410 428891 1005413
rect 432873 1005410 432939 1005413
rect 428628 1005408 428891 1005410
rect 428628 1005352 428830 1005408
rect 428886 1005352 428891 1005408
rect 428628 1005350 428891 1005352
rect 432676 1005408 432939 1005410
rect 432676 1005352 432878 1005408
rect 432934 1005352 432939 1005408
rect 432676 1005350 432939 1005352
rect 428825 1005347 428891 1005350
rect 432873 1005347 432939 1005350
rect 432505 1005274 432571 1005277
rect 432308 1005272 432571 1005274
rect 432308 1005216 432510 1005272
rect 432566 1005216 432571 1005272
rect 432308 1005214 432571 1005216
rect 432505 1005211 432571 1005214
rect 421465 1002010 421531 1002013
rect 424317 1002010 424383 1002013
rect 421465 1002008 421636 1002010
rect 421465 1001952 421470 1002008
rect 421526 1001952 421636 1002008
rect 421465 1001950 421636 1001952
rect 424120 1002008 424383 1002010
rect 424120 1001952 424322 1002008
rect 424378 1001952 424383 1002008
rect 424120 1001950 424383 1001952
rect 421465 1001947 421531 1001950
rect 424317 1001947 424383 1001950
rect 426341 1002010 426407 1002013
rect 426341 1002008 426604 1002010
rect 426341 1001952 426346 1002008
rect 426402 1001952 426604 1002008
rect 426341 1001950 426604 1001952
rect 426341 1001947 426407 1001950
rect 372337 998338 372403 998341
rect 383469 998338 383535 998341
rect 372337 998336 383535 998338
rect 372337 998280 372342 998336
rect 372398 998280 383474 998336
rect 383530 998280 383535 998336
rect 372337 998278 383535 998280
rect 372337 998275 372403 998278
rect 383469 998275 383535 998278
rect 430849 998202 430915 998205
rect 430652 998200 430915 998202
rect 430652 998144 430854 998200
rect 430910 998144 430915 998200
rect 430652 998142 430915 998144
rect 430849 998139 430915 998142
rect 429653 998066 429719 998069
rect 429456 998064 429719 998066
rect 429456 998008 429658 998064
rect 429714 998008 429719 998064
rect 429456 998006 429719 998008
rect 429653 998003 429719 998006
rect 430849 998066 430915 998069
rect 431677 998066 431743 998069
rect 430849 998064 431020 998066
rect 430849 998008 430854 998064
rect 430910 998008 431020 998064
rect 430849 998006 431020 998008
rect 431480 998064 431743 998066
rect 431480 998008 431682 998064
rect 431738 998008 431743 998064
rect 431480 998006 431743 998008
rect 430849 998003 430915 998006
rect 431677 998003 431743 998006
rect 429193 997930 429259 997933
rect 430389 997930 430455 997933
rect 432045 997930 432111 997933
rect 428996 997928 429259 997930
rect 428996 997872 429198 997928
rect 429254 997872 429259 997928
rect 428996 997870 429259 997872
rect 430284 997928 430455 997930
rect 430284 997872 430394 997928
rect 430450 997872 430455 997928
rect 430284 997870 430455 997872
rect 431940 997928 432111 997930
rect 431940 997872 432050 997928
rect 432106 997872 432111 997928
rect 431940 997870 432111 997872
rect 429193 997867 429259 997870
rect 430389 997867 430455 997870
rect 432045 997867 432111 997870
rect 383561 997794 383627 997797
rect 383694 997794 383700 997796
rect 383561 997792 383700 997794
rect 383561 997736 383566 997792
rect 383622 997736 383700 997792
rect 383561 997734 383700 997736
rect 383561 997731 383627 997734
rect 383694 997732 383700 997734
rect 383764 997732 383770 997796
rect 435357 997794 435423 997797
rect 433136 997792 435423 997794
rect 433136 997736 435362 997792
rect 435418 997736 435423 997792
rect 433136 997734 435423 997736
rect 435357 997731 435423 997734
rect 433977 997386 434043 997389
rect 436553 997386 436619 997389
rect 433977 997384 436619 997386
rect 433977 997328 433982 997384
rect 434038 997328 436558 997384
rect 436614 997328 436619 997384
rect 433977 997326 436619 997328
rect 433977 997323 434043 997326
rect 436553 997323 436619 997326
rect 372337 997250 372403 997253
rect 399937 997250 400003 997253
rect 372337 997248 400003 997250
rect 372337 997192 372342 997248
rect 372398 997192 399942 997248
rect 399998 997192 400003 997248
rect 372337 997190 400003 997192
rect 372337 997187 372403 997190
rect 399937 997187 400003 997190
rect 372337 996978 372403 996981
rect 400029 996978 400095 996981
rect 372337 996976 400095 996978
rect 372337 996920 372342 996976
rect 372398 996920 400034 996976
rect 400090 996920 400095 996976
rect 372337 996918 400095 996920
rect 372337 996915 372403 996918
rect 400029 996915 400095 996918
rect 436782 996677 437982 1029666
rect 372337 996298 372403 996301
rect 387558 996298 387564 996300
rect 372337 996296 387564 996298
rect 372337 996240 372342 996296
rect 372398 996240 387564 996296
rect 372337 996238 387564 996240
rect 372337 996235 372403 996238
rect 387558 996236 387564 996238
rect 387628 996236 387634 996300
rect 377397 996162 377463 996165
rect 390318 996162 390324 996164
rect 377397 996160 390324 996162
rect 377397 996104 377402 996160
rect 377458 996104 390324 996160
rect 377397 996102 390324 996104
rect 377397 996099 377463 996102
rect 390318 996100 390324 996102
rect 390388 996100 390394 996164
rect 383694 995964 383700 996028
rect 383764 996026 383770 996028
rect 383764 995966 389282 996026
rect 383764 995964 383770 995966
rect 374637 995890 374703 995893
rect 389030 995890 389036 995892
rect 374637 995888 389036 995890
rect 374637 995832 374642 995888
rect 374698 995832 389036 995888
rect 374637 995830 389036 995832
rect 374637 995827 374703 995830
rect 389030 995828 389036 995830
rect 389100 995828 389106 995892
rect 378317 995754 378383 995757
rect 388621 995754 388687 995757
rect 378317 995752 388687 995754
rect 378317 995696 378322 995752
rect 378378 995696 388626 995752
rect 388682 995696 388687 995752
rect 378317 995694 388687 995696
rect 389222 995754 389282 995966
rect 389398 995828 389404 995892
rect 389468 995890 389474 995892
rect 389468 995830 393330 995890
rect 389468 995828 389474 995830
rect 389357 995754 389423 995757
rect 389222 995752 389423 995754
rect 389222 995696 389362 995752
rect 389418 995696 389423 995752
rect 389222 995694 389423 995696
rect 378317 995691 378383 995694
rect 388621 995691 388687 995694
rect 389357 995691 389423 995694
rect 390318 995692 390324 995756
rect 390388 995754 390394 995756
rect 392393 995754 392459 995757
rect 390388 995752 392459 995754
rect 390388 995696 392398 995752
rect 392454 995696 392459 995752
rect 390388 995694 392459 995696
rect 393270 995754 393330 995830
rect 393405 995754 393471 995757
rect 393270 995752 393471 995754
rect 393270 995696 393410 995752
rect 393466 995696 393471 995752
rect 393270 995694 393471 995696
rect 390388 995692 390394 995694
rect 392393 995691 392459 995694
rect 393405 995691 393471 995694
rect 372429 995618 372495 995621
rect 391933 995618 391999 995621
rect 372429 995616 391999 995618
rect 372429 995560 372434 995616
rect 372490 995560 391938 995616
rect 391994 995560 391999 995616
rect 372429 995558 391999 995560
rect 372429 995555 372495 995558
rect 391933 995555 391999 995558
rect 436782 995573 436827 996677
rect 437931 995573 437982 996677
rect 436782 995502 437982 995573
rect 372337 995482 372403 995485
rect 396717 995482 396783 995485
rect 372337 995480 396783 995482
rect 372337 995424 372342 995480
rect 372398 995424 396722 995480
rect 396778 995424 396783 995480
rect 372337 995422 396783 995424
rect 372337 995419 372403 995422
rect 396717 995419 396783 995422
rect 372337 995346 372403 995349
rect 395153 995346 395219 995349
rect 372337 995344 395219 995346
rect 372337 995288 372342 995344
rect 372398 995288 395158 995344
rect 395214 995288 395219 995344
rect 372337 995286 395219 995288
rect 372337 995283 372403 995286
rect 395153 995283 395219 995286
rect 372337 995210 372403 995213
rect 387793 995210 387859 995213
rect 372337 995208 387859 995210
rect 372337 995152 372342 995208
rect 372398 995152 387798 995208
rect 387854 995152 387859 995208
rect 372337 995150 387859 995152
rect 372337 995147 372403 995150
rect 387793 995147 387859 995150
rect 370982 993979 371045 995083
rect 372149 993979 372182 995083
rect 438382 995083 439582 1030864
rect 515382 1031568 516582 1031696
rect 515382 1030864 515409 1031568
rect 516553 1030864 516582 1031568
rect 513782 1030370 514982 1030482
rect 513782 1029666 513813 1030370
rect 514957 1029666 514982 1030370
rect 508681 1006498 508747 1006501
rect 508484 1006496 508747 1006498
rect 508484 1006440 508686 1006496
rect 508742 1006440 508747 1006496
rect 508484 1006438 508747 1006440
rect 508681 1006435 508747 1006438
rect 501321 1006362 501387 1006365
rect 501124 1006360 501387 1006362
rect 501124 1006304 501326 1006360
rect 501382 1006304 501387 1006360
rect 501124 1006302 501387 1006304
rect 501321 1006299 501387 1006302
rect 505829 1006226 505895 1006229
rect 505632 1006224 505895 1006226
rect 505632 1006168 505834 1006224
rect 505890 1006168 505895 1006224
rect 505632 1006166 505895 1006168
rect 505829 1006163 505895 1006166
rect 499665 1006090 499731 1006093
rect 504541 1006090 504607 1006093
rect 505369 1006090 505435 1006093
rect 499100 1006030 499468 1006090
rect 499665 1006088 499928 1006090
rect 499665 1006032 499670 1006088
rect 499726 1006032 499928 1006088
rect 499665 1006030 499928 1006032
rect 504436 1006088 504607 1006090
rect 504436 1006032 504546 1006088
rect 504602 1006032 504607 1006088
rect 504436 1006030 504607 1006032
rect 505172 1006088 505435 1006090
rect 505172 1006032 505374 1006088
rect 505430 1006032 505435 1006088
rect 505172 1006030 505435 1006032
rect 499665 1006027 499731 1006030
rect 504541 1006027 504607 1006030
rect 505369 1006027 505435 1006030
rect 509877 1005410 509943 1005413
rect 509680 1005408 509943 1005410
rect 509680 1005352 509882 1005408
rect 509938 1005352 509943 1005408
rect 509680 1005350 509943 1005352
rect 509877 1005347 509943 1005350
rect 502885 1005274 502951 1005277
rect 502780 1005272 502951 1005274
rect 502780 1005216 502890 1005272
rect 502946 1005216 502951 1005272
rect 502780 1005214 502951 1005216
rect 502885 1005211 502951 1005214
rect 501689 1004866 501755 1004869
rect 501689 1004864 501952 1004866
rect 501689 1004808 501694 1004864
rect 501750 1004808 501952 1004864
rect 501689 1004806 501952 1004808
rect 501689 1004803 501755 1004806
rect 500493 1004730 500559 1004733
rect 500296 1004728 500559 1004730
rect 500296 1004672 500498 1004728
rect 500554 1004672 500559 1004728
rect 500296 1004670 500559 1004672
rect 500493 1004667 500559 1004670
rect 500493 1004594 500559 1004597
rect 501321 1004594 501387 1004597
rect 500493 1004592 500756 1004594
rect 500493 1004536 500498 1004592
rect 500554 1004536 500756 1004592
rect 500493 1004534 500756 1004536
rect 501321 1004592 501492 1004594
rect 501321 1004536 501326 1004592
rect 501382 1004536 501492 1004592
rect 501321 1004534 501492 1004536
rect 500493 1004531 500559 1004534
rect 501321 1004531 501387 1004534
rect 502517 1002146 502583 1002149
rect 502412 1002144 502583 1002146
rect 502412 1002088 502522 1002144
rect 502578 1002088 502583 1002144
rect 502412 1002086 502583 1002088
rect 502517 1002083 502583 1002086
rect 498469 1002010 498535 1002013
rect 502885 1002010 502951 1002013
rect 503345 1002010 503411 1002013
rect 505001 1002010 505067 1002013
rect 498469 1002008 498732 1002010
rect 498469 1001952 498474 1002008
rect 498530 1001952 498732 1002008
rect 498469 1001950 498732 1001952
rect 502885 1002008 503148 1002010
rect 502885 1001952 502890 1002008
rect 502946 1001952 503148 1002008
rect 502885 1001950 503148 1001952
rect 503345 1002008 503608 1002010
rect 503345 1001952 503350 1002008
rect 503406 1001952 503608 1002008
rect 503345 1001950 503608 1001952
rect 504804 1002008 505067 1002010
rect 504804 1001952 505006 1002008
rect 505062 1001952 505067 1002008
rect 504804 1001950 505067 1001952
rect 498469 1001947 498535 1001950
rect 502885 1001947 502951 1001950
rect 503345 1001947 503411 1001950
rect 505001 1001947 505067 1001950
rect 443637 998338 443703 998341
rect 472709 998338 472775 998341
rect 443637 998336 472775 998338
rect 443637 998280 443642 998336
rect 443698 998280 472714 998336
rect 472770 998280 472775 998336
rect 443637 998278 472775 998280
rect 443637 998275 443703 998278
rect 472709 998275 472775 998278
rect 507025 998066 507091 998069
rect 508221 998066 508287 998069
rect 506828 998064 507091 998066
rect 506828 998008 507030 998064
rect 507086 998008 507091 998064
rect 506828 998006 507091 998008
rect 508116 998064 508287 998066
rect 508116 998008 508226 998064
rect 508282 998008 508287 998064
rect 508116 998006 508287 998008
rect 507025 998003 507091 998006
rect 508221 998003 508287 998006
rect 506197 997930 506263 997933
rect 507853 997930 507919 997933
rect 509049 997930 509115 997933
rect 506000 997928 506263 997930
rect 506000 997872 506202 997928
rect 506258 997872 506263 997928
rect 506000 997870 506263 997872
rect 507656 997928 507919 997930
rect 507656 997872 507858 997928
rect 507914 997872 507919 997928
rect 507656 997870 507919 997872
rect 508852 997928 509115 997930
rect 508852 997872 509054 997928
rect 509110 997872 509115 997928
rect 508852 997870 509115 997872
rect 506197 997867 506263 997870
rect 507853 997867 507919 997870
rect 509049 997867 509115 997870
rect 506565 997794 506631 997797
rect 507393 997794 507459 997797
rect 509509 997794 509575 997797
rect 512637 997794 512703 997797
rect 506460 997792 506631 997794
rect 506460 997736 506570 997792
rect 506626 997736 506631 997792
rect 506460 997734 506631 997736
rect 507196 997792 507459 997794
rect 507196 997736 507398 997792
rect 507454 997736 507459 997792
rect 507196 997734 507459 997736
rect 509312 997792 509575 997794
rect 509312 997736 509514 997792
rect 509570 997736 509575 997792
rect 509312 997734 509575 997736
rect 510140 997792 512703 997794
rect 510140 997736 512642 997792
rect 512698 997736 512703 997792
rect 510140 997734 512703 997736
rect 506565 997731 506631 997734
rect 507393 997731 507459 997734
rect 509509 997731 509575 997734
rect 512637 997731 512703 997734
rect 439681 997250 439747 997253
rect 488901 997250 488967 997253
rect 439681 997248 488967 997250
rect 439681 997192 439686 997248
rect 439742 997192 488906 997248
rect 488962 997192 488967 997248
rect 439681 997190 488967 997192
rect 439681 997187 439747 997190
rect 488901 997187 488967 997190
rect 513782 996677 514982 1029666
rect 448605 996298 448671 996301
rect 448605 996296 480270 996298
rect 448605 996240 448610 996296
rect 448666 996240 480270 996296
rect 448605 996238 480270 996240
rect 448605 996235 448671 996238
rect 454677 996162 454743 996165
rect 454677 996160 470610 996162
rect 454677 996104 454682 996160
rect 454738 996104 470610 996160
rect 454677 996102 470610 996104
rect 454677 996099 454743 996102
rect 470550 995754 470610 996102
rect 480210 995890 480270 996238
rect 480210 995830 482570 995890
rect 481541 995754 481607 995757
rect 470550 995752 481607 995754
rect 470550 995696 481546 995752
rect 481602 995696 481607 995752
rect 470550 995694 481607 995696
rect 482510 995754 482570 995830
rect 482645 995754 482711 995757
rect 485589 995756 485655 995757
rect 485589 995754 485636 995756
rect 482510 995752 482711 995754
rect 482510 995696 482650 995752
rect 482706 995696 482711 995752
rect 482510 995694 482711 995696
rect 485544 995752 485636 995754
rect 485544 995696 485594 995752
rect 485544 995694 485636 995696
rect 481541 995691 481607 995694
rect 482645 995691 482711 995694
rect 485589 995692 485636 995694
rect 485700 995692 485706 995756
rect 485589 995691 485655 995692
rect 469857 995618 469923 995621
rect 483749 995618 483815 995621
rect 469857 995616 483815 995618
rect 469857 995560 469862 995616
rect 469918 995560 483754 995616
rect 483810 995560 483815 995616
rect 469857 995558 483815 995560
rect 469857 995555 469923 995558
rect 483749 995555 483815 995558
rect 451917 995482 451983 995485
rect 476941 995482 477007 995485
rect 451917 995480 477007 995482
rect 451917 995424 451922 995480
rect 451978 995424 476946 995480
rect 477002 995424 477007 995480
rect 451917 995422 477007 995424
rect 451917 995419 451983 995422
rect 476941 995419 477007 995422
rect 439681 995346 439747 995349
rect 478597 995346 478663 995349
rect 439681 995344 478663 995346
rect 439681 995288 439686 995344
rect 439742 995288 478602 995344
rect 478658 995288 478663 995344
rect 439681 995286 478663 995288
rect 503946 995346 504006 996132
rect 506422 995828 506428 995892
rect 506492 995890 506498 995892
rect 511073 995890 511139 995893
rect 506492 995888 511139 995890
rect 506492 995832 511078 995888
rect 511134 995832 511139 995888
rect 506492 995830 511139 995832
rect 506492 995828 506498 995830
rect 511073 995827 511139 995830
rect 513782 995573 513827 996677
rect 514931 995573 514982 996677
rect 513782 995502 514982 995573
rect 515213 995346 515279 995349
rect 503946 995344 515279 995346
rect 503946 995288 515218 995344
rect 515274 995288 515279 995344
rect 503946 995286 515279 995288
rect 439681 995283 439747 995286
rect 478597 995283 478663 995286
rect 515213 995283 515279 995286
rect 440877 995210 440943 995213
rect 481081 995210 481147 995213
rect 440877 995208 481147 995210
rect 440877 995152 440882 995208
rect 440938 995152 481086 995208
rect 481142 995152 481147 995208
rect 440877 995150 481147 995152
rect 440877 995147 440943 995150
rect 481081 995147 481147 995150
rect 500953 995210 501019 995213
rect 515213 995210 515279 995213
rect 500953 995208 515279 995210
rect 500953 995152 500958 995208
rect 501014 995152 515218 995208
rect 515274 995152 515279 995208
rect 500953 995150 515279 995152
rect 500953 995147 501019 995150
rect 515213 995147 515279 995150
rect 387558 995012 387564 995076
rect 387628 995074 387634 995076
rect 388069 995074 388135 995077
rect 387628 995072 388135 995074
rect 387628 995016 388074 995072
rect 388130 995016 388135 995072
rect 387628 995014 388135 995016
rect 387628 995012 387634 995014
rect 388069 995011 388135 995014
rect 370982 993858 372182 993979
rect 438382 993979 438445 995083
rect 439549 993979 439582 995083
rect 515382 995083 516582 1030864
rect 566782 1031568 567982 1031696
rect 566782 1030864 566809 1031568
rect 567953 1030864 567982 1031568
rect 565182 1030370 566382 1030482
rect 565182 1029666 565213 1030370
rect 566357 1029666 566382 1030370
rect 551921 1006362 551987 1006365
rect 553945 1006362 554011 1006365
rect 551724 1006360 551987 1006362
rect 551724 1006304 551926 1006360
rect 551982 1006304 551987 1006360
rect 551724 1006302 551987 1006304
rect 553748 1006360 554011 1006362
rect 553748 1006304 553950 1006360
rect 554006 1006304 554011 1006360
rect 553748 1006302 554011 1006304
rect 551921 1006299 551987 1006302
rect 553945 1006299 554011 1006302
rect 555969 1006226 556035 1006229
rect 557165 1006226 557231 1006229
rect 555772 1006224 556035 1006226
rect 555772 1006168 555974 1006224
rect 556030 1006168 556035 1006224
rect 555772 1006166 556035 1006168
rect 557060 1006224 557231 1006226
rect 557060 1006168 557170 1006224
rect 557226 1006168 557231 1006224
rect 557060 1006166 557231 1006168
rect 555969 1006163 556035 1006166
rect 557165 1006163 557231 1006166
rect 550265 1006090 550331 1006093
rect 551093 1006090 551159 1006093
rect 553117 1006090 553183 1006093
rect 556797 1006090 556863 1006093
rect 564341 1006090 564407 1006093
rect 550068 1006088 550331 1006090
rect 550068 1006032 550270 1006088
rect 550326 1006032 550331 1006088
rect 550068 1006030 550331 1006032
rect 550436 1006030 550896 1006090
rect 551093 1006088 551356 1006090
rect 551093 1006032 551098 1006088
rect 551154 1006032 551356 1006088
rect 551093 1006030 551356 1006032
rect 552920 1006088 553183 1006090
rect 552920 1006032 553122 1006088
rect 553178 1006032 553183 1006088
rect 552920 1006030 553183 1006032
rect 556600 1006088 556863 1006090
rect 556600 1006032 556802 1006088
rect 556858 1006032 556863 1006088
rect 556600 1006030 556863 1006032
rect 561476 1006088 564407 1006090
rect 561476 1006032 564346 1006088
rect 564402 1006032 564407 1006088
rect 561476 1006030 564407 1006032
rect 550265 1006027 550331 1006030
rect 551093 1006027 551159 1006030
rect 553117 1006027 553183 1006030
rect 556797 1006027 556863 1006030
rect 564341 1006027 564407 1006030
rect 556337 1004730 556403 1004733
rect 557625 1004730 557691 1004733
rect 556232 1004728 556403 1004730
rect 556232 1004672 556342 1004728
rect 556398 1004672 556403 1004728
rect 556232 1004670 556403 1004672
rect 557428 1004728 557691 1004730
rect 557428 1004672 557630 1004728
rect 557686 1004672 557691 1004728
rect 557428 1004670 557691 1004672
rect 556337 1004667 556403 1004670
rect 557625 1004667 557691 1004670
rect 552749 1002690 552815 1002693
rect 552552 1002688 552815 1002690
rect 552552 1002632 552754 1002688
rect 552810 1002632 552815 1002688
rect 552552 1002630 552815 1002632
rect 552749 1002627 552815 1002630
rect 552289 1002554 552355 1002557
rect 552092 1002552 552355 1002554
rect 552092 1002496 552294 1002552
rect 552350 1002496 552355 1002552
rect 552092 1002494 552355 1002496
rect 552289 1002491 552355 1002494
rect 559189 1002282 559255 1002285
rect 559649 1002282 559715 1002285
rect 559084 1002280 559255 1002282
rect 559084 1002224 559194 1002280
rect 559250 1002224 559255 1002280
rect 559084 1002222 559255 1002224
rect 559452 1002280 559715 1002282
rect 559452 1002224 559654 1002280
rect 559710 1002224 559715 1002280
rect 559452 1002222 559715 1002224
rect 559189 1002219 559255 1002222
rect 559649 1002219 559715 1002222
rect 554773 1002146 554839 1002149
rect 558453 1002146 558519 1002149
rect 560017 1002146 560083 1002149
rect 561305 1002146 561371 1002149
rect 554773 1002144 555036 1002146
rect 554773 1002088 554778 1002144
rect 554834 1002088 555036 1002144
rect 554773 1002086 555036 1002088
rect 558256 1002144 558519 1002146
rect 558256 1002088 558458 1002144
rect 558514 1002088 558519 1002144
rect 558256 1002086 558519 1002088
rect 559820 1002144 560083 1002146
rect 559820 1002088 560022 1002144
rect 560078 1002088 560083 1002144
rect 559820 1002086 560083 1002088
rect 561108 1002144 561371 1002146
rect 561108 1002088 561310 1002144
rect 561366 1002088 561371 1002144
rect 561108 1002086 561371 1002088
rect 554773 1002083 554839 1002086
rect 558453 1002083 558519 1002086
rect 560017 1002083 560083 1002086
rect 561305 1002083 561371 1002086
rect 553117 1002010 553183 1002013
rect 553945 1002010 554011 1002013
rect 554313 1002010 554379 1002013
rect 555141 1002010 555207 1002013
rect 557993 1002010 558059 1002013
rect 558821 1002010 558887 1002013
rect 560477 1002010 560543 1002013
rect 560845 1002010 560911 1002013
rect 553117 1002008 553380 1002010
rect 553117 1001952 553122 1002008
rect 553178 1001952 553380 1002008
rect 553117 1001950 553380 1001952
rect 553945 1002008 554116 1002010
rect 553945 1001952 553950 1002008
rect 554006 1001952 554116 1002008
rect 553945 1001950 554116 1001952
rect 554313 1002008 554576 1002010
rect 554313 1001952 554318 1002008
rect 554374 1001952 554576 1002008
rect 554313 1001950 554576 1001952
rect 555141 1002008 555404 1002010
rect 555141 1001952 555146 1002008
rect 555202 1001952 555404 1002008
rect 555141 1001950 555404 1001952
rect 557796 1002008 558059 1002010
rect 557796 1001952 557998 1002008
rect 558054 1001952 558059 1002008
rect 557796 1001950 558059 1001952
rect 558624 1002008 558887 1002010
rect 558624 1001952 558826 1002008
rect 558882 1001952 558887 1002008
rect 558624 1001950 558887 1001952
rect 560280 1002008 560543 1002010
rect 560280 1001952 560482 1002008
rect 560538 1001952 560543 1002008
rect 560280 1001950 560543 1001952
rect 560740 1002008 560911 1002010
rect 560740 1001952 560850 1002008
rect 560906 1001952 560911 1002008
rect 560740 1001950 560911 1001952
rect 553117 1001947 553183 1001950
rect 553945 1001947 554011 1001950
rect 554313 1001947 554379 1001950
rect 555141 1001947 555207 1001950
rect 557993 1001947 558059 1001950
rect 558821 1001947 558887 1001950
rect 560477 1001947 560543 1001950
rect 560845 1001947 560911 1001950
rect 517973 998474 518039 998477
rect 523953 998474 524019 998477
rect 517973 998472 524019 998474
rect 517973 998416 517978 998472
rect 518034 998416 523958 998472
rect 524014 998416 524019 998472
rect 517973 998414 524019 998416
rect 517973 998411 518039 998414
rect 523953 998411 524019 998414
rect 516685 998338 516751 998341
rect 524045 998338 524111 998341
rect 516685 998336 524111 998338
rect 516685 998280 516690 998336
rect 516746 998280 524050 998336
rect 524106 998280 524111 998336
rect 516685 998278 524111 998280
rect 516685 998275 516751 998278
rect 524045 998275 524111 998278
rect 561673 997386 561739 997389
rect 564985 997386 565051 997389
rect 561673 997384 565051 997386
rect 561673 997328 561678 997384
rect 561734 997328 564990 997384
rect 565046 997328 565051 997384
rect 561673 997326 565051 997328
rect 561673 997323 561739 997326
rect 564985 997323 565051 997326
rect 516685 997250 516751 997253
rect 540881 997250 540947 997253
rect 516685 997248 540947 997250
rect 516685 997192 516690 997248
rect 516746 997192 540886 997248
rect 540942 997192 540947 997248
rect 516685 997190 540947 997192
rect 516685 997187 516751 997190
rect 540881 997187 540947 997190
rect 561673 996978 561739 996981
rect 564985 996978 565051 996981
rect 561673 996976 565051 996978
rect 561673 996920 561678 996976
rect 561734 996920 564990 996976
rect 565046 996920 565051 996976
rect 561673 996918 565051 996920
rect 561673 996915 561739 996918
rect 564985 996915 565051 996918
rect 565182 996677 566382 1029666
rect 523953 996434 524019 996437
rect 523953 996432 526178 996434
rect 523953 996376 523958 996432
rect 524014 996376 526178 996432
rect 523953 996374 526178 996376
rect 523953 996371 524019 996374
rect 526118 995757 526178 996374
rect 516685 995754 516751 995757
rect 525333 995754 525399 995757
rect 516685 995752 525399 995754
rect 516685 995696 516690 995752
rect 516746 995696 525338 995752
rect 525394 995696 525399 995752
rect 516685 995694 525399 995696
rect 526118 995752 526227 995757
rect 526118 995696 526166 995752
rect 526222 995696 526227 995752
rect 526118 995694 526227 995696
rect 516685 995691 516751 995694
rect 525333 995691 525399 995694
rect 526161 995691 526227 995694
rect 516685 995618 516751 995621
rect 529013 995618 529079 995621
rect 516685 995616 529079 995618
rect 516685 995560 516690 995616
rect 516746 995560 529018 995616
rect 529074 995560 529079 995616
rect 516685 995558 529079 995560
rect 516685 995555 516751 995558
rect 529013 995555 529079 995558
rect 565182 995573 565227 996677
rect 566331 995573 566382 996677
rect 565182 995502 566382 995573
rect 516685 995482 516751 995485
rect 538949 995482 539015 995485
rect 516685 995480 539015 995482
rect 516685 995424 516690 995480
rect 516746 995424 538954 995480
rect 539010 995424 539015 995480
rect 516685 995422 539015 995424
rect 516685 995419 516751 995422
rect 538949 995419 539015 995422
rect 516685 995346 516751 995349
rect 532141 995346 532207 995349
rect 516685 995344 532207 995346
rect 516685 995288 516690 995344
rect 516746 995288 532146 995344
rect 532202 995288 532207 995344
rect 516685 995286 532207 995288
rect 516685 995283 516751 995286
rect 532141 995283 532207 995286
rect 516685 995210 516751 995213
rect 532601 995210 532667 995213
rect 516685 995208 532667 995210
rect 516685 995152 516690 995208
rect 516746 995152 532606 995208
rect 532662 995152 532667 995208
rect 516685 995150 532667 995152
rect 516685 995147 516751 995150
rect 532601 995147 532667 995150
rect 446305 995074 446371 995077
rect 487797 995074 487863 995077
rect 446305 995072 487863 995074
rect 446305 995016 446310 995072
rect 446366 995016 487802 995072
rect 487858 995016 487863 995072
rect 446305 995014 487863 995016
rect 446305 995011 446371 995014
rect 487797 995011 487863 995014
rect 438382 993858 439582 993979
rect 515382 993979 515445 995083
rect 516549 993979 516582 995083
rect 515382 993858 516582 993979
rect 566782 995083 567982 1030864
rect 568113 997250 568179 997253
rect 575197 997250 575263 997253
rect 568113 997248 575263 997250
rect 568113 997192 568118 997248
rect 568174 997192 575202 997248
rect 575258 997192 575263 997248
rect 568113 997190 575263 997192
rect 568113 997187 568179 997190
rect 575197 997187 575263 997190
rect 575700 997067 580479 997678
rect 580901 997250 580967 997253
rect 585133 997250 585199 997253
rect 580901 997248 585199 997250
rect 580901 997192 580906 997248
rect 580962 997192 585138 997248
rect 585194 997192 585199 997248
rect 580901 997190 585199 997192
rect 580901 997187 580967 997190
rect 585133 997187 585199 997190
rect 568113 996842 568179 996845
rect 575473 996842 575539 996845
rect 568113 996840 575539 996842
rect 568113 996784 568118 996840
rect 568174 996784 575478 996840
rect 575534 996784 575539 996840
rect 568113 996782 575539 996784
rect 568113 996779 568179 996782
rect 575473 996779 575539 996782
rect 566782 993979 566845 995083
rect 567949 993979 567982 995083
rect 575700 995123 575774 997067
rect 580398 995123 580479 997067
rect 585678 997073 590458 997678
rect 590929 997250 590995 997253
rect 590929 997248 605850 997250
rect 590929 997192 590934 997248
rect 590990 997192 605850 997248
rect 590929 997190 605850 997192
rect 590929 997187 590995 997190
rect 580717 996842 580783 996845
rect 585501 996842 585567 996845
rect 580717 996840 585567 996842
rect 580717 996784 580722 996840
rect 580778 996784 585506 996840
rect 585562 996784 585567 996840
rect 580717 996782 585567 996784
rect 580717 996779 580783 996782
rect 585501 996779 585567 996782
rect 575700 995032 580479 995123
rect 585678 995129 585744 997073
rect 590368 995129 590458 997073
rect 605790 997114 605850 997190
rect 605790 997054 634830 997114
rect 590561 996842 590627 996845
rect 590561 996840 634002 996842
rect 590561 996784 590566 996840
rect 590622 996784 634002 996840
rect 590561 996782 634002 996784
rect 590561 996779 590627 996782
rect 623681 996706 623747 996709
rect 625889 996706 625955 996709
rect 623681 996704 625955 996706
rect 623681 996648 623686 996704
rect 623742 996648 625894 996704
rect 625950 996648 625955 996704
rect 623681 996646 625955 996648
rect 623681 996643 623747 996646
rect 625889 996643 625955 996646
rect 605925 996298 605991 996301
rect 605925 996296 625170 996298
rect 605925 996240 605930 996296
rect 605986 996240 625170 996296
rect 605925 996238 625170 996240
rect 605925 996235 605991 996238
rect 625110 995618 625170 996238
rect 633942 995757 634002 996782
rect 634770 996434 634830 997054
rect 634770 996374 640810 996434
rect 640750 995757 640810 996374
rect 633942 995752 634051 995757
rect 633942 995696 633990 995752
rect 634046 995696 634051 995752
rect 633942 995694 634051 995696
rect 640750 995752 640859 995757
rect 640750 995696 640798 995752
rect 640854 995696 640859 995752
rect 640750 995694 640859 995696
rect 633985 995691 634051 995694
rect 640793 995691 640859 995694
rect 635181 995618 635247 995621
rect 625110 995616 635247 995618
rect 625110 995560 635186 995616
rect 635242 995560 635247 995616
rect 625110 995558 635247 995560
rect 635181 995555 635247 995558
rect 585678 995032 590458 995129
rect 622393 995074 622459 995077
rect 629661 995074 629727 995077
rect 622393 995072 629727 995074
rect 622393 995016 622398 995072
rect 622454 995016 629666 995072
rect 629722 995016 629727 995072
rect 622393 995014 629727 995016
rect 622393 995011 622459 995014
rect 629661 995011 629727 995014
rect 638953 994938 639019 994941
rect 640793 994938 640859 994941
rect 638953 994936 640859 994938
rect 638953 994880 638958 994936
rect 639014 994880 640798 994936
rect 640854 994880 640859 994936
rect 638953 994878 640859 994880
rect 638953 994875 639019 994878
rect 640793 994875 640859 994878
rect 566782 993858 567982 993979
rect 114502 990932 114508 990996
rect 114572 990994 114578 990996
rect 122097 990994 122163 990997
rect 114572 990992 122163 990994
rect 114572 990936 122102 990992
rect 122158 990936 122163 990992
rect 114572 990934 122163 990936
rect 114572 990932 114578 990934
rect 122097 990931 122163 990934
rect 62113 976034 62179 976037
rect 62113 976032 64492 976034
rect 62113 975976 62118 976032
rect 62174 975976 64492 976032
rect 62113 975974 64492 975976
rect 62113 975971 62179 975974
rect 651649 975898 651715 975901
rect 650164 975896 651715 975898
rect 650164 975840 651654 975896
rect 651710 975840 651715 975896
rect 650164 975838 651715 975840
rect 651649 975835 651715 975838
rect 40534 968764 40540 968828
rect 40604 968826 40610 968828
rect 41781 968826 41847 968829
rect 40604 968824 41847 968826
rect 40604 968768 41786 968824
rect 41842 968768 41847 968824
rect 40604 968766 41847 968768
rect 40604 968764 40610 968766
rect 41781 968763 41847 968766
rect 40718 967268 40724 967332
rect 40788 967330 40794 967332
rect 41781 967330 41847 967333
rect 40788 967328 41847 967330
rect 40788 967272 41786 967328
rect 41842 967272 41847 967328
rect 40788 967270 41847 967272
rect 40788 967268 40794 967270
rect 41781 967267 41847 967270
rect 675753 966514 675819 966517
rect 676438 966514 676444 966516
rect 675753 966512 676444 966514
rect 675753 966456 675758 966512
rect 675814 966456 676444 966512
rect 675753 966454 676444 966456
rect 675753 966451 675819 966454
rect 676438 966452 676444 966454
rect 676508 966452 676514 966516
rect 675753 966242 675819 966245
rect 676254 966242 676260 966244
rect 675753 966240 676260 966242
rect 675753 966184 675758 966240
rect 675814 966184 676260 966240
rect 675753 966182 676260 966184
rect 675753 966179 675819 966182
rect 676254 966180 676260 966182
rect 676324 966180 676330 966244
rect 41638 965092 41644 965156
rect 41708 965154 41714 965156
rect 41781 965154 41847 965157
rect 41708 965152 41847 965154
rect 41708 965096 41786 965152
rect 41842 965096 41847 965152
rect 41708 965094 41847 965096
rect 41708 965092 41714 965094
rect 41781 965091 41847 965094
rect 675753 965018 675819 965021
rect 676622 965018 676628 965020
rect 675753 965016 676628 965018
rect 675753 964960 675758 965016
rect 675814 964960 676628 965016
rect 675753 964958 676628 964960
rect 675753 964955 675819 964958
rect 676622 964956 676628 964958
rect 676692 964956 676698 965020
rect 40902 963460 40908 963524
rect 40972 963522 40978 963524
rect 41781 963522 41847 963525
rect 40972 963520 41847 963522
rect 40972 963464 41786 963520
rect 41842 963464 41847 963520
rect 40972 963462 41847 963464
rect 40972 963460 40978 963462
rect 41781 963459 41847 963462
rect 675753 963386 675819 963389
rect 676070 963386 676076 963388
rect 675753 963384 676076 963386
rect 675753 963328 675758 963384
rect 675814 963328 676076 963384
rect 675753 963326 676076 963328
rect 675753 963323 675819 963326
rect 676070 963324 676076 963326
rect 676140 963324 676146 963388
rect 62113 962978 62179 962981
rect 62113 962976 64492 962978
rect 62113 962920 62118 962976
rect 62174 962920 64492 962976
rect 62113 962918 64492 962920
rect 62113 962915 62179 962918
rect 675661 962844 675727 962845
rect 675661 962840 675708 962844
rect 675772 962842 675778 962844
rect 675661 962784 675666 962840
rect 675661 962780 675708 962784
rect 675772 962782 675818 962842
rect 675772 962780 675778 962782
rect 675661 962779 675727 962780
rect 652017 962570 652083 962573
rect 650164 962568 652083 962570
rect 650164 962512 652022 962568
rect 652078 962512 652083 962568
rect 650164 962510 652083 962512
rect 652017 962507 652083 962510
rect 41781 962164 41847 962165
rect 41781 962160 41828 962164
rect 41892 962162 41898 962164
rect 41781 962104 41786 962160
rect 41781 962100 41828 962104
rect 41892 962102 41938 962162
rect 41892 962100 41898 962102
rect 41781 962099 41847 962100
rect 675477 961892 675543 961893
rect 675477 961888 675524 961892
rect 675588 961890 675594 961892
rect 675477 961832 675482 961888
rect 675477 961828 675524 961832
rect 675588 961830 675634 961890
rect 675588 961828 675594 961830
rect 675477 961827 675543 961828
rect 675753 959170 675819 959173
rect 675886 959170 675892 959172
rect 675753 959168 675892 959170
rect 675753 959112 675758 959168
rect 675814 959112 675892 959168
rect 675753 959110 675892 959112
rect 675753 959107 675819 959110
rect 675886 959108 675892 959110
rect 675956 959108 675962 959172
rect 42057 958492 42123 958493
rect 42006 958490 42012 958492
rect 41966 958430 42012 958490
rect 42076 958488 42123 958492
rect 42118 958432 42123 958488
rect 42006 958428 42012 958430
rect 42076 958428 42123 958432
rect 42057 958427 42123 958428
rect 675017 957946 675083 957949
rect 676806 957946 676812 957948
rect 675017 957944 676812 957946
rect 675017 957888 675022 957944
rect 675078 957888 676812 957944
rect 675017 957886 676812 957888
rect 675017 957883 675083 957886
rect 676806 957884 676812 957886
rect 676876 957884 676882 957948
rect 41454 957748 41460 957812
rect 41524 957810 41530 957812
rect 41781 957810 41847 957813
rect 41524 957808 41847 957810
rect 41524 957752 41786 957808
rect 41842 957752 41847 957808
rect 41524 957750 41847 957752
rect 41524 957748 41530 957750
rect 41781 957747 41847 957750
rect 675753 957808 675819 957813
rect 675753 957752 675758 957808
rect 675814 957752 675819 957808
rect 675753 957747 675819 957752
rect 675756 957674 675816 957747
rect 676990 957674 676996 957676
rect 675756 957614 676996 957674
rect 676990 957612 676996 957614
rect 677060 957612 677066 957676
rect 675385 954004 675451 954005
rect 675334 954002 675340 954004
rect 675294 953942 675340 954002
rect 675404 954000 675451 954004
rect 675446 953944 675451 954000
rect 675334 953940 675340 953942
rect 675404 953940 675451 953944
rect 675385 953939 675451 953940
rect 31017 952914 31083 952917
rect 41822 952914 41828 952916
rect 31017 952912 41828 952914
rect 31017 952856 31022 952912
rect 31078 952856 41828 952912
rect 31017 952854 41828 952856
rect 31017 952851 31083 952854
rect 41822 952852 41828 952854
rect 41892 952852 41898 952916
rect 36721 952370 36787 952373
rect 42006 952370 42012 952372
rect 36721 952368 42012 952370
rect 36721 952312 36726 952368
rect 36782 952312 42012 952368
rect 36721 952310 42012 952312
rect 36721 952307 36787 952310
rect 42006 952308 42012 952310
rect 42076 952308 42082 952372
rect 36537 952234 36603 952237
rect 41638 952234 41644 952236
rect 36537 952232 41644 952234
rect 36537 952176 36542 952232
rect 36598 952176 41644 952232
rect 36537 952174 41644 952176
rect 36537 952171 36603 952174
rect 41638 952172 41644 952174
rect 41708 952172 41714 952236
rect 6022 949953 58218 949982
rect 6022 948809 6150 949953
rect 6854 949949 58218 949953
rect 6854 948845 54235 949949
rect 55339 949682 58218 949949
rect 62113 949922 62179 949925
rect 62113 949920 64492 949922
rect 62113 949864 62118 949920
rect 62174 949864 64492 949920
rect 62113 949862 64492 949864
rect 62113 949859 62179 949862
rect 675702 949724 675708 949788
rect 675772 949786 675778 949788
rect 679801 949786 679867 949789
rect 675772 949784 679867 949786
rect 675772 949728 679806 949784
rect 679862 949728 679867 949784
rect 675772 949726 679867 949728
rect 675772 949724 675778 949726
rect 679801 949723 679867 949726
rect 55339 949629 63922 949682
rect 55339 948845 63339 949629
rect 6854 948809 63339 948845
rect 6022 948782 63339 948809
rect 57038 948525 63339 948782
rect 63883 948525 63922 949629
rect 675518 949588 675524 949652
rect 675588 949650 675594 949652
rect 679617 949650 679683 949653
rect 675588 949648 679683 949650
rect 675588 949592 679622 949648
rect 679678 949592 679683 949648
rect 675588 949590 679683 949592
rect 675588 949588 675594 949590
rect 679617 949587 679683 949590
rect 675334 949452 675340 949516
rect 675404 949514 675410 949516
rect 676857 949514 676923 949517
rect 675404 949512 676923 949514
rect 675404 949456 676862 949512
rect 676918 949456 676923 949512
rect 675404 949454 676923 949456
rect 675404 949452 675410 949454
rect 676857 949451 676923 949454
rect 651557 949378 651623 949381
rect 650164 949376 651623 949378
rect 650164 949320 651562 949376
rect 651618 949320 651623 949376
rect 650164 949318 651623 949320
rect 651557 949315 651623 949318
rect 57038 948482 63922 948525
rect 7236 948357 56610 948382
rect 7236 947213 7348 948357
rect 8052 948331 56610 948357
rect 8052 947227 52641 948331
rect 53745 948182 56610 948331
rect 53745 948121 62944 948182
rect 53745 947227 62371 948121
rect 8052 947213 62371 947227
rect 7236 947182 62371 947213
rect 55432 947017 62371 947182
rect 62915 947017 62944 948121
rect 55432 946982 62944 947017
rect 27613 943802 27679 943805
rect 27613 943800 27722 943802
rect 27613 943744 27618 943800
rect 27674 943744 27722 943800
rect 27613 943739 27722 943744
rect 40718 943740 40724 943804
rect 40788 943802 40794 943804
rect 41965 943802 42031 943805
rect 40788 943800 42031 943802
rect 40788 943744 41970 943800
rect 42026 943744 42031 943800
rect 40788 943742 42031 943744
rect 40788 943740 40794 943742
rect 41965 943739 42031 943742
rect 27662 943500 27722 943739
rect 35801 943122 35867 943125
rect 35788 943120 35867 943122
rect 35788 943064 35806 943120
rect 35862 943064 35867 943120
rect 35788 943062 35867 943064
rect 35801 943059 35867 943062
rect 35709 942714 35775 942717
rect 35709 942712 35788 942714
rect 35709 942656 35714 942712
rect 35770 942656 35788 942712
rect 35709 942654 35788 942656
rect 35709 942651 35775 942654
rect 46197 942306 46263 942309
rect 41492 942304 46263 942306
rect 41492 942248 46202 942304
rect 46258 942248 46263 942304
rect 41492 942246 46263 942248
rect 46197 942243 46263 942246
rect 41781 941898 41847 941901
rect 41492 941896 41847 941898
rect 41492 941840 41786 941896
rect 41842 941840 41847 941896
rect 41492 941838 41847 941840
rect 41781 941835 41847 941838
rect 47577 941490 47643 941493
rect 41492 941488 47643 941490
rect 41492 941432 47582 941488
rect 47638 941432 47643 941488
rect 41492 941430 47643 941432
rect 47577 941427 47643 941430
rect 41781 941082 41847 941085
rect 41492 941080 41847 941082
rect 41492 941024 41786 941080
rect 41842 941024 41847 941080
rect 41492 941022 41847 941024
rect 41781 941019 41847 941022
rect 44817 940674 44883 940677
rect 41492 940672 44883 940674
rect 41492 940616 44822 940672
rect 44878 940616 44883 940672
rect 41492 940614 44883 940616
rect 44817 940611 44883 940614
rect 41873 940266 41939 940269
rect 41492 940264 41939 940266
rect 41492 940208 41878 940264
rect 41934 940208 41939 940264
rect 41492 940206 41939 940208
rect 41873 940203 41939 940206
rect 676029 939994 676095 939997
rect 676029 939992 676292 939994
rect 676029 939936 676034 939992
rect 676090 939936 676292 939992
rect 676029 939934 676292 939936
rect 676029 939931 676095 939934
rect 55857 939858 55923 939861
rect 41492 939856 55923 939858
rect 41492 939800 55862 939856
rect 55918 939800 55923 939856
rect 41492 939798 55923 939800
rect 55857 939795 55923 939798
rect 41492 939390 41890 939450
rect 41689 939314 41755 939317
rect 41830 939314 41890 939390
rect 676262 939317 676322 939556
rect 41689 939312 41890 939314
rect 41689 939256 41694 939312
rect 41750 939256 41890 939312
rect 41689 939254 41890 939256
rect 676213 939312 676322 939317
rect 676213 939256 676218 939312
rect 676274 939256 676322 939312
rect 676213 939254 676322 939256
rect 41689 939251 41755 939254
rect 676213 939251 676279 939254
rect 676029 939178 676095 939181
rect 676029 939176 676292 939178
rect 676029 939120 676034 939176
rect 676090 939120 676292 939176
rect 676029 939118 676292 939120
rect 676029 939115 676095 939118
rect 42149 939042 42215 939045
rect 41492 939040 42215 939042
rect 41492 938984 42154 939040
rect 42210 938984 42215 939040
rect 41492 938982 42215 938984
rect 42149 938979 42215 938982
rect 676029 938770 676095 938773
rect 676029 938768 676292 938770
rect 676029 938712 676034 938768
rect 676090 938712 676292 938768
rect 676029 938710 676292 938712
rect 676029 938707 676095 938710
rect 41965 938634 42031 938637
rect 41492 938632 42031 938634
rect 41492 938576 41970 938632
rect 42026 938576 42031 938632
rect 41492 938574 42031 938576
rect 41965 938571 42031 938574
rect 676029 938362 676095 938365
rect 676029 938360 676292 938362
rect 676029 938304 676034 938360
rect 676090 938304 676292 938360
rect 676029 938302 676292 938304
rect 676029 938299 676095 938302
rect 32397 938226 32463 938229
rect 32397 938224 32476 938226
rect 32397 938168 32402 938224
rect 32458 938168 32476 938224
rect 32397 938166 32476 938168
rect 32397 938163 32463 938166
rect 42006 937818 42012 937820
rect 41492 937758 42012 937818
rect 42006 937756 42012 937758
rect 42076 937756 42082 937820
rect 676262 937685 676322 937924
rect 676213 937680 676322 937685
rect 676213 937624 676218 937680
rect 676274 937624 676322 937680
rect 676213 937622 676322 937624
rect 676213 937619 676279 937622
rect 676029 937546 676095 937549
rect 676029 937544 676292 937546
rect 676029 937488 676034 937544
rect 676090 937488 676292 937544
rect 676029 937486 676292 937488
rect 676029 937483 676095 937486
rect 31017 937410 31083 937413
rect 31004 937408 31083 937410
rect 31004 937352 31022 937408
rect 31078 937352 31083 937408
rect 31004 937350 31083 937352
rect 31017 937347 31083 937350
rect 676213 937274 676279 937277
rect 676213 937272 676322 937274
rect 676213 937216 676218 937272
rect 676274 937216 676322 937272
rect 676213 937211 676322 937216
rect 676262 937108 676322 937211
rect 62113 937002 62179 937005
rect 41492 936942 41890 937002
rect 41830 936868 41890 936942
rect 62113 937000 64492 937002
rect 62113 936944 62118 937000
rect 62174 936944 64492 937000
rect 62113 936942 64492 936944
rect 62113 936939 62179 936942
rect 41822 936804 41828 936868
rect 41892 936804 41898 936868
rect 37917 936594 37983 936597
rect 37917 936592 37996 936594
rect 37917 936536 37922 936592
rect 37978 936536 37996 936592
rect 37917 936534 37996 936536
rect 37917 936531 37983 936534
rect 676121 936458 676187 936461
rect 676262 936458 676322 936700
rect 676121 936456 676322 936458
rect 676121 936400 676126 936456
rect 676182 936400 676322 936456
rect 676121 936398 676322 936400
rect 676121 936395 676187 936398
rect 36721 936186 36787 936189
rect 651557 936186 651623 936189
rect 36708 936184 36787 936186
rect 36708 936128 36726 936184
rect 36782 936128 36787 936184
rect 36708 936126 36787 936128
rect 650164 936184 651623 936186
rect 650164 936128 651562 936184
rect 651618 936128 651623 936184
rect 650164 936126 651623 936128
rect 36721 936123 36787 936126
rect 651557 936123 651623 936126
rect 676262 936053 676322 936292
rect 676213 936048 676322 936053
rect 676213 935992 676218 936048
rect 676274 935992 676322 936048
rect 676213 935990 676322 935992
rect 676213 935987 676279 935990
rect 676029 935914 676095 935917
rect 676029 935912 676292 935914
rect 676029 935856 676034 935912
rect 676090 935856 676292 935912
rect 676029 935854 676292 935856
rect 676029 935851 676095 935854
rect 42977 935778 43043 935781
rect 41492 935776 43043 935778
rect 41492 935720 42982 935776
rect 43038 935720 43043 935776
rect 41492 935718 43043 935720
rect 42977 935715 43043 935718
rect 676622 935580 676628 935644
rect 676692 935580 676698 935644
rect 676630 935476 676690 935580
rect 36537 935370 36603 935373
rect 36524 935368 36603 935370
rect 36524 935312 36542 935368
rect 36598 935312 36603 935368
rect 36524 935310 36603 935312
rect 36537 935307 36603 935310
rect 676857 935234 676923 935237
rect 676814 935232 676923 935234
rect 676814 935176 676862 935232
rect 676918 935176 676923 935232
rect 676814 935171 676923 935176
rect 676814 935068 676874 935171
rect 42006 934962 42012 934964
rect 41492 934902 42012 934962
rect 42006 934900 42012 934902
rect 42076 934900 42082 934964
rect 676438 934764 676444 934828
rect 676508 934764 676514 934828
rect 676446 934660 676506 934764
rect 44173 934554 44239 934557
rect 41492 934552 44239 934554
rect 41492 934496 44178 934552
rect 44234 934496 44239 934552
rect 41492 934494 44239 934496
rect 44173 934491 44239 934494
rect 42885 934146 42951 934149
rect 41492 934144 42951 934146
rect 41492 934088 42890 934144
rect 42946 934088 42951 934144
rect 41492 934086 42951 934088
rect 42885 934083 42951 934086
rect 676070 933948 676076 934012
rect 676140 934010 676146 934012
rect 676262 934010 676322 934252
rect 676140 933950 676322 934010
rect 676140 933948 676146 933950
rect 675886 933812 675892 933876
rect 675956 933874 675962 933876
rect 675956 933814 676292 933874
rect 675956 933812 675962 933814
rect 42793 933738 42859 933741
rect 41492 933736 42859 933738
rect 41492 933680 42798 933736
rect 42854 933680 42859 933736
rect 41492 933678 42859 933680
rect 42793 933675 42859 933678
rect 678237 933602 678303 933605
rect 678237 933600 678346 933602
rect 678237 933544 678242 933600
rect 678298 933544 678346 933600
rect 678237 933539 678346 933544
rect 678286 933436 678346 933539
rect 39941 933330 40007 933333
rect 39941 933328 40020 933330
rect 39941 933272 39946 933328
rect 40002 933272 40020 933328
rect 39941 933270 40020 933272
rect 39941 933267 40007 933270
rect 676622 933132 676628 933196
rect 676692 933132 676698 933196
rect 676630 933028 676690 933132
rect 21774 932484 21834 932910
rect 679801 932786 679867 932789
rect 679758 932784 679867 932786
rect 679758 932728 679806 932784
rect 679862 932728 679867 932784
rect 679758 932723 679867 932728
rect 679758 932620 679818 932723
rect 679617 932378 679683 932381
rect 679574 932376 679683 932378
rect 679574 932320 679622 932376
rect 679678 932320 679683 932376
rect 679574 932315 679683 932320
rect 41689 932242 41755 932245
rect 41689 932240 41890 932242
rect 41689 932184 41694 932240
rect 41750 932184 41890 932240
rect 679574 932212 679634 932315
rect 41689 932182 41890 932184
rect 41689 932179 41755 932182
rect 41830 932106 41890 932182
rect 41492 932046 41890 932106
rect 676029 931834 676095 931837
rect 676029 931832 676292 931834
rect 676029 931776 676034 931832
rect 676090 931776 676292 931832
rect 676029 931774 676292 931776
rect 676029 931771 676095 931774
rect 676990 931500 676996 931564
rect 677060 931500 677066 931564
rect 676998 931396 677058 931500
rect 676806 931092 676812 931156
rect 676876 931092 676882 931156
rect 676814 930988 676874 931092
rect 676213 930746 676279 930749
rect 676213 930744 676322 930746
rect 676213 930688 676218 930744
rect 676274 930688 676322 930744
rect 676213 930683 676322 930688
rect 676262 930580 676322 930683
rect 676213 930338 676279 930341
rect 676213 930336 676322 930338
rect 676213 930280 676218 930336
rect 676274 930280 676322 930336
rect 676213 930275 676322 930280
rect 676262 930172 676322 930275
rect 683070 929525 683130 929764
rect 683070 929520 683179 929525
rect 683070 929464 683118 929520
rect 683174 929464 683179 929520
rect 683070 929462 683179 929464
rect 683113 929459 683179 929462
rect 685830 928948 685890 929356
rect 683113 928706 683179 928709
rect 683070 928704 683179 928706
rect 683070 928648 683118 928704
rect 683174 928648 683179 928704
rect 683070 928643 683179 928648
rect 683070 928540 683130 928643
rect 62113 923810 62179 923813
rect 62113 923808 64492 923810
rect 62113 923752 62118 923808
rect 62174 923752 64492 923808
rect 62113 923750 64492 923752
rect 62113 923747 62179 923750
rect 651557 922722 651623 922725
rect 650164 922720 651623 922722
rect 650164 922664 651562 922720
rect 651618 922664 651623 922720
rect 650164 922662 651623 922664
rect 651557 922659 651623 922662
rect 62113 910754 62179 910757
rect 62113 910752 64492 910754
rect 62113 910696 62118 910752
rect 62174 910696 64492 910752
rect 62113 910694 64492 910696
rect 62113 910691 62179 910694
rect 651557 909530 651623 909533
rect 650164 909528 651623 909530
rect 650164 909472 651562 909528
rect 651618 909472 651623 909528
rect 650164 909470 651623 909472
rect 651557 909467 651623 909470
rect 62113 897834 62179 897837
rect 62113 897832 64492 897834
rect 62113 897776 62118 897832
rect 62174 897776 64492 897832
rect 62113 897774 64492 897776
rect 62113 897771 62179 897774
rect 651557 896202 651623 896205
rect 650164 896200 651623 896202
rect 650164 896144 651562 896200
rect 651618 896144 651623 896200
rect 650164 896142 651623 896144
rect 651557 896139 651623 896142
rect 62113 884778 62179 884781
rect 62113 884776 64492 884778
rect 62113 884720 62118 884776
rect 62174 884720 64492 884776
rect 62113 884718 64492 884720
rect 62113 884715 62179 884718
rect 652017 882874 652083 882877
rect 650164 882872 652083 882874
rect 650164 882816 652022 882872
rect 652078 882816 652083 882872
rect 650164 882814 652083 882816
rect 652017 882811 652083 882814
rect 675150 877236 675156 877300
rect 675220 877298 675226 877300
rect 675385 877298 675451 877301
rect 675220 877296 675451 877298
rect 675220 877240 675390 877296
rect 675446 877240 675451 877296
rect 675220 877238 675451 877240
rect 675220 877236 675226 877238
rect 675385 877235 675451 877238
rect 675753 876618 675819 876621
rect 676254 876618 676260 876620
rect 675753 876616 676260 876618
rect 675753 876560 675758 876616
rect 675814 876560 676260 876616
rect 675753 876558 676260 876560
rect 675753 876555 675819 876558
rect 676254 876556 676260 876558
rect 676324 876556 676330 876620
rect 675753 875938 675819 875941
rect 676070 875938 676076 875940
rect 675753 875936 676076 875938
rect 675753 875880 675758 875936
rect 675814 875880 676076 875936
rect 675753 875878 676076 875880
rect 675753 875875 675819 875878
rect 676070 875876 676076 875878
rect 676140 875876 676146 875940
rect 675753 874034 675819 874037
rect 675886 874034 675892 874036
rect 675753 874032 675892 874034
rect 675753 873976 675758 874032
rect 675814 873976 675892 874032
rect 675753 873974 675892 873976
rect 675753 873971 675819 873974
rect 675886 873972 675892 873974
rect 675956 873972 675962 874036
rect 62113 871722 62179 871725
rect 62113 871720 64492 871722
rect 62113 871664 62118 871720
rect 62174 871664 64492 871720
rect 62113 871662 64492 871664
rect 62113 871659 62179 871662
rect 651557 869682 651623 869685
rect 650164 869680 651623 869682
rect 650164 869624 651562 869680
rect 651618 869624 651623 869680
rect 650164 869622 651623 869624
rect 651557 869619 651623 869622
rect 675753 866826 675819 866829
rect 676438 866826 676444 866828
rect 675753 866824 676444 866826
rect 675753 866768 675758 866824
rect 675814 866768 676444 866824
rect 675753 866766 676444 866768
rect 675753 866763 675819 866766
rect 676438 866764 676444 866766
rect 676508 866764 676514 866828
rect 675753 864788 675819 864789
rect 675702 864786 675708 864788
rect 675662 864726 675708 864786
rect 675772 864784 675819 864788
rect 675814 864728 675819 864784
rect 675702 864724 675708 864726
rect 675772 864724 675819 864728
rect 675753 864723 675819 864724
rect 62113 858666 62179 858669
rect 62113 858664 64492 858666
rect 62113 858608 62118 858664
rect 62174 858608 64492 858664
rect 62113 858606 64492 858608
rect 62113 858603 62179 858606
rect 651557 856354 651623 856357
rect 650164 856352 651623 856354
rect 650164 856296 651562 856352
rect 651618 856296 651623 856352
rect 650164 856294 651623 856296
rect 651557 856291 651623 856294
rect 62113 845610 62179 845613
rect 62113 845608 64492 845610
rect 62113 845552 62118 845608
rect 62174 845552 64492 845608
rect 62113 845550 64492 845552
rect 62113 845547 62179 845550
rect 651557 843026 651623 843029
rect 650164 843024 651623 843026
rect 650164 842968 651562 843024
rect 651618 842968 651623 843024
rect 650164 842966 651623 842968
rect 651557 842963 651623 842966
rect 39852 842334 50002 842458
rect 39852 837790 47909 842334
rect 49693 837790 50002 842334
rect 39852 837678 50002 837790
rect 667172 833210 677818 833301
rect 62113 832554 62179 832557
rect 62113 832552 64492 832554
rect 62113 832496 62118 832552
rect 62174 832496 64492 832552
rect 62113 832494 64492 832496
rect 62113 832491 62179 832494
rect 39852 832402 50002 832479
rect 39852 827858 47909 832402
rect 49693 827858 50002 832402
rect 651557 829834 651623 829837
rect 650164 829832 651623 829834
rect 650164 829776 651562 829832
rect 651618 829776 651623 829832
rect 650164 829774 651623 829776
rect 651557 829771 651623 829774
rect 667172 828626 667276 833210
rect 669740 828626 677818 833210
rect 667172 828521 677818 828626
rect 39852 827699 50002 827858
rect 6022 824153 63922 824182
rect 6022 823009 6150 824153
rect 6854 824149 63922 824153
rect 6854 823045 54235 824149
rect 55339 824129 63922 824149
rect 55339 823045 63339 824129
rect 6854 823025 63339 823045
rect 63883 823025 63922 824129
rect 6854 823009 63922 823025
rect 6022 822982 63922 823009
rect 667172 823216 677818 823322
rect 7236 822557 62944 822582
rect 7236 821413 7348 822557
rect 8052 822531 62944 822557
rect 8052 821427 52641 822531
rect 53745 822521 62944 822531
rect 53745 821427 62371 822521
rect 8052 821417 62371 821427
rect 62915 821417 62944 822521
rect 8052 821413 62944 821417
rect 7236 821382 62944 821413
rect 62113 819498 62179 819501
rect 62113 819496 64492 819498
rect 62113 819440 62118 819496
rect 62174 819440 64492 819496
rect 62113 819438 64492 819440
rect 62113 819435 62179 819438
rect 667172 818632 667262 823216
rect 669726 818632 677818 823216
rect 667172 818542 677818 818632
rect 41229 818002 41295 818005
rect 41229 818000 41338 818002
rect 41229 817944 41234 818000
rect 41290 817944 41338 818000
rect 41229 817939 41338 817944
rect 41278 817700 41338 817939
rect 41321 817322 41387 817325
rect 41308 817320 41387 817322
rect 41308 817264 41326 817320
rect 41382 817264 41387 817320
rect 41308 817262 41387 817264
rect 41321 817259 41387 817262
rect 54477 816914 54543 816917
rect 41492 816912 54543 816914
rect 41492 816856 54482 816912
rect 54538 816856 54543 816912
rect 41492 816854 54543 816856
rect 54477 816851 54543 816854
rect 41689 816642 41755 816645
rect 41689 816640 41890 816642
rect 41689 816584 41694 816640
rect 41750 816584 41890 816640
rect 41689 816582 41890 816584
rect 41689 816579 41755 816582
rect 41830 816506 41890 816582
rect 651557 816506 651623 816509
rect 41492 816446 41890 816506
rect 650164 816504 651623 816506
rect 650164 816448 651562 816504
rect 651618 816448 651623 816504
rect 650164 816446 651623 816448
rect 651557 816443 651623 816446
rect 42006 816098 42012 816100
rect 41492 816038 42012 816098
rect 42006 816036 42012 816038
rect 42076 816036 42082 816100
rect 41873 815690 41939 815693
rect 41492 815688 41939 815690
rect 41492 815632 41878 815688
rect 41934 815632 41939 815688
rect 41492 815630 41939 815632
rect 41873 815627 41939 815630
rect 44265 815282 44331 815285
rect 41492 815280 44331 815282
rect 41492 815224 44270 815280
rect 44326 815224 44331 815280
rect 41492 815222 44331 815224
rect 44265 815219 44331 815222
rect 41965 814874 42031 814877
rect 41492 814872 42031 814874
rect 41492 814816 41970 814872
rect 42026 814816 42031 814872
rect 41492 814814 42031 814816
rect 41965 814811 42031 814814
rect 41822 814466 41828 814468
rect 41492 814406 41828 814466
rect 41822 814404 41828 814406
rect 41892 814404 41898 814468
rect 41781 814058 41847 814061
rect 41492 814056 41847 814058
rect 41492 814000 41786 814056
rect 41842 814000 41847 814056
rect 41492 813998 41847 814000
rect 41781 813995 41847 813998
rect 44173 813650 44239 813653
rect 41492 813648 44239 813650
rect 41492 813592 44178 813648
rect 44234 813592 44239 813648
rect 41492 813590 44239 813592
rect 44173 813587 44239 813590
rect 40677 813242 40743 813245
rect 40677 813240 40756 813242
rect 40677 813184 40682 813240
rect 40738 813184 40756 813240
rect 40677 813182 40756 813184
rect 40677 813179 40743 813182
rect 42149 812834 42215 812837
rect 41492 812832 42215 812834
rect 41492 812776 42154 812832
rect 42210 812776 42215 812832
rect 41492 812774 42215 812776
rect 42149 812771 42215 812774
rect 33777 812426 33843 812429
rect 33764 812424 33843 812426
rect 33764 812368 33782 812424
rect 33838 812368 33843 812424
rect 33764 812366 33843 812368
rect 33777 812363 33843 812366
rect 42190 812018 42196 812020
rect 41492 811958 42196 812018
rect 42190 811956 42196 811958
rect 42260 811956 42266 812020
rect 41781 811610 41847 811613
rect 41492 811608 41847 811610
rect 41492 811552 41786 811608
rect 41842 811552 41847 811608
rect 41492 811550 41847 811552
rect 41781 811547 41847 811550
rect 42333 811202 42399 811205
rect 41492 811200 42399 811202
rect 41492 811144 42338 811200
rect 42394 811144 42399 811200
rect 41492 811142 42399 811144
rect 42333 811139 42399 811142
rect 34421 810794 34487 810797
rect 34421 810792 34500 810794
rect 34421 810736 34426 810792
rect 34482 810736 34500 810792
rect 34421 810734 34500 810736
rect 34421 810731 34487 810734
rect 33041 810386 33107 810389
rect 33028 810384 33107 810386
rect 33028 810328 33046 810384
rect 33102 810328 33107 810384
rect 33028 810326 33107 810328
rect 33041 810323 33107 810326
rect 42793 809978 42859 809981
rect 41492 809976 42859 809978
rect 41492 809920 42798 809976
rect 42854 809920 42859 809976
rect 41492 809918 42859 809920
rect 42793 809915 42859 809918
rect 42057 809570 42123 809573
rect 41492 809568 42123 809570
rect 41492 809512 42062 809568
rect 42118 809512 42123 809568
rect 41492 809510 42123 809512
rect 42057 809507 42123 809510
rect 32397 809162 32463 809165
rect 32397 809160 32476 809162
rect 32397 809104 32402 809160
rect 32458 809104 32476 809160
rect 32397 809102 32476 809104
rect 32397 809099 32463 809102
rect 35157 808754 35223 808757
rect 35157 808752 35236 808754
rect 35157 808696 35162 808752
rect 35218 808696 35236 808752
rect 35157 808694 35236 808696
rect 35157 808691 35223 808694
rect 44357 808346 44423 808349
rect 41492 808344 44423 808346
rect 41492 808288 44362 808344
rect 44418 808288 44423 808344
rect 41492 808286 44423 808288
rect 44357 808283 44423 808286
rect 41822 807938 41828 807940
rect 41492 807878 41828 807938
rect 41822 807876 41828 807878
rect 41892 807876 41898 807940
rect 39806 807333 39866 807500
rect 39806 807328 39915 807333
rect 39806 807272 39854 807328
rect 39910 807272 39915 807328
rect 39806 807270 39915 807272
rect 39849 807267 39915 807270
rect 24902 806684 24962 807092
rect 62113 806578 62179 806581
rect 62113 806576 64492 806578
rect 62113 806520 62118 806576
rect 62174 806520 64492 806576
rect 62113 806518 64492 806520
rect 62113 806515 62179 806518
rect 41781 806306 41847 806309
rect 43437 806306 43503 806309
rect 41492 806304 43503 806306
rect 41492 806248 41786 806304
rect 41842 806248 43442 806304
rect 43498 806248 43503 806304
rect 41492 806246 43503 806248
rect 41781 806243 41847 806246
rect 43437 806243 43503 806246
rect 651557 803314 651623 803317
rect 650164 803312 651623 803314
rect 650164 803256 651562 803312
rect 651618 803256 651623 803312
rect 650164 803254 651623 803256
rect 651557 803251 651623 803254
rect 34421 802634 34487 802637
rect 41638 802634 41644 802636
rect 34421 802632 41644 802634
rect 34421 802576 34426 802632
rect 34482 802576 41644 802632
rect 34421 802574 41644 802576
rect 34421 802571 34487 802574
rect 41638 802572 41644 802574
rect 41708 802572 41714 802636
rect 33041 802498 33107 802501
rect 42006 802498 42012 802500
rect 33041 802496 42012 802498
rect 33041 802440 33046 802496
rect 33102 802440 42012 802496
rect 33041 802438 42012 802440
rect 33041 802435 33107 802438
rect 42006 802436 42012 802438
rect 42076 802436 42082 802500
rect 40677 801682 40743 801685
rect 41822 801682 41828 801684
rect 40677 801680 41828 801682
rect 40677 801624 40682 801680
rect 40738 801624 41828 801680
rect 40677 801622 41828 801624
rect 40677 801619 40743 801622
rect 41822 801620 41828 801622
rect 41892 801620 41898 801684
rect 33777 801002 33843 801005
rect 41454 801002 41460 801004
rect 33777 801000 41460 801002
rect 33777 800944 33782 801000
rect 33838 800944 41460 801000
rect 33777 800942 41460 800944
rect 33777 800939 33843 800942
rect 41454 800940 41460 800942
rect 41524 800940 41530 801004
rect 40534 796724 40540 796788
rect 40604 796786 40610 796788
rect 42425 796786 42491 796789
rect 40604 796784 42491 796786
rect 40604 796728 42430 796784
rect 42486 796728 42491 796784
rect 40604 796726 42491 796728
rect 40604 796724 40610 796726
rect 42425 796723 42491 796726
rect 62113 793658 62179 793661
rect 62113 793656 64492 793658
rect 62113 793600 62118 793656
rect 62174 793600 64492 793656
rect 62113 793598 64492 793600
rect 62113 793595 62179 793598
rect 42006 791964 42012 792028
rect 42076 792026 42082 792028
rect 42333 792026 42399 792029
rect 42076 792024 42399 792026
rect 42076 791968 42338 792024
rect 42394 791968 42399 792024
rect 42076 791966 42399 791968
rect 42076 791964 42082 791966
rect 42333 791963 42399 791966
rect 42190 791828 42196 791892
rect 42260 791890 42266 791892
rect 42701 791890 42767 791893
rect 42260 791888 42767 791890
rect 42260 791832 42706 791888
rect 42762 791832 42767 791888
rect 42260 791830 42767 791832
rect 42260 791828 42266 791830
rect 42701 791827 42767 791830
rect 651649 789986 651715 789989
rect 650164 789984 651715 789986
rect 650164 789928 651654 789984
rect 651710 789928 651715 789984
rect 650164 789926 651715 789928
rect 651649 789923 651715 789926
rect 41454 788156 41460 788220
rect 41524 788218 41530 788220
rect 42701 788218 42767 788221
rect 41524 788216 42767 788218
rect 41524 788160 42706 788216
rect 42762 788160 42767 788216
rect 41524 788158 42767 788160
rect 41524 788156 41530 788158
rect 42701 788155 42767 788158
rect 41822 788020 41828 788084
rect 41892 788082 41898 788084
rect 42425 788082 42491 788085
rect 41892 788080 42491 788082
rect 41892 788024 42430 788080
rect 42486 788024 42491 788080
rect 41892 788022 42491 788024
rect 41892 788020 41898 788022
rect 42425 788019 42491 788022
rect 41638 786116 41644 786180
rect 41708 786178 41714 786180
rect 41781 786178 41847 786181
rect 41708 786176 41847 786178
rect 41708 786120 41786 786176
rect 41842 786120 41847 786176
rect 41708 786118 41847 786120
rect 41708 786116 41714 786118
rect 41781 786115 41847 786118
rect 675702 785164 675708 785228
rect 675772 785164 675778 785228
rect 675710 784954 675770 785164
rect 675886 784954 675892 784956
rect 675710 784894 675892 784954
rect 675886 784892 675892 784894
rect 675956 784892 675962 784956
rect 675477 784820 675543 784821
rect 675477 784816 675524 784820
rect 675588 784818 675594 784820
rect 675477 784760 675482 784816
rect 675477 784756 675524 784760
rect 675588 784758 675634 784818
rect 675588 784756 675594 784758
rect 675477 784755 675543 784756
rect 675150 784212 675156 784276
rect 675220 784274 675226 784276
rect 675702 784274 675708 784276
rect 675220 784214 675708 784274
rect 675220 784212 675226 784214
rect 675702 784212 675708 784214
rect 675772 784212 675778 784276
rect 675753 784138 675819 784141
rect 676622 784138 676628 784140
rect 675753 784136 676628 784138
rect 675753 784080 675758 784136
rect 675814 784080 676628 784136
rect 675753 784078 676628 784080
rect 675753 784075 675819 784078
rect 676622 784076 676628 784078
rect 676692 784076 676698 784140
rect 56078 782129 63922 782182
rect 56078 781025 63339 782129
rect 63883 781025 63922 782129
rect 56078 780982 63922 781025
rect 6022 780953 57370 780982
rect 6022 779809 6150 780953
rect 6854 780949 57370 780953
rect 6854 779845 54235 780949
rect 55339 779845 57370 780949
rect 62113 780466 62179 780469
rect 62113 780464 64492 780466
rect 62113 780408 62118 780464
rect 62174 780408 64492 780464
rect 62113 780406 64492 780408
rect 62113 780403 62179 780406
rect 675385 779922 675451 779925
rect 677174 779922 677180 779924
rect 675385 779920 677180 779922
rect 675385 779864 675390 779920
rect 675446 779864 677180 779920
rect 675385 779862 677180 779864
rect 675385 779859 675451 779862
rect 677174 779860 677180 779862
rect 677244 779860 677250 779924
rect 6854 779809 57370 779845
rect 6022 779782 57370 779809
rect 7236 779357 62944 779382
rect 7236 778213 7348 779357
rect 8052 779331 62944 779357
rect 8052 778227 52641 779331
rect 53745 779321 62944 779331
rect 53745 778227 62371 779321
rect 8052 778217 62371 778227
rect 62915 778217 62944 779321
rect 8052 778213 62944 778217
rect 7236 778182 62944 778213
rect 651557 776658 651623 776661
rect 650164 776656 651623 776658
rect 650164 776600 651562 776656
rect 651618 776600 651623 776656
rect 650164 776598 651623 776600
rect 651557 776595 651623 776598
rect 675150 775644 675156 775708
rect 675220 775706 675226 775708
rect 675385 775706 675451 775709
rect 675220 775704 675451 775706
rect 675220 775648 675390 775704
rect 675446 775648 675451 775704
rect 675220 775646 675451 775648
rect 675220 775644 675226 775646
rect 675385 775643 675451 775646
rect 675334 774828 675340 774892
rect 675404 774890 675410 774892
rect 676806 774890 676812 774892
rect 675404 774830 676812 774890
rect 675404 774828 675410 774830
rect 676806 774828 676812 774830
rect 676876 774828 676882 774892
rect 35758 774349 35818 774452
rect 35758 774344 35867 774349
rect 35758 774288 35806 774344
rect 35862 774288 35867 774344
rect 35758 774286 35867 774288
rect 35801 774283 35867 774286
rect 41462 773938 41522 774044
rect 50337 773938 50403 773941
rect 41462 773936 50403 773938
rect 41462 773880 50342 773936
rect 50398 773880 50403 773936
rect 41462 773878 50403 773880
rect 50337 773875 50403 773878
rect 43621 773666 43687 773669
rect 41492 773664 43687 773666
rect 41492 773608 43626 773664
rect 43682 773608 43687 773664
rect 41492 773606 43687 773608
rect 43621 773603 43687 773606
rect 40166 773468 40172 773532
rect 40236 773468 40242 773532
rect 40174 773228 40234 773468
rect 675753 773396 675819 773397
rect 675702 773394 675708 773396
rect 675662 773334 675708 773394
rect 675772 773392 675819 773396
rect 675814 773336 675819 773392
rect 675702 773332 675708 773334
rect 675772 773332 675819 773336
rect 675753 773331 675819 773332
rect 44725 772850 44791 772853
rect 41492 772848 44791 772850
rect 41492 772792 44730 772848
rect 44786 772792 44791 772848
rect 41492 772790 44791 772792
rect 44725 772787 44791 772790
rect 675886 772652 675892 772716
rect 675956 772714 675962 772716
rect 679617 772714 679683 772717
rect 675956 772712 679683 772714
rect 675956 772656 679622 772712
rect 679678 772656 679683 772712
rect 675956 772654 679683 772656
rect 675956 772652 675962 772654
rect 679617 772651 679683 772654
rect 44265 772442 44331 772445
rect 41492 772440 44331 772442
rect 41492 772384 44270 772440
rect 44326 772384 44331 772440
rect 41492 772382 44331 772384
rect 44265 772379 44331 772382
rect 42793 772034 42859 772037
rect 41492 772032 42859 772034
rect 41492 771976 42798 772032
rect 42854 771976 42859 772032
rect 41492 771974 42859 771976
rect 42793 771971 42859 771974
rect 39982 771836 39988 771900
rect 40052 771836 40058 771900
rect 39990 771596 40050 771836
rect 39990 771084 40050 771188
rect 39982 771020 39988 771084
rect 40052 771020 40058 771084
rect 44173 770810 44239 770813
rect 41492 770808 44239 770810
rect 41492 770752 44178 770808
rect 44234 770752 44239 770808
rect 41492 770750 44239 770752
rect 44173 770747 44239 770750
rect 44633 770402 44699 770405
rect 41492 770400 44699 770402
rect 41492 770344 44638 770400
rect 44694 770344 44699 770400
rect 41492 770342 44699 770344
rect 44633 770339 44699 770342
rect 44357 769994 44423 769997
rect 41492 769992 44423 769994
rect 41492 769936 44362 769992
rect 44418 769936 44423 769992
rect 41492 769934 44423 769936
rect 44357 769931 44423 769934
rect 33734 769453 33794 769556
rect 33734 769448 33843 769453
rect 33734 769392 33782 769448
rect 33838 769392 33843 769448
rect 33734 769390 33843 769392
rect 33777 769387 33843 769390
rect 40726 769045 40786 769148
rect 40677 769040 40786 769045
rect 40677 768984 40682 769040
rect 40738 768984 40786 769040
rect 40677 768982 40786 768984
rect 40677 768979 40743 768982
rect 32446 768637 32506 768740
rect 32397 768632 32506 768637
rect 32397 768576 32402 768632
rect 32458 768576 32506 768632
rect 32397 768574 32506 768576
rect 32397 768571 32463 768574
rect 44449 768362 44515 768365
rect 41492 768360 44515 768362
rect 41492 768304 44454 768360
rect 44510 768304 44515 768360
rect 41492 768302 44515 768304
rect 44449 768299 44515 768302
rect 30974 767821 31034 767924
rect 30974 767816 31083 767821
rect 30974 767760 31022 767816
rect 31078 767760 31083 767816
rect 30974 767758 31083 767760
rect 31017 767755 31083 767758
rect 35206 767413 35266 767516
rect 35157 767408 35266 767413
rect 35157 767352 35162 767408
rect 35218 767352 35266 767408
rect 35157 767350 35266 767352
rect 62113 767410 62179 767413
rect 62113 767408 64492 767410
rect 62113 767352 62118 767408
rect 62174 767352 64492 767408
rect 62113 767350 64492 767352
rect 35157 767347 35223 767350
rect 62113 767347 62179 767350
rect 42885 767138 42951 767141
rect 41492 767136 42951 767138
rect 41492 767080 42890 767136
rect 42946 767080 42951 767136
rect 41492 767078 42951 767080
rect 42885 767075 42951 767078
rect 32446 766597 32506 766700
rect 32446 766592 32555 766597
rect 32446 766536 32494 766592
rect 32550 766536 32555 766592
rect 32446 766534 32555 766536
rect 32489 766531 32555 766534
rect 40910 766188 40970 766292
rect 40902 766124 40908 766188
rect 40972 766124 40978 766188
rect 42977 765914 43043 765917
rect 41492 765912 43043 765914
rect 41492 765856 42982 765912
rect 43038 765856 43043 765912
rect 41492 765854 43043 765856
rect 42977 765851 43043 765854
rect 44541 765506 44607 765509
rect 41492 765504 44607 765506
rect 41492 765448 44546 765504
rect 44602 765448 44607 765504
rect 41492 765446 44607 765448
rect 44541 765443 44607 765446
rect 40542 764964 40602 765068
rect 40534 764900 40540 764964
rect 40604 764900 40610 764964
rect 40726 764556 40786 764660
rect 40718 764492 40724 764556
rect 40788 764492 40794 764556
rect 30422 764149 30482 764252
rect 30373 764144 30482 764149
rect 30373 764088 30378 764144
rect 30434 764088 30482 764144
rect 30373 764086 30482 764088
rect 30373 764083 30439 764086
rect 30422 763436 30482 763844
rect 30373 763330 30439 763333
rect 651557 763330 651623 763333
rect 30373 763328 30482 763330
rect 30373 763272 30378 763328
rect 30434 763272 30482 763328
rect 30373 763267 30482 763272
rect 650164 763328 651623 763330
rect 650164 763272 651562 763328
rect 651618 763272 651623 763328
rect 650164 763270 651623 763272
rect 651557 763267 651623 763270
rect 30422 763028 30482 763267
rect 41462 762925 41522 763028
rect 41462 762920 41571 762925
rect 41462 762864 41510 762920
rect 41566 762864 41571 762920
rect 41462 762862 41571 762864
rect 41505 762859 41571 762862
rect 676121 761290 676187 761293
rect 676262 761290 676322 761532
rect 676121 761288 676322 761290
rect 676121 761232 676126 761288
rect 676182 761232 676322 761288
rect 676121 761230 676322 761232
rect 676121 761227 676187 761230
rect 676262 760885 676322 761124
rect 676213 760880 676322 760885
rect 676213 760824 676218 760880
rect 676274 760824 676322 760880
rect 676213 760822 676322 760824
rect 676213 760819 676279 760822
rect 676029 760746 676095 760749
rect 676029 760744 676292 760746
rect 676029 760688 676034 760744
rect 676090 760688 676292 760744
rect 676029 760686 676292 760688
rect 676029 760683 676095 760686
rect 676029 760338 676095 760341
rect 676029 760336 676292 760338
rect 676029 760280 676034 760336
rect 676090 760280 676292 760336
rect 676029 760278 676292 760280
rect 676029 760275 676095 760278
rect 676262 759661 676322 759900
rect 676213 759656 676322 759661
rect 676213 759600 676218 759656
rect 676274 759600 676322 759656
rect 676213 759598 676322 759600
rect 676213 759595 676279 759598
rect 676029 759522 676095 759525
rect 676029 759520 676292 759522
rect 676029 759464 676034 759520
rect 676090 759464 676292 759520
rect 676029 759462 676292 759464
rect 676029 759459 676095 759462
rect 672349 759114 672415 759117
rect 672758 759114 672764 759116
rect 672349 759112 672764 759114
rect 672349 759056 672354 759112
rect 672410 759056 672764 759112
rect 672349 759054 672764 759056
rect 672349 759051 672415 759054
rect 672758 759052 672764 759054
rect 672828 759052 672834 759116
rect 676029 759114 676095 759117
rect 676029 759112 676292 759114
rect 676029 759056 676034 759112
rect 676090 759056 676292 759112
rect 676029 759054 676292 759056
rect 676029 759051 676095 759054
rect 672809 758434 672875 758437
rect 676262 758434 676322 758676
rect 672809 758432 676322 758434
rect 672809 758376 672814 758432
rect 672870 758376 676322 758432
rect 672809 758374 676322 758376
rect 672809 758371 672875 758374
rect 35157 758298 35223 758301
rect 41638 758298 41644 758300
rect 35157 758296 41644 758298
rect 35157 758240 35162 758296
rect 35218 758240 41644 758296
rect 35157 758238 41644 758240
rect 35157 758235 35223 758238
rect 41638 758236 41644 758238
rect 41708 758236 41714 758300
rect 676029 758298 676095 758301
rect 676029 758296 676292 758298
rect 676029 758240 676034 758296
rect 676090 758240 676292 758296
rect 676029 758238 676292 758240
rect 676029 758235 676095 758238
rect 672758 757828 672764 757892
rect 672828 757890 672834 757892
rect 672828 757830 676292 757890
rect 672828 757828 672834 757830
rect 40677 757754 40743 757757
rect 41454 757754 41460 757756
rect 40677 757752 41460 757754
rect 40677 757696 40682 757752
rect 40738 757696 41460 757752
rect 40677 757694 41460 757696
rect 40677 757691 40743 757694
rect 41454 757692 41460 757694
rect 41524 757692 41530 757756
rect 674741 757482 674807 757485
rect 674741 757480 676292 757482
rect 674741 757424 674746 757480
rect 674802 757424 676292 757480
rect 674741 757422 676292 757424
rect 674741 757419 674807 757422
rect 676070 757148 676076 757212
rect 676140 757210 676146 757212
rect 676140 757150 676322 757210
rect 676140 757148 676146 757150
rect 676262 757044 676322 757150
rect 679617 756802 679683 756805
rect 679574 756800 679683 756802
rect 679574 756744 679622 756800
rect 679678 756744 679683 756800
rect 679574 756739 679683 756744
rect 679574 756636 679634 756739
rect 42701 756532 42767 756533
rect 42701 756530 42748 756532
rect 42656 756528 42748 756530
rect 42656 756472 42706 756528
rect 42656 756470 42748 756472
rect 42701 756468 42748 756470
rect 42812 756468 42818 756532
rect 42701 756467 42767 756468
rect 675753 756258 675819 756261
rect 675753 756256 676292 756258
rect 675753 756200 675758 756256
rect 675814 756200 676292 756256
rect 675753 756198 676292 756200
rect 675753 756195 675819 756198
rect 676806 755924 676812 755988
rect 676876 755924 676882 755988
rect 676814 755820 676874 755924
rect 676213 755578 676279 755581
rect 676213 755576 676322 755578
rect 676213 755520 676218 755576
rect 676274 755520 676322 755576
rect 676213 755515 676322 755520
rect 676262 755412 676322 755515
rect 40902 755244 40908 755308
rect 40972 755306 40978 755308
rect 41822 755306 41828 755308
rect 40972 755246 41828 755306
rect 40972 755244 40978 755246
rect 41822 755244 41828 755246
rect 41892 755244 41898 755308
rect 676029 755034 676095 755037
rect 676029 755032 676292 755034
rect 676029 754976 676034 755032
rect 676090 754976 676292 755032
rect 676029 754974 676292 754976
rect 676029 754971 676095 754974
rect 676254 754700 676260 754764
rect 676324 754700 676330 754764
rect 676262 754596 676322 754700
rect 62113 754354 62179 754357
rect 676213 754354 676279 754357
rect 62113 754352 64492 754354
rect 62113 754296 62118 754352
rect 62174 754296 64492 754352
rect 62113 754294 64492 754296
rect 676213 754352 676322 754354
rect 676213 754296 676218 754352
rect 676274 754296 676322 754352
rect 62113 754291 62179 754294
rect 676213 754291 676322 754296
rect 676262 754188 676322 754291
rect 676029 753810 676095 753813
rect 676029 753808 676292 753810
rect 676029 753752 676034 753808
rect 676090 753752 676292 753808
rect 676029 753750 676292 753752
rect 676029 753747 676095 753750
rect 676438 753476 676444 753540
rect 676508 753476 676514 753540
rect 676446 753372 676506 753476
rect 41781 753132 41847 753133
rect 41781 753128 41828 753132
rect 41892 753130 41898 753132
rect 676213 753130 676279 753133
rect 41781 753072 41786 753128
rect 41781 753068 41828 753072
rect 41892 753070 41938 753130
rect 676213 753128 676322 753130
rect 676213 753072 676218 753128
rect 676274 753072 676322 753128
rect 41892 753068 41898 753070
rect 41781 753067 41847 753068
rect 676213 753067 676322 753072
rect 676262 752964 676322 753067
rect 676213 752722 676279 752725
rect 676213 752720 676322 752722
rect 676213 752664 676218 752720
rect 676274 752664 676322 752720
rect 676213 752659 676322 752664
rect 676262 752556 676322 752659
rect 676213 752314 676279 752317
rect 676213 752312 676322 752314
rect 676213 752256 676218 752312
rect 676274 752256 676322 752312
rect 676213 752251 676322 752256
rect 676262 752148 676322 752251
rect 40718 751708 40724 751772
rect 40788 751770 40794 751772
rect 41781 751770 41847 751773
rect 40788 751768 41847 751770
rect 40788 751712 41786 751768
rect 41842 751712 41847 751768
rect 40788 751710 41847 751712
rect 40788 751708 40794 751710
rect 41781 751707 41847 751710
rect 676262 751501 676322 751740
rect 676213 751496 676322 751501
rect 676213 751440 676218 751496
rect 676274 751440 676322 751496
rect 676213 751438 676322 751440
rect 676213 751435 676279 751438
rect 683070 751093 683130 751332
rect 683070 751088 683179 751093
rect 683070 751032 683118 751088
rect 683174 751032 683179 751088
rect 683070 751030 683179 751032
rect 683113 751027 683179 751030
rect 683070 750516 683130 750924
rect 40534 750348 40540 750412
rect 40604 750410 40610 750412
rect 41781 750410 41847 750413
rect 40604 750408 41847 750410
rect 40604 750352 41786 750408
rect 41842 750352 41847 750408
rect 40604 750350 41847 750352
rect 40604 750348 40610 750350
rect 41781 750347 41847 750350
rect 683113 750274 683179 750277
rect 683070 750272 683179 750274
rect 683070 750216 683118 750272
rect 683174 750216 683179 750272
rect 683070 750211 683179 750216
rect 651557 750138 651623 750141
rect 650164 750136 651623 750138
rect 650164 750080 651562 750136
rect 651618 750080 651623 750136
rect 683070 750108 683130 750211
rect 650164 750078 651623 750080
rect 651557 750075 651623 750078
rect 42701 749324 42767 749325
rect 42701 749322 42748 749324
rect 42656 749320 42748 749322
rect 42656 749264 42706 749320
rect 42656 749262 42748 749264
rect 42701 749260 42748 749262
rect 42812 749260 42818 749324
rect 42701 749259 42767 749260
rect 41638 746540 41644 746604
rect 41708 746602 41714 746604
rect 42609 746602 42675 746605
rect 41708 746600 42675 746602
rect 41708 746544 42614 746600
rect 42670 746544 42675 746600
rect 41708 746542 42675 746544
rect 41708 746540 41714 746542
rect 42609 746539 42675 746542
rect 41454 742324 41460 742388
rect 41524 742386 41530 742388
rect 41781 742386 41847 742389
rect 41524 742384 41847 742386
rect 41524 742328 41786 742384
rect 41842 742328 41847 742384
rect 41524 742326 41847 742328
rect 41524 742324 41530 742326
rect 41781 742323 41847 742326
rect 675334 741644 675340 741708
rect 675404 741706 675410 741708
rect 675477 741706 675543 741709
rect 675404 741704 675543 741706
rect 675404 741648 675482 741704
rect 675538 741648 675543 741704
rect 675404 741646 675543 741648
rect 675404 741644 675410 741646
rect 675477 741643 675543 741646
rect 62113 741298 62179 741301
rect 62113 741296 64492 741298
rect 62113 741240 62118 741296
rect 62174 741240 64492 741296
rect 62113 741238 64492 741240
rect 62113 741235 62179 741238
rect 675753 739938 675819 739941
rect 675886 739938 675892 739940
rect 675753 739936 675892 739938
rect 675753 739880 675758 739936
rect 675814 739880 675892 739936
rect 675753 739878 675892 739880
rect 675753 739875 675819 739878
rect 675886 739876 675892 739878
rect 675956 739876 675962 739940
rect 675661 739260 675727 739261
rect 675661 739256 675708 739260
rect 675772 739258 675778 739260
rect 675661 739200 675666 739256
rect 675661 739196 675708 739200
rect 675772 739198 675818 739258
rect 675772 739196 675778 739198
rect 675661 739195 675727 739196
rect 6022 737753 63922 737782
rect 6022 736609 6150 737753
rect 6854 737749 63922 737753
rect 6854 736645 54235 737749
rect 55339 737729 63922 737749
rect 55339 736645 63339 737729
rect 6854 736625 63339 736645
rect 63883 736625 63922 737729
rect 651557 736810 651623 736813
rect 650164 736808 651623 736810
rect 650164 736752 651562 736808
rect 651618 736752 651623 736808
rect 650164 736750 651623 736752
rect 651557 736747 651623 736750
rect 6854 736609 63922 736625
rect 6022 736582 63922 736609
rect 7236 736157 62944 736182
rect 7236 735013 7348 736157
rect 8052 736131 62944 736157
rect 8052 735027 52641 736131
rect 53745 736121 62944 736131
rect 53745 735027 62371 736121
rect 8052 735017 62371 735027
rect 62915 735017 62944 736121
rect 8052 735013 62944 735017
rect 7236 734982 62944 735013
rect 675753 734362 675819 734365
rect 676806 734362 676812 734364
rect 675753 734360 676812 734362
rect 675753 734304 675758 734360
rect 675814 734304 676812 734360
rect 675753 734302 676812 734304
rect 675753 734299 675819 734302
rect 676806 734300 676812 734302
rect 676876 734300 676882 734364
rect 675753 733002 675819 733005
rect 676990 733002 676996 733004
rect 675753 733000 676996 733002
rect 675753 732944 675758 733000
rect 675814 732944 676996 733000
rect 675753 732942 676996 732944
rect 675753 732939 675819 732942
rect 676990 732940 676996 732942
rect 677060 732940 677066 733004
rect 31526 731101 31586 731340
rect 31477 731096 31586 731101
rect 31477 731040 31482 731096
rect 31538 731040 31586 731096
rect 31477 731038 31586 731040
rect 31661 731098 31727 731101
rect 31661 731096 31770 731098
rect 31661 731040 31666 731096
rect 31722 731040 31770 731096
rect 31477 731035 31543 731038
rect 31661 731035 31770 731040
rect 31710 730932 31770 731035
rect 31569 730690 31635 730693
rect 31526 730688 31635 730690
rect 31526 730632 31574 730688
rect 31630 730632 31635 730688
rect 31526 730627 31635 730632
rect 31526 730524 31586 730627
rect 31385 730282 31451 730285
rect 31342 730280 31451 730282
rect 31342 730224 31390 730280
rect 31446 730224 31451 730280
rect 31342 730219 31451 730224
rect 31342 730116 31402 730219
rect 40174 729468 40234 729708
rect 40166 729404 40172 729468
rect 40236 729404 40242 729468
rect 42793 729330 42859 729333
rect 41492 729328 42859 729330
rect 41492 729272 42798 729328
rect 42854 729272 42859 729328
rect 41492 729270 42859 729272
rect 42793 729267 42859 729270
rect 44173 728922 44239 728925
rect 41492 728920 44239 728922
rect 41492 728864 44178 728920
rect 44234 728864 44239 728920
rect 41492 728862 44239 728864
rect 44173 728859 44239 728862
rect 39982 728588 39988 728652
rect 40052 728588 40058 728652
rect 39990 728484 40050 728588
rect 62113 728242 62179 728245
rect 62113 728240 64492 728242
rect 62113 728184 62118 728240
rect 62174 728184 64492 728240
rect 62113 728182 64492 728184
rect 62113 728179 62179 728182
rect 39990 727836 40050 728076
rect 39982 727772 39988 727836
rect 40052 727772 40058 727836
rect 44633 727698 44699 727701
rect 41492 727696 44699 727698
rect 41492 727640 44638 727696
rect 44694 727640 44699 727696
rect 41492 727638 44699 727640
rect 44633 727635 44699 727638
rect 42793 727290 42859 727293
rect 41492 727288 42859 727290
rect 41492 727232 42798 727288
rect 42854 727232 42859 727288
rect 41492 727230 42859 727232
rect 42793 727227 42859 727230
rect 675150 727228 675156 727292
rect 675220 727290 675226 727292
rect 678237 727290 678303 727293
rect 675220 727288 678303 727290
rect 675220 727232 678242 727288
rect 678298 727232 678303 727288
rect 675220 727230 678303 727232
rect 675220 727228 675226 727230
rect 678237 727227 678303 727230
rect 30974 726613 31034 726852
rect 30974 726608 31083 726613
rect 30974 726552 31022 726608
rect 31078 726552 31083 726608
rect 30974 726550 31083 726552
rect 31017 726547 31083 726550
rect 40726 726205 40786 726444
rect 40677 726200 40786 726205
rect 40677 726144 40682 726200
rect 40738 726144 40786 726200
rect 40677 726142 40786 726144
rect 40677 726139 40743 726142
rect 41454 726140 41460 726204
rect 41524 726140 41530 726204
rect 41462 726036 41522 726140
rect 33734 725389 33794 725628
rect 33734 725384 33843 725389
rect 33734 725328 33782 725384
rect 33838 725328 33843 725384
rect 33734 725326 33843 725328
rect 33777 725323 33843 725326
rect 42149 725250 42215 725253
rect 41492 725248 42215 725250
rect 41492 725192 42154 725248
rect 42210 725192 42215 725248
rect 41492 725190 42215 725192
rect 42149 725187 42215 725190
rect 40910 724573 40970 724812
rect 40861 724568 40970 724573
rect 40861 724512 40866 724568
rect 40922 724512 40970 724568
rect 40861 724510 40970 724512
rect 40861 724507 40927 724510
rect 42885 724434 42951 724437
rect 41492 724432 42951 724434
rect 41492 724376 42890 724432
rect 42946 724376 42951 724432
rect 41492 724374 42951 724376
rect 42885 724371 42951 724374
rect 42057 724026 42123 724029
rect 41492 724024 42123 724026
rect 41492 723968 42062 724024
rect 42118 723968 42123 724024
rect 41492 723966 42123 723968
rect 42057 723963 42123 723966
rect 34470 723349 34530 723588
rect 652017 723482 652083 723485
rect 650164 723480 652083 723482
rect 650164 723424 652022 723480
rect 652078 723424 652083 723480
rect 650164 723422 652083 723424
rect 652017 723419 652083 723422
rect 34421 723344 34530 723349
rect 40769 723346 40835 723349
rect 34421 723288 34426 723344
rect 34482 723288 34530 723344
rect 34421 723286 34530 723288
rect 40726 723344 40835 723346
rect 40726 723288 40774 723344
rect 40830 723288 40835 723344
rect 34421 723283 34487 723286
rect 40726 723283 40835 723288
rect 40726 723180 40786 723283
rect 44541 722802 44607 722805
rect 41492 722800 44607 722802
rect 41492 722744 44546 722800
rect 44602 722744 44607 722800
rect 41492 722742 44607 722744
rect 44541 722739 44607 722742
rect 42977 722394 43043 722397
rect 41492 722392 43043 722394
rect 41492 722336 42982 722392
rect 43038 722336 43043 722392
rect 41492 722334 43043 722336
rect 42977 722331 43043 722334
rect 44357 721986 44423 721989
rect 41492 721984 44423 721986
rect 41492 721928 44362 721984
rect 44418 721928 44423 721984
rect 41492 721926 44423 721928
rect 44357 721923 44423 721926
rect 40542 721308 40602 721548
rect 40534 721244 40540 721308
rect 40604 721244 40610 721308
rect 41462 720901 41522 721140
rect 41462 720896 41571 720901
rect 41462 720840 41510 720896
rect 41566 720840 41571 720896
rect 41462 720838 41571 720840
rect 41505 720835 41571 720838
rect 27662 720324 27722 720732
rect 41462 719677 41522 719916
rect 41462 719672 41571 719677
rect 41462 719616 41510 719672
rect 41566 719616 41571 719672
rect 41462 719614 41571 719616
rect 41505 719611 41571 719614
rect 676029 716546 676095 716549
rect 676029 716544 676292 716546
rect 676029 716488 676034 716544
rect 676090 716488 676292 716544
rect 676029 716486 676292 716488
rect 676029 716483 676095 716486
rect 676029 716138 676095 716141
rect 676029 716136 676292 716138
rect 676029 716080 676034 716136
rect 676090 716080 676292 716136
rect 676029 716078 676292 716080
rect 676029 716075 676095 716078
rect 676029 715730 676095 715733
rect 676029 715728 676292 715730
rect 676029 715672 676034 715728
rect 676090 715672 676292 715728
rect 676029 715670 676292 715672
rect 676029 715667 676095 715670
rect 33777 715594 33843 715597
rect 41822 715594 41828 715596
rect 33777 715592 41828 715594
rect 33777 715536 33782 715592
rect 33838 715536 41828 715592
rect 33777 715534 41828 715536
rect 33777 715531 33843 715534
rect 41822 715532 41828 715534
rect 41892 715532 41898 715596
rect 31017 715458 31083 715461
rect 41638 715458 41644 715460
rect 31017 715456 41644 715458
rect 31017 715400 31022 715456
rect 31078 715400 41644 715456
rect 31017 715398 41644 715400
rect 31017 715395 31083 715398
rect 41638 715396 41644 715398
rect 41708 715396 41714 715460
rect 62113 715322 62179 715325
rect 675937 715322 676003 715325
rect 62113 715320 64492 715322
rect 62113 715264 62118 715320
rect 62174 715264 64492 715320
rect 62113 715262 64492 715264
rect 675937 715320 676292 715322
rect 675937 715264 675942 715320
rect 675998 715264 676292 715320
rect 675937 715262 676292 715264
rect 62113 715259 62179 715262
rect 675937 715259 676003 715262
rect 676029 714914 676095 714917
rect 676029 714912 676292 714914
rect 676029 714856 676034 714912
rect 676090 714856 676292 714912
rect 676029 714854 676292 714856
rect 676029 714851 676095 714854
rect 676029 714506 676095 714509
rect 676029 714504 676292 714506
rect 676029 714448 676034 714504
rect 676090 714448 676292 714504
rect 676029 714446 676292 714448
rect 676029 714443 676095 714446
rect 40769 714098 40835 714101
rect 40902 714098 40908 714100
rect 40769 714096 40908 714098
rect 40769 714040 40774 714096
rect 40830 714040 40908 714096
rect 40769 714038 40908 714040
rect 40769 714035 40835 714038
rect 40902 714036 40908 714038
rect 40972 714036 40978 714100
rect 676029 714098 676095 714101
rect 676029 714096 676292 714098
rect 676029 714040 676034 714096
rect 676090 714040 676292 714096
rect 676029 714038 676292 714040
rect 676029 714035 676095 714038
rect 42057 713828 42123 713829
rect 42006 713826 42012 713828
rect 41966 713766 42012 713826
rect 42076 713824 42123 713828
rect 42118 713768 42123 713824
rect 42006 713764 42012 713766
rect 42076 713764 42123 713768
rect 42057 713763 42123 713764
rect 676029 713690 676095 713693
rect 676029 713688 676292 713690
rect 676029 713632 676034 713688
rect 676090 713632 676292 713688
rect 676029 713630 676292 713632
rect 676029 713627 676095 713630
rect 677317 713492 677383 713493
rect 677317 713488 677364 713492
rect 677428 713490 677434 713492
rect 677317 713432 677322 713488
rect 677317 713428 677364 713432
rect 677428 713430 677474 713490
rect 677428 713428 677434 713430
rect 677317 713427 677383 713428
rect 42190 713220 42196 713284
rect 42260 713282 42266 713284
rect 42425 713282 42491 713285
rect 42260 713280 42491 713282
rect 42260 713224 42430 713280
rect 42486 713224 42491 713280
rect 42260 713222 42491 713224
rect 42260 713220 42266 713222
rect 42425 713219 42491 713222
rect 676029 713282 676095 713285
rect 676029 713280 676292 713282
rect 676029 713224 676034 713280
rect 676090 713224 676292 713280
rect 676029 713222 676292 713224
rect 676029 713219 676095 713222
rect 674741 712874 674807 712877
rect 674741 712872 676292 712874
rect 674741 712816 674746 712872
rect 674802 712816 676292 712872
rect 674741 712814 676292 712816
rect 674741 712811 674807 712814
rect 676029 712466 676095 712469
rect 676029 712464 676292 712466
rect 676029 712408 676034 712464
rect 676090 712408 676292 712464
rect 676029 712406 676292 712408
rect 676029 712403 676095 712406
rect 42374 712268 42380 712332
rect 42444 712330 42450 712332
rect 42517 712330 42583 712333
rect 42444 712328 42583 712330
rect 42444 712272 42522 712328
rect 42578 712272 42583 712328
rect 42444 712270 42583 712272
rect 42444 712268 42450 712270
rect 42517 712267 42583 712270
rect 676029 712058 676095 712061
rect 676029 712056 676292 712058
rect 676029 712000 676034 712056
rect 676090 712000 676292 712056
rect 676029 711998 676292 712000
rect 676029 711995 676095 711998
rect 42149 711788 42215 711789
rect 42149 711786 42196 711788
rect 42104 711784 42196 711786
rect 42104 711728 42154 711784
rect 42104 711726 42196 711728
rect 42149 711724 42196 711726
rect 42260 711724 42266 711788
rect 42149 711723 42215 711724
rect 678237 711650 678303 711653
rect 678237 711648 678316 711650
rect 678237 711592 678242 711648
rect 678298 711592 678316 711648
rect 678237 711590 678316 711592
rect 678237 711587 678303 711590
rect 676029 711242 676095 711245
rect 676029 711240 676292 711242
rect 676029 711184 676034 711240
rect 676090 711184 676292 711240
rect 676029 711182 676292 711184
rect 676029 711179 676095 711182
rect 675937 711106 676003 711109
rect 676070 711106 676076 711108
rect 675937 711104 676076 711106
rect 675937 711048 675942 711104
rect 675998 711048 676076 711104
rect 675937 711046 676076 711048
rect 675937 711043 676003 711046
rect 676070 711044 676076 711046
rect 676140 711044 676146 711108
rect 40534 710772 40540 710836
rect 40604 710834 40610 710836
rect 42517 710834 42583 710837
rect 40604 710832 42583 710834
rect 40604 710776 42522 710832
rect 42578 710776 42583 710832
rect 40604 710774 42583 710776
rect 40604 710772 40610 710774
rect 42517 710771 42583 710774
rect 675518 710772 675524 710836
rect 675588 710834 675594 710836
rect 675588 710774 676292 710834
rect 675588 710772 675594 710774
rect 676029 710426 676095 710429
rect 676029 710424 676292 710426
rect 676029 710368 676034 710424
rect 676090 710368 676292 710424
rect 676029 710366 676292 710368
rect 676029 710363 676095 710366
rect 651557 710290 651623 710293
rect 650164 710288 651623 710290
rect 650164 710232 651562 710288
rect 651618 710232 651623 710288
rect 650164 710230 651623 710232
rect 651557 710227 651623 710230
rect 676029 710018 676095 710021
rect 676029 710016 676292 710018
rect 676029 709960 676034 710016
rect 676090 709960 676292 710016
rect 676029 709958 676292 709960
rect 676029 709955 676095 709958
rect 40902 709820 40908 709884
rect 40972 709882 40978 709884
rect 41781 709882 41847 709885
rect 40972 709880 41847 709882
rect 40972 709824 41786 709880
rect 41842 709824 41847 709880
rect 40972 709822 41847 709824
rect 40972 709820 40978 709822
rect 41781 709819 41847 709822
rect 676029 709610 676095 709613
rect 676029 709608 676292 709610
rect 676029 709552 676034 709608
rect 676090 709552 676292 709608
rect 676029 709550 676292 709552
rect 676029 709547 676095 709550
rect 676029 709202 676095 709205
rect 676029 709200 676292 709202
rect 676029 709144 676034 709200
rect 676090 709144 676292 709200
rect 676029 709142 676292 709144
rect 676029 709139 676095 709142
rect 676070 708868 676076 708932
rect 676140 708868 676146 708932
rect 676078 708794 676138 708868
rect 676078 708734 676292 708794
rect 42374 708460 42380 708524
rect 42444 708522 42450 708524
rect 42517 708522 42583 708525
rect 42444 708520 42583 708522
rect 42444 708464 42522 708520
rect 42578 708464 42583 708520
rect 42444 708462 42583 708464
rect 42444 708460 42450 708462
rect 42517 708459 42583 708462
rect 676029 708386 676095 708389
rect 676029 708384 676292 708386
rect 676029 708328 676034 708384
rect 676090 708328 676292 708384
rect 676029 708326 676292 708328
rect 676029 708323 676095 708326
rect 676029 707978 676095 707981
rect 676029 707976 676292 707978
rect 676029 707920 676034 707976
rect 676090 707920 676292 707976
rect 676029 707918 676292 707920
rect 676029 707915 676095 707918
rect 676029 707570 676095 707573
rect 676029 707568 676292 707570
rect 676029 707512 676034 707568
rect 676090 707512 676292 707568
rect 676029 707510 676292 707512
rect 676029 707507 676095 707510
rect 676029 707162 676095 707165
rect 676029 707160 676292 707162
rect 676029 707104 676034 707160
rect 676090 707104 676292 707160
rect 676029 707102 676292 707104
rect 676029 707099 676095 707102
rect 676029 706754 676095 706757
rect 676029 706752 676292 706754
rect 676029 706696 676034 706752
rect 676090 706696 676292 706752
rect 676029 706694 676292 706696
rect 676029 706691 676095 706694
rect 42006 706556 42012 706620
rect 42076 706618 42082 706620
rect 42517 706618 42583 706621
rect 42076 706616 42583 706618
rect 42076 706560 42522 706616
rect 42578 706560 42583 706616
rect 42076 706558 42583 706560
rect 42076 706556 42082 706558
rect 42517 706555 42583 706558
rect 676029 706346 676095 706349
rect 676029 706344 676292 706346
rect 676029 706288 676034 706344
rect 676090 706288 676292 706344
rect 676029 706286 676292 706288
rect 676029 706283 676095 706286
rect 685830 705500 685890 705908
rect 676029 705122 676095 705125
rect 676029 705120 676292 705122
rect 676029 705064 676034 705120
rect 676090 705064 676292 705120
rect 676029 705062 676292 705064
rect 676029 705059 676095 705062
rect 41822 704924 41828 704988
rect 41892 704986 41898 704988
rect 42241 704986 42307 704989
rect 41892 704984 42307 704986
rect 41892 704928 42246 704984
rect 42302 704928 42307 704984
rect 41892 704926 42307 704928
rect 41892 704924 41898 704926
rect 42241 704923 42307 704926
rect 675937 704442 676003 704445
rect 676254 704442 676260 704444
rect 675937 704440 676260 704442
rect 675937 704384 675942 704440
rect 675998 704384 676260 704440
rect 675937 704382 676260 704384
rect 675937 704379 676003 704382
rect 676254 704380 676260 704382
rect 676324 704380 676330 704444
rect 41638 702884 41644 702948
rect 41708 702946 41714 702948
rect 42425 702946 42491 702949
rect 41708 702944 42491 702946
rect 41708 702888 42430 702944
rect 42486 702888 42491 702944
rect 41708 702886 42491 702888
rect 41708 702884 41714 702886
rect 42425 702883 42491 702886
rect 62757 702266 62823 702269
rect 62757 702264 64492 702266
rect 62757 702208 62762 702264
rect 62818 702208 64492 702264
rect 62757 702206 64492 702208
rect 62757 702203 62823 702206
rect 41454 699348 41460 699412
rect 41524 699410 41530 699412
rect 41781 699410 41847 699413
rect 41524 699408 41847 699410
rect 41524 699352 41786 699408
rect 41842 699352 41847 699408
rect 41524 699350 41847 699352
rect 41524 699348 41530 699350
rect 41781 699347 41847 699350
rect 674598 697308 674604 697372
rect 674668 697370 674674 697372
rect 675385 697370 675451 697373
rect 674668 697368 675451 697370
rect 674668 697312 675390 697368
rect 675446 697312 675451 697368
rect 674668 697310 675451 697312
rect 674668 697308 674674 697310
rect 675385 697307 675451 697310
rect 652017 696962 652083 696965
rect 650164 696960 652083 696962
rect 650164 696904 652022 696960
rect 652078 696904 652083 696960
rect 650164 696902 652083 696904
rect 652017 696899 652083 696902
rect 675661 696964 675727 696965
rect 675661 696960 675708 696964
rect 675772 696962 675778 696964
rect 675661 696904 675666 696960
rect 675661 696900 675708 696904
rect 675772 696902 675818 696962
rect 675772 696900 675778 696902
rect 675661 696899 675727 696900
rect 675753 695058 675819 695061
rect 676070 695058 676076 695060
rect 675753 695056 676076 695058
rect 675753 695000 675758 695056
rect 675814 695000 676076 695056
rect 675753 694998 676076 695000
rect 675753 694995 675819 694998
rect 676070 694996 676076 694998
rect 676140 694996 676146 695060
rect 6022 694553 63922 694582
rect 6022 693409 6150 694553
rect 6854 694549 63922 694553
rect 6854 693445 54235 694549
rect 55339 694529 63922 694549
rect 55339 693445 63339 694529
rect 6854 693425 63339 693445
rect 63883 693425 63922 694529
rect 675753 694242 675819 694245
rect 676438 694242 676444 694244
rect 675753 694240 676444 694242
rect 675753 694184 675758 694240
rect 675814 694184 676444 694240
rect 675753 694182 676444 694184
rect 675753 694179 675819 694182
rect 676438 694180 676444 694182
rect 676508 694180 676514 694244
rect 6854 693409 63922 693425
rect 6022 693382 63922 693409
rect 7236 692957 62944 692982
rect 7236 691813 7348 692957
rect 8052 692931 62944 692957
rect 8052 691827 52641 692931
rect 53745 692921 62944 692931
rect 53745 691827 62371 692921
rect 8052 691817 62371 691827
rect 62915 691817 62944 692921
rect 8052 691813 62944 691817
rect 7236 691782 62944 691813
rect 62113 689210 62179 689213
rect 62113 689208 64492 689210
rect 62113 689152 62118 689208
rect 62174 689152 64492 689208
rect 62113 689150 64492 689152
rect 62113 689147 62179 689150
rect 35617 688394 35683 688397
rect 35574 688392 35683 688394
rect 35574 688336 35622 688392
rect 35678 688336 35683 688392
rect 35574 688331 35683 688336
rect 35574 688092 35634 688331
rect 35801 687714 35867 687717
rect 35788 687712 35867 687714
rect 35788 687656 35806 687712
rect 35862 687656 35867 687712
rect 35788 687654 35867 687656
rect 35801 687651 35867 687654
rect 35709 687306 35775 687309
rect 35709 687304 35788 687306
rect 35709 687248 35714 687304
rect 35770 687248 35788 687304
rect 35709 687246 35788 687248
rect 35709 687243 35775 687246
rect 40166 687108 40172 687172
rect 40236 687108 40242 687172
rect 40174 686868 40234 687108
rect 44265 686490 44331 686493
rect 41492 686488 44331 686490
rect 41492 686432 44270 686488
rect 44326 686432 44331 686488
rect 41492 686430 44331 686432
rect 44265 686427 44331 686430
rect 44173 686082 44239 686085
rect 41492 686080 44239 686082
rect 41492 686024 44178 686080
rect 44234 686024 44239 686080
rect 41492 686022 44239 686024
rect 44173 686019 44239 686022
rect 44173 685674 44239 685677
rect 41492 685672 44239 685674
rect 41492 685616 44178 685672
rect 44234 685616 44239 685672
rect 41492 685614 44239 685616
rect 44173 685611 44239 685614
rect 39982 685476 39988 685540
rect 40052 685476 40058 685540
rect 39990 685236 40050 685476
rect 39990 684724 40050 684828
rect 39982 684660 39988 684724
rect 40052 684660 40058 684724
rect 42793 684450 42859 684453
rect 41492 684448 42859 684450
rect 41492 684392 42798 684448
rect 42854 684392 42859 684448
rect 41492 684390 42859 684392
rect 42793 684387 42859 684390
rect 42793 684042 42859 684045
rect 41492 684040 42859 684042
rect 41492 683984 42798 684040
rect 42854 683984 42859 684040
rect 41492 683982 42859 683984
rect 42793 683979 42859 683982
rect 39297 683634 39363 683637
rect 651833 683634 651899 683637
rect 39284 683632 39363 683634
rect 39284 683576 39302 683632
rect 39358 683576 39363 683632
rect 39284 683574 39363 683576
rect 650164 683632 651899 683634
rect 650164 683576 651838 683632
rect 651894 683576 651899 683632
rect 650164 683574 651899 683576
rect 39297 683571 39363 683574
rect 651833 683571 651899 683574
rect 41462 683090 41522 683196
rect 41689 683090 41755 683093
rect 41462 683088 41755 683090
rect 41462 683032 41694 683088
rect 41750 683032 41755 683088
rect 41462 683030 41755 683032
rect 41689 683027 41755 683030
rect 32397 682818 32463 682821
rect 32397 682816 32476 682818
rect 32397 682760 32402 682816
rect 32458 682760 32476 682816
rect 32397 682758 32476 682760
rect 32397 682755 32463 682758
rect 41462 682276 41522 682380
rect 41454 682212 41460 682276
rect 41524 682212 41530 682276
rect 41462 681866 41522 681972
rect 41689 681866 41755 681869
rect 41462 681864 41755 681866
rect 41462 681808 41694 681864
rect 41750 681808 41755 681864
rect 41462 681806 41755 681808
rect 41689 681803 41755 681806
rect 31017 681594 31083 681597
rect 31004 681592 31083 681594
rect 31004 681536 31022 681592
rect 31078 681536 31083 681592
rect 31004 681534 31083 681536
rect 31017 681531 31083 681534
rect 44357 681186 44423 681189
rect 41492 681184 44423 681186
rect 41492 681128 44362 681184
rect 44418 681128 44423 681184
rect 41492 681126 44423 681128
rect 44357 681123 44423 681126
rect 41965 680778 42031 680781
rect 41492 680776 42031 680778
rect 41492 680720 41970 680776
rect 42026 680720 42031 680776
rect 41492 680718 42031 680720
rect 41965 680715 42031 680718
rect 35157 680370 35223 680373
rect 35157 680368 35236 680370
rect 35157 680312 35162 680368
rect 35218 680312 35236 680368
rect 35157 680310 35236 680312
rect 35157 680307 35223 680310
rect 44449 679962 44515 679965
rect 41492 679960 44515 679962
rect 41492 679904 44454 679960
rect 44510 679904 44515 679960
rect 41492 679902 44515 679904
rect 44449 679899 44515 679902
rect 40542 679420 40602 679524
rect 40534 679356 40540 679420
rect 40604 679356 40610 679420
rect 42885 679146 42951 679149
rect 41492 679144 42951 679146
rect 41492 679088 42890 679144
rect 42946 679088 42951 679144
rect 41492 679086 42951 679088
rect 42885 679083 42951 679086
rect 675334 678948 675340 679012
rect 675404 679010 675410 679012
rect 678237 679010 678303 679013
rect 675404 679008 678303 679010
rect 675404 678952 678242 679008
rect 678298 678952 678303 679008
rect 675404 678950 678303 678952
rect 675404 678948 675410 678950
rect 678237 678947 678303 678950
rect 42977 678738 43043 678741
rect 41492 678736 43043 678738
rect 41492 678680 42982 678736
rect 43038 678680 43043 678736
rect 41492 678678 43043 678680
rect 42977 678675 43043 678678
rect 40726 678196 40786 678300
rect 40718 678132 40724 678196
rect 40788 678132 40794 678196
rect 30606 677788 30666 677892
rect 30598 677724 30604 677788
rect 30668 677724 30674 677788
rect 27662 677076 27722 677484
rect 30465 676868 30531 676871
rect 30422 676866 30531 676868
rect 30422 676810 30470 676866
rect 30526 676810 30531 676866
rect 30422 676805 30531 676810
rect 30422 676698 30482 676805
rect 30422 676668 30636 676698
rect 30452 676638 30666 676668
rect 30606 676564 30666 676638
rect 30598 676500 30604 676564
rect 30668 676500 30674 676564
rect 62113 676154 62179 676157
rect 62113 676152 64492 676154
rect 62113 676096 62118 676152
rect 62174 676096 64492 676152
rect 62113 676094 64492 676096
rect 62113 676091 62179 676094
rect 32397 671394 32463 671397
rect 41638 671394 41644 671396
rect 32397 671392 41644 671394
rect 32397 671336 32402 671392
rect 32458 671336 41644 671392
rect 32397 671334 41644 671336
rect 32397 671331 32463 671334
rect 41638 671332 41644 671334
rect 41708 671332 41714 671396
rect 676262 671125 676322 671364
rect 676213 671120 676322 671125
rect 676213 671064 676218 671120
rect 676274 671064 676322 671120
rect 676213 671062 676322 671064
rect 676213 671059 676279 671062
rect 39297 670986 39363 670989
rect 41822 670986 41828 670988
rect 39297 670984 41828 670986
rect 39297 670928 39302 670984
rect 39358 670928 41828 670984
rect 39297 670926 41828 670928
rect 39297 670923 39363 670926
rect 41822 670924 41828 670926
rect 41892 670924 41898 670988
rect 676029 670986 676095 670989
rect 676029 670984 676292 670986
rect 676029 670928 676034 670984
rect 676090 670928 676292 670984
rect 676029 670926 676292 670928
rect 676029 670923 676095 670926
rect 42057 670716 42123 670717
rect 42006 670652 42012 670716
rect 42076 670714 42123 670716
rect 42076 670712 42168 670714
rect 42118 670656 42168 670712
rect 42076 670654 42168 670656
rect 42076 670652 42123 670654
rect 42057 670651 42123 670652
rect 651557 670442 651623 670445
rect 650164 670440 651623 670442
rect 650164 670384 651562 670440
rect 651618 670384 651623 670440
rect 650164 670382 651623 670384
rect 651557 670379 651623 670382
rect 676262 670309 676322 670548
rect 676262 670304 676371 670309
rect 676262 670248 676310 670304
rect 676366 670248 676371 670304
rect 676262 670246 676371 670248
rect 676305 670243 676371 670246
rect 42190 670108 42196 670172
rect 42260 670170 42266 670172
rect 42425 670170 42491 670173
rect 42260 670168 42491 670170
rect 42260 670112 42430 670168
rect 42486 670112 42491 670168
rect 42260 670110 42491 670112
rect 42260 670108 42266 670110
rect 42425 670107 42491 670110
rect 676121 669898 676187 669901
rect 676262 669898 676322 670140
rect 676121 669896 676322 669898
rect 676121 669840 676126 669896
rect 676182 669840 676322 669896
rect 676121 669838 676322 669840
rect 676121 669835 676187 669838
rect 674741 669762 674807 669765
rect 674741 669760 676292 669762
rect 674741 669704 674746 669760
rect 674802 669704 676292 669760
rect 674741 669702 676292 669704
rect 674741 669699 674807 669702
rect 42701 669490 42767 669493
rect 42566 669488 42767 669490
rect 42566 669432 42706 669488
rect 42762 669432 42767 669488
rect 42566 669430 42767 669432
rect 42057 668538 42123 668541
rect 42566 668538 42626 669430
rect 42701 669427 42767 669430
rect 676213 669490 676279 669493
rect 676213 669488 676322 669490
rect 676213 669432 676218 669488
rect 676274 669432 676322 669488
rect 676213 669427 676322 669432
rect 676262 669324 676322 669427
rect 676029 668946 676095 668949
rect 676029 668944 676292 668946
rect 676029 668888 676034 668944
rect 676090 668888 676292 668944
rect 676029 668886 676292 668888
rect 676029 668883 676095 668886
rect 676213 668674 676279 668677
rect 676213 668672 676322 668674
rect 676213 668616 676218 668672
rect 676274 668616 676322 668672
rect 676213 668611 676322 668616
rect 42057 668536 42626 668538
rect 42057 668480 42062 668536
rect 42118 668480 42626 668536
rect 676262 668508 676322 668611
rect 42057 668478 42626 668480
rect 42057 668475 42123 668478
rect 676029 668130 676095 668133
rect 676029 668128 676292 668130
rect 676029 668072 676034 668128
rect 676090 668072 676292 668128
rect 676029 668070 676292 668072
rect 676029 668067 676095 668070
rect 676213 667858 676279 667861
rect 676213 667856 676322 667858
rect 676213 667800 676218 667856
rect 676274 667800 676322 667856
rect 676213 667795 676322 667800
rect 676262 667692 676322 667795
rect 676262 667045 676322 667284
rect 676213 667040 676322 667045
rect 676213 666984 676218 667040
rect 676274 666984 676322 667040
rect 676213 666982 676322 666984
rect 678237 667042 678303 667045
rect 678237 667040 678346 667042
rect 678237 666984 678242 667040
rect 678298 666984 678346 667040
rect 676213 666979 676279 666982
rect 678237 666979 678346 666984
rect 678286 666876 678346 666979
rect 676029 666498 676095 666501
rect 676029 666496 676292 666498
rect 676029 666440 676034 666496
rect 676090 666440 676292 666496
rect 676029 666438 676292 666440
rect 676029 666435 676095 666438
rect 676262 665821 676322 666060
rect 676213 665816 676322 665821
rect 676213 665760 676218 665816
rect 676274 665760 676322 665816
rect 676213 665758 676322 665760
rect 676213 665755 676279 665758
rect 675886 665620 675892 665684
rect 675956 665682 675962 665684
rect 675956 665622 676292 665682
rect 675956 665620 675962 665622
rect 40718 665348 40724 665412
rect 40788 665410 40794 665412
rect 41781 665410 41847 665413
rect 40788 665408 41847 665410
rect 40788 665352 41786 665408
rect 41842 665352 41847 665408
rect 40788 665350 41847 665352
rect 40788 665348 40794 665350
rect 41781 665347 41847 665350
rect 676029 665274 676095 665277
rect 676029 665272 676292 665274
rect 676029 665216 676034 665272
rect 676090 665216 676292 665272
rect 676029 665214 676292 665216
rect 676029 665211 676095 665214
rect 676213 665002 676279 665005
rect 676213 665000 676322 665002
rect 676213 664944 676218 665000
rect 676274 664944 676322 665000
rect 676213 664939 676322 664944
rect 676262 664836 676322 664939
rect 40534 664532 40540 664596
rect 40604 664594 40610 664596
rect 41781 664594 41847 664597
rect 40604 664592 41847 664594
rect 40604 664536 41786 664592
rect 41842 664536 41847 664592
rect 40604 664534 41847 664536
rect 40604 664532 40610 664534
rect 41781 664531 41847 664534
rect 676262 664189 676322 664428
rect 676213 664184 676322 664189
rect 676213 664128 676218 664184
rect 676274 664128 676322 664184
rect 676213 664126 676322 664128
rect 676213 664123 676279 664126
rect 676262 663781 676322 664020
rect 676213 663776 676322 663781
rect 676213 663720 676218 663776
rect 676274 663720 676322 663776
rect 676213 663718 676322 663720
rect 676213 663715 676279 663718
rect 42057 663372 42123 663373
rect 676262 663372 676322 663612
rect 42006 663370 42012 663372
rect 41966 663310 42012 663370
rect 42076 663368 42123 663372
rect 42118 663312 42123 663368
rect 42006 663308 42012 663310
rect 42076 663308 42123 663312
rect 676254 663308 676260 663372
rect 676324 663308 676330 663372
rect 676990 663308 676996 663372
rect 677060 663308 677066 663372
rect 42057 663307 42123 663308
rect 676998 663204 677058 663308
rect 62113 663098 62179 663101
rect 62113 663096 64492 663098
rect 62113 663040 62118 663096
rect 62174 663040 64492 663096
rect 62113 663038 64492 663040
rect 62113 663035 62179 663038
rect 676806 662900 676812 662964
rect 676876 662900 676882 662964
rect 676814 662796 676874 662900
rect 676029 662418 676095 662421
rect 676029 662416 676292 662418
rect 676029 662360 676034 662416
rect 676090 662360 676292 662416
rect 676029 662358 676292 662360
rect 676029 662355 676095 662358
rect 676262 661741 676322 661980
rect 676213 661736 676322 661741
rect 676213 661680 676218 661736
rect 676274 661680 676322 661736
rect 676213 661678 676322 661680
rect 676213 661675 676279 661678
rect 676029 661602 676095 661605
rect 676029 661600 676292 661602
rect 676029 661544 676034 661600
rect 676090 661544 676292 661600
rect 676029 661542 676292 661544
rect 676029 661539 676095 661542
rect 41454 661268 41460 661332
rect 41524 661330 41530 661332
rect 42701 661330 42767 661333
rect 41524 661328 42767 661330
rect 41524 661272 42706 661328
rect 42762 661272 42767 661328
rect 41524 661270 42767 661272
rect 41524 661268 41530 661270
rect 42701 661267 42767 661270
rect 683070 660925 683130 661164
rect 683070 660920 683179 660925
rect 683070 660864 683118 660920
rect 683174 660864 683179 660920
rect 683070 660862 683179 660864
rect 683113 660859 683179 660862
rect 42149 660516 42215 660517
rect 42149 660514 42196 660516
rect 42104 660512 42196 660514
rect 42104 660456 42154 660512
rect 42104 660454 42196 660456
rect 42149 660452 42196 660454
rect 42260 660452 42266 660516
rect 42149 660451 42215 660452
rect 41822 660316 41828 660380
rect 41892 660378 41898 660380
rect 42517 660378 42583 660381
rect 41892 660376 42583 660378
rect 41892 660320 42522 660376
rect 42578 660320 42583 660376
rect 685830 660348 685890 660756
rect 41892 660318 42583 660320
rect 41892 660316 41898 660318
rect 42517 660315 42583 660318
rect 683113 660106 683179 660109
rect 683070 660104 683179 660106
rect 683070 660048 683118 660104
rect 683174 660048 683179 660104
rect 683070 660043 683179 660048
rect 673862 659908 673868 659972
rect 673932 659970 673938 659972
rect 683070 659970 683130 660043
rect 673932 659940 683130 659970
rect 673932 659910 683100 659940
rect 673932 659908 673938 659910
rect 41638 658276 41644 658340
rect 41708 658338 41714 658340
rect 42333 658338 42399 658341
rect 41708 658336 42399 658338
rect 41708 658280 42338 658336
rect 42394 658280 42399 658336
rect 41708 658278 42399 658280
rect 41708 658276 41714 658278
rect 42333 658275 42399 658278
rect 651557 657114 651623 657117
rect 650164 657112 651623 657114
rect 650164 657056 651562 657112
rect 651618 657056 651623 657112
rect 650164 657054 651623 657056
rect 651557 657051 651623 657054
rect 674414 652156 674420 652220
rect 674484 652218 674490 652220
rect 675477 652218 675543 652221
rect 674484 652216 675543 652218
rect 674484 652160 675482 652216
rect 675538 652160 675543 652216
rect 674484 652158 675543 652160
rect 674484 652156 674490 652158
rect 675477 652155 675543 652158
rect 675753 651538 675819 651541
rect 675886 651538 675892 651540
rect 675753 651536 675892 651538
rect 675753 651480 675758 651536
rect 675814 651480 675892 651536
rect 675753 651478 675892 651480
rect 675753 651475 675819 651478
rect 675886 651476 675892 651478
rect 675956 651476 675962 651540
rect 6022 651353 63922 651382
rect 6022 650209 6150 651353
rect 6854 651349 63922 651353
rect 6854 650245 54235 651349
rect 55339 651329 63922 651349
rect 55339 650245 63339 651329
rect 6854 650225 63339 650245
rect 63883 650225 63922 651329
rect 6854 650209 63922 650225
rect 6022 650182 63922 650209
rect 62113 650042 62179 650045
rect 62113 650040 64492 650042
rect 62113 649984 62118 650040
rect 62174 649984 64492 650040
rect 62113 649982 64492 649984
rect 62113 649979 62179 649982
rect 7236 649757 62944 649782
rect 7236 648613 7348 649757
rect 8052 649731 62944 649757
rect 8052 648627 52641 649731
rect 53745 649721 62944 649731
rect 53745 648627 62371 649721
rect 8052 648617 62371 648627
rect 62915 648617 62944 649721
rect 673310 649164 673316 649228
rect 673380 649226 673386 649228
rect 675385 649226 675451 649229
rect 673380 649224 675451 649226
rect 673380 649168 675390 649224
rect 675446 649168 675451 649224
rect 673380 649166 675451 649168
rect 673380 649164 673386 649166
rect 675385 649163 675451 649166
rect 675753 648682 675819 648685
rect 676254 648682 676260 648684
rect 675753 648680 676260 648682
rect 675753 648624 675758 648680
rect 675814 648624 676260 648680
rect 675753 648622 676260 648624
rect 675753 648619 675819 648622
rect 676254 648620 676260 648622
rect 676324 648620 676330 648684
rect 8052 648613 62944 648617
rect 7236 648582 62944 648613
rect 35574 644741 35634 644912
rect 35574 644736 35683 644741
rect 35801 644738 35867 644741
rect 35574 644680 35622 644736
rect 35678 644680 35683 644736
rect 35574 644678 35683 644680
rect 35617 644675 35683 644678
rect 35758 644736 35867 644738
rect 35758 644680 35806 644736
rect 35862 644680 35867 644736
rect 35758 644675 35867 644680
rect 675753 644738 675819 644741
rect 676622 644738 676628 644740
rect 675753 644736 676628 644738
rect 675753 644680 675758 644736
rect 675814 644680 676628 644736
rect 675753 644678 676628 644680
rect 675753 644675 675819 644678
rect 676622 644676 676628 644678
rect 676692 644676 676698 644740
rect 35758 644504 35818 644675
rect 676990 644602 676996 644604
rect 675710 644542 676996 644602
rect 41462 643922 41522 644096
rect 41462 643862 45570 643922
rect 44265 643786 44331 643789
rect 41462 643784 44331 643786
rect 41462 643728 44270 643784
rect 44326 643728 44331 643784
rect 41462 643726 44331 643728
rect 41462 643688 41522 643726
rect 44265 643723 44331 643726
rect 45510 643514 45570 643862
rect 651557 643786 651623 643789
rect 650164 643784 651623 643786
rect 650164 643728 651562 643784
rect 651618 643728 651623 643784
rect 650164 643726 651623 643728
rect 651557 643723 651623 643726
rect 62757 643514 62823 643517
rect 45510 643512 62823 643514
rect 45510 643456 62762 643512
rect 62818 643456 62823 643512
rect 45510 643454 62823 643456
rect 62757 643451 62823 643454
rect 41462 643242 41522 643280
rect 44357 643242 44423 643245
rect 41462 643240 44423 643242
rect 41462 643184 44362 643240
rect 44418 643184 44423 643240
rect 41462 643182 44423 643184
rect 44357 643179 44423 643182
rect 675710 643109 675770 644542
rect 676990 644540 676996 644542
rect 677060 644540 677066 644604
rect 44173 643106 44239 643109
rect 41462 643104 44239 643106
rect 41462 643048 44178 643104
rect 44234 643048 44239 643104
rect 41462 643046 44239 643048
rect 41462 642872 41522 643046
rect 44173 643043 44239 643046
rect 675661 643104 675770 643109
rect 675661 643048 675666 643104
rect 675722 643048 675770 643104
rect 675661 643046 675770 643048
rect 675661 643043 675727 643046
rect 39982 642228 39988 642292
rect 40052 642228 40058 642292
rect 41462 642290 41522 642464
rect 44173 642290 44239 642293
rect 41462 642288 44239 642290
rect 41462 642232 44178 642288
rect 44234 642232 44239 642288
rect 41462 642230 44239 642232
rect 39990 642056 40050 642228
rect 44173 642227 44239 642230
rect 39990 641476 40050 641648
rect 39982 641412 39988 641476
rect 40052 641412 40058 641476
rect 42793 641474 42859 641477
rect 41462 641472 42859 641474
rect 41462 641416 42798 641472
rect 42854 641416 42859 641472
rect 41462 641414 42859 641416
rect 41462 641240 41522 641414
rect 42793 641411 42859 641414
rect 41462 640794 41522 640832
rect 44265 640794 44331 640797
rect 41462 640792 44331 640794
rect 41462 640736 44270 640792
rect 44326 640736 44331 640792
rect 41462 640734 44331 640736
rect 44265 640731 44331 640734
rect 41454 640596 41460 640660
rect 41524 640596 41530 640660
rect 41462 640424 41522 640596
rect 675477 640388 675543 640389
rect 675477 640384 675524 640388
rect 675588 640386 675594 640388
rect 675477 640328 675482 640384
rect 675477 640324 675524 640328
rect 675588 640326 675634 640386
rect 675588 640324 675594 640326
rect 675477 640323 675543 640324
rect 33734 639845 33794 640016
rect 33734 639840 33843 639845
rect 33734 639784 33782 639840
rect 33838 639784 33843 639840
rect 33734 639782 33843 639784
rect 33777 639779 33843 639782
rect 40726 639437 40786 639608
rect 40677 639432 40786 639437
rect 40677 639376 40682 639432
rect 40738 639376 40786 639432
rect 40677 639374 40786 639376
rect 40677 639371 40743 639374
rect 40910 639029 40970 639200
rect 40861 639024 40970 639029
rect 40861 638968 40866 639024
rect 40922 638968 40970 639024
rect 40861 638966 40970 638968
rect 40861 638963 40927 638966
rect 41462 638618 41522 638792
rect 42793 638618 42859 638621
rect 41462 638616 42859 638618
rect 41462 638560 42798 638616
rect 42854 638560 42859 638616
rect 41462 638558 42859 638560
rect 42793 638555 42859 638558
rect 32446 638213 32506 638384
rect 32397 638208 32506 638213
rect 32397 638152 32402 638208
rect 32458 638152 32506 638208
rect 32397 638150 32506 638152
rect 32397 638147 32463 638150
rect 675518 638148 675524 638212
rect 675588 638210 675594 638212
rect 675661 638210 675727 638213
rect 675588 638208 675727 638210
rect 675588 638152 675666 638208
rect 675722 638152 675727 638208
rect 675588 638150 675727 638152
rect 675588 638148 675594 638150
rect 675661 638147 675727 638150
rect 35206 637805 35266 637976
rect 35157 637800 35266 637805
rect 35157 637744 35162 637800
rect 35218 637744 35266 637800
rect 35157 637742 35266 637744
rect 35157 637739 35223 637742
rect 41094 637397 41154 637568
rect 41045 637392 41154 637397
rect 41045 637336 41050 637392
rect 41106 637336 41154 637392
rect 41045 637334 41154 637336
rect 41045 637331 41111 637334
rect 41462 636986 41522 637160
rect 62113 637122 62179 637125
rect 62113 637120 64492 637122
rect 62113 637064 62118 637120
rect 62174 637064 64492 637120
rect 62113 637062 64492 637064
rect 62113 637059 62179 637062
rect 44449 636986 44515 636989
rect 41462 636984 44515 636986
rect 41462 636928 44454 636984
rect 44510 636928 44515 636984
rect 41462 636926 44515 636928
rect 44449 636923 44515 636926
rect 40910 636580 40970 636752
rect 40902 636516 40908 636580
rect 40972 636516 40978 636580
rect 40542 636172 40602 636344
rect 40534 636108 40540 636172
rect 40604 636108 40610 636172
rect 41462 635762 41522 635936
rect 42885 635762 42951 635765
rect 41462 635760 42951 635762
rect 41462 635704 42890 635760
rect 42946 635704 42951 635760
rect 41462 635702 42951 635704
rect 42885 635699 42951 635702
rect 41462 635354 41522 635528
rect 43069 635354 43135 635357
rect 41462 635352 43135 635354
rect 41462 635296 43074 635352
rect 43130 635296 43135 635352
rect 41462 635294 43135 635296
rect 43069 635291 43135 635294
rect 40726 634948 40786 635120
rect 40718 634884 40724 634948
rect 40788 634884 40794 634948
rect 41462 634538 41522 634712
rect 41462 634478 41890 634538
rect 30422 633896 30482 634304
rect 41830 633722 41890 634478
rect 41462 633662 41890 633722
rect 41462 633450 41522 633662
rect 53097 633450 53163 633453
rect 41462 633448 53163 633450
rect 41462 633392 53102 633448
rect 53158 633392 53163 633448
rect 41462 633390 53163 633392
rect 53097 633387 53163 633390
rect 675702 633388 675708 633452
rect 675772 633450 675778 633452
rect 678237 633450 678303 633453
rect 675772 633448 678303 633450
rect 675772 633392 678242 633448
rect 678298 633392 678303 633448
rect 675772 633390 678303 633392
rect 675772 633388 675778 633390
rect 678237 633387 678303 633390
rect 651557 630594 651623 630597
rect 650164 630592 651623 630594
rect 650164 630536 651562 630592
rect 651618 630536 651623 630592
rect 650164 630534 651623 630536
rect 651557 630531 651623 630534
rect 35157 629914 35223 629917
rect 41822 629914 41828 629916
rect 35157 629912 41828 629914
rect 35157 629856 35162 629912
rect 35218 629856 41828 629912
rect 35157 629854 41828 629856
rect 35157 629851 35223 629854
rect 41822 629852 41828 629854
rect 41892 629852 41898 629916
rect 41045 629234 41111 629237
rect 42006 629234 42012 629236
rect 41045 629232 42012 629234
rect 41045 629176 41050 629232
rect 41106 629176 42012 629232
rect 41045 629174 42012 629176
rect 41045 629171 41111 629174
rect 42006 629172 42012 629174
rect 42076 629172 42082 629236
rect 40677 629098 40743 629101
rect 41638 629098 41644 629100
rect 40677 629096 41644 629098
rect 40677 629040 40682 629096
rect 40738 629040 41644 629096
rect 40677 629038 41644 629040
rect 40677 629035 40743 629038
rect 41638 629036 41644 629038
rect 41708 629036 41714 629100
rect 40861 628962 40927 628965
rect 42190 628962 42196 628964
rect 40861 628960 42196 628962
rect 40861 628904 40866 628960
rect 40922 628904 42196 628960
rect 40861 628902 42196 628904
rect 40861 628899 40927 628902
rect 42190 628900 42196 628902
rect 42260 628900 42266 628964
rect 676121 626106 676187 626109
rect 676262 626106 676322 626348
rect 676121 626104 676322 626106
rect 676121 626048 676126 626104
rect 676182 626048 676322 626104
rect 676121 626046 676322 626048
rect 676121 626043 676187 626046
rect 676262 625701 676322 625940
rect 676213 625696 676322 625701
rect 676213 625640 676218 625696
rect 676274 625640 676322 625696
rect 676213 625638 676322 625640
rect 676213 625635 676279 625638
rect 676262 625293 676322 625532
rect 40902 625228 40908 625292
rect 40972 625290 40978 625292
rect 40972 625230 42442 625290
rect 40972 625228 40978 625230
rect 42382 625154 42442 625230
rect 676213 625288 676322 625293
rect 676213 625232 676218 625288
rect 676274 625232 676322 625288
rect 676213 625230 676322 625232
rect 676213 625227 676279 625230
rect 42517 625154 42583 625157
rect 42382 625152 42583 625154
rect 42382 625096 42522 625152
rect 42578 625096 42583 625152
rect 42382 625094 42583 625096
rect 42517 625091 42583 625094
rect 674741 625154 674807 625157
rect 674741 625152 676292 625154
rect 674741 625096 674746 625152
rect 674802 625096 676292 625152
rect 674741 625094 676292 625096
rect 674741 625091 674807 625094
rect 676262 624477 676322 624716
rect 676213 624472 676322 624477
rect 676213 624416 676218 624472
rect 676274 624416 676322 624472
rect 676213 624414 676322 624416
rect 676213 624411 676279 624414
rect 676029 624338 676095 624341
rect 676029 624336 676292 624338
rect 676029 624280 676034 624336
rect 676090 624280 676292 624336
rect 676029 624278 676292 624280
rect 676029 624275 676095 624278
rect 62113 624066 62179 624069
rect 62113 624064 64492 624066
rect 62113 624008 62118 624064
rect 62174 624008 64492 624064
rect 62113 624006 64492 624008
rect 62113 624003 62179 624006
rect 676029 623930 676095 623933
rect 676029 623928 676292 623930
rect 676029 623872 676034 623928
rect 676090 623872 676292 623928
rect 676029 623870 676292 623872
rect 676029 623867 676095 623870
rect 40718 623732 40724 623796
rect 40788 623794 40794 623796
rect 42517 623794 42583 623797
rect 40788 623792 42583 623794
rect 40788 623736 42522 623792
rect 42578 623736 42583 623792
rect 40788 623734 42583 623736
rect 40788 623732 40794 623734
rect 42517 623731 42583 623734
rect 676121 623250 676187 623253
rect 676262 623250 676322 623492
rect 676121 623248 676322 623250
rect 676121 623192 676126 623248
rect 676182 623192 676322 623248
rect 676121 623190 676322 623192
rect 676121 623187 676187 623190
rect 676262 622845 676322 623084
rect 676213 622840 676322 622845
rect 676213 622784 676218 622840
rect 676274 622784 676322 622840
rect 676213 622782 676322 622784
rect 676213 622779 676279 622782
rect 676029 622706 676095 622709
rect 676029 622704 676292 622706
rect 676029 622648 676034 622704
rect 676090 622648 676292 622704
rect 676029 622646 676292 622648
rect 676029 622643 676095 622646
rect 676029 622298 676095 622301
rect 676029 622296 676292 622298
rect 676029 622240 676034 622296
rect 676090 622240 676292 622296
rect 676029 622238 676292 622240
rect 676029 622235 676095 622238
rect 678237 622026 678303 622029
rect 678237 622024 678346 622026
rect 678237 621968 678242 622024
rect 678298 621968 678346 622024
rect 678237 621963 678346 621968
rect 678286 621860 678346 621963
rect 40534 621420 40540 621484
rect 40604 621482 40610 621484
rect 41781 621482 41847 621485
rect 40604 621480 41847 621482
rect 40604 621424 41786 621480
rect 41842 621424 41847 621480
rect 40604 621422 41847 621424
rect 40604 621420 40610 621422
rect 41781 621419 41847 621422
rect 676029 621482 676095 621485
rect 676029 621480 676292 621482
rect 676029 621424 676034 621480
rect 676090 621424 676292 621480
rect 676029 621422 676292 621424
rect 676029 621419 676095 621422
rect 676213 621210 676279 621213
rect 676213 621208 676322 621210
rect 676213 621152 676218 621208
rect 676274 621152 676322 621208
rect 676213 621147 676322 621152
rect 676262 621044 676322 621147
rect 676070 620740 676076 620804
rect 676140 620802 676146 620804
rect 676140 620742 676322 620802
rect 676140 620740 676146 620742
rect 676262 620636 676322 620742
rect 676262 619989 676322 620228
rect 676213 619984 676322 619989
rect 676213 619928 676218 619984
rect 676274 619928 676322 619984
rect 676213 619926 676322 619928
rect 676213 619923 676279 619926
rect 676029 619850 676095 619853
rect 676029 619848 676292 619850
rect 676029 619792 676034 619848
rect 676090 619792 676292 619848
rect 676029 619790 676292 619792
rect 676029 619787 676095 619790
rect 674598 619380 674604 619444
rect 674668 619442 674674 619444
rect 674668 619382 676292 619442
rect 674668 619380 674674 619382
rect 676213 619170 676279 619173
rect 676213 619168 676322 619170
rect 676213 619112 676218 619168
rect 676274 619112 676322 619168
rect 676213 619107 676322 619112
rect 42006 618972 42012 619036
rect 42076 619034 42082 619036
rect 42241 619034 42307 619037
rect 42076 619032 42307 619034
rect 42076 618976 42246 619032
rect 42302 618976 42307 619032
rect 676262 619004 676322 619107
rect 42076 618974 42307 618976
rect 42076 618972 42082 618974
rect 42241 618971 42307 618974
rect 676438 618700 676444 618764
rect 676508 618700 676514 618764
rect 676446 618596 676506 618700
rect 676121 617946 676187 617949
rect 676262 617946 676322 618188
rect 676121 617944 676322 617946
rect 676121 617888 676126 617944
rect 676182 617888 676322 617944
rect 676121 617886 676322 617888
rect 676121 617883 676187 617886
rect 676029 617810 676095 617813
rect 676029 617808 676292 617810
rect 676029 617752 676034 617808
rect 676090 617752 676292 617808
rect 676029 617750 676292 617752
rect 676029 617747 676095 617750
rect 652385 617266 652451 617269
rect 650164 617264 652451 617266
rect 650164 617208 652390 617264
rect 652446 617208 652451 617264
rect 650164 617206 652451 617208
rect 652385 617203 652451 617206
rect 676262 617133 676322 617372
rect 676213 617128 676322 617133
rect 676213 617072 676218 617128
rect 676274 617072 676322 617128
rect 676213 617070 676322 617072
rect 676213 617067 676279 617070
rect 676029 616994 676095 616997
rect 676029 616992 676292 616994
rect 676029 616936 676034 616992
rect 676090 616936 676292 616992
rect 676029 616934 676292 616936
rect 676029 616931 676095 616934
rect 41822 616796 41828 616860
rect 41892 616858 41898 616860
rect 42517 616858 42583 616861
rect 41892 616856 42583 616858
rect 41892 616800 42522 616856
rect 42578 616800 42583 616856
rect 41892 616798 42583 616800
rect 41892 616796 41898 616798
rect 42517 616795 42583 616798
rect 676262 616317 676322 616556
rect 676213 616312 676322 616317
rect 676213 616256 676218 616312
rect 676274 616256 676322 616312
rect 676213 616254 676322 616256
rect 676213 616251 676279 616254
rect 42241 616044 42307 616045
rect 42190 615980 42196 616044
rect 42260 616042 42307 616044
rect 42260 616040 42352 616042
rect 42302 615984 42352 616040
rect 42260 615982 42352 615984
rect 42260 615980 42307 615982
rect 42241 615979 42307 615980
rect 683070 615909 683130 616148
rect 683070 615904 683179 615909
rect 683070 615848 683118 615904
rect 683174 615848 683179 615904
rect 683070 615846 683179 615848
rect 683113 615843 683179 615846
rect 683070 615332 683130 615740
rect 683113 615090 683179 615093
rect 683070 615088 683179 615090
rect 683070 615032 683118 615088
rect 683174 615032 683179 615088
rect 683070 615027 683179 615032
rect 683070 614924 683130 615027
rect 41454 614076 41460 614140
rect 41524 614138 41530 614140
rect 41873 614138 41939 614141
rect 41524 614136 41939 614138
rect 41524 614080 41878 614136
rect 41934 614080 41939 614136
rect 41524 614078 41939 614080
rect 41524 614076 41530 614078
rect 41873 614075 41939 614078
rect 41638 612716 41644 612780
rect 41708 612778 41714 612780
rect 41781 612778 41847 612781
rect 41708 612776 41847 612778
rect 41708 612720 41786 612776
rect 41842 612720 41847 612776
rect 41708 612718 41847 612720
rect 41708 612716 41714 612718
rect 41781 612715 41847 612718
rect 62113 611010 62179 611013
rect 62113 611008 64492 611010
rect 62113 610952 62118 611008
rect 62174 610952 64492 611008
rect 62113 610950 64492 610952
rect 62113 610947 62179 610950
rect 6022 608153 63922 608182
rect 6022 607009 6150 608153
rect 6854 608149 63922 608153
rect 6854 607045 54235 608149
rect 55339 608129 63922 608149
rect 55339 607045 63339 608129
rect 6854 607025 63339 607045
rect 63883 607025 63922 608129
rect 675477 607884 675543 607885
rect 675477 607880 675524 607884
rect 675588 607882 675594 607884
rect 675477 607824 675482 607880
rect 675477 607820 675524 607824
rect 675588 607822 675634 607882
rect 675588 607820 675594 607822
rect 675477 607819 675543 607820
rect 6854 607009 63922 607025
rect 6022 606982 63922 607009
rect 7236 606557 62944 606582
rect 7236 605413 7348 606557
rect 8052 606531 62944 606557
rect 8052 605427 52641 606531
rect 53745 606521 62944 606531
rect 675385 606524 675451 606525
rect 675334 606522 675340 606524
rect 53745 605427 62371 606521
rect 8052 605417 62371 605427
rect 62915 605417 62944 606521
rect 675294 606462 675340 606522
rect 675404 606520 675451 606524
rect 675446 606464 675451 606520
rect 675334 606460 675340 606462
rect 675404 606460 675451 606464
rect 675385 606459 675451 606460
rect 675334 605780 675340 605844
rect 675404 605842 675410 605844
rect 675702 605842 675708 605844
rect 675404 605782 675708 605842
rect 675404 605780 675410 605782
rect 675702 605780 675708 605782
rect 675772 605780 675778 605844
rect 8052 605413 62944 605417
rect 7236 605382 62944 605413
rect 651557 603938 651623 603941
rect 650164 603936 651623 603938
rect 650164 603880 651562 603936
rect 651618 603880 651623 603936
rect 650164 603878 651623 603880
rect 651557 603875 651623 603878
rect 35801 601898 35867 601901
rect 35758 601896 35867 601898
rect 35758 601840 35806 601896
rect 35862 601840 35867 601896
rect 35758 601835 35867 601840
rect 35758 601732 35818 601835
rect 35801 601490 35867 601493
rect 35758 601488 35867 601490
rect 35758 601432 35806 601488
rect 35862 601432 35867 601488
rect 35758 601427 35867 601432
rect 35758 601324 35818 601427
rect 35801 601082 35867 601085
rect 35758 601080 35867 601082
rect 35758 601024 35806 601080
rect 35862 601024 35867 601080
rect 35758 601019 35867 601024
rect 35758 600916 35818 601019
rect 675201 600946 675267 600949
rect 675702 600946 675708 600948
rect 675201 600944 675708 600946
rect 675201 600888 675206 600944
rect 675262 600888 675708 600944
rect 675201 600886 675708 600888
rect 675201 600883 675267 600886
rect 675702 600884 675708 600886
rect 675772 600884 675778 600948
rect 35709 600674 35775 600677
rect 35709 600672 35818 600674
rect 35709 600616 35714 600672
rect 35770 600616 35818 600672
rect 35709 600611 35818 600616
rect 35758 600508 35818 600611
rect 675569 600268 675635 600269
rect 675518 600266 675524 600268
rect 675478 600206 675524 600266
rect 675588 600264 675635 600268
rect 675630 600208 675635 600264
rect 675518 600204 675524 600206
rect 675588 600204 675635 600208
rect 675569 600203 675635 600204
rect 41462 599858 41522 600100
rect 44081 599858 44147 599861
rect 41462 599856 44147 599858
rect 41462 599800 44086 599856
rect 44142 599800 44147 599856
rect 41462 599798 44147 599800
rect 44081 599795 44147 599798
rect 44173 599722 44239 599725
rect 41492 599720 44239 599722
rect 41492 599664 44178 599720
rect 44234 599664 44239 599720
rect 41492 599662 44239 599664
rect 44173 599659 44239 599662
rect 44541 599314 44607 599317
rect 41492 599312 44607 599314
rect 41492 599256 44546 599312
rect 44602 599256 44607 599312
rect 41492 599254 44607 599256
rect 44541 599251 44607 599254
rect 39982 598980 39988 599044
rect 40052 598980 40058 599044
rect 675753 599042 675819 599045
rect 676438 599042 676444 599044
rect 675753 599040 676444 599042
rect 675753 598984 675758 599040
rect 675814 598984 676444 599040
rect 675753 598982 676444 598984
rect 39990 598876 40050 598980
rect 675753 598979 675819 598982
rect 676438 598980 676444 598982
rect 676508 598980 676514 599044
rect 39990 598228 40050 598468
rect 39982 598164 39988 598228
rect 40052 598164 40058 598228
rect 44265 598090 44331 598093
rect 41492 598088 44331 598090
rect 41492 598032 44270 598088
rect 44326 598032 44331 598088
rect 41492 598030 44331 598032
rect 44265 598027 44331 598030
rect 62113 597954 62179 597957
rect 62113 597952 64492 597954
rect 62113 597896 62118 597952
rect 62174 597896 64492 597952
rect 62113 597894 64492 597896
rect 62113 597891 62179 597894
rect 675753 597818 675819 597821
rect 676806 597818 676812 597820
rect 675753 597816 676812 597818
rect 675753 597760 675758 597816
rect 675814 597760 676812 597816
rect 675753 597758 676812 597760
rect 675753 597755 675819 597758
rect 676806 597756 676812 597758
rect 676876 597756 676882 597820
rect 42793 597682 42859 597685
rect 41492 597680 42859 597682
rect 41492 597624 42798 597680
rect 42854 597624 42859 597680
rect 41492 597622 42859 597624
rect 42793 597619 42859 597622
rect 39254 597005 39314 597244
rect 39254 597000 39363 597005
rect 39254 596944 39302 597000
rect 39358 596944 39363 597000
rect 39254 596942 39363 596944
rect 39297 596939 39363 596942
rect 40726 596597 40786 596836
rect 40677 596592 40786 596597
rect 40677 596536 40682 596592
rect 40738 596536 40786 596592
rect 40677 596534 40786 596536
rect 40677 596531 40743 596534
rect 41454 596532 41460 596596
rect 41524 596532 41530 596596
rect 41462 596428 41522 596532
rect 40726 595781 40786 596020
rect 40726 595776 40835 595781
rect 40726 595720 40774 595776
rect 40830 595720 40835 595776
rect 40726 595718 40835 595720
rect 40769 595715 40835 595718
rect 44357 595642 44423 595645
rect 41492 595640 44423 595642
rect 41492 595584 44362 595640
rect 44418 595584 44423 595640
rect 41492 595582 44423 595584
rect 44357 595579 44423 595582
rect 33734 594965 33794 595204
rect 33734 594960 33843 594965
rect 41638 594962 41644 594964
rect 33734 594904 33782 594960
rect 33838 594904 33843 594960
rect 33734 594902 33843 594904
rect 33777 594899 33843 594902
rect 41462 594902 41644 594962
rect 41462 594796 41522 594902
rect 41638 594900 41644 594902
rect 41708 594900 41714 594964
rect 42885 594418 42951 594421
rect 41492 594416 42951 594418
rect 41492 594360 42890 594416
rect 42946 594360 42951 594416
rect 41492 594358 42951 594360
rect 42885 594355 42951 594358
rect 42057 594010 42123 594013
rect 41492 594008 42123 594010
rect 41492 593952 42062 594008
rect 42118 593952 42123 594008
rect 41492 593950 42123 593952
rect 42057 593947 42123 593950
rect 32446 593333 32506 593572
rect 32397 593328 32506 593333
rect 32397 593272 32402 593328
rect 32458 593272 32506 593328
rect 32397 593270 32506 593272
rect 32397 593267 32463 593270
rect 44449 593194 44515 593197
rect 675477 593196 675543 593197
rect 675661 593196 675727 593197
rect 675477 593194 675524 593196
rect 41492 593192 44515 593194
rect 41492 593136 44454 593192
rect 44510 593136 44515 593192
rect 41492 593134 44515 593136
rect 675432 593192 675524 593194
rect 675432 593136 675482 593192
rect 675432 593134 675524 593136
rect 44449 593131 44515 593134
rect 675477 593132 675524 593134
rect 675588 593132 675594 593196
rect 675661 593192 675708 593196
rect 675772 593194 675778 593196
rect 675661 593136 675666 593192
rect 675661 593132 675708 593136
rect 675772 593134 675818 593194
rect 675772 593132 675778 593134
rect 675477 593131 675543 593132
rect 675661 593131 675727 593132
rect 42977 592786 43043 592789
rect 41492 592784 43043 592786
rect 41492 592728 42982 592784
rect 43038 592728 43043 592784
rect 41492 592726 43043 592728
rect 42977 592723 43043 592726
rect 40542 592108 40602 592348
rect 40534 592044 40540 592108
rect 40604 592044 40610 592108
rect 40726 591700 40786 591940
rect 40718 591636 40724 591700
rect 40788 591636 40794 591700
rect 41462 591293 41522 591532
rect 41462 591288 41571 591293
rect 41462 591232 41510 591288
rect 41566 591232 41571 591288
rect 41462 591230 41571 591232
rect 41505 591227 41571 591230
rect 30422 590716 30482 591124
rect 651557 590746 651623 590749
rect 650164 590744 651623 590746
rect 650164 590688 651562 590744
rect 651618 590688 651623 590744
rect 650164 590686 651623 590688
rect 651557 590683 651623 590686
rect 41462 590069 41522 590308
rect 41462 590064 41571 590069
rect 41462 590008 41510 590064
rect 41566 590008 41571 590064
rect 41462 590006 41571 590008
rect 41505 590003 41571 590006
rect 676070 589188 676076 589252
rect 676140 589250 676146 589252
rect 678237 589250 678303 589253
rect 676140 589248 678303 589250
rect 676140 589192 678242 589248
rect 678298 589192 678303 589248
rect 676140 589190 678303 589192
rect 676140 589188 676146 589190
rect 678237 589187 678303 589190
rect 39297 585170 39363 585173
rect 42374 585170 42380 585172
rect 39297 585168 42380 585170
rect 39297 585112 39302 585168
rect 39358 585112 42380 585168
rect 39297 585110 42380 585112
rect 39297 585107 39363 585110
rect 42374 585108 42380 585110
rect 42444 585108 42450 585172
rect 62113 584898 62179 584901
rect 62113 584896 64492 584898
rect 62113 584840 62118 584896
rect 62174 584840 64492 584896
rect 62113 584838 64492 584840
rect 62113 584835 62179 584838
rect 41781 584220 41847 584221
rect 41965 584220 42031 584221
rect 41781 584218 41828 584220
rect 41736 584216 41828 584218
rect 41736 584160 41786 584216
rect 41736 584158 41828 584160
rect 41781 584156 41828 584158
rect 41892 584156 41898 584220
rect 41965 584216 42012 584220
rect 42076 584218 42082 584220
rect 41965 584160 41970 584216
rect 41965 584156 42012 584160
rect 42076 584158 42122 584218
rect 42076 584156 42082 584158
rect 41781 584155 41847 584156
rect 41965 584155 42031 584156
rect 42425 583674 42491 583677
rect 42558 583674 42564 583676
rect 42425 583672 42564 583674
rect 42425 583616 42430 583672
rect 42486 583616 42564 583672
rect 42425 583614 42564 583616
rect 42425 583611 42491 583614
rect 42558 583612 42564 583614
rect 42628 583612 42634 583676
rect 41965 582180 42031 582181
rect 41965 582176 42012 582180
rect 42076 582178 42082 582180
rect 41965 582120 41970 582176
rect 41965 582116 42012 582120
rect 42076 582118 42122 582178
rect 42076 582116 42082 582118
rect 41965 582115 42031 582116
rect 676029 581090 676095 581093
rect 676029 581088 676292 581090
rect 676029 581032 676034 581088
rect 676090 581032 676292 581088
rect 676029 581030 676292 581032
rect 676029 581027 676095 581030
rect 676121 580546 676187 580549
rect 676262 580546 676322 580652
rect 676121 580544 676322 580546
rect 676121 580488 676126 580544
rect 676182 580488 676322 580544
rect 676121 580486 676322 580488
rect 676121 580483 676187 580486
rect 41781 580276 41847 580277
rect 41781 580272 41828 580276
rect 41892 580274 41898 580276
rect 676029 580274 676095 580277
rect 41781 580216 41786 580272
rect 41781 580212 41828 580216
rect 41892 580214 41938 580274
rect 676029 580272 676292 580274
rect 676029 580216 676034 580272
rect 676090 580216 676292 580272
rect 676029 580214 676292 580216
rect 41892 580212 41898 580214
rect 41781 580211 41847 580212
rect 676029 580211 676095 580214
rect 676213 580138 676279 580141
rect 676213 580136 676322 580138
rect 676213 580080 676218 580136
rect 676274 580080 676322 580136
rect 676213 580075 676322 580080
rect 676262 579836 676322 580075
rect 676262 579325 676322 579428
rect 676213 579320 676322 579325
rect 676213 579264 676218 579320
rect 676274 579264 676322 579320
rect 676213 579262 676322 579264
rect 676213 579259 676279 579262
rect 40718 578988 40724 579052
rect 40788 579050 40794 579052
rect 41781 579050 41847 579053
rect 40788 579048 41847 579050
rect 40788 578992 41786 579048
rect 41842 578992 41847 579048
rect 40788 578990 41847 578992
rect 40788 578988 40794 578990
rect 41781 578987 41847 578990
rect 676262 578917 676322 579020
rect 676213 578912 676322 578917
rect 676213 578856 676218 578912
rect 676274 578856 676322 578912
rect 676213 578854 676322 578856
rect 676213 578851 676279 578854
rect 676029 578642 676095 578645
rect 676029 578640 676292 578642
rect 676029 578584 676034 578640
rect 676090 578584 676292 578640
rect 676029 578582 676292 578584
rect 676029 578579 676095 578582
rect 676262 578101 676322 578204
rect 676213 578096 676322 578101
rect 676213 578040 676218 578096
rect 676274 578040 676322 578096
rect 676213 578038 676322 578040
rect 676213 578035 676279 578038
rect 676121 577690 676187 577693
rect 676262 577690 676322 577796
rect 676121 577688 676322 577690
rect 676121 577632 676126 577688
rect 676182 577632 676322 577688
rect 676121 577630 676322 577632
rect 676121 577627 676187 577630
rect 40534 577492 40540 577556
rect 40604 577554 40610 577556
rect 41781 577554 41847 577557
rect 40604 577552 41847 577554
rect 40604 577496 41786 577552
rect 41842 577496 41847 577552
rect 40604 577494 41847 577496
rect 40604 577492 40610 577494
rect 41781 577491 41847 577494
rect 651557 577418 651623 577421
rect 650164 577416 651623 577418
rect 650164 577360 651562 577416
rect 651618 577360 651623 577416
rect 650164 577358 651623 577360
rect 651557 577355 651623 577358
rect 676029 577418 676095 577421
rect 676029 577416 676292 577418
rect 676029 577360 676034 577416
rect 676090 577360 676292 577416
rect 676029 577358 676292 577360
rect 676029 577355 676095 577358
rect 676029 577010 676095 577013
rect 676029 577008 676292 577010
rect 676029 576952 676034 577008
rect 676090 576952 676292 577008
rect 676029 576950 676292 576952
rect 676029 576947 676095 576950
rect 42190 576812 42196 576876
rect 42260 576874 42266 576876
rect 42701 576874 42767 576877
rect 42260 576872 42767 576874
rect 42260 576816 42706 576872
rect 42762 576816 42767 576872
rect 42260 576814 42767 576816
rect 42260 576812 42266 576814
rect 42701 576811 42767 576814
rect 678237 576874 678303 576877
rect 678237 576872 678346 576874
rect 678237 576816 678242 576872
rect 678298 576816 678346 576872
rect 678237 576811 678346 576816
rect 678286 576572 678346 576811
rect 675661 576194 675727 576197
rect 675661 576192 676292 576194
rect 675661 576136 675666 576192
rect 675722 576136 676292 576192
rect 675661 576134 676292 576136
rect 675661 576131 675727 576134
rect 42190 575860 42196 575924
rect 42260 575922 42266 575924
rect 42333 575922 42399 575925
rect 42260 575920 42399 575922
rect 42260 575864 42338 575920
rect 42394 575864 42399 575920
rect 42260 575862 42399 575864
rect 42260 575860 42266 575862
rect 42333 575859 42399 575862
rect 676262 575653 676322 575756
rect 676213 575648 676322 575653
rect 676213 575592 676218 575648
rect 676274 575592 676322 575648
rect 676213 575590 676322 575592
rect 676213 575587 676279 575590
rect 676029 575378 676095 575381
rect 676029 575376 676292 575378
rect 676029 575320 676034 575376
rect 676090 575320 676292 575376
rect 676029 575318 676292 575320
rect 676029 575315 676095 575318
rect 676262 574837 676322 574940
rect 676213 574832 676322 574837
rect 676213 574776 676218 574832
rect 676274 574776 676322 574832
rect 676213 574774 676322 574776
rect 676213 574771 676279 574774
rect 676029 574562 676095 574565
rect 676029 574560 676292 574562
rect 676029 574504 676034 574560
rect 676090 574504 676292 574560
rect 676029 574502 676292 574504
rect 676029 574499 676095 574502
rect 674414 574092 674420 574156
rect 674484 574154 674490 574156
rect 674484 574094 676292 574154
rect 674484 574092 674490 574094
rect 41822 573684 41828 573748
rect 41892 573746 41898 573748
rect 42333 573746 42399 573749
rect 41892 573744 42399 573746
rect 41892 573688 42338 573744
rect 42394 573688 42399 573744
rect 41892 573686 42399 573688
rect 41892 573684 41898 573686
rect 42333 573683 42399 573686
rect 676262 573610 676322 573716
rect 674790 573550 676322 573610
rect 41965 572796 42031 572797
rect 41965 572792 42012 572796
rect 42076 572794 42082 572796
rect 41965 572736 41970 572792
rect 41965 572732 42012 572736
rect 42076 572734 42122 572794
rect 42076 572732 42082 572734
rect 673310 572732 673316 572796
rect 673380 572794 673386 572796
rect 674790 572794 674850 573550
rect 676262 573204 676322 573308
rect 676254 573140 676260 573204
rect 676324 573140 676330 573204
rect 676990 573140 676996 573204
rect 677060 573140 677066 573204
rect 676998 572900 677058 573140
rect 673380 572734 674850 572794
rect 673380 572732 673386 572734
rect 676622 572732 676628 572796
rect 676692 572732 676698 572796
rect 41965 572731 42031 572732
rect 676630 572492 676690 572732
rect 676262 571981 676322 572084
rect 676213 571976 676322 571981
rect 676213 571920 676218 571976
rect 676274 571920 676322 571976
rect 676213 571918 676322 571920
rect 676213 571915 676279 571918
rect 62113 571842 62179 571845
rect 62113 571840 64492 571842
rect 62113 571784 62118 571840
rect 62174 571784 64492 571840
rect 62113 571782 64492 571784
rect 62113 571779 62179 571782
rect 676029 571706 676095 571709
rect 676029 571704 676292 571706
rect 676029 571648 676034 571704
rect 676090 571648 676292 571704
rect 676029 571646 676292 571648
rect 676029 571643 676095 571646
rect 41454 571508 41460 571572
rect 41524 571570 41530 571572
rect 42701 571570 42767 571573
rect 41524 571568 42767 571570
rect 41524 571512 42706 571568
rect 42762 571512 42767 571568
rect 41524 571510 42767 571512
rect 41524 571508 41530 571510
rect 42701 571507 42767 571510
rect 676262 571165 676322 571268
rect 676213 571160 676322 571165
rect 676213 571104 676218 571160
rect 676274 571104 676322 571160
rect 676213 571102 676322 571104
rect 676213 571099 676279 571102
rect 683070 570757 683130 570860
rect 683070 570752 683179 570757
rect 683070 570696 683118 570752
rect 683174 570696 683179 570752
rect 683070 570694 683179 570696
rect 683113 570691 683179 570694
rect 41638 570420 41644 570484
rect 41708 570482 41714 570484
rect 42149 570482 42215 570485
rect 41708 570480 42215 570482
rect 41708 570424 42154 570480
rect 42210 570424 42215 570480
rect 41708 570422 42215 570424
rect 41708 570420 41714 570422
rect 42149 570419 42215 570422
rect 685830 570044 685890 570452
rect 683113 569938 683179 569941
rect 683070 569936 683179 569938
rect 683070 569880 683118 569936
rect 683174 569880 683179 569936
rect 683070 569875 683179 569880
rect 683070 569636 683130 569875
rect 675477 568578 675543 568581
rect 676990 568578 676996 568580
rect 675477 568576 676996 568578
rect 675477 568520 675482 568576
rect 675538 568520 676996 568576
rect 675477 568518 676996 568520
rect 675477 568515 675543 568518
rect 676990 568516 676996 568518
rect 677060 568516 677066 568580
rect 6022 564953 63922 564982
rect 6022 563809 6150 564953
rect 6854 564949 63922 564953
rect 6854 563845 54235 564949
rect 55339 564929 63922 564949
rect 55339 563845 63339 564929
rect 6854 563825 63339 563845
rect 63883 563825 63922 564929
rect 652109 564090 652175 564093
rect 650164 564088 652175 564090
rect 650164 564032 652114 564088
rect 652170 564032 652175 564088
rect 650164 564030 652175 564032
rect 652109 564027 652175 564030
rect 6854 563809 63922 563825
rect 6022 563782 63922 563809
rect 7236 563357 62944 563382
rect 7236 562213 7348 563357
rect 8052 563331 62944 563357
rect 8052 562227 52641 563331
rect 53745 563321 62944 563331
rect 53745 562227 62371 563321
rect 8052 562217 62371 562227
rect 62915 562217 62944 563321
rect 675753 562730 675819 562733
rect 675886 562730 675892 562732
rect 675753 562728 675892 562730
rect 675753 562672 675758 562728
rect 675814 562672 675892 562728
rect 675753 562670 675892 562672
rect 675753 562667 675819 562670
rect 675886 562668 675892 562670
rect 675956 562668 675962 562732
rect 8052 562213 62944 562217
rect 7236 562182 62944 562213
rect 675753 561234 675819 561237
rect 676070 561234 676076 561236
rect 675753 561232 676076 561234
rect 675753 561176 675758 561232
rect 675814 561176 676076 561232
rect 675753 561174 676076 561176
rect 675753 561171 675819 561174
rect 676070 561172 676076 561174
rect 676140 561172 676146 561236
rect 675334 559540 675340 559604
rect 675404 559602 675410 559604
rect 675477 559602 675543 559605
rect 675404 559600 675543 559602
rect 675404 559544 675482 559600
rect 675538 559544 675543 559600
rect 675404 559542 675543 559544
rect 675404 559540 675410 559542
rect 675477 559539 675543 559542
rect 62113 558786 62179 558789
rect 62113 558784 64492 558786
rect 62113 558728 62118 558784
rect 62174 558728 64492 558784
rect 62113 558726 64492 558728
rect 62113 558723 62179 558726
rect 35758 558381 35818 558484
rect 35617 558378 35683 558381
rect 35574 558376 35683 558378
rect 35574 558320 35622 558376
rect 35678 558320 35683 558376
rect 35574 558315 35683 558320
rect 35758 558376 35867 558381
rect 35758 558320 35806 558376
rect 35862 558320 35867 558376
rect 35758 558318 35867 558320
rect 35801 558315 35867 558318
rect 675753 558378 675819 558381
rect 676254 558378 676260 558380
rect 675753 558376 676260 558378
rect 675753 558320 675758 558376
rect 675814 558320 676260 558376
rect 675753 558318 676260 558320
rect 675753 558315 675819 558318
rect 676254 558316 676260 558318
rect 676324 558316 676330 558380
rect 35574 558076 35634 558315
rect 35709 557970 35775 557973
rect 35709 557968 35818 557970
rect 35709 557912 35714 557968
rect 35770 557912 35818 557968
rect 35709 557907 35818 557912
rect 35758 557668 35818 557907
rect 44173 557290 44239 557293
rect 41492 557288 44239 557290
rect 41492 557232 44178 557288
rect 44234 557232 44239 557288
rect 41492 557230 44239 557232
rect 44173 557227 44239 557230
rect 42977 556882 43043 556885
rect 41492 556880 43043 556882
rect 41492 556824 42982 556880
rect 43038 556824 43043 556880
rect 41492 556822 43043 556824
rect 42977 556819 43043 556822
rect 44541 556474 44607 556477
rect 41492 556472 44607 556474
rect 41492 556416 44546 556472
rect 44602 556416 44607 556472
rect 41492 556414 44607 556416
rect 44541 556411 44607 556414
rect 42885 556066 42951 556069
rect 41492 556064 42951 556066
rect 41492 556008 42890 556064
rect 42946 556008 42951 556064
rect 41492 556006 42951 556008
rect 42885 556003 42951 556006
rect 39982 555868 39988 555932
rect 40052 555868 40058 555932
rect 39990 555628 40050 555868
rect 44173 555250 44239 555253
rect 41492 555248 44239 555250
rect 41492 555192 44178 555248
rect 44234 555192 44239 555248
rect 41492 555190 44239 555192
rect 44173 555187 44239 555190
rect 42793 554842 42859 554845
rect 41492 554840 42859 554842
rect 41492 554784 42798 554840
rect 42854 554784 42859 554840
rect 41492 554782 42859 554784
rect 42793 554779 42859 554782
rect 44633 554434 44699 554437
rect 41492 554432 44699 554434
rect 41492 554376 44638 554432
rect 44694 554376 44699 554432
rect 41492 554374 44699 554376
rect 44633 554371 44699 554374
rect 40910 553893 40970 553996
rect 40861 553888 40970 553893
rect 40861 553832 40866 553888
rect 40922 553832 40970 553888
rect 40861 553830 40970 553832
rect 40861 553827 40927 553830
rect 40726 553485 40786 553588
rect 40677 553480 40786 553485
rect 40677 553424 40682 553480
rect 40738 553424 40786 553480
rect 40677 553422 40786 553424
rect 40677 553419 40743 553422
rect 40910 553077 40970 553180
rect 40910 553072 41019 553077
rect 40910 553016 40958 553072
rect 41014 553016 41019 553072
rect 40910 553014 41019 553016
rect 40953 553011 41019 553014
rect 32446 552669 32506 552772
rect 32397 552664 32506 552669
rect 32397 552608 32402 552664
rect 32458 552608 32506 552664
rect 32397 552606 32506 552608
rect 32397 552603 32463 552606
rect 40726 552261 40786 552364
rect 40726 552256 40835 552261
rect 40726 552200 40774 552256
rect 40830 552200 40835 552256
rect 40726 552198 40835 552200
rect 40769 552195 40835 552198
rect 675753 551986 675819 551989
rect 676622 551986 676628 551988
rect 675753 551984 676628 551986
rect 30974 551853 31034 551956
rect 675753 551928 675758 551984
rect 675814 551928 676628 551984
rect 675753 551926 676628 551928
rect 675753 551923 675819 551926
rect 676622 551924 676628 551926
rect 676692 551924 676698 551988
rect 30974 551848 31083 551853
rect 30974 551792 31022 551848
rect 31078 551792 31083 551848
rect 30974 551790 31083 551792
rect 31017 551787 31083 551790
rect 44357 551578 44423 551581
rect 41492 551576 44423 551578
rect 41492 551520 44362 551576
rect 44418 551520 44423 551576
rect 41492 551518 44423 551520
rect 44357 551515 44423 551518
rect 42977 551170 43043 551173
rect 41492 551168 43043 551170
rect 41492 551112 42982 551168
rect 43038 551112 43043 551168
rect 41492 551110 43043 551112
rect 42977 551107 43043 551110
rect 651557 550898 651623 550901
rect 650164 550896 651623 550898
rect 650164 550840 651562 550896
rect 651618 550840 651623 550896
rect 650164 550838 651623 550840
rect 651557 550835 651623 550838
rect 40542 550628 40602 550732
rect 40534 550564 40540 550628
rect 40604 550564 40610 550628
rect 44541 550354 44607 550357
rect 41492 550352 44607 550354
rect 41492 550296 44546 550352
rect 44602 550296 44607 550352
rect 41492 550294 44607 550296
rect 44541 550291 44607 550294
rect 43069 549946 43135 549949
rect 41492 549944 43135 549946
rect 41492 549888 43074 549944
rect 43130 549888 43135 549944
rect 41492 549886 43135 549888
rect 43069 549883 43135 549886
rect 40726 549404 40786 549508
rect 40718 549340 40724 549404
rect 40788 549340 40794 549404
rect 40910 548996 40970 549100
rect 40902 548932 40908 548996
rect 40972 548932 40978 548996
rect 44449 548722 44515 548725
rect 41492 548720 44515 548722
rect 41492 548664 44454 548720
rect 44510 548664 44515 548720
rect 41492 548662 44515 548664
rect 44449 548659 44515 548662
rect 31710 548181 31770 548284
rect 31661 548176 31770 548181
rect 31661 548120 31666 548176
rect 31722 548120 31770 548176
rect 31661 548118 31770 548120
rect 31661 548115 31727 548118
rect 27662 547468 27722 547890
rect 35758 546957 35818 547060
rect 35758 546952 35867 546957
rect 35758 546896 35806 546952
rect 35862 546896 35867 546952
rect 35758 546894 35867 546896
rect 35801 546891 35867 546894
rect 675518 546484 675524 546548
rect 675588 546546 675594 546548
rect 680997 546546 681063 546549
rect 675588 546544 681063 546546
rect 675588 546488 681002 546544
rect 681058 546488 681063 546544
rect 675588 546486 681063 546488
rect 675588 546484 675594 546486
rect 680997 546483 681063 546486
rect 62757 545866 62823 545869
rect 62757 545864 64492 545866
rect 62757 545808 62762 545864
rect 62818 545808 64492 545864
rect 62757 545806 64492 545808
rect 62757 545803 62823 545806
rect 40861 545186 40927 545189
rect 41454 545186 41460 545188
rect 40861 545184 41460 545186
rect 40861 545128 40866 545184
rect 40922 545128 41460 545184
rect 40861 545126 41460 545128
rect 40861 545123 40927 545126
rect 41454 545124 41460 545126
rect 41524 545124 41530 545188
rect 675702 543764 675708 543828
rect 675772 543826 675778 543828
rect 678237 543826 678303 543829
rect 675772 543824 678303 543826
rect 675772 543768 678242 543824
rect 678298 543768 678303 543824
rect 675772 543766 678303 543768
rect 675772 543764 675778 543766
rect 678237 543763 678303 543766
rect 40953 543010 41019 543013
rect 41638 543010 41644 543012
rect 40953 543008 41644 543010
rect 40953 542952 40958 543008
rect 41014 542952 41644 543008
rect 40953 542950 41644 542952
rect 40953 542947 41019 542950
rect 41638 542948 41644 542950
rect 41708 542948 41714 543012
rect 32397 542874 32463 542877
rect 41822 542874 41828 542876
rect 32397 542872 41828 542874
rect 32397 542816 32402 542872
rect 32458 542816 41828 542872
rect 32397 542814 41828 542816
rect 32397 542811 32463 542814
rect 41822 542812 41828 542814
rect 41892 542812 41898 542876
rect 40769 542330 40835 542333
rect 42006 542330 42012 542332
rect 40769 542328 42012 542330
rect 40769 542272 40774 542328
rect 40830 542272 42012 542328
rect 40769 542270 42012 542272
rect 40769 542267 40835 542270
rect 42006 542268 42012 542270
rect 42076 542268 42082 542332
rect 651557 537570 651623 537573
rect 650164 537568 651623 537570
rect 650164 537512 651562 537568
rect 651618 537512 651623 537568
rect 650164 537510 651623 537512
rect 651557 537507 651623 537510
rect 676262 535941 676322 536112
rect 42006 535876 42012 535940
rect 42076 535938 42082 535940
rect 42609 535938 42675 535941
rect 42076 535936 42675 535938
rect 42076 535880 42614 535936
rect 42670 535880 42675 535936
rect 42076 535878 42675 535880
rect 42076 535876 42082 535878
rect 42609 535875 42675 535878
rect 676213 535936 676322 535941
rect 676213 535880 676218 535936
rect 676274 535880 676322 535936
rect 676213 535878 676322 535880
rect 676213 535875 676279 535878
rect 676029 535734 676095 535737
rect 676029 535732 676292 535734
rect 676029 535676 676034 535732
rect 676090 535676 676292 535732
rect 676029 535674 676292 535676
rect 676029 535671 676095 535674
rect 676262 535125 676322 535296
rect 676213 535120 676322 535125
rect 676213 535064 676218 535120
rect 676274 535064 676322 535120
rect 676213 535062 676322 535064
rect 676213 535059 676279 535062
rect 676029 534918 676095 534921
rect 676029 534916 676292 534918
rect 676029 534860 676034 534916
rect 676090 534860 676292 534916
rect 676029 534858 676292 534860
rect 676029 534855 676095 534858
rect 40902 534516 40908 534580
rect 40972 534578 40978 534580
rect 41781 534578 41847 534581
rect 40972 534576 41847 534578
rect 40972 534520 41786 534576
rect 41842 534520 41847 534576
rect 40972 534518 41847 534520
rect 40972 534516 40978 534518
rect 41781 534515 41847 534518
rect 683254 534309 683314 534480
rect 683254 534304 683363 534309
rect 683254 534248 683302 534304
rect 683358 534248 683363 534304
rect 683254 534246 683363 534248
rect 683297 534243 683363 534246
rect 676029 534102 676095 534105
rect 676029 534100 676292 534102
rect 676029 534044 676034 534100
rect 676090 534044 676292 534100
rect 676029 534042 676292 534044
rect 676029 534039 676095 534042
rect 40718 533836 40724 533900
rect 40788 533898 40794 533900
rect 42609 533898 42675 533901
rect 40788 533896 42675 533898
rect 40788 533840 42614 533896
rect 42670 533840 42675 533896
rect 40788 533838 42675 533840
rect 40788 533836 40794 533838
rect 42609 533835 42675 533838
rect 683622 533493 683682 533664
rect 683622 533488 683731 533493
rect 683622 533432 683670 533488
rect 683726 533432 683731 533488
rect 683622 533430 683731 533432
rect 683665 533427 683731 533430
rect 676262 533085 676322 533256
rect 676213 533080 676322 533085
rect 676213 533024 676218 533080
rect 676274 533024 676322 533080
rect 676213 533022 676322 533024
rect 676213 533019 676279 533022
rect 62113 532810 62179 532813
rect 62113 532808 64492 532810
rect 62113 532752 62118 532808
rect 62174 532752 64492 532808
rect 62113 532750 64492 532752
rect 62113 532747 62179 532750
rect 677366 532677 677426 532848
rect 41822 532612 41828 532676
rect 41892 532674 41898 532676
rect 42333 532674 42399 532677
rect 41892 532672 42399 532674
rect 41892 532616 42338 532672
rect 42394 532616 42399 532672
rect 41892 532614 42399 532616
rect 41892 532612 41898 532614
rect 42333 532611 42399 532614
rect 677317 532672 677426 532677
rect 677317 532616 677322 532672
rect 677378 532616 677426 532672
rect 677317 532614 677426 532616
rect 677317 532611 677383 532614
rect 676262 532269 676322 532440
rect 676213 532264 676322 532269
rect 676213 532208 676218 532264
rect 676274 532208 676322 532264
rect 676213 532206 676322 532208
rect 676213 532203 676279 532206
rect 677550 531861 677610 532032
rect 677501 531856 677610 531861
rect 677501 531800 677506 531856
rect 677562 531800 677610 531856
rect 677501 531798 677610 531800
rect 678237 531858 678303 531861
rect 678237 531856 678346 531858
rect 678237 531800 678242 531856
rect 678298 531800 678346 531856
rect 677501 531795 677567 531798
rect 678237 531795 678346 531800
rect 678286 531624 678346 531795
rect 676262 531045 676322 531216
rect 676213 531040 676322 531045
rect 676213 530984 676218 531040
rect 676274 530984 676322 531040
rect 676213 530982 676322 530984
rect 680997 531042 681063 531045
rect 680997 531040 681106 531042
rect 680997 530984 681002 531040
rect 681058 530984 681106 531040
rect 676213 530979 676279 530982
rect 680997 530979 681106 530984
rect 681046 530808 681106 530979
rect 40534 530708 40540 530772
rect 40604 530770 40610 530772
rect 41781 530770 41847 530773
rect 40604 530768 41847 530770
rect 40604 530712 41786 530768
rect 41842 530712 41847 530768
rect 40604 530710 41847 530712
rect 40604 530708 40610 530710
rect 41781 530707 41847 530710
rect 676029 530430 676095 530433
rect 676029 530428 676292 530430
rect 676029 530372 676034 530428
rect 676090 530372 676292 530428
rect 676029 530370 676292 530372
rect 676029 530367 676095 530370
rect 676990 530164 676996 530228
rect 677060 530164 677066 530228
rect 676998 529992 677058 530164
rect 41454 529892 41460 529956
rect 41524 529954 41530 529956
rect 41524 529894 42258 529954
rect 41524 529892 41530 529894
rect 42198 529546 42258 529894
rect 42333 529546 42399 529549
rect 42198 529544 42399 529546
rect 42198 529488 42338 529544
rect 42394 529488 42399 529544
rect 42198 529486 42399 529488
rect 42333 529483 42399 529486
rect 41638 529348 41644 529412
rect 41708 529410 41714 529412
rect 42609 529410 42675 529413
rect 41708 529408 42675 529410
rect 41708 529352 42614 529408
rect 42670 529352 42675 529408
rect 41708 529350 42675 529352
rect 41708 529348 41714 529350
rect 42609 529347 42675 529350
rect 676121 529410 676187 529413
rect 676262 529410 676322 529584
rect 676121 529408 676322 529410
rect 676121 529352 676126 529408
rect 676182 529352 676322 529408
rect 676121 529350 676322 529352
rect 676121 529347 676187 529350
rect 676262 529005 676322 529176
rect 676213 529000 676322 529005
rect 676213 528944 676218 529000
rect 676274 528944 676322 529000
rect 676213 528942 676322 528944
rect 676213 528939 676279 528942
rect 676029 528798 676095 528801
rect 676029 528796 676292 528798
rect 676029 528740 676034 528796
rect 676090 528740 676292 528796
rect 676029 528738 676292 528740
rect 676029 528735 676095 528738
rect 676029 528390 676095 528393
rect 676029 528388 676292 528390
rect 676029 528332 676034 528388
rect 676090 528332 676292 528388
rect 676029 528330 676292 528332
rect 676029 528327 676095 528330
rect 676806 528124 676812 528188
rect 676876 528124 676882 528188
rect 676814 527952 676874 528124
rect 676438 527716 676444 527780
rect 676508 527716 676514 527780
rect 676446 527544 676506 527716
rect 676262 526965 676322 527136
rect 676213 526960 676322 526965
rect 676213 526904 676218 526960
rect 676274 526904 676322 526960
rect 676213 526902 676322 526904
rect 676213 526899 676279 526902
rect 676029 526758 676095 526761
rect 676029 526756 676292 526758
rect 676029 526700 676034 526756
rect 676090 526700 676292 526756
rect 676029 526698 676292 526700
rect 676029 526695 676095 526698
rect 676029 526350 676095 526353
rect 676029 526348 676292 526350
rect 676029 526292 676034 526348
rect 676090 526292 676292 526348
rect 676029 526290 676292 526292
rect 676029 526287 676095 526290
rect 683070 525741 683130 525912
rect 683070 525736 683179 525741
rect 683070 525680 683118 525736
rect 683174 525680 683179 525736
rect 683070 525678 683179 525680
rect 683113 525675 683179 525678
rect 685830 525096 685890 525504
rect 683113 524922 683179 524925
rect 683070 524920 683179 524922
rect 683070 524864 683118 524920
rect 683174 524864 683179 524920
rect 683070 524859 683179 524864
rect 683070 524688 683130 524859
rect 651557 524242 651623 524245
rect 650164 524240 651623 524242
rect 650164 524184 651562 524240
rect 651618 524184 651623 524240
rect 650164 524182 651623 524184
rect 651557 524179 651623 524182
rect 62113 519754 62179 519757
rect 62113 519752 64492 519754
rect 62113 519696 62118 519752
rect 62174 519696 64492 519752
rect 62113 519694 64492 519696
rect 62113 519691 62179 519694
rect 667062 518591 677700 518701
rect 667062 514047 667329 518591
rect 669713 514047 677700 518591
rect 667062 513921 677700 514047
rect 651557 511050 651623 511053
rect 650164 511048 651623 511050
rect 650164 510992 651562 511048
rect 651618 510992 651623 511048
rect 650164 510990 651623 510992
rect 651557 510987 651623 510990
rect 667062 508601 677700 508722
rect 62113 506698 62179 506701
rect 62113 506696 64492 506698
rect 62113 506640 62118 506696
rect 62174 506640 64492 506696
rect 62113 506638 64492 506640
rect 62113 506635 62179 506638
rect 667062 504057 667343 508601
rect 669727 504057 677700 508601
rect 667062 503942 677700 504057
rect 675886 503644 675892 503708
rect 675956 503706 675962 503708
rect 679617 503706 679683 503709
rect 675956 503704 679683 503706
rect 675956 503648 679622 503704
rect 679678 503648 679683 503704
rect 675956 503646 679683 503648
rect 675956 503644 675962 503646
rect 679617 503643 679683 503646
rect 675334 503508 675340 503572
rect 675404 503570 675410 503572
rect 679801 503570 679867 503573
rect 675404 503568 679867 503570
rect 675404 503512 679806 503568
rect 679862 503512 679867 503568
rect 675404 503510 679867 503512
rect 675404 503508 675410 503510
rect 679801 503507 679867 503510
rect 39924 497743 52292 497858
rect 39924 493239 50356 497743
rect 52100 493239 52292 497743
rect 651557 497722 651623 497725
rect 650164 497720 651623 497722
rect 650164 497664 651562 497720
rect 651618 497664 651623 497720
rect 650164 497662 651623 497664
rect 651557 497659 651623 497662
rect 62113 493642 62179 493645
rect 62113 493640 64492 493642
rect 62113 493584 62118 493640
rect 62174 493584 64492 493640
rect 62113 493582 64492 493584
rect 62113 493579 62179 493582
rect 39924 493078 52292 493239
rect 675937 492146 676003 492149
rect 675937 492144 676292 492146
rect 675937 492088 675942 492144
rect 675998 492088 676292 492144
rect 675937 492086 676292 492088
rect 675937 492083 676003 492086
rect 676029 491738 676095 491741
rect 676029 491736 676292 491738
rect 676029 491680 676034 491736
rect 676090 491680 676292 491736
rect 676029 491678 676292 491680
rect 676029 491675 676095 491678
rect 676029 491330 676095 491333
rect 676029 491328 676292 491330
rect 676029 491272 676034 491328
rect 676090 491272 676292 491328
rect 676029 491270 676292 491272
rect 676029 491267 676095 491270
rect 676029 490922 676095 490925
rect 676029 490920 676292 490922
rect 676029 490864 676034 490920
rect 676090 490864 676292 490920
rect 676029 490862 676292 490864
rect 676029 490859 676095 490862
rect 676029 490514 676095 490517
rect 676029 490512 676292 490514
rect 676029 490456 676034 490512
rect 676090 490456 676292 490512
rect 676029 490454 676292 490456
rect 676029 490451 676095 490454
rect 675845 490106 675911 490109
rect 675845 490104 676292 490106
rect 675845 490048 675850 490104
rect 675906 490048 676292 490104
rect 675845 490046 676292 490048
rect 675845 490043 675911 490046
rect 677409 489930 677475 489933
rect 677366 489928 677475 489930
rect 677366 489872 677414 489928
rect 677470 489872 677475 489928
rect 677366 489867 677475 489872
rect 677366 489668 677426 489867
rect 675937 489290 676003 489293
rect 675937 489288 676292 489290
rect 675937 489232 675942 489288
rect 675998 489232 676292 489288
rect 675937 489230 676292 489232
rect 675937 489227 676003 489230
rect 675937 488882 676003 488885
rect 675937 488880 676292 488882
rect 675937 488824 675942 488880
rect 675998 488824 676292 488880
rect 675937 488822 676292 488824
rect 675937 488819 676003 488822
rect 675937 488474 676003 488477
rect 675937 488472 676292 488474
rect 675937 488416 675942 488472
rect 675998 488416 676292 488472
rect 675937 488414 676292 488416
rect 675937 488411 676003 488414
rect 675845 488066 675911 488069
rect 675845 488064 676292 488066
rect 675845 488008 675850 488064
rect 675906 488008 676292 488064
rect 675845 488006 676292 488008
rect 675845 488003 675911 488006
rect 39924 487753 52292 487879
rect 39924 483249 50344 487753
rect 52088 483249 52292 487753
rect 676070 487732 676076 487796
rect 676140 487732 676146 487796
rect 676078 487658 676138 487732
rect 676078 487598 676292 487658
rect 675937 487250 676003 487253
rect 675937 487248 676292 487250
rect 675937 487192 675942 487248
rect 675998 487192 676292 487248
rect 675937 487190 676292 487192
rect 675937 487187 676003 487190
rect 679617 486842 679683 486845
rect 679604 486840 679683 486842
rect 679604 486784 679622 486840
rect 679678 486784 679683 486840
rect 679604 486782 679683 486784
rect 679617 486779 679683 486782
rect 679801 486434 679867 486437
rect 679788 486432 679867 486434
rect 679788 486376 679806 486432
rect 679862 486376 679867 486432
rect 679788 486374 679867 486376
rect 679801 486371 679867 486374
rect 675937 486026 676003 486029
rect 675937 486024 676292 486026
rect 675937 485968 675942 486024
rect 675998 485968 676292 486024
rect 675937 485966 676292 485968
rect 675937 485963 676003 485966
rect 674741 485618 674807 485621
rect 674741 485616 676292 485618
rect 674741 485560 674746 485616
rect 674802 485560 676292 485616
rect 674741 485558 676292 485560
rect 674741 485555 674807 485558
rect 675845 485210 675911 485213
rect 675845 485208 676292 485210
rect 675845 485152 675850 485208
rect 675906 485152 676292 485208
rect 675845 485150 676292 485152
rect 675845 485147 675911 485150
rect 675937 484802 676003 484805
rect 675937 484800 676292 484802
rect 675937 484744 675942 484800
rect 675998 484744 676292 484800
rect 675937 484742 676292 484744
rect 675937 484739 676003 484742
rect 676254 484570 676260 484634
rect 676324 484570 676330 484634
rect 651557 484530 651623 484533
rect 650164 484528 651623 484530
rect 650164 484472 651562 484528
rect 651618 484472 651623 484528
rect 650164 484470 651623 484472
rect 651557 484467 651623 484470
rect 676262 484364 676322 484570
rect 676078 483926 676292 483986
rect 676078 483852 676138 483926
rect 676070 483788 676076 483852
rect 676140 483788 676146 483852
rect 675937 483578 676003 483581
rect 675937 483576 676292 483578
rect 675937 483520 675942 483576
rect 675998 483520 676292 483576
rect 675937 483518 676292 483520
rect 675937 483515 676003 483518
rect 39924 483099 52292 483249
rect 675937 483170 676003 483173
rect 675937 483168 676292 483170
rect 675937 483112 675942 483168
rect 675998 483112 676292 483168
rect 675937 483110 676292 483112
rect 675937 483107 676003 483110
rect 675845 482762 675911 482765
rect 675845 482760 676292 482762
rect 675845 482704 675850 482760
rect 675906 482704 676292 482760
rect 675845 482702 676292 482704
rect 675845 482699 675911 482702
rect 675937 482354 676003 482357
rect 675937 482352 676292 482354
rect 675937 482296 675942 482352
rect 675998 482296 676292 482352
rect 675937 482294 676292 482296
rect 675937 482291 676003 482294
rect 676078 481886 676292 481946
rect 676078 480722 676138 481886
rect 685830 481100 685890 481508
rect 678973 480722 679039 480725
rect 676078 480720 679166 480722
rect 676078 480664 678978 480720
rect 679034 480664 679166 480720
rect 676078 480662 679166 480664
rect 678973 480659 679039 480662
rect 62113 480586 62179 480589
rect 62113 480584 64492 480586
rect 62113 480528 62118 480584
rect 62174 480528 64492 480584
rect 62113 480526 64492 480528
rect 62113 480523 62179 480526
rect 651649 471202 651715 471205
rect 650164 471200 651715 471202
rect 650164 471144 651654 471200
rect 651710 471144 651715 471200
rect 650164 471142 651715 471144
rect 651649 471139 651715 471142
rect 62113 467530 62179 467533
rect 62113 467528 64492 467530
rect 62113 467472 62118 467528
rect 62174 467472 64492 467528
rect 62113 467470 64492 467472
rect 62113 467467 62179 467470
rect 651557 457874 651623 457877
rect 650164 457872 651623 457874
rect 650164 457816 651562 457872
rect 651618 457816 651623 457872
rect 650164 457814 651623 457816
rect 651557 457811 651623 457814
rect 62113 454610 62179 454613
rect 62113 454608 64492 454610
rect 62113 454552 62118 454608
rect 62174 454552 64492 454608
rect 62113 454550 64492 454552
rect 62113 454547 62179 454550
rect 651557 444546 651623 444549
rect 650164 444544 651623 444546
rect 650164 444488 651562 444544
rect 651618 444488 651623 444544
rect 650164 444486 651623 444488
rect 651557 444483 651623 444486
rect 62113 441554 62179 441557
rect 62113 441552 64492 441554
rect 62113 441496 62118 441552
rect 62174 441496 64492 441552
rect 62113 441494 64492 441496
rect 62113 441491 62179 441494
rect 6022 437353 63922 437382
rect 6022 436209 6150 437353
rect 6854 437349 63922 437353
rect 6854 436245 54235 437349
rect 55339 437329 63922 437349
rect 55339 436245 63339 437329
rect 6854 436225 63339 436245
rect 63883 436225 63922 437329
rect 6854 436209 63922 436225
rect 6022 436182 63922 436209
rect 7236 435757 62944 435782
rect 7236 434613 7348 435757
rect 8052 435731 62944 435757
rect 8052 434627 52641 435731
rect 53745 435721 62944 435731
rect 53745 434627 62371 435721
rect 8052 434617 62371 434627
rect 62915 434617 62944 435721
rect 8052 434613 62944 434617
rect 7236 434582 62944 434613
rect 651557 431354 651623 431357
rect 650164 431352 651623 431354
rect 650164 431296 651562 431352
rect 651618 431296 651623 431352
rect 650164 431294 651623 431296
rect 651557 431291 651623 431294
rect 43345 430946 43411 430949
rect 41492 430944 43411 430946
rect 41492 430888 43350 430944
rect 43406 430888 43411 430944
rect 41492 430886 43411 430888
rect 43345 430883 43411 430886
rect 41781 430538 41847 430541
rect 41492 430536 41847 430538
rect 41492 430480 41786 430536
rect 41842 430480 41847 430536
rect 41492 430478 41847 430480
rect 41781 430475 41847 430478
rect 663914 430389 677712 430501
rect 41781 430130 41847 430133
rect 41492 430128 41847 430130
rect 41492 430072 41786 430128
rect 41842 430072 41847 430128
rect 41492 430070 41847 430072
rect 41781 430067 41847 430070
rect 42885 429722 42951 429725
rect 41492 429720 42951 429722
rect 41492 429664 42890 429720
rect 42946 429664 42951 429720
rect 41492 429662 42951 429664
rect 42885 429659 42951 429662
rect 44357 429314 44423 429317
rect 41492 429312 44423 429314
rect 41492 429256 44362 429312
rect 44418 429256 44423 429312
rect 41492 429254 44423 429256
rect 44357 429251 44423 429254
rect 42793 428906 42859 428909
rect 41492 428904 42859 428906
rect 41492 428848 42798 428904
rect 42854 428848 42859 428904
rect 41492 428846 42859 428848
rect 42793 428843 42859 428846
rect 44265 428498 44331 428501
rect 41492 428496 44331 428498
rect 41492 428440 44270 428496
rect 44326 428440 44331 428496
rect 41492 428438 44331 428440
rect 44265 428435 44331 428438
rect 62113 428498 62179 428501
rect 62113 428496 64492 428498
rect 62113 428440 62118 428496
rect 62174 428440 64492 428496
rect 62113 428438 64492 428440
rect 62113 428435 62179 428438
rect 44173 428090 44239 428093
rect 41492 428088 44239 428090
rect 41492 428032 44178 428088
rect 44234 428032 44239 428088
rect 41492 428030 44239 428032
rect 44173 428027 44239 428030
rect 43161 427682 43227 427685
rect 41492 427680 43227 427682
rect 41492 427624 43166 427680
rect 43222 427624 43227 427680
rect 41492 427622 43227 427624
rect 43161 427619 43227 427622
rect 44633 427274 44699 427277
rect 41492 427272 44699 427274
rect 41492 427216 44638 427272
rect 44694 427216 44699 427272
rect 41492 427214 44699 427216
rect 44633 427211 44699 427214
rect 42885 426866 42951 426869
rect 41492 426864 42951 426866
rect 41492 426808 42890 426864
rect 42946 426808 42951 426864
rect 41492 426806 42951 426808
rect 42885 426803 42951 426806
rect 41781 426458 41847 426461
rect 41492 426456 41847 426458
rect 41492 426400 41786 426456
rect 41842 426400 41847 426456
rect 41492 426398 41847 426400
rect 41781 426395 41847 426398
rect 42190 426050 42196 426052
rect 41492 425990 42196 426050
rect 42190 425988 42196 425990
rect 42260 425988 42266 426052
rect 663914 425685 664125 430389
rect 666549 425748 677712 430389
rect 666549 425685 667110 425748
rect 41822 425642 41828 425644
rect 41492 425582 41828 425642
rect 41822 425580 41828 425582
rect 41892 425580 41898 425644
rect 663914 425562 667110 425685
rect 35157 425234 35223 425237
rect 35157 425232 35236 425234
rect 35157 425176 35162 425232
rect 35218 425176 35236 425232
rect 35157 425174 35236 425176
rect 35157 425171 35223 425174
rect 40769 425072 40835 425073
rect 40718 425070 40724 425072
rect 40678 425010 40724 425070
rect 40788 425068 40835 425072
rect 41321 425070 41387 425073
rect 40830 425012 40835 425068
rect 40718 425008 40724 425010
rect 40788 425008 40835 425012
rect 40769 425007 40835 425008
rect 41278 425068 41387 425070
rect 41278 425012 41326 425068
rect 41382 425012 41387 425068
rect 41278 425007 41387 425012
rect 41278 424796 41338 425007
rect 32397 424418 32463 424421
rect 32397 424416 32476 424418
rect 32397 424360 32402 424416
rect 32458 424360 32476 424416
rect 32397 424358 32476 424360
rect 32397 424355 32463 424358
rect 41822 424010 41828 424012
rect 41492 423950 41828 424010
rect 41822 423948 41828 423950
rect 41892 423948 41898 424012
rect 42006 423602 42012 423604
rect 41492 423542 42012 423602
rect 42006 423540 42012 423542
rect 42076 423540 42082 423604
rect 44357 423194 44423 423197
rect 41492 423192 44423 423194
rect 41492 423136 44362 423192
rect 44418 423136 44423 423192
rect 41492 423134 44423 423136
rect 44357 423131 44423 423134
rect 41822 422786 41828 422788
rect 41492 422726 41828 422786
rect 41822 422724 41828 422726
rect 41892 422724 41898 422788
rect 31017 422378 31083 422381
rect 31004 422376 31083 422378
rect 31004 422320 31022 422376
rect 31078 422320 31083 422376
rect 31004 422318 31083 422320
rect 31017 422315 31083 422318
rect 42793 421970 42859 421973
rect 41492 421968 42859 421970
rect 41492 421912 42798 421968
rect 42854 421912 42859 421968
rect 41492 421910 42859 421912
rect 42793 421907 42859 421910
rect 44449 421562 44515 421565
rect 41492 421560 44515 421562
rect 41492 421504 44454 421560
rect 44510 421504 44515 421560
rect 41492 421502 44515 421504
rect 44449 421499 44515 421502
rect 43069 421154 43135 421157
rect 41492 421152 43135 421154
rect 41492 421096 43074 421152
rect 43130 421096 43135 421152
rect 41492 421094 43135 421096
rect 43069 421091 43135 421094
rect 30598 420868 30604 420932
rect 30668 420868 30674 420932
rect 30606 420716 30666 420868
rect 663914 420471 677712 420522
rect 21774 419900 21834 420308
rect 41781 419522 41847 419525
rect 41492 419520 41847 419522
rect 21774 419386 21834 419492
rect 41492 419464 41786 419520
rect 41842 419464 41847 419520
rect 41492 419462 41847 419464
rect 41781 419459 41847 419462
rect 21406 419326 21834 419386
rect 21406 418842 21466 419326
rect 30598 418842 30604 418844
rect 21406 418782 30604 418842
rect 30598 418780 30604 418782
rect 30668 418780 30674 418844
rect 41321 418026 41387 418029
rect 41638 418026 41644 418028
rect 41321 418024 41644 418026
rect 41321 417968 41326 418024
rect 41382 417968 41644 418024
rect 41321 417966 41644 417968
rect 41321 417963 41387 417966
rect 41638 417964 41644 417966
rect 41708 417964 41714 418028
rect 651557 418026 651623 418029
rect 650164 418024 651623 418026
rect 650164 417968 651562 418024
rect 651618 417968 651623 418024
rect 650164 417966 651623 417968
rect 651557 417963 651623 417966
rect 663914 415847 664108 420471
rect 666532 415847 677712 420471
rect 663914 415742 677712 415847
rect 62113 415442 62179 415445
rect 62113 415440 64492 415442
rect 62113 415384 62118 415440
rect 62174 415384 64492 415440
rect 62113 415382 64492 415384
rect 62113 415379 62179 415382
rect 35157 414626 35223 414629
rect 41822 414626 41828 414628
rect 35157 414624 41828 414626
rect 35157 414568 35162 414624
rect 35218 414568 41828 414624
rect 35157 414566 41828 414568
rect 35157 414563 35223 414566
rect 41822 414564 41828 414566
rect 41892 414564 41898 414628
rect 42149 411226 42215 411229
rect 42374 411226 42380 411228
rect 42149 411224 42380 411226
rect 42149 411168 42154 411224
rect 42210 411168 42380 411224
rect 42149 411166 42380 411168
rect 42149 411163 42215 411166
rect 42374 411164 42380 411166
rect 42444 411164 42450 411228
rect 41086 409396 41092 409460
rect 41156 409458 41162 409460
rect 41781 409458 41847 409461
rect 41156 409456 41847 409458
rect 41156 409400 41786 409456
rect 41842 409400 41847 409456
rect 41156 409398 41847 409400
rect 41156 409396 41162 409398
rect 41781 409395 41847 409398
rect 41638 406268 41644 406332
rect 41708 406330 41714 406332
rect 41781 406330 41847 406333
rect 41708 406328 41847 406330
rect 41708 406272 41786 406328
rect 41842 406272 41847 406328
rect 41708 406270 41847 406272
rect 41708 406268 41714 406270
rect 41781 406267 41847 406270
rect 652017 404698 652083 404701
rect 650164 404696 652083 404698
rect 650164 404640 652022 404696
rect 652078 404640 652083 404696
rect 650164 404638 652083 404640
rect 652017 404635 652083 404638
rect 676262 403749 676322 403852
rect 676213 403744 676322 403749
rect 676213 403688 676218 403744
rect 676274 403688 676322 403744
rect 676213 403686 676322 403688
rect 676213 403683 676279 403686
rect 676446 403341 676506 403444
rect 676213 403338 676279 403341
rect 676213 403336 676322 403338
rect 676213 403280 676218 403336
rect 676274 403280 676322 403336
rect 676213 403275 676322 403280
rect 676397 403336 676506 403341
rect 676397 403280 676402 403336
rect 676458 403280 676506 403336
rect 676397 403278 676506 403280
rect 676397 403275 676463 403278
rect 676262 403036 676322 403275
rect 676029 402658 676095 402661
rect 676029 402656 676292 402658
rect 676029 402600 676034 402656
rect 676090 402600 676292 402656
rect 676029 402598 676292 402600
rect 676029 402595 676095 402598
rect 41454 402460 41460 402524
rect 41524 402522 41530 402524
rect 41781 402522 41847 402525
rect 41524 402520 41847 402522
rect 41524 402464 41786 402520
rect 41842 402464 41847 402520
rect 41524 402462 41847 402464
rect 41524 402460 41530 402462
rect 41781 402459 41847 402462
rect 62113 402386 62179 402389
rect 62113 402384 64492 402386
rect 62113 402328 62118 402384
rect 62174 402328 64492 402384
rect 62113 402326 64492 402328
rect 62113 402323 62179 402326
rect 676262 402117 676322 402220
rect 676213 402112 676322 402117
rect 676213 402056 676218 402112
rect 676274 402056 676322 402112
rect 676213 402054 676322 402056
rect 677317 402114 677383 402117
rect 677317 402112 677426 402114
rect 677317 402056 677322 402112
rect 677378 402056 677426 402112
rect 676213 402051 676279 402054
rect 677317 402051 677426 402056
rect 41965 401844 42031 401845
rect 41965 401840 42012 401844
rect 42076 401842 42082 401844
rect 41965 401784 41970 401840
rect 41965 401780 42012 401784
rect 42076 401782 42122 401842
rect 677366 401812 677426 402051
rect 42076 401780 42082 401782
rect 41965 401779 42031 401780
rect 676121 401298 676187 401301
rect 676262 401298 676322 401404
rect 676121 401296 676322 401298
rect 676121 401240 676126 401296
rect 676182 401240 676322 401296
rect 676121 401238 676322 401240
rect 676121 401235 676187 401238
rect 676029 401026 676095 401029
rect 676029 401024 676292 401026
rect 676029 400968 676034 401024
rect 676090 400968 676292 401024
rect 676029 400966 676292 400968
rect 676029 400963 676095 400966
rect 676262 400485 676322 400588
rect 676213 400480 676322 400485
rect 677225 400482 677291 400485
rect 676213 400424 676218 400480
rect 676274 400424 676322 400480
rect 676213 400422 676322 400424
rect 677182 400480 677291 400482
rect 677182 400424 677230 400480
rect 677286 400424 677291 400480
rect 676213 400419 676279 400422
rect 677182 400419 677291 400424
rect 677182 400180 677242 400419
rect 40718 400012 40724 400076
rect 40788 400074 40794 400076
rect 41781 400074 41847 400077
rect 40788 400072 41847 400074
rect 40788 400016 41786 400072
rect 41842 400016 41847 400072
rect 40788 400014 41847 400016
rect 40788 400012 40794 400014
rect 41781 400011 41847 400014
rect 676262 399669 676322 399772
rect 40902 399604 40908 399668
rect 40972 399666 40978 399668
rect 41781 399666 41847 399669
rect 40972 399664 41847 399666
rect 40972 399608 41786 399664
rect 41842 399608 41847 399664
rect 40972 399606 41847 399608
rect 40972 399604 40978 399606
rect 41781 399603 41847 399606
rect 676213 399664 676322 399669
rect 676213 399608 676218 399664
rect 676274 399608 676322 399664
rect 676213 399606 676322 399608
rect 676213 399603 676279 399606
rect 675702 399332 675708 399396
rect 675772 399394 675778 399396
rect 675772 399334 676292 399394
rect 675772 399332 675778 399334
rect 40534 398788 40540 398852
rect 40604 398850 40610 398852
rect 41781 398850 41847 398853
rect 676262 398852 676322 398956
rect 40604 398848 41847 398850
rect 40604 398792 41786 398848
rect 41842 398792 41847 398848
rect 40604 398790 41847 398792
rect 40604 398788 40610 398790
rect 41781 398787 41847 398790
rect 676254 398788 676260 398852
rect 676324 398788 676330 398852
rect 676029 398578 676095 398581
rect 676029 398576 676292 398578
rect 676029 398520 676034 398576
rect 676090 398520 676292 398576
rect 676029 398518 676292 398520
rect 676029 398515 676095 398518
rect 676029 398170 676095 398173
rect 676029 398168 676292 398170
rect 676029 398112 676034 398168
rect 676090 398112 676292 398168
rect 676029 398110 676292 398112
rect 676029 398107 676095 398110
rect 676814 397629 676874 397732
rect 676814 397624 676923 397629
rect 676814 397568 676862 397624
rect 676918 397568 676923 397624
rect 676814 397566 676923 397568
rect 676857 397563 676923 397566
rect 676446 397220 676506 397324
rect 676438 397156 676444 397220
rect 676508 397156 676514 397220
rect 676998 396813 677058 396916
rect 676949 396808 677058 396813
rect 676949 396752 676954 396808
rect 677010 396752 677058 396808
rect 676949 396750 677058 396752
rect 676949 396747 677015 396750
rect 679574 396405 679634 396508
rect 679574 396400 679683 396405
rect 679574 396344 679622 396400
rect 679678 396344 679683 396400
rect 679574 396342 679683 396344
rect 679617 396339 679683 396342
rect 678286 395997 678346 396100
rect 678237 395992 678346 395997
rect 678237 395936 678242 395992
rect 678298 395936 678346 395992
rect 678237 395934 678346 395936
rect 678237 395931 678303 395934
rect 676070 395524 676076 395588
rect 676140 395586 676146 395588
rect 676262 395586 676322 395692
rect 676140 395526 676322 395586
rect 676140 395524 676146 395526
rect 675886 395252 675892 395316
rect 675956 395314 675962 395316
rect 675956 395254 676292 395314
rect 675956 395252 675962 395254
rect 676446 394773 676506 394876
rect 676446 394768 676555 394773
rect 676446 394712 676494 394768
rect 676550 394712 676555 394768
rect 676446 394710 676555 394712
rect 676489 394707 676555 394710
rect 676262 394365 676322 394468
rect 676213 394360 676322 394365
rect 676213 394304 676218 394360
rect 676274 394304 676322 394360
rect 676213 394302 676322 394304
rect 676213 394299 676279 394302
rect 6022 394153 63922 394182
rect 6022 393009 6150 394153
rect 6854 394149 63922 394153
rect 6854 393045 54235 394149
rect 55339 394129 63922 394149
rect 55339 393045 63339 394129
rect 6854 393025 63339 393045
rect 63883 393025 63922 394129
rect 676029 394090 676095 394093
rect 676029 394088 676292 394090
rect 676029 394032 676034 394088
rect 676090 394032 676292 394088
rect 676029 394030 676292 394032
rect 676029 394027 676095 394030
rect 683070 393549 683130 393652
rect 683070 393544 683179 393549
rect 683070 393488 683118 393544
rect 683174 393488 683179 393544
rect 683070 393486 683179 393488
rect 683113 393483 683179 393486
rect 6854 393009 63922 393025
rect 6022 392982 63922 393009
rect 685830 392836 685890 393244
rect 7236 392557 62944 392582
rect 7236 391413 7348 392557
rect 8052 392531 62944 392557
rect 8052 391427 52641 392531
rect 53745 392521 62944 392531
rect 53745 391427 62371 392521
rect 8052 391417 62371 391427
rect 62915 391417 62944 392521
rect 683070 392325 683130 392428
rect 683070 392320 683179 392325
rect 683070 392264 683118 392320
rect 683174 392264 683179 392320
rect 683070 392262 683179 392264
rect 683113 392259 683179 392262
rect 651557 391506 651623 391509
rect 650164 391504 651623 391506
rect 650164 391448 651562 391504
rect 651618 391448 651623 391504
rect 650164 391446 651623 391448
rect 651557 391443 651623 391446
rect 8052 391413 62944 391417
rect 7236 391382 62944 391413
rect 62113 389330 62179 389333
rect 62113 389328 64492 389330
rect 62113 389272 62118 389328
rect 62174 389272 64492 389328
rect 62113 389270 64492 389272
rect 62113 389267 62179 389270
rect 675518 388452 675524 388516
rect 675588 388514 675594 388516
rect 676857 388514 676923 388517
rect 675588 388512 676923 388514
rect 675588 388456 676862 388512
rect 676918 388456 676923 388512
rect 675588 388454 676923 388456
rect 675588 388452 675594 388454
rect 676857 388451 676923 388454
rect 675334 388180 675340 388244
rect 675404 388242 675410 388244
rect 679617 388242 679683 388245
rect 675404 388240 679683 388242
rect 675404 388184 679622 388240
rect 679678 388184 679683 388240
rect 675404 388182 679683 388184
rect 675404 388180 675410 388182
rect 679617 388179 679683 388182
rect 35758 387565 35818 387668
rect 35758 387560 35867 387565
rect 35758 387504 35806 387560
rect 35862 387504 35867 387560
rect 35758 387502 35867 387504
rect 35801 387499 35867 387502
rect 35758 387157 35818 387260
rect 35617 387154 35683 387157
rect 35574 387152 35683 387154
rect 35574 387096 35622 387152
rect 35678 387096 35683 387152
rect 35574 387091 35683 387096
rect 35758 387152 35867 387157
rect 35758 387096 35806 387152
rect 35862 387096 35867 387152
rect 35758 387094 35867 387096
rect 35801 387091 35867 387094
rect 35574 386852 35634 387091
rect 35709 386746 35775 386749
rect 35709 386744 35818 386746
rect 35709 386688 35714 386744
rect 35770 386688 35818 386744
rect 35709 386683 35818 386688
rect 35758 386444 35818 386683
rect 44265 386066 44331 386069
rect 41492 386064 44331 386066
rect 41492 386008 44270 386064
rect 44326 386008 44331 386064
rect 41492 386006 44331 386008
rect 44265 386003 44331 386006
rect 44173 385658 44239 385661
rect 41492 385656 44239 385658
rect 41492 385600 44178 385656
rect 44234 385600 44239 385656
rect 41492 385598 44239 385600
rect 44173 385595 44239 385598
rect 44633 385250 44699 385253
rect 41492 385248 44699 385250
rect 41492 385192 44638 385248
rect 44694 385192 44699 385248
rect 41492 385190 44699 385192
rect 44633 385187 44699 385190
rect 675753 384980 675819 384981
rect 675702 384978 675708 384980
rect 675662 384918 675708 384978
rect 675772 384976 675819 384980
rect 675814 384920 675819 384976
rect 675702 384916 675708 384918
rect 675772 384916 675819 384920
rect 675753 384915 675819 384916
rect 43161 384842 43227 384845
rect 41492 384840 43227 384842
rect 41492 384784 43166 384840
rect 43222 384784 43227 384840
rect 41492 384782 43227 384784
rect 43161 384779 43227 384782
rect 44173 384434 44239 384437
rect 41492 384432 44239 384434
rect 41492 384376 44178 384432
rect 44234 384376 44239 384432
rect 41492 384374 44239 384376
rect 44173 384371 44239 384374
rect 42885 384026 42951 384029
rect 41492 384024 42951 384026
rect 41492 383968 42890 384024
rect 42946 383968 42951 384024
rect 41492 383966 42951 383968
rect 42885 383963 42951 383966
rect 42793 383618 42859 383621
rect 41492 383616 42859 383618
rect 41492 383560 42798 383616
rect 42854 383560 42859 383616
rect 41492 383558 42859 383560
rect 42793 383555 42859 383558
rect 40726 383076 40786 383180
rect 40718 383012 40724 383076
rect 40788 383012 40794 383076
rect 40910 382669 40970 382772
rect 40861 382664 40970 382669
rect 40861 382608 40866 382664
rect 40922 382608 40970 382664
rect 40861 382606 40970 382608
rect 40861 382603 40927 382606
rect 40542 382260 40602 382364
rect 675385 382260 675451 382261
rect 40534 382196 40540 382260
rect 40604 382196 40610 382260
rect 675334 382258 675340 382260
rect 675294 382198 675340 382258
rect 675404 382256 675451 382260
rect 675446 382200 675451 382256
rect 675334 382196 675340 382198
rect 675404 382196 675451 382200
rect 675385 382195 675451 382196
rect 41462 381852 41522 381956
rect 41454 381788 41460 381852
rect 41524 381788 41530 381852
rect 37966 381445 38026 381548
rect 37917 381440 38026 381445
rect 37917 381384 37922 381440
rect 37978 381384 38026 381440
rect 37917 381382 38026 381384
rect 37917 381379 37983 381382
rect 30974 381037 31034 381140
rect 30974 381032 31083 381037
rect 30974 380976 31022 381032
rect 31078 380976 31083 381032
rect 30974 380974 31083 380976
rect 31017 380971 31083 380974
rect 44449 380762 44515 380765
rect 41492 380760 44515 380762
rect 41492 380704 44454 380760
rect 44510 380704 44515 380760
rect 41492 380702 44515 380704
rect 44449 380699 44515 380702
rect 42885 380354 42951 380357
rect 41492 380352 42951 380354
rect 41492 380296 42890 380352
rect 42946 380296 42951 380352
rect 41492 380294 42951 380296
rect 42885 380291 42951 380294
rect 40910 379812 40970 379916
rect 40902 379748 40908 379812
rect 40972 379748 40978 379812
rect 40726 379405 40786 379508
rect 40677 379400 40786 379405
rect 40677 379344 40682 379400
rect 40738 379344 40786 379400
rect 40677 379342 40786 379344
rect 40677 379339 40743 379342
rect 44541 379130 44607 379133
rect 41492 379128 44607 379130
rect 41492 379072 44546 379128
rect 44602 379072 44607 379128
rect 41492 379070 44607 379072
rect 44541 379067 44607 379070
rect 42977 378722 43043 378725
rect 41492 378720 43043 378722
rect 41492 378664 42982 378720
rect 43038 378664 43043 378720
rect 41492 378662 43043 378664
rect 42977 378659 43043 378662
rect 675477 378724 675543 378725
rect 675477 378720 675524 378724
rect 675588 378722 675594 378724
rect 675477 378664 675482 378720
rect 675477 378660 675524 378664
rect 675588 378662 675634 378722
rect 675588 378660 675594 378662
rect 675477 378659 675543 378660
rect 33734 378181 33794 378284
rect 33734 378176 33843 378181
rect 651557 378178 651623 378181
rect 33734 378120 33782 378176
rect 33838 378120 33843 378176
rect 33734 378118 33843 378120
rect 650164 378176 651623 378178
rect 650164 378120 651562 378176
rect 651618 378120 651623 378176
rect 650164 378118 651623 378120
rect 33777 378115 33843 378118
rect 651557 378115 651623 378118
rect 43069 377906 43135 377909
rect 41492 377904 43135 377906
rect 41492 377848 43074 377904
rect 43130 377848 43135 377904
rect 41492 377846 43135 377848
rect 43069 377843 43135 377846
rect 35758 377365 35818 377468
rect 35758 377360 35867 377365
rect 35758 377304 35806 377360
rect 35862 377304 35867 377360
rect 35758 377302 35867 377304
rect 35801 377299 35867 377302
rect 675753 377362 675819 377365
rect 675886 377362 675892 377364
rect 675753 377360 675892 377362
rect 675753 377304 675758 377360
rect 675814 377304 675892 377360
rect 675753 377302 675892 377304
rect 675753 377299 675819 377302
rect 675886 377300 675892 377302
rect 675956 377300 675962 377364
rect 27662 376652 27722 377060
rect 62113 376274 62179 376277
rect 62113 376272 64492 376274
rect 41462 376141 41522 376244
rect 62113 376216 62118 376272
rect 62174 376216 64492 376272
rect 62113 376214 64492 376216
rect 62113 376211 62179 376214
rect 41462 376136 41571 376141
rect 41462 376080 41510 376136
rect 41566 376080 41571 376136
rect 41462 376078 41571 376080
rect 41505 376075 41571 376078
rect 675753 375050 675819 375053
rect 676070 375050 676076 375052
rect 675753 375048 676076 375050
rect 675753 374992 675758 375048
rect 675814 374992 676076 375048
rect 675753 374990 676076 374992
rect 675753 374987 675819 374990
rect 676070 374988 676076 374990
rect 676140 374988 676146 375052
rect 675753 373690 675819 373693
rect 676254 373690 676260 373692
rect 675753 373688 676260 373690
rect 675753 373632 675758 373688
rect 675814 373632 676260 373688
rect 675753 373630 676260 373632
rect 675753 373627 675819 373630
rect 676254 373628 676260 373630
rect 676324 373628 676330 373692
rect 675753 372058 675819 372061
rect 676438 372058 676444 372060
rect 675753 372056 676444 372058
rect 675753 372000 675758 372056
rect 675814 372000 676444 372056
rect 675753 371998 676444 372000
rect 675753 371995 675819 371998
rect 676438 371996 676444 371998
rect 676508 371996 676514 372060
rect 33777 371922 33843 371925
rect 42006 371922 42012 371924
rect 33777 371920 42012 371922
rect 33777 371864 33782 371920
rect 33838 371864 42012 371920
rect 33777 371862 42012 371864
rect 33777 371859 33843 371862
rect 42006 371860 42012 371862
rect 42076 371860 42082 371924
rect 37917 371378 37983 371381
rect 41638 371378 41644 371380
rect 37917 371376 41644 371378
rect 37917 371320 37922 371376
rect 37978 371320 41644 371376
rect 37917 371318 41644 371320
rect 37917 371315 37983 371318
rect 41638 371316 41644 371318
rect 41708 371316 41714 371380
rect 41781 370292 41847 370293
rect 41781 370290 41828 370292
rect 41736 370288 41828 370290
rect 41736 370232 41786 370288
rect 41736 370230 41828 370232
rect 41781 370228 41828 370230
rect 41892 370228 41898 370292
rect 41781 370227 41847 370228
rect 41873 366348 41939 366349
rect 41822 366346 41828 366348
rect 41782 366286 41828 366346
rect 41892 366344 41939 366348
rect 41934 366288 41939 366344
rect 41822 366284 41828 366286
rect 41892 366284 41939 366288
rect 41873 366283 41939 366284
rect 652017 364850 652083 364853
rect 650164 364848 652083 364850
rect 650164 364792 652022 364848
rect 652078 364792 652083 364848
rect 650164 364790 652083 364792
rect 652017 364787 652083 364790
rect 41965 363764 42031 363765
rect 41965 363760 42012 363764
rect 42076 363762 42082 363764
rect 41965 363704 41970 363760
rect 41965 363700 42012 363704
rect 42076 363702 42122 363762
rect 42076 363700 42082 363702
rect 41965 363699 42031 363700
rect 62113 363354 62179 363357
rect 62113 363352 64492 363354
rect 62113 363296 62118 363352
rect 62174 363296 64492 363352
rect 62113 363294 64492 363296
rect 62113 363291 62179 363294
rect 41638 362884 41644 362948
rect 41708 362946 41714 362948
rect 41781 362946 41847 362949
rect 41708 362944 41847 362946
rect 41708 362888 41786 362944
rect 41842 362888 41847 362944
rect 41708 362886 41847 362888
rect 41708 362884 41714 362886
rect 41781 362883 41847 362886
rect 40902 360164 40908 360228
rect 40972 360226 40978 360228
rect 40972 360166 41706 360226
rect 40972 360164 40978 360166
rect 41646 360090 41706 360166
rect 41781 360090 41847 360093
rect 41646 360088 41847 360090
rect 41646 360032 41786 360088
rect 41842 360032 41847 360088
rect 41646 360030 41847 360032
rect 41781 360027 41847 360030
rect 41454 358668 41460 358732
rect 41524 358730 41530 358732
rect 41781 358730 41847 358733
rect 41524 358728 41847 358730
rect 41524 358672 41786 358728
rect 41842 358672 41847 358728
rect 41524 358670 41847 358672
rect 41524 358668 41530 358670
rect 41781 358667 41847 358670
rect 675845 358730 675911 358733
rect 675845 358728 676292 358730
rect 675845 358672 675850 358728
rect 675906 358672 676292 358728
rect 675845 358670 676292 358672
rect 675845 358667 675911 358670
rect 675937 358322 676003 358325
rect 675937 358320 676292 358322
rect 675937 358264 675942 358320
rect 675998 358264 676292 358320
rect 675937 358262 676292 358264
rect 675937 358259 676003 358262
rect 676029 357914 676095 357917
rect 676029 357912 676292 357914
rect 676029 357856 676034 357912
rect 676090 357856 676292 357912
rect 676029 357854 676292 357856
rect 676029 357851 676095 357854
rect 676029 357506 676095 357509
rect 676029 357504 676292 357506
rect 676029 357448 676034 357504
rect 676090 357448 676292 357504
rect 676029 357446 676292 357448
rect 676029 357443 676095 357446
rect 676029 357098 676095 357101
rect 676029 357096 676292 357098
rect 676029 357040 676034 357096
rect 676090 357040 676292 357096
rect 676029 357038 676292 357040
rect 676029 357035 676095 357038
rect 40718 356900 40724 356964
rect 40788 356962 40794 356964
rect 41781 356962 41847 356965
rect 40788 356960 41847 356962
rect 40788 356904 41786 356960
rect 41842 356904 41847 356960
rect 40788 356902 41847 356904
rect 40788 356900 40794 356902
rect 41781 356899 41847 356902
rect 676029 356690 676095 356693
rect 676029 356688 676292 356690
rect 676029 356632 676034 356688
rect 676090 356632 676292 356688
rect 676029 356630 676292 356632
rect 676029 356627 676095 356630
rect 676029 356282 676095 356285
rect 676029 356280 676292 356282
rect 676029 356224 676034 356280
rect 676090 356224 676292 356280
rect 676029 356222 676292 356224
rect 676029 356219 676095 356222
rect 676029 355874 676095 355877
rect 676029 355872 676292 355874
rect 676029 355816 676034 355872
rect 676090 355816 676292 355872
rect 676029 355814 676292 355816
rect 676029 355811 676095 355814
rect 40534 355676 40540 355740
rect 40604 355738 40610 355740
rect 41781 355738 41847 355741
rect 40604 355736 41847 355738
rect 40604 355680 41786 355736
rect 41842 355680 41847 355736
rect 40604 355678 41847 355680
rect 40604 355676 40610 355678
rect 41781 355675 41847 355678
rect 676029 355466 676095 355469
rect 676029 355464 676292 355466
rect 676029 355408 676034 355464
rect 676090 355408 676292 355464
rect 676029 355406 676292 355408
rect 676029 355403 676095 355406
rect 674741 355058 674807 355061
rect 674741 355056 676292 355058
rect 674741 355000 674746 355056
rect 674802 355000 676292 355056
rect 674741 354998 676292 355000
rect 674741 354995 674807 354998
rect 676029 354650 676095 354653
rect 676029 354648 676292 354650
rect 676029 354592 676034 354648
rect 676090 354592 676292 354648
rect 676029 354590 676292 354592
rect 676029 354587 676095 354590
rect 675886 354180 675892 354244
rect 675956 354242 675962 354244
rect 675956 354182 676292 354242
rect 675956 354180 675962 354182
rect 676078 353774 676292 353834
rect 676078 353700 676138 353774
rect 676070 353636 676076 353700
rect 676140 353636 676146 353700
rect 675702 353364 675708 353428
rect 675772 353426 675778 353428
rect 675772 353366 676292 353426
rect 675772 353364 675778 353366
rect 675334 352956 675340 353020
rect 675404 353018 675410 353020
rect 675404 352958 676292 353018
rect 675404 352956 675410 352958
rect 679617 352610 679683 352613
rect 679604 352608 679683 352610
rect 679604 352552 679622 352608
rect 679678 352552 679683 352608
rect 679604 352550 679683 352552
rect 679617 352547 679683 352550
rect 676078 352142 676292 352202
rect 676078 352068 676138 352142
rect 676070 352004 676076 352068
rect 676140 352004 676146 352068
rect 679801 351794 679867 351797
rect 679788 351792 679867 351794
rect 55968 351729 63922 351782
rect 679788 351736 679806 351792
rect 679862 351736 679867 351792
rect 679788 351734 679867 351736
rect 679801 351731 679867 351734
rect 55968 350982 63339 351729
rect 6022 350953 63339 350982
rect 6022 349809 6150 350953
rect 6854 350949 63339 350953
rect 6854 349845 54235 350949
rect 55339 350625 63339 350949
rect 63883 350625 63922 351729
rect 651557 351658 651623 351661
rect 650164 351656 651623 351658
rect 650164 351600 651562 351656
rect 651618 351600 651623 351656
rect 650164 351598 651623 351600
rect 651557 351595 651623 351598
rect 676029 351386 676095 351389
rect 676029 351384 676292 351386
rect 676029 351328 676034 351384
rect 676090 351328 676292 351384
rect 676029 351326 676292 351328
rect 676029 351323 676095 351326
rect 676029 350978 676095 350981
rect 676029 350976 676292 350978
rect 676029 350920 676034 350976
rect 676090 350920 676292 350976
rect 676029 350918 676292 350920
rect 676029 350915 676095 350918
rect 55339 350582 63922 350625
rect 55339 349845 57264 350582
rect 676029 350570 676095 350573
rect 676029 350568 676292 350570
rect 676029 350512 676034 350568
rect 676090 350512 676292 350568
rect 676029 350510 676292 350512
rect 676029 350507 676095 350510
rect 62113 350298 62179 350301
rect 62113 350296 64492 350298
rect 62113 350240 62118 350296
rect 62174 350240 64492 350296
rect 62113 350238 64492 350240
rect 62113 350235 62179 350238
rect 676029 350162 676095 350165
rect 676029 350160 676292 350162
rect 676029 350104 676034 350160
rect 676090 350104 676292 350160
rect 676029 350102 676292 350104
rect 676029 350099 676095 350102
rect 6854 349809 57264 349845
rect 6022 349782 57264 349809
rect 675937 349754 676003 349757
rect 675937 349752 676292 349754
rect 675937 349696 675942 349752
rect 675998 349696 676292 349752
rect 675937 349694 676292 349696
rect 675937 349691 676003 349694
rect 7236 349357 62944 349382
rect 7236 348213 7348 349357
rect 8052 349331 62944 349357
rect 8052 348227 52641 349331
rect 53745 349321 62944 349331
rect 53745 348227 62371 349321
rect 8052 348217 62371 348227
rect 62915 348217 62944 349321
rect 676029 349346 676095 349349
rect 676029 349344 676292 349346
rect 676029 349288 676034 349344
rect 676090 349288 676292 349344
rect 676029 349286 676292 349288
rect 676029 349283 676095 349286
rect 676029 348938 676095 348941
rect 676029 348936 676292 348938
rect 676029 348880 676034 348936
rect 676090 348880 676292 348936
rect 676029 348878 676292 348880
rect 676029 348875 676095 348878
rect 676029 348530 676095 348533
rect 676029 348528 676292 348530
rect 676029 348472 676034 348528
rect 676090 348472 676292 348528
rect 676029 348470 676292 348472
rect 676029 348467 676095 348470
rect 8052 348213 62944 348217
rect 7236 348182 62944 348213
rect 676262 347684 676322 348092
rect 676029 347306 676095 347309
rect 676029 347304 676292 347306
rect 676029 347248 676034 347304
rect 676090 347248 676292 347304
rect 676029 347246 676292 347248
rect 676029 347243 676095 347246
rect 675937 346626 676003 346629
rect 676990 346626 676996 346628
rect 675937 346624 676996 346626
rect 675937 346568 675942 346624
rect 675998 346568 676996 346624
rect 675937 346566 676996 346568
rect 675937 346563 676003 346566
rect 676990 346564 676996 346566
rect 677060 346564 677066 346628
rect 676121 346490 676187 346493
rect 676765 346492 676831 346493
rect 676622 346490 676628 346492
rect 676121 346488 676628 346490
rect 676121 346432 676126 346488
rect 676182 346432 676628 346488
rect 676121 346430 676628 346432
rect 676121 346427 676187 346430
rect 676622 346428 676628 346430
rect 676692 346428 676698 346492
rect 676765 346488 676812 346492
rect 676876 346490 676882 346492
rect 676765 346432 676770 346488
rect 676765 346428 676812 346432
rect 676876 346430 676922 346490
rect 676876 346428 676882 346430
rect 676765 346427 676831 346428
rect 35574 344317 35634 344556
rect 35574 344312 35683 344317
rect 35801 344314 35867 344317
rect 35574 344256 35622 344312
rect 35678 344256 35683 344312
rect 35574 344254 35683 344256
rect 35617 344251 35683 344254
rect 35758 344312 35867 344314
rect 35758 344256 35806 344312
rect 35862 344256 35867 344312
rect 35758 344251 35867 344256
rect 35758 344148 35818 344251
rect 35709 343906 35775 343909
rect 35709 343904 35818 343906
rect 35709 343848 35714 343904
rect 35770 343848 35818 343904
rect 35709 343843 35818 343848
rect 35758 343740 35818 343843
rect 44265 343362 44331 343365
rect 41492 343360 44331 343362
rect 41492 343304 44270 343360
rect 44326 343304 44331 343360
rect 41492 343302 44331 343304
rect 44265 343299 44331 343302
rect 44357 342954 44423 342957
rect 41492 342952 44423 342954
rect 41492 342896 44362 342952
rect 44418 342896 44423 342952
rect 41492 342894 44423 342896
rect 44357 342891 44423 342894
rect 44633 342546 44699 342549
rect 41492 342544 44699 342546
rect 41492 342488 44638 342544
rect 44694 342488 44699 342544
rect 41492 342486 44699 342488
rect 44633 342483 44699 342486
rect 676070 342348 676076 342412
rect 676140 342410 676146 342412
rect 679617 342410 679683 342413
rect 676140 342408 679683 342410
rect 676140 342352 679622 342408
rect 679678 342352 679683 342408
rect 676140 342350 679683 342352
rect 676140 342348 676146 342350
rect 679617 342347 679683 342350
rect 675293 342274 675359 342277
rect 679801 342274 679867 342277
rect 675293 342272 679867 342274
rect 675293 342216 675298 342272
rect 675354 342216 679806 342272
rect 679862 342216 679867 342272
rect 675293 342214 679867 342216
rect 675293 342211 675359 342214
rect 679801 342211 679867 342214
rect 44265 342138 44331 342141
rect 41492 342136 44331 342138
rect 41492 342080 44270 342136
rect 44326 342080 44331 342136
rect 41492 342078 44331 342080
rect 44265 342075 44331 342078
rect 44173 341730 44239 341733
rect 41492 341728 44239 341730
rect 41492 341672 44178 341728
rect 44234 341672 44239 341728
rect 41492 341670 44239 341672
rect 44173 341667 44239 341670
rect 44357 341322 44423 341325
rect 41492 341320 44423 341322
rect 41492 341264 44362 341320
rect 44418 341264 44423 341320
rect 41492 341262 44423 341264
rect 44357 341259 44423 341262
rect 42793 340914 42859 340917
rect 41492 340912 42859 340914
rect 41492 340856 42798 340912
rect 42854 340856 42859 340912
rect 41492 340854 42859 340856
rect 42793 340851 42859 340854
rect 675661 340780 675727 340781
rect 675661 340776 675708 340780
rect 675772 340778 675778 340780
rect 675661 340720 675666 340776
rect 675661 340716 675708 340720
rect 675772 340718 675818 340778
rect 675772 340716 675778 340718
rect 675661 340715 675727 340716
rect 42793 340506 42859 340509
rect 41492 340504 42859 340506
rect 41492 340448 42798 340504
rect 42854 340448 42859 340504
rect 41492 340446 42859 340448
rect 42793 340443 42859 340446
rect 40726 339828 40786 340068
rect 40718 339764 40724 339828
rect 40788 339764 40794 339828
rect 40910 339421 40970 339660
rect 40861 339416 40970 339421
rect 40861 339360 40866 339416
rect 40922 339360 40970 339416
rect 40861 339358 40970 339360
rect 675753 339418 675819 339421
rect 675886 339418 675892 339420
rect 675753 339416 675892 339418
rect 675753 339360 675758 339416
rect 675814 339360 675892 339416
rect 675753 339358 675892 339360
rect 40861 339355 40927 339358
rect 675753 339355 675819 339358
rect 675886 339356 675892 339358
rect 675956 339356 675962 339420
rect 40542 339012 40602 339252
rect 40534 338948 40540 339012
rect 40604 338948 40610 339012
rect 41462 338604 41522 338844
rect 41454 338540 41460 338604
rect 41524 338540 41530 338604
rect 40726 338197 40786 338436
rect 651649 338330 651715 338333
rect 650164 338328 651715 338330
rect 650164 338272 651654 338328
rect 651710 338272 651715 338328
rect 650164 338270 651715 338272
rect 651649 338267 651715 338270
rect 40677 338192 40786 338197
rect 40677 338136 40682 338192
rect 40738 338136 40786 338192
rect 40677 338134 40786 338136
rect 40677 338131 40743 338134
rect 43069 338058 43135 338061
rect 41492 338056 43135 338058
rect 41492 338000 43074 338056
rect 43130 338000 43135 338056
rect 41492 337998 43135 338000
rect 43069 337995 43135 337998
rect 675334 337860 675340 337924
rect 675404 337922 675410 337924
rect 675477 337922 675543 337925
rect 675404 337920 675543 337922
rect 675404 337864 675482 337920
rect 675538 337864 675543 337920
rect 675404 337862 675543 337864
rect 675404 337860 675410 337862
rect 675477 337859 675543 337862
rect 40910 337380 40970 337620
rect 40902 337316 40908 337380
rect 40972 337316 40978 337380
rect 62113 337242 62179 337245
rect 62113 337240 64492 337242
rect 41462 336970 41522 337212
rect 62113 337184 62118 337240
rect 62174 337184 64492 337240
rect 62113 337182 64492 337184
rect 62113 337179 62179 337182
rect 41638 336970 41644 336972
rect 41462 336910 41644 336970
rect 41638 336908 41644 336910
rect 41708 336908 41714 336972
rect 44449 336834 44515 336837
rect 41492 336832 44515 336834
rect 41492 336776 44454 336832
rect 44510 336776 44515 336832
rect 41492 336774 44515 336776
rect 44449 336771 44515 336774
rect 42977 336426 43043 336429
rect 41492 336424 43043 336426
rect 41492 336368 42982 336424
rect 43038 336368 43043 336424
rect 41492 336366 43043 336368
rect 42977 336363 43043 336366
rect 41278 335748 41338 335988
rect 675753 335882 675819 335885
rect 676990 335882 676996 335884
rect 675753 335880 676996 335882
rect 675753 335824 675758 335880
rect 675814 335824 676996 335880
rect 675753 335822 676996 335824
rect 675753 335819 675819 335822
rect 676990 335820 676996 335822
rect 677060 335820 677066 335884
rect 41270 335684 41276 335748
rect 41340 335684 41346 335748
rect 41094 335340 41154 335580
rect 41086 335276 41092 335340
rect 41156 335276 41162 335340
rect 674833 335338 674899 335341
rect 676806 335338 676812 335340
rect 674833 335336 676812 335338
rect 674833 335280 674838 335336
rect 674894 335280 676812 335336
rect 674833 335278 676812 335280
rect 674833 335275 674899 335278
rect 676806 335276 676812 335278
rect 676876 335276 676882 335340
rect 44541 335202 44607 335205
rect 41492 335200 44607 335202
rect 41492 335144 44546 335200
rect 44602 335144 44607 335200
rect 41492 335142 44607 335144
rect 44541 335139 44607 335142
rect 42885 334794 42951 334797
rect 41492 334792 42951 334794
rect 41492 334736 42890 334792
rect 42946 334736 42951 334792
rect 41492 334734 42951 334736
rect 42885 334731 42951 334734
rect 30422 334117 30482 334356
rect 30373 334112 30482 334117
rect 30373 334056 30378 334112
rect 30434 334056 30482 334112
rect 30373 334054 30482 334056
rect 40861 334114 40927 334117
rect 41822 334114 41828 334116
rect 40861 334112 41828 334114
rect 40861 334056 40866 334112
rect 40922 334056 41828 334112
rect 40861 334054 41828 334056
rect 30373 334051 30439 334054
rect 40861 334051 40927 334054
rect 41822 334052 41828 334054
rect 41892 334052 41898 334116
rect 30422 333540 30482 333948
rect 675753 333570 675819 333573
rect 676070 333570 676076 333572
rect 675753 333568 676076 333570
rect 675753 333512 675758 333568
rect 675814 333512 676076 333568
rect 675753 333510 676076 333512
rect 675753 333507 675819 333510
rect 676070 333508 676076 333510
rect 676140 333508 676146 333572
rect 30373 333298 30439 333301
rect 30373 333296 30482 333298
rect 30373 333240 30378 333296
rect 30434 333240 30482 333296
rect 30373 333235 30482 333240
rect 30422 333132 30482 333235
rect 676622 332618 676628 332620
rect 675710 332558 676628 332618
rect 675710 332213 675770 332558
rect 676622 332556 676628 332558
rect 676692 332556 676698 332620
rect 675710 332208 675819 332213
rect 675710 332152 675758 332208
rect 675814 332152 675819 332208
rect 675710 332150 675819 332152
rect 675753 332147 675819 332150
rect 40677 328402 40743 328405
rect 42006 328402 42012 328404
rect 40677 328400 42012 328402
rect 40677 328344 40682 328400
rect 40738 328344 42012 328400
rect 40677 328342 42012 328344
rect 40677 328339 40743 328342
rect 42006 328340 42012 328342
rect 42076 328340 42082 328404
rect 675109 325682 675175 325685
rect 676438 325682 676444 325684
rect 675109 325680 676444 325682
rect 675109 325624 675114 325680
rect 675170 325624 676444 325680
rect 675109 325622 676444 325624
rect 675109 325619 675175 325622
rect 676438 325620 676444 325622
rect 676508 325620 676514 325684
rect 675753 325546 675819 325549
rect 676254 325546 676260 325548
rect 675753 325544 676260 325546
rect 675753 325488 675758 325544
rect 675814 325488 676260 325544
rect 675753 325486 676260 325488
rect 675753 325483 675819 325486
rect 676254 325484 676260 325486
rect 676324 325484 676330 325548
rect 651557 325002 651623 325005
rect 650164 325000 651623 325002
rect 650164 324944 651562 325000
rect 651618 324944 651623 325000
rect 650164 324942 651623 324944
rect 651557 324939 651623 324942
rect 41781 324868 41847 324869
rect 41781 324864 41828 324868
rect 41892 324866 41898 324868
rect 41781 324808 41786 324864
rect 41781 324804 41828 324808
rect 41892 324806 41938 324866
rect 41892 324804 41898 324806
rect 41781 324803 41847 324804
rect 62113 324186 62179 324189
rect 62113 324184 64492 324186
rect 62113 324128 62118 324184
rect 62174 324128 64492 324184
rect 62113 324126 64492 324128
rect 62113 324123 62179 324126
rect 41270 321132 41276 321196
rect 41340 321194 41346 321196
rect 41781 321194 41847 321197
rect 41340 321192 41847 321194
rect 41340 321136 41786 321192
rect 41842 321136 41847 321192
rect 41340 321134 41847 321136
rect 41340 321132 41346 321134
rect 41781 321131 41847 321134
rect 41965 319972 42031 319973
rect 41965 319968 42012 319972
rect 42076 319970 42082 319972
rect 41965 319912 41970 319968
rect 41965 319908 42012 319912
rect 42076 319910 42122 319970
rect 42076 319908 42082 319910
rect 41965 319907 42031 319908
rect 41086 317324 41092 317388
rect 41156 317386 41162 317388
rect 41781 317386 41847 317389
rect 41156 317384 41847 317386
rect 41156 317328 41786 317384
rect 41842 317328 41847 317384
rect 41156 317326 41847 317328
rect 41156 317324 41162 317326
rect 41781 317323 41847 317326
rect 41638 315828 41644 315892
rect 41708 315890 41714 315892
rect 41781 315890 41847 315893
rect 41708 315888 41847 315890
rect 41708 315832 41786 315888
rect 41842 315832 41847 315888
rect 41708 315830 41847 315832
rect 41708 315828 41714 315830
rect 41781 315827 41847 315830
rect 41454 315420 41460 315484
rect 41524 315482 41530 315484
rect 41781 315482 41847 315485
rect 41524 315480 41847 315482
rect 41524 315424 41786 315480
rect 41842 315424 41847 315480
rect 41524 315422 41847 315424
rect 41524 315420 41530 315422
rect 41781 315419 41847 315422
rect 40718 313788 40724 313852
rect 40788 313850 40794 313852
rect 41873 313850 41939 313853
rect 40788 313848 41939 313850
rect 40788 313792 41878 313848
rect 41934 313792 41939 313848
rect 40788 313790 41939 313792
rect 40788 313788 40794 313790
rect 41873 313787 41939 313790
rect 676262 313581 676322 313684
rect 676213 313576 676322 313581
rect 676213 313520 676218 313576
rect 676274 313520 676322 313576
rect 676213 313518 676322 313520
rect 676213 313515 676279 313518
rect 676029 313306 676095 313309
rect 676029 313304 676292 313306
rect 676029 313248 676034 313304
rect 676090 313248 676292 313304
rect 676029 313246 676292 313248
rect 676029 313243 676095 313246
rect 40902 313108 40908 313172
rect 40972 313170 40978 313172
rect 41781 313170 41847 313173
rect 40972 313168 41847 313170
rect 40972 313112 41786 313168
rect 41842 313112 41847 313168
rect 40972 313110 41847 313112
rect 40972 313108 40978 313110
rect 41781 313107 41847 313110
rect 676262 312765 676322 312868
rect 676213 312760 676322 312765
rect 676213 312704 676218 312760
rect 676274 312704 676322 312760
rect 676213 312702 676322 312704
rect 676213 312699 676279 312702
rect 676029 312490 676095 312493
rect 676029 312488 676292 312490
rect 676029 312432 676034 312488
rect 676090 312432 676292 312488
rect 676029 312430 676292 312432
rect 676029 312427 676095 312430
rect 40534 312292 40540 312356
rect 40604 312354 40610 312356
rect 41781 312354 41847 312357
rect 40604 312352 41847 312354
rect 40604 312296 41786 312352
rect 41842 312296 41847 312352
rect 40604 312294 41847 312296
rect 40604 312292 40610 312294
rect 41781 312291 41847 312294
rect 676262 311949 676322 312052
rect 676213 311944 676322 311949
rect 676213 311888 676218 311944
rect 676274 311888 676322 311944
rect 676213 311886 676322 311888
rect 676213 311883 676279 311886
rect 652385 311810 652451 311813
rect 650164 311808 652451 311810
rect 650164 311752 652390 311808
rect 652446 311752 652451 311808
rect 650164 311750 652451 311752
rect 652385 311747 652451 311750
rect 676029 311674 676095 311677
rect 676029 311672 676292 311674
rect 676029 311616 676034 311672
rect 676090 311616 676292 311672
rect 676029 311614 676292 311616
rect 676029 311611 676095 311614
rect 676262 311133 676322 311236
rect 62113 311130 62179 311133
rect 62113 311128 64492 311130
rect 62113 311072 62118 311128
rect 62174 311072 64492 311128
rect 62113 311070 64492 311072
rect 676213 311128 676322 311133
rect 676213 311072 676218 311128
rect 676274 311072 676322 311128
rect 676213 311070 676322 311072
rect 62113 311067 62179 311070
rect 676213 311067 676279 311070
rect 676262 310725 676322 310828
rect 676213 310720 676322 310725
rect 676213 310664 676218 310720
rect 676274 310664 676322 310720
rect 676213 310662 676322 310664
rect 676213 310659 676279 310662
rect 676262 310317 676322 310420
rect 676262 310312 676371 310317
rect 676262 310256 676310 310312
rect 676366 310256 676371 310312
rect 676262 310254 676371 310256
rect 676305 310251 676371 310254
rect 676121 309906 676187 309909
rect 676262 309906 676322 310012
rect 676121 309904 676322 309906
rect 676121 309848 676126 309904
rect 676182 309848 676322 309904
rect 676121 309846 676322 309848
rect 676121 309843 676187 309846
rect 676262 309501 676322 309604
rect 676213 309496 676322 309501
rect 676213 309440 676218 309496
rect 676274 309440 676322 309496
rect 676213 309438 676322 309440
rect 676213 309435 676279 309438
rect 681046 309093 681106 309196
rect 680997 309088 681106 309093
rect 680997 309032 681002 309088
rect 681058 309032 681106 309088
rect 680997 309030 681106 309032
rect 680997 309027 681063 309030
rect 676446 308684 676506 308788
rect 676438 308620 676444 308684
rect 676508 308620 676514 308684
rect 679758 308277 679818 308380
rect 679709 308272 679818 308277
rect 679709 308216 679714 308272
rect 679770 308216 679818 308272
rect 679709 308214 679818 308216
rect 679709 308211 679775 308214
rect 679574 307869 679634 307972
rect 679574 307864 679683 307869
rect 679574 307808 679622 307864
rect 679678 307808 679683 307864
rect 679574 307806 679683 307808
rect 679617 307803 679683 307806
rect 6022 307753 63922 307782
rect 6022 306609 6150 307753
rect 6854 307749 63922 307753
rect 6854 306645 54235 307749
rect 55339 307729 63922 307749
rect 55339 306645 63339 307729
rect 6854 306625 63339 306645
rect 63883 306625 63922 307729
rect 676070 307396 676076 307460
rect 676140 307458 676146 307460
rect 676262 307458 676322 307564
rect 676140 307398 676322 307458
rect 676140 307396 676146 307398
rect 676262 307052 676322 307156
rect 676254 306988 676260 307052
rect 676324 306988 676330 307052
rect 6854 306609 63922 306625
rect 6022 306582 63922 306609
rect 676814 306645 676874 306748
rect 676814 306640 676923 306645
rect 676814 306584 676862 306640
rect 676918 306584 676923 306640
rect 676814 306582 676923 306584
rect 676857 306579 676923 306582
rect 676262 306237 676322 306340
rect 676262 306232 676371 306237
rect 7236 306157 62944 306182
rect 676262 306176 676310 306232
rect 676366 306176 676371 306232
rect 676262 306174 676371 306176
rect 676305 306171 676371 306174
rect 7236 305013 7348 306157
rect 8052 306131 62944 306157
rect 8052 305027 52641 306131
rect 53745 306121 62944 306131
rect 53745 305027 62371 306121
rect 8052 305017 62371 305027
rect 62915 305017 62944 306121
rect 676446 305829 676506 305932
rect 676397 305824 676506 305829
rect 676397 305768 676402 305824
rect 676458 305768 676506 305824
rect 676397 305766 676506 305768
rect 676397 305763 676463 305766
rect 677550 305421 677610 305524
rect 677550 305416 677659 305421
rect 677550 305360 677598 305416
rect 677654 305360 677659 305416
rect 677550 305358 677659 305360
rect 677593 305355 677659 305358
rect 8052 305013 62944 305017
rect 7236 304982 62944 305013
rect 676630 305012 676690 305116
rect 676622 304948 676628 305012
rect 676692 304948 676698 305012
rect 676262 304605 676322 304708
rect 676213 304600 676322 304605
rect 676213 304544 676218 304600
rect 676274 304544 676322 304600
rect 676213 304542 676322 304544
rect 676213 304539 676279 304542
rect 676121 304194 676187 304197
rect 676262 304194 676322 304300
rect 676121 304192 676322 304194
rect 676121 304136 676126 304192
rect 676182 304136 676322 304192
rect 676121 304134 676322 304136
rect 676121 304131 676187 304134
rect 676262 303789 676322 303892
rect 676213 303784 676322 303789
rect 676213 303728 676218 303784
rect 676274 303728 676322 303784
rect 676213 303726 676322 303728
rect 676213 303723 676279 303726
rect 683070 303381 683130 303484
rect 683070 303376 683179 303381
rect 683070 303320 683118 303376
rect 683174 303320 683179 303376
rect 683070 303318 683179 303320
rect 683113 303315 683179 303318
rect 685830 302668 685890 303076
rect 683113 302562 683179 302565
rect 683070 302560 683179 302562
rect 683070 302504 683118 302560
rect 683174 302504 683179 302560
rect 683070 302499 683179 302504
rect 683070 302260 683130 302499
rect 42057 301338 42123 301341
rect 41492 301336 42123 301338
rect 41492 301280 42062 301336
rect 42118 301280 42123 301336
rect 41492 301278 42123 301280
rect 42057 301275 42123 301278
rect 41965 300930 42031 300933
rect 41492 300928 42031 300930
rect 41492 300872 41970 300928
rect 42026 300872 42031 300928
rect 41492 300870 42031 300872
rect 41965 300867 42031 300870
rect 43621 300522 43687 300525
rect 41492 300520 43687 300522
rect 41492 300464 43626 300520
rect 43682 300464 43687 300520
rect 41492 300462 43687 300464
rect 43621 300459 43687 300462
rect 44265 300114 44331 300117
rect 41492 300112 44331 300114
rect 41492 300056 44270 300112
rect 44326 300056 44331 300112
rect 41492 300054 44331 300056
rect 44265 300051 44331 300054
rect 44725 299706 44791 299709
rect 41492 299704 44791 299706
rect 41492 299648 44730 299704
rect 44786 299648 44791 299704
rect 41492 299646 44791 299648
rect 44725 299643 44791 299646
rect 675886 299372 675892 299436
rect 675956 299434 675962 299436
rect 680997 299434 681063 299437
rect 675956 299432 681063 299434
rect 675956 299376 681002 299432
rect 681058 299376 681063 299432
rect 675956 299374 681063 299376
rect 675956 299372 675962 299374
rect 680997 299371 681063 299374
rect 44173 299298 44239 299301
rect 41492 299296 44239 299298
rect 41492 299240 44178 299296
rect 44234 299240 44239 299296
rect 41492 299238 44239 299240
rect 44173 299235 44239 299238
rect 43069 298890 43135 298893
rect 41492 298888 43135 298890
rect 41492 298832 43074 298888
rect 43130 298832 43135 298888
rect 41492 298830 43135 298832
rect 43069 298827 43135 298830
rect 44357 298482 44423 298485
rect 652017 298482 652083 298485
rect 41492 298480 44423 298482
rect 41492 298424 44362 298480
rect 44418 298424 44423 298480
rect 41492 298422 44423 298424
rect 650164 298480 652083 298482
rect 650164 298424 652022 298480
rect 652078 298424 652083 298480
rect 650164 298422 652083 298424
rect 44357 298419 44423 298422
rect 652017 298419 652083 298422
rect 62113 298210 62179 298213
rect 62113 298208 64492 298210
rect 62113 298152 62118 298208
rect 62174 298152 64492 298208
rect 62113 298150 64492 298152
rect 62113 298147 62179 298150
rect 44265 298074 44331 298077
rect 41492 298072 44331 298074
rect 41492 298016 44270 298072
rect 44326 298016 44331 298072
rect 41492 298014 44331 298016
rect 44265 298011 44331 298014
rect 675702 297740 675708 297804
rect 675772 297802 675778 297804
rect 679617 297802 679683 297805
rect 675772 297800 679683 297802
rect 675772 297744 679622 297800
rect 679678 297744 679683 297800
rect 675772 297742 679683 297744
rect 675772 297740 675778 297742
rect 679617 297739 679683 297742
rect 42793 297666 42859 297669
rect 41492 297664 42859 297666
rect 41492 297608 42798 297664
rect 42854 297608 42859 297664
rect 41492 297606 42859 297608
rect 42793 297603 42859 297606
rect 675334 297468 675340 297532
rect 675404 297530 675410 297532
rect 677593 297530 677659 297533
rect 675404 297528 677659 297530
rect 675404 297472 677598 297528
rect 677654 297472 677659 297528
rect 675404 297470 677659 297472
rect 675404 297468 675410 297470
rect 677593 297467 677659 297470
rect 675518 297332 675524 297396
rect 675588 297394 675594 297396
rect 676305 297394 676371 297397
rect 675588 297392 676371 297394
rect 675588 297336 676310 297392
rect 676366 297336 676371 297392
rect 675588 297334 676371 297336
rect 675588 297332 675594 297334
rect 676305 297331 676371 297334
rect 44633 297258 44699 297261
rect 41492 297256 44699 297258
rect 41492 297200 44638 297256
rect 44694 297200 44699 297256
rect 41492 297198 44699 297200
rect 44633 297195 44699 297198
rect 42374 296850 42380 296852
rect 41492 296790 42380 296850
rect 42374 296788 42380 296790
rect 42444 296788 42450 296852
rect 33777 296442 33843 296445
rect 33764 296440 33843 296442
rect 33764 296384 33782 296440
rect 33838 296384 33843 296440
rect 33764 296382 33843 296384
rect 33777 296379 33843 296382
rect 41822 296034 41828 296036
rect 41492 295974 41828 296034
rect 41822 295972 41828 295974
rect 41892 295972 41898 296036
rect 42190 295626 42196 295628
rect 41492 295566 42196 295626
rect 42190 295564 42196 295566
rect 42260 295564 42266 295628
rect 42006 295218 42012 295220
rect 41492 295158 42012 295218
rect 42006 295156 42012 295158
rect 42076 295156 42082 295220
rect 42425 294810 42491 294813
rect 41492 294808 42491 294810
rect 41492 294752 42430 294808
rect 42486 294752 42491 294808
rect 41492 294750 42491 294752
rect 42425 294747 42491 294750
rect 675753 294810 675819 294813
rect 675886 294810 675892 294812
rect 675753 294808 675892 294810
rect 675753 294752 675758 294808
rect 675814 294752 675892 294808
rect 675753 294750 675892 294752
rect 675753 294747 675819 294750
rect 675886 294748 675892 294750
rect 675956 294748 675962 294812
rect 41822 294402 41828 294404
rect 41492 294342 41828 294402
rect 41822 294340 41828 294342
rect 41892 294340 41898 294404
rect 41822 293994 41828 293996
rect 41492 293934 41828 293994
rect 41822 293932 41828 293934
rect 41892 293932 41898 293996
rect 44449 293586 44515 293589
rect 41492 293584 44515 293586
rect 41492 293528 44454 293584
rect 44510 293528 44515 293584
rect 41492 293526 44515 293528
rect 44449 293523 44515 293526
rect 42977 293178 43043 293181
rect 41492 293176 43043 293178
rect 41492 293120 42982 293176
rect 43038 293120 43043 293176
rect 41492 293118 43043 293120
rect 42977 293115 43043 293118
rect 41462 292592 41522 292740
rect 675661 292636 675727 292637
rect 675661 292634 675708 292636
rect 675616 292632 675708 292634
rect 41454 292528 41460 292592
rect 41524 292528 41530 292592
rect 675616 292576 675666 292632
rect 675616 292574 675708 292576
rect 675661 292572 675708 292574
rect 675772 292572 675778 292636
rect 675661 292571 675727 292572
rect 44541 292362 44607 292365
rect 41492 292360 44607 292362
rect 41492 292304 44546 292360
rect 44602 292304 44607 292360
rect 41492 292302 44607 292304
rect 44541 292299 44607 292302
rect 675477 292092 675543 292093
rect 675477 292088 675524 292092
rect 675588 292090 675594 292092
rect 675477 292032 675482 292088
rect 675477 292028 675524 292032
rect 675588 292030 675634 292090
rect 675588 292028 675594 292030
rect 675477 292027 675543 292028
rect 42885 291954 42951 291957
rect 41492 291952 42951 291954
rect 41492 291896 42890 291952
rect 42946 291896 42951 291952
rect 41492 291894 42951 291896
rect 42885 291891 42951 291894
rect 44173 291546 44239 291549
rect 41492 291544 44239 291546
rect 41492 291488 44178 291544
rect 44234 291488 44239 291544
rect 41492 291486 44239 291488
rect 44173 291483 44239 291486
rect 43989 291138 44055 291141
rect 41492 291136 44055 291138
rect 41492 291080 43994 291136
rect 44050 291080 44055 291136
rect 41492 291078 44055 291080
rect 43989 291075 44055 291078
rect 43805 290730 43871 290733
rect 41492 290728 43871 290730
rect 41492 290672 43810 290728
rect 43866 290672 43871 290728
rect 41492 290670 43871 290672
rect 43805 290667 43871 290670
rect 45001 289914 45067 289917
rect 41492 289912 45067 289914
rect 41492 289856 45006 289912
rect 45062 289856 45067 289912
rect 41492 289854 45067 289856
rect 45001 289851 45067 289854
rect 675753 288418 675819 288421
rect 676070 288418 676076 288420
rect 675753 288416 676076 288418
rect 675753 288360 675758 288416
rect 675814 288360 676076 288416
rect 675753 288358 676076 288360
rect 675753 288355 675819 288358
rect 676070 288356 676076 288358
rect 676140 288356 676146 288420
rect 41822 288084 41828 288148
rect 41892 288084 41898 288148
rect 41830 287876 41890 288084
rect 41822 287812 41828 287876
rect 41892 287812 41898 287876
rect 675753 287330 675819 287333
rect 676622 287330 676628 287332
rect 675753 287328 676628 287330
rect 675753 287272 675758 287328
rect 675814 287272 676628 287328
rect 675753 287270 676628 287272
rect 675753 287267 675819 287270
rect 676622 287268 676628 287270
rect 676692 287268 676698 287332
rect 675334 285500 675340 285564
rect 675404 285562 675410 285564
rect 675477 285562 675543 285565
rect 675404 285560 675543 285562
rect 675404 285504 675482 285560
rect 675538 285504 675543 285560
rect 675404 285502 675543 285504
rect 675404 285500 675410 285502
rect 675477 285499 675543 285502
rect 651557 285290 651623 285293
rect 650164 285288 651623 285290
rect 650164 285232 651562 285288
rect 651618 285232 651623 285288
rect 650164 285230 651623 285232
rect 651557 285227 651623 285230
rect 62113 285154 62179 285157
rect 62113 285152 64492 285154
rect 62113 285096 62118 285152
rect 62174 285096 64492 285152
rect 62113 285094 64492 285096
rect 62113 285091 62179 285094
rect 41638 284956 41644 285020
rect 41708 285018 41714 285020
rect 42006 285018 42012 285020
rect 41708 284958 42012 285018
rect 41708 284956 41714 284958
rect 42006 284956 42012 284958
rect 42076 284956 42082 285020
rect 33777 284882 33843 284885
rect 41454 284882 41460 284884
rect 33777 284880 41460 284882
rect 33777 284824 33782 284880
rect 33838 284824 41460 284880
rect 33777 284822 41460 284824
rect 33777 284819 33843 284822
rect 41454 284820 41460 284822
rect 41524 284820 41530 284884
rect 675753 283658 675819 283661
rect 676438 283658 676444 283660
rect 675753 283656 676444 283658
rect 675753 283600 675758 283656
rect 675814 283600 676444 283656
rect 675753 283598 676444 283600
rect 675753 283595 675819 283598
rect 676438 283596 676444 283598
rect 676508 283596 676514 283660
rect 41454 281420 41460 281484
rect 41524 281482 41530 281484
rect 41781 281482 41847 281485
rect 41524 281480 41847 281482
rect 41524 281424 41786 281480
rect 41842 281424 41847 281480
rect 41524 281422 41847 281424
rect 41524 281420 41530 281422
rect 41781 281419 41847 281422
rect 675753 281482 675819 281485
rect 676254 281482 676260 281484
rect 675753 281480 676260 281482
rect 675753 281424 675758 281480
rect 675814 281424 676260 281480
rect 675753 281422 676260 281424
rect 675753 281419 675819 281422
rect 676254 281420 676260 281422
rect 676324 281420 676330 281484
rect 40902 278700 40908 278764
rect 40972 278762 40978 278764
rect 42701 278762 42767 278765
rect 40972 278760 42767 278762
rect 40972 278704 42706 278760
rect 42762 278704 42767 278760
rect 40972 278702 42767 278704
rect 40972 278700 40978 278702
rect 42701 278699 42767 278702
rect 40902 277340 40908 277404
rect 40972 277402 40978 277404
rect 41781 277402 41847 277405
rect 40972 277400 41847 277402
rect 40972 277344 41786 277400
rect 41842 277344 41847 277400
rect 40972 277342 41847 277344
rect 40972 277340 40978 277342
rect 41781 277339 41847 277342
rect 41781 276724 41847 276725
rect 41781 276720 41828 276724
rect 41892 276722 41898 276724
rect 41781 276664 41786 276720
rect 41781 276660 41828 276664
rect 41892 276662 41938 276722
rect 41892 276660 41898 276662
rect 41781 276659 41847 276660
rect 368381 275498 368447 275501
rect 530485 275498 530551 275501
rect 368381 275496 530551 275498
rect 368381 275440 368386 275496
rect 368442 275440 530490 275496
rect 530546 275440 530551 275496
rect 368381 275438 530551 275440
rect 368381 275435 368447 275438
rect 530485 275435 530551 275438
rect 371141 275362 371207 275365
rect 537569 275362 537635 275365
rect 371141 275360 537635 275362
rect 371141 275304 371146 275360
rect 371202 275304 537574 275360
rect 537630 275304 537635 275360
rect 371141 275302 537635 275304
rect 371141 275299 371207 275302
rect 537569 275299 537635 275302
rect 373901 275226 373967 275229
rect 544653 275226 544719 275229
rect 373901 275224 544719 275226
rect 373901 275168 373906 275224
rect 373962 275168 544658 275224
rect 544714 275168 544719 275224
rect 373901 275166 544719 275168
rect 373901 275163 373967 275166
rect 544653 275163 544719 275166
rect 411069 274002 411135 274005
rect 419533 274002 419599 274005
rect 411069 274000 419599 274002
rect 411069 273944 411074 274000
rect 411130 273944 419538 274000
rect 419594 273944 419599 274000
rect 411069 273942 419599 273944
rect 411069 273939 411135 273942
rect 419533 273939 419599 273942
rect 386229 273866 386295 273869
rect 580073 273866 580139 273869
rect 386229 273864 580139 273866
rect 386229 273808 386234 273864
rect 386290 273808 580078 273864
rect 580134 273808 580139 273864
rect 386229 273806 580139 273808
rect 386229 273803 386295 273806
rect 580073 273803 580139 273806
rect 404261 272778 404327 272781
rect 628557 272778 628623 272781
rect 404261 272776 628623 272778
rect 404261 272720 404266 272776
rect 404322 272720 628562 272776
rect 628618 272720 628623 272776
rect 404261 272718 628623 272720
rect 404261 272715 404327 272718
rect 628557 272715 628623 272718
rect 406929 272642 406995 272645
rect 635641 272642 635707 272645
rect 406929 272640 635707 272642
rect 406929 272584 406934 272640
rect 406990 272584 635646 272640
rect 635702 272584 635707 272640
rect 406929 272582 635707 272584
rect 406929 272579 406995 272582
rect 635641 272579 635707 272582
rect 408309 272506 408375 272509
rect 639229 272506 639295 272509
rect 408309 272504 639295 272506
rect 408309 272448 408314 272504
rect 408370 272448 639234 272504
rect 639290 272448 639295 272504
rect 408309 272446 639295 272448
rect 408309 272443 408375 272446
rect 639229 272443 639295 272446
rect 41638 272308 41644 272372
rect 41708 272370 41714 272372
rect 41781 272370 41847 272373
rect 41708 272368 41847 272370
rect 41708 272312 41786 272368
rect 41842 272312 41847 272368
rect 41708 272310 41847 272312
rect 41708 272308 41714 272310
rect 41781 272307 41847 272310
rect 379237 271418 379303 271421
rect 561213 271418 561279 271421
rect 379237 271416 561279 271418
rect 379237 271360 379242 271416
rect 379298 271360 561218 271416
rect 561274 271360 561279 271416
rect 379237 271358 561279 271360
rect 379237 271355 379303 271358
rect 561213 271355 561279 271358
rect 382089 271282 382155 271285
rect 568297 271282 568363 271285
rect 382089 271280 568363 271282
rect 382089 271224 382094 271280
rect 382150 271224 568302 271280
rect 568358 271224 568363 271280
rect 382089 271222 568363 271224
rect 382089 271219 382155 271222
rect 568297 271219 568363 271222
rect 383285 271146 383351 271149
rect 571793 271146 571859 271149
rect 383285 271144 571859 271146
rect 383285 271088 383290 271144
rect 383346 271088 571798 271144
rect 571854 271088 571859 271144
rect 383285 271086 571859 271088
rect 383285 271083 383351 271086
rect 571793 271083 571859 271086
rect 41965 270468 42031 270469
rect 41965 270464 42012 270468
rect 42076 270466 42082 270468
rect 41965 270408 41970 270464
rect 41965 270404 42012 270408
rect 42076 270406 42122 270466
rect 42076 270404 42082 270406
rect 41965 270403 42031 270404
rect 350257 270194 350323 270197
rect 484393 270194 484459 270197
rect 350257 270192 484459 270194
rect 350257 270136 350262 270192
rect 350318 270136 484398 270192
rect 484454 270136 484459 270192
rect 350257 270134 484459 270136
rect 350257 270131 350323 270134
rect 484393 270131 484459 270134
rect 383377 270058 383443 270061
rect 572713 270058 572779 270061
rect 383377 270056 572779 270058
rect 383377 270000 383382 270056
rect 383438 270000 572718 270056
rect 572774 270000 572779 270056
rect 383377 269998 572779 270000
rect 383377 269995 383443 269998
rect 572713 269995 572779 269998
rect 388253 269922 388319 269925
rect 585133 269922 585199 269925
rect 388253 269920 585199 269922
rect 388253 269864 388258 269920
rect 388314 269864 585138 269920
rect 585194 269864 585199 269920
rect 388253 269862 585199 269864
rect 388253 269859 388319 269862
rect 585133 269859 585199 269862
rect 40718 269724 40724 269788
rect 40788 269786 40794 269788
rect 41781 269786 41847 269789
rect 40788 269784 41847 269786
rect 40788 269728 41786 269784
rect 41842 269728 41847 269784
rect 40788 269726 41847 269728
rect 40788 269724 40794 269726
rect 41781 269723 41847 269726
rect 401593 269786 401659 269789
rect 618253 269786 618319 269789
rect 401593 269784 618319 269786
rect 401593 269728 401598 269784
rect 401654 269728 618258 269784
rect 618314 269728 618319 269784
rect 401593 269726 618319 269728
rect 401593 269723 401659 269726
rect 618253 269723 618319 269726
rect 40534 269044 40540 269108
rect 40604 269106 40610 269108
rect 41781 269106 41847 269109
rect 40604 269104 41847 269106
rect 40604 269048 41786 269104
rect 41842 269048 41847 269104
rect 40604 269046 41847 269048
rect 40604 269044 40610 269046
rect 41781 269043 41847 269046
rect 350349 268970 350415 268973
rect 433333 268970 433399 268973
rect 350349 268968 433399 268970
rect 350349 268912 350354 268968
rect 350410 268912 433338 268968
rect 433394 268912 433399 268968
rect 350349 268910 433399 268912
rect 350349 268907 350415 268910
rect 433333 268907 433399 268910
rect 368197 268834 368263 268837
rect 532693 268834 532759 268837
rect 368197 268832 532759 268834
rect 368197 268776 368202 268832
rect 368258 268776 532698 268832
rect 532754 268776 532759 268832
rect 368197 268774 532759 268776
rect 368197 268771 368263 268774
rect 532693 268771 532759 268774
rect 398465 268698 398531 268701
rect 612733 268698 612799 268701
rect 398465 268696 612799 268698
rect 398465 268640 398470 268696
rect 398526 268640 612738 268696
rect 612794 268640 612799 268696
rect 398465 268638 612799 268640
rect 398465 268635 398531 268638
rect 612733 268635 612799 268638
rect 676262 268565 676322 268668
rect 402513 268562 402579 268565
rect 623773 268562 623839 268565
rect 402513 268560 623839 268562
rect 402513 268504 402518 268560
rect 402574 268504 623778 268560
rect 623834 268504 623839 268560
rect 402513 268502 623839 268504
rect 402513 268499 402579 268502
rect 623773 268499 623839 268502
rect 676213 268560 676322 268565
rect 676213 268504 676218 268560
rect 676274 268504 676322 268560
rect 676213 268502 676322 268504
rect 676213 268499 676279 268502
rect 405181 268426 405247 268429
rect 630673 268426 630739 268429
rect 405181 268424 630739 268426
rect 405181 268368 405186 268424
rect 405242 268368 630678 268424
rect 630734 268368 630739 268424
rect 405181 268366 630739 268368
rect 405181 268363 405247 268366
rect 630673 268363 630739 268366
rect 676121 268154 676187 268157
rect 676262 268154 676322 268260
rect 676121 268152 676322 268154
rect 676121 268096 676126 268152
rect 676182 268096 676322 268152
rect 676121 268094 676322 268096
rect 676121 268091 676187 268094
rect 676262 267749 676322 267852
rect 397637 267746 397703 267749
rect 411897 267746 411963 267749
rect 397637 267744 411963 267746
rect 397637 267688 397642 267744
rect 397698 267688 411902 267744
rect 411958 267688 411963 267744
rect 397637 267686 411963 267688
rect 397637 267683 397703 267686
rect 411897 267683 411963 267686
rect 676213 267744 676322 267749
rect 676213 267688 676218 267744
rect 676274 267688 676322 267744
rect 676213 267686 676322 267688
rect 676213 267683 676279 267686
rect 403433 267610 403499 267613
rect 469305 267610 469371 267613
rect 403433 267608 469371 267610
rect 403433 267552 403438 267608
rect 403494 267552 469310 267608
rect 469366 267552 469371 267608
rect 403433 267550 469371 267552
rect 403433 267547 403499 267550
rect 469305 267547 469371 267550
rect 357985 267474 358051 267477
rect 493317 267474 493383 267477
rect 357985 267472 493383 267474
rect 357985 267416 357990 267472
rect 358046 267416 493322 267472
rect 493378 267416 493383 267472
rect 357985 267414 493383 267416
rect 357985 267411 358051 267414
rect 493317 267411 493383 267414
rect 674741 267474 674807 267477
rect 674741 267472 676292 267474
rect 674741 267416 674746 267472
rect 674802 267416 676292 267472
rect 674741 267414 676292 267416
rect 674741 267411 674807 267414
rect 365989 267338 366055 267341
rect 518985 267338 519051 267341
rect 365989 267336 519051 267338
rect 365989 267280 365994 267336
rect 366050 267280 518990 267336
rect 519046 267280 519051 267336
rect 365989 267278 519051 267280
rect 365989 267275 366055 267278
rect 518985 267275 519051 267278
rect 411437 267202 411503 267205
rect 647233 267202 647299 267205
rect 411437 267200 647299 267202
rect 411437 267144 411442 267200
rect 411498 267144 647238 267200
rect 647294 267144 647299 267200
rect 411437 267142 647299 267144
rect 411437 267139 411503 267142
rect 647233 267139 647299 267142
rect 380709 267066 380775 267069
rect 388437 267066 388503 267069
rect 380709 267064 388503 267066
rect 380709 267008 380714 267064
rect 380770 267008 388442 267064
rect 388498 267008 388503 267064
rect 380709 267006 388503 267008
rect 380709 267003 380775 267006
rect 388437 267003 388503 267006
rect 411897 267066 411963 267069
rect 648613 267066 648679 267069
rect 411897 267064 648679 267066
rect 411897 267008 411902 267064
rect 411958 267008 648618 267064
rect 648674 267008 648679 267064
rect 411897 267006 648679 267008
rect 411897 267003 411963 267006
rect 648613 267003 648679 267006
rect 676262 266933 676322 267036
rect 676213 266928 676322 266933
rect 676213 266872 676218 266928
rect 676274 266872 676322 266928
rect 676213 266870 676322 266872
rect 676213 266867 676279 266870
rect 676029 266658 676095 266661
rect 676029 266656 676292 266658
rect 676029 266600 676034 266656
rect 676090 266600 676292 266656
rect 676029 266598 676292 266600
rect 676029 266595 676095 266598
rect 391381 266386 391447 266389
rect 392577 266386 392643 266389
rect 391381 266384 392643 266386
rect 391381 266328 391386 266384
rect 391442 266328 392582 266384
rect 392638 266328 392643 266384
rect 391381 266326 392643 266328
rect 391381 266323 391447 266326
rect 392577 266323 392643 266326
rect 407389 266386 407455 266389
rect 410425 266386 410491 266389
rect 407389 266384 410491 266386
rect 407389 266328 407394 266384
rect 407450 266328 410430 266384
rect 410486 266328 410491 266384
rect 407389 266326 410491 266328
rect 407389 266323 407455 266326
rect 410425 266323 410491 266326
rect 676262 266117 676322 266220
rect 676213 266112 676322 266117
rect 676213 266056 676218 266112
rect 676274 266056 676322 266112
rect 676213 266054 676322 266056
rect 676213 266051 676279 266054
rect 389633 265978 389699 265981
rect 589273 265978 589339 265981
rect 389633 265976 589339 265978
rect 389633 265920 389638 265976
rect 389694 265920 589278 265976
rect 589334 265920 589339 265976
rect 389633 265918 589339 265920
rect 389633 265915 389699 265918
rect 589273 265915 589339 265918
rect 392301 265842 392367 265845
rect 596173 265842 596239 265845
rect 392301 265840 596239 265842
rect 392301 265784 392306 265840
rect 392362 265784 596178 265840
rect 596234 265784 596239 265840
rect 392301 265782 596239 265784
rect 392301 265779 392367 265782
rect 596173 265779 596239 265782
rect 676262 265709 676322 265812
rect 406561 265706 406627 265709
rect 633433 265706 633499 265709
rect 406561 265704 633499 265706
rect 406561 265648 406566 265704
rect 406622 265648 633438 265704
rect 633494 265648 633499 265704
rect 406561 265646 633499 265648
rect 406561 265643 406627 265646
rect 633433 265643 633499 265646
rect 676213 265704 676322 265709
rect 676213 265648 676218 265704
rect 676274 265648 676322 265704
rect 676213 265646 676322 265648
rect 676213 265643 676279 265646
rect 409229 265570 409295 265573
rect 640517 265570 640583 265573
rect 409229 265568 640583 265570
rect 409229 265512 409234 265568
rect 409290 265512 640522 265568
rect 640578 265512 640583 265568
rect 409229 265510 640583 265512
rect 409229 265507 409295 265510
rect 640517 265507 640583 265510
rect 676121 265298 676187 265301
rect 676262 265298 676322 265404
rect 676121 265296 676322 265298
rect 676121 265240 676126 265296
rect 676182 265240 676322 265296
rect 676121 265238 676322 265240
rect 676121 265235 676187 265238
rect 676029 265026 676095 265029
rect 676029 265024 676292 265026
rect 676029 264968 676034 265024
rect 676090 264968 676292 265024
rect 676029 264966 676292 264968
rect 676029 264963 676095 264966
rect 6022 264553 55460 264582
rect 6022 263409 6150 264553
rect 6854 264549 55460 264553
rect 6854 263445 54235 264549
rect 55339 263445 55460 264549
rect 676262 264485 676322 264588
rect 676213 264480 676322 264485
rect 676213 264424 676218 264480
rect 676274 264424 676322 264480
rect 676213 264422 676322 264424
rect 676213 264419 676279 264422
rect 396993 264210 397059 264213
rect 401225 264210 401291 264213
rect 396993 264208 401291 264210
rect 396993 264152 396998 264208
rect 397054 264152 401230 264208
rect 401286 264152 401291 264208
rect 396993 264150 401291 264152
rect 396993 264147 397059 264150
rect 401225 264147 401291 264150
rect 675886 264148 675892 264212
rect 675956 264210 675962 264212
rect 675956 264150 676292 264210
rect 675956 264148 675962 264150
rect 676998 263634 677058 263772
rect 676990 263570 676996 263634
rect 677060 263570 677066 263634
rect 6854 263409 55460 263445
rect 6022 263382 55460 263409
rect 678286 263261 678346 263364
rect 678237 263256 678346 263261
rect 678237 263200 678242 263256
rect 678298 263200 678346 263256
rect 678237 263198 678346 263200
rect 678237 263195 678303 263198
rect 7236 262957 53816 262982
rect 7236 261813 7348 262957
rect 8052 262931 53816 262957
rect 8052 261827 52641 262931
rect 53745 261827 53816 262931
rect 675702 262924 675708 262988
rect 675772 262986 675778 262988
rect 675772 262926 676292 262986
rect 675772 262924 675778 262926
rect 678286 262445 678346 262548
rect 678286 262440 678395 262445
rect 678286 262384 678334 262440
rect 678390 262384 678395 262440
rect 678286 262382 678395 262384
rect 678329 262379 678395 262382
rect 415301 262306 415367 262309
rect 412436 262304 415367 262306
rect 412436 262248 415306 262304
rect 415362 262248 415367 262304
rect 412436 262246 415367 262248
rect 415301 262243 415367 262246
rect 677182 262036 677242 262140
rect 677174 261972 677180 262036
rect 677244 261972 677250 262036
rect 8052 261813 53816 261827
rect 7236 261782 53816 261813
rect 677366 261628 677426 261732
rect 677358 261564 677364 261628
rect 677428 261564 677434 261628
rect 676814 261221 676874 261324
rect 676814 261216 676923 261221
rect 676814 261160 676862 261216
rect 676918 261160 676923 261216
rect 676814 261158 676923 261160
rect 676857 261155 676923 261158
rect 676998 260813 677058 260916
rect 676949 260808 677058 260813
rect 676949 260752 676954 260808
rect 677010 260752 677058 260808
rect 676949 260750 677058 260752
rect 676949 260747 677015 260750
rect 676070 260340 676076 260404
rect 676140 260402 676146 260404
rect 676262 260402 676322 260508
rect 676140 260342 676322 260402
rect 676140 260340 676146 260342
rect 676446 259997 676506 260100
rect 676397 259992 676506 259997
rect 676397 259936 676402 259992
rect 676458 259936 676506 259992
rect 676397 259934 676506 259936
rect 676397 259931 676463 259934
rect 676446 259589 676506 259692
rect 676446 259584 676555 259589
rect 676446 259528 676494 259584
rect 676550 259528 676555 259584
rect 676446 259526 676555 259528
rect 676489 259523 676555 259526
rect 676262 259181 676322 259284
rect 414197 259178 414263 259181
rect 412436 259176 414263 259178
rect 412436 259120 414202 259176
rect 414258 259120 414263 259176
rect 412436 259118 414263 259120
rect 414197 259115 414263 259118
rect 676213 259176 676322 259181
rect 676213 259120 676218 259176
rect 676274 259120 676322 259176
rect 676213 259118 676322 259120
rect 676213 259115 676279 259118
rect 676262 258773 676322 258876
rect 676213 258768 676322 258773
rect 676213 258712 676218 258768
rect 676274 258712 676322 258768
rect 676213 258710 676322 258712
rect 676213 258707 676279 258710
rect 189073 258634 189139 258637
rect 189073 258632 191820 258634
rect 189073 258576 189078 258632
rect 189134 258576 191820 258632
rect 189073 258574 191820 258576
rect 189073 258571 189139 258574
rect 683070 258365 683130 258468
rect 35801 258362 35867 258365
rect 35758 258360 35867 258362
rect 35758 258304 35806 258360
rect 35862 258304 35867 258360
rect 35758 258299 35867 258304
rect 683070 258360 683179 258365
rect 683070 258304 683118 258360
rect 683174 258304 683179 258360
rect 683070 258302 683179 258304
rect 683113 258299 683179 258302
rect 35758 258060 35818 258299
rect 31661 257954 31727 257957
rect 31661 257952 31770 257954
rect 31661 257896 31666 257952
rect 31722 257896 31770 257952
rect 31661 257891 31770 257896
rect 31710 257652 31770 257891
rect 683070 257652 683130 258060
rect 31661 257546 31727 257549
rect 683113 257546 683179 257549
rect 31661 257544 31770 257546
rect 31661 257488 31666 257544
rect 31722 257488 31770 257544
rect 31661 257483 31770 257488
rect 31710 257244 31770 257483
rect 683070 257544 683179 257546
rect 683070 257488 683118 257544
rect 683174 257488 683179 257544
rect 683070 257483 683179 257488
rect 683070 257244 683130 257483
rect 31569 257138 31635 257141
rect 31526 257136 31635 257138
rect 31526 257080 31574 257136
rect 31630 257080 31635 257136
rect 31526 257075 31635 257080
rect 31526 256836 31586 257075
rect 42885 256458 42951 256461
rect 41492 256456 42951 256458
rect 41492 256400 42890 256456
rect 42946 256400 42951 256456
rect 41492 256398 42951 256400
rect 42885 256395 42951 256398
rect 43069 256050 43135 256053
rect 41492 256048 43135 256050
rect 41492 255992 43074 256048
rect 43130 255992 43135 256048
rect 41492 255990 43135 255992
rect 43069 255987 43135 255990
rect 415301 255914 415367 255917
rect 412436 255912 415367 255914
rect 412436 255856 415306 255912
rect 415362 255856 415367 255912
rect 412436 255854 415367 255856
rect 415301 255851 415367 255854
rect 43069 255642 43135 255645
rect 41492 255640 43135 255642
rect 41492 255584 43074 255640
rect 43130 255584 43135 255640
rect 41492 255582 43135 255584
rect 43069 255579 43135 255582
rect 44265 255234 44331 255237
rect 41492 255232 44331 255234
rect 41492 255176 44270 255232
rect 44326 255176 44331 255232
rect 41492 255174 44331 255176
rect 44265 255171 44331 255174
rect 44541 254826 44607 254829
rect 41492 254824 44607 254826
rect 41492 254768 44546 254824
rect 44602 254768 44607 254824
rect 41492 254766 44607 254768
rect 44541 254763 44607 254766
rect 44633 254418 44699 254421
rect 41492 254416 44699 254418
rect 41492 254360 44638 254416
rect 44694 254360 44699 254416
rect 41492 254358 44699 254360
rect 44633 254355 44699 254358
rect 44265 254010 44331 254013
rect 41492 254008 44331 254010
rect 41492 253952 44270 254008
rect 44326 253952 44331 254008
rect 41492 253950 44331 253952
rect 44265 253947 44331 253950
rect 42190 253602 42196 253604
rect 41492 253542 42196 253602
rect 42190 253540 42196 253542
rect 42260 253540 42266 253604
rect 41822 253194 41828 253196
rect 41492 253134 41828 253194
rect 41822 253132 41828 253134
rect 41892 253132 41898 253196
rect 414381 252786 414447 252789
rect 412436 252784 414447 252786
rect 40542 252652 40602 252756
rect 412436 252728 414386 252784
rect 414442 252728 414447 252784
rect 412436 252726 414447 252728
rect 414381 252723 414447 252726
rect 40534 252588 40540 252652
rect 40604 252588 40610 252652
rect 674782 252588 674788 252652
rect 674852 252650 674858 252652
rect 678329 252650 678395 252653
rect 674852 252648 678395 252650
rect 674852 252592 678334 252648
rect 678390 252592 678395 252648
rect 674852 252590 678395 252592
rect 674852 252588 674858 252590
rect 678329 252587 678395 252590
rect 41462 252242 41522 252348
rect 41638 252242 41644 252244
rect 41462 252182 41644 252242
rect 41638 252180 41644 252182
rect 41708 252180 41714 252244
rect 30974 251837 31034 251940
rect 30974 251832 31083 251837
rect 30974 251776 31022 251832
rect 31078 251776 31083 251832
rect 30974 251774 31083 251776
rect 31017 251771 31083 251774
rect 673913 251698 673979 251701
rect 676397 251698 676463 251701
rect 673913 251696 676463 251698
rect 673913 251640 673918 251696
rect 673974 251640 676402 251696
rect 676458 251640 676463 251696
rect 673913 251638 676463 251640
rect 673913 251635 673979 251638
rect 676397 251635 676463 251638
rect 42701 251562 42767 251565
rect 41492 251560 42767 251562
rect 41492 251504 42706 251560
rect 42762 251504 42767 251560
rect 41492 251502 42767 251504
rect 42701 251499 42767 251502
rect 676438 251500 676444 251564
rect 676508 251562 676514 251564
rect 677358 251562 677364 251564
rect 676508 251502 677364 251562
rect 676508 251500 676514 251502
rect 677358 251500 677364 251502
rect 677428 251500 677434 251564
rect 44357 251154 44423 251157
rect 41492 251152 44423 251154
rect 41492 251096 44362 251152
rect 44418 251096 44423 251152
rect 41492 251094 44423 251096
rect 44357 251091 44423 251094
rect 39990 250613 40050 250716
rect 39941 250608 40050 250613
rect 39941 250552 39946 250608
rect 40002 250552 40050 250608
rect 39941 250550 40050 250552
rect 39941 250547 40007 250550
rect 42977 250338 43043 250341
rect 41492 250336 43043 250338
rect 41492 250280 42982 250336
rect 43038 250280 43043 250336
rect 41492 250278 43043 250280
rect 42977 250275 43043 250278
rect 675753 250338 675819 250341
rect 676438 250338 676444 250340
rect 675753 250336 676444 250338
rect 675753 250280 675758 250336
rect 675814 250280 676444 250336
rect 675753 250278 676444 250280
rect 675753 250275 675819 250278
rect 676438 250276 676444 250278
rect 676508 250276 676514 250340
rect 40174 249796 40234 249900
rect 40166 249732 40172 249796
rect 40236 249732 40242 249796
rect 673729 249794 673795 249797
rect 674782 249794 674788 249796
rect 673729 249792 674788 249794
rect 673729 249736 673734 249792
rect 673790 249736 674788 249792
rect 673729 249734 674788 249736
rect 673729 249731 673795 249734
rect 674782 249732 674788 249734
rect 674852 249732 674858 249796
rect 675753 249794 675819 249797
rect 675886 249794 675892 249796
rect 675753 249792 675892 249794
rect 675753 249736 675758 249792
rect 675814 249736 675892 249792
rect 675753 249734 675892 249736
rect 675753 249731 675819 249734
rect 675886 249732 675892 249734
rect 675956 249732 675962 249796
rect 673821 249660 673887 249661
rect 673821 249658 673868 249660
rect 673776 249656 673868 249658
rect 673776 249600 673826 249656
rect 673776 249598 673868 249600
rect 673821 249596 673868 249598
rect 673932 249596 673938 249660
rect 675017 249658 675083 249661
rect 675702 249658 675708 249660
rect 675017 249656 675708 249658
rect 675017 249600 675022 249656
rect 675078 249600 675708 249656
rect 675017 249598 675708 249600
rect 673821 249595 673887 249596
rect 675017 249595 675083 249598
rect 675702 249596 675708 249598
rect 675772 249596 675778 249660
rect 676070 249596 676076 249660
rect 676140 249596 676146 249660
rect 414197 249522 414263 249525
rect 412436 249520 414263 249522
rect 40358 249388 40418 249492
rect 412436 249464 414202 249520
rect 414258 249464 414263 249520
rect 412436 249462 414263 249464
rect 414197 249459 414263 249462
rect 675201 249522 675267 249525
rect 676078 249522 676138 249596
rect 675201 249520 676138 249522
rect 675201 249464 675206 249520
rect 675262 249464 676138 249520
rect 675201 249462 676138 249464
rect 675201 249459 675267 249462
rect 40350 249324 40356 249388
rect 40420 249324 40426 249388
rect 39990 248980 40050 249084
rect 39982 248916 39988 248980
rect 40052 248916 40058 248980
rect 44449 248706 44515 248709
rect 41492 248704 44515 248706
rect 41492 248648 44454 248704
rect 44510 248648 44515 248704
rect 41492 248646 44515 248648
rect 44449 248643 44515 248646
rect 44541 248298 44607 248301
rect 41492 248296 44607 248298
rect 41492 248240 44546 248296
rect 44602 248240 44607 248296
rect 41492 248238 44607 248240
rect 44541 248235 44607 248238
rect 190361 248026 190427 248029
rect 190361 248024 191820 248026
rect 190361 247968 190366 248024
rect 190422 247968 191820 248024
rect 190361 247966 191820 247968
rect 190361 247963 190427 247966
rect 41462 247754 41522 247860
rect 41462 247694 55230 247754
rect 41462 247346 41522 247452
rect 55170 247346 55230 247694
rect 85021 247346 85087 247349
rect 41462 247286 45570 247346
rect 55170 247344 85087 247346
rect 55170 247288 85026 247344
rect 85082 247288 85087 247344
rect 55170 247286 85087 247288
rect 45510 247210 45570 247286
rect 85021 247283 85087 247286
rect 84837 247210 84903 247213
rect 45510 247208 84903 247210
rect 45510 247152 84842 247208
rect 84898 247152 84903 247208
rect 45510 247150 84903 247152
rect 84837 247147 84903 247150
rect 35758 246533 35818 246636
rect 35758 246528 35867 246533
rect 35758 246472 35806 246528
rect 35862 246472 35867 246528
rect 35758 246470 35867 246472
rect 35801 246467 35867 246470
rect 415301 246394 415367 246397
rect 412436 246392 415367 246394
rect 412436 246336 415306 246392
rect 415362 246336 415367 246392
rect 412436 246334 415367 246336
rect 415301 246331 415367 246334
rect 673913 246258 673979 246261
rect 674966 246258 674972 246260
rect 673913 246256 674972 246258
rect 673913 246200 673918 246256
rect 673974 246200 674972 246256
rect 673913 246198 674972 246200
rect 673913 246195 673979 246198
rect 674966 246196 674972 246198
rect 675036 246196 675042 246260
rect 675201 246258 675267 246261
rect 675334 246258 675340 246260
rect 675201 246256 675340 246258
rect 675201 246200 675206 246256
rect 675262 246200 675340 246256
rect 675201 246198 675340 246200
rect 675201 246195 675267 246198
rect 675334 246196 675340 246198
rect 675404 246196 675410 246260
rect 673821 246124 673887 246125
rect 673821 246120 673868 246124
rect 673932 246122 673938 246124
rect 673821 246064 673826 246120
rect 673821 246060 673868 246064
rect 673932 246062 673978 246122
rect 673932 246060 673938 246062
rect 673821 246059 673887 246060
rect 42190 245788 42196 245852
rect 42260 245850 42266 245852
rect 42793 245850 42859 245853
rect 42260 245848 42859 245850
rect 42260 245792 42798 245848
rect 42854 245792 42859 245848
rect 42260 245790 42859 245792
rect 42260 245788 42266 245790
rect 42793 245787 42859 245790
rect 41822 245652 41828 245716
rect 41892 245714 41898 245716
rect 42701 245714 42767 245717
rect 41892 245712 42767 245714
rect 41892 245656 42706 245712
rect 42762 245656 42767 245712
rect 41892 245654 42767 245656
rect 41892 245652 41898 245654
rect 42701 245651 42767 245654
rect 40033 244628 40099 244629
rect 39982 244626 39988 244628
rect 39942 244566 39988 244626
rect 40052 244624 40099 244628
rect 40094 244568 40099 244624
rect 39982 244564 39988 244566
rect 40052 244564 40099 244568
rect 40033 244563 40099 244564
rect 40033 244218 40099 244221
rect 40166 244218 40172 244220
rect 40033 244216 40172 244218
rect 40033 244160 40038 244216
rect 40094 244160 40172 244216
rect 40033 244158 40172 244160
rect 40033 244155 40099 244158
rect 40166 244156 40172 244158
rect 40236 244156 40242 244220
rect 31017 243538 31083 243541
rect 40493 243538 40559 243541
rect 31017 243536 40559 243538
rect 31017 243480 31022 243536
rect 31078 243480 40498 243536
rect 40554 243480 40559 243536
rect 31017 243478 40559 243480
rect 31017 243475 31083 243478
rect 40493 243475 40559 243478
rect 414381 243130 414447 243133
rect 412436 243128 414447 243130
rect 412436 243072 414386 243128
rect 414442 243072 414447 243128
rect 412436 243070 414447 243072
rect 414381 243067 414447 243070
rect 674966 241844 674972 241908
rect 675036 241906 675042 241908
rect 675293 241906 675359 241909
rect 675036 241904 675359 241906
rect 675036 241848 675298 241904
rect 675354 241848 675359 241904
rect 675036 241846 675359 241848
rect 675036 241844 675042 241846
rect 675293 241843 675359 241846
rect 39941 241634 40007 241637
rect 43161 241634 43227 241637
rect 39941 241632 43227 241634
rect 39941 241576 39946 241632
rect 40002 241576 43166 241632
rect 43222 241576 43227 241632
rect 39941 241574 43227 241576
rect 39941 241571 40007 241574
rect 43161 241571 43227 241574
rect 40493 240954 40559 240957
rect 40493 240952 40602 240954
rect 40493 240896 40498 240952
rect 40554 240896 40602 240952
rect 40493 240891 40602 240896
rect 40542 238914 40602 240891
rect 675385 240276 675451 240277
rect 675334 240274 675340 240276
rect 675294 240214 675340 240274
rect 675404 240272 675451 240276
rect 675446 240216 675451 240272
rect 675334 240212 675340 240214
rect 675404 240212 675451 240216
rect 675385 240211 675451 240212
rect 414289 240002 414355 240005
rect 412436 240000 414355 240002
rect 412436 239944 414294 240000
rect 414350 239944 414355 240000
rect 412436 239942 414355 239944
rect 414289 239939 414355 239942
rect 40718 238988 40724 239052
rect 40788 239050 40794 239052
rect 40788 238990 41706 239050
rect 40788 238988 40794 238990
rect 40542 238854 41430 238914
rect 41370 238778 41430 238854
rect 41370 238718 41522 238778
rect 40350 238444 40356 238508
rect 40420 238506 40426 238508
rect 40420 238446 41338 238506
rect 40420 238444 40426 238446
rect 40534 238172 40540 238236
rect 40604 238234 40610 238236
rect 40604 238174 41154 238234
rect 40604 238172 40610 238174
rect 41094 238100 41154 238174
rect 41278 238100 41338 238446
rect 41462 238100 41522 238718
rect 41646 238100 41706 238990
rect 42701 238914 42767 238917
rect 41830 238912 42767 238914
rect 41830 238856 42706 238912
rect 42762 238856 42767 238912
rect 41830 238854 42767 238856
rect 41830 238509 41890 238854
rect 42701 238851 42767 238854
rect 41830 238504 41939 238509
rect 41830 238448 41878 238504
rect 41934 238448 41939 238504
rect 41830 238446 41939 238448
rect 41873 238443 41939 238446
rect 675753 238506 675819 238509
rect 676990 238506 676996 238508
rect 675753 238504 676996 238506
rect 675753 238448 675758 238504
rect 675814 238448 676996 238504
rect 675753 238446 676996 238448
rect 675753 238443 675819 238446
rect 676990 238444 676996 238446
rect 677060 238444 677066 238508
rect 41086 238036 41092 238100
rect 41156 238036 41162 238100
rect 41270 238036 41276 238100
rect 41340 238036 41346 238100
rect 41454 238036 41460 238100
rect 41524 238036 41530 238100
rect 41638 238036 41644 238100
rect 41708 238036 41714 238100
rect 42190 238036 42196 238100
rect 42260 238098 42266 238100
rect 42793 238098 42859 238101
rect 42260 238096 42859 238098
rect 42260 238040 42798 238096
rect 42854 238040 42859 238096
rect 42260 238038 42859 238040
rect 42260 238036 42266 238038
rect 42793 238035 42859 238038
rect 42558 237900 42564 237964
rect 42628 237962 42634 237964
rect 42701 237962 42767 237965
rect 42628 237960 42767 237962
rect 42628 237904 42706 237960
rect 42762 237904 42767 237960
rect 42628 237902 42767 237904
rect 42628 237900 42634 237902
rect 42701 237899 42767 237902
rect 189073 237418 189139 237421
rect 189073 237416 191820 237418
rect 189073 237360 189078 237416
rect 189134 237360 191820 237416
rect 189073 237358 191820 237360
rect 189073 237355 189139 237358
rect 675753 236874 675819 236877
rect 677174 236874 677180 236876
rect 675753 236872 677180 236874
rect 675753 236816 675758 236872
rect 675814 236816 677180 236872
rect 675753 236814 677180 236816
rect 675753 236811 675819 236814
rect 677174 236812 677180 236814
rect 677244 236812 677250 236876
rect 40534 236676 40540 236740
rect 40604 236738 40610 236740
rect 41781 236738 41847 236741
rect 414933 236738 414999 236741
rect 40604 236736 41847 236738
rect 40604 236680 41786 236736
rect 41842 236680 41847 236736
rect 40604 236678 41847 236680
rect 412436 236736 414999 236738
rect 412436 236680 414938 236736
rect 414994 236680 414999 236736
rect 412436 236678 414999 236680
rect 40604 236676 40610 236678
rect 41781 236675 41847 236678
rect 414933 236675 414999 236678
rect 41270 234772 41276 234836
rect 41340 234834 41346 234836
rect 41781 234834 41847 234837
rect 41340 234832 41847 234834
rect 41340 234776 41786 234832
rect 41842 234776 41847 234832
rect 41340 234774 41847 234776
rect 41340 234772 41346 234774
rect 41781 234771 41847 234774
rect 414197 233610 414263 233613
rect 412436 233608 414263 233610
rect 412436 233552 414202 233608
rect 414258 233552 414263 233608
rect 412436 233550 414263 233552
rect 414197 233547 414263 233550
rect 41454 233276 41460 233340
rect 41524 233338 41530 233340
rect 41781 233338 41847 233341
rect 41524 233336 41847 233338
rect 41524 233280 41786 233336
rect 41842 233280 41847 233336
rect 41524 233278 41847 233280
rect 41524 233276 41530 233278
rect 41781 233275 41847 233278
rect 40718 230420 40724 230484
rect 40788 230482 40794 230484
rect 41781 230482 41847 230485
rect 40788 230480 41847 230482
rect 40788 230424 41786 230480
rect 41842 230424 41847 230480
rect 40788 230422 41847 230424
rect 40788 230420 40794 230422
rect 41781 230419 41847 230422
rect 647325 230482 647391 230485
rect 647734 230482 647740 230484
rect 647325 230480 647740 230482
rect 647325 230424 647330 230480
rect 647386 230424 647740 230480
rect 647325 230422 647740 230424
rect 647325 230419 647391 230422
rect 647734 230420 647740 230422
rect 647804 230420 647810 230484
rect 196617 230346 196683 230349
rect 199009 230346 199075 230349
rect 196617 230344 199075 230346
rect 196617 230288 196622 230344
rect 196678 230288 199014 230344
rect 199070 230288 199075 230344
rect 196617 230286 199075 230288
rect 196617 230283 196683 230286
rect 199009 230283 199075 230286
rect 376937 230346 377003 230349
rect 428641 230346 428707 230349
rect 376937 230344 428707 230346
rect 376937 230288 376942 230344
rect 376998 230288 428646 230344
rect 428702 230288 428707 230344
rect 376937 230286 428707 230288
rect 376937 230283 377003 230286
rect 428641 230283 428707 230286
rect 377305 230210 377371 230213
rect 478137 230210 478203 230213
rect 377305 230208 478203 230210
rect 377305 230152 377310 230208
rect 377366 230152 478142 230208
rect 478198 230152 478203 230208
rect 377305 230150 478203 230152
rect 377305 230147 377371 230150
rect 478137 230147 478203 230150
rect 375833 230074 375899 230077
rect 486417 230074 486483 230077
rect 375833 230072 486483 230074
rect 375833 230016 375838 230072
rect 375894 230016 486422 230072
rect 486478 230016 486483 230072
rect 375833 230014 486483 230016
rect 375833 230011 375899 230014
rect 486417 230011 486483 230014
rect 42149 229938 42215 229941
rect 42558 229938 42564 229940
rect 42149 229936 42564 229938
rect 42149 229880 42154 229936
rect 42210 229880 42564 229936
rect 42149 229878 42564 229880
rect 42149 229875 42215 229878
rect 42558 229876 42564 229878
rect 42628 229876 42634 229940
rect 66897 229938 66963 229941
rect 196157 229938 196223 229941
rect 66897 229936 196223 229938
rect 66897 229880 66902 229936
rect 66958 229880 196162 229936
rect 196218 229880 196223 229936
rect 66897 229878 196223 229880
rect 66897 229875 66963 229878
rect 196157 229875 196223 229878
rect 378685 229938 378751 229941
rect 493317 229938 493383 229941
rect 378685 229936 493383 229938
rect 378685 229880 378690 229936
rect 378746 229880 493322 229936
rect 493378 229880 493383 229936
rect 378685 229878 493383 229880
rect 378685 229875 378751 229878
rect 493317 229875 493383 229878
rect 58617 229802 58683 229805
rect 194777 229802 194843 229805
rect 58617 229800 194843 229802
rect 58617 229744 58622 229800
rect 58678 229744 194782 229800
rect 194838 229744 194843 229800
rect 58617 229742 194843 229744
rect 58617 229739 58683 229742
rect 194777 229739 194843 229742
rect 380157 229802 380223 229805
rect 496077 229802 496143 229805
rect 380157 229800 496143 229802
rect 380157 229744 380162 229800
rect 380218 229744 496082 229800
rect 496138 229744 496143 229800
rect 380157 229742 496143 229744
rect 380157 229739 380223 229742
rect 496077 229739 496143 229742
rect 41638 228924 41644 228988
rect 41708 228986 41714 228988
rect 41781 228986 41847 228989
rect 41708 228984 41847 228986
rect 41708 228928 41786 228984
rect 41842 228928 41847 228984
rect 41708 228926 41847 228928
rect 41708 228924 41714 228926
rect 41781 228923 41847 228926
rect 387241 228714 387307 228717
rect 513373 228714 513439 228717
rect 387241 228712 513439 228714
rect 387241 228656 387246 228712
rect 387302 228656 513378 228712
rect 513434 228656 513439 228712
rect 387241 228654 513439 228656
rect 387241 228651 387307 228654
rect 513373 228651 513439 228654
rect 399385 228578 399451 228581
rect 541525 228578 541591 228581
rect 399385 228576 541591 228578
rect 399385 228520 399390 228576
rect 399446 228520 541530 228576
rect 541586 228520 541591 228576
rect 399385 228518 541591 228520
rect 399385 228515 399451 228518
rect 541525 228515 541591 228518
rect 90541 228442 90607 228445
rect 207933 228442 207999 228445
rect 90541 228440 207999 228442
rect 90541 228384 90546 228440
rect 90602 228384 207938 228440
rect 207994 228384 207999 228440
rect 90541 228382 207999 228384
rect 90541 228379 90607 228382
rect 207933 228379 207999 228382
rect 402605 228442 402671 228445
rect 549253 228442 549319 228445
rect 402605 228440 549319 228442
rect 402605 228384 402610 228440
rect 402666 228384 549258 228440
rect 549314 228384 549319 228440
rect 402605 228382 549319 228384
rect 402605 228379 402671 228382
rect 549253 228379 549319 228382
rect 86861 228306 86927 228309
rect 206553 228306 206619 228309
rect 86861 228304 206619 228306
rect 86861 228248 86866 228304
rect 86922 228248 206558 228304
rect 206614 228248 206619 228304
rect 86861 228246 206619 228248
rect 86861 228243 86927 228246
rect 206553 228243 206619 228246
rect 411161 228306 411227 228309
rect 564433 228306 564499 228309
rect 411161 228304 564499 228306
rect 411161 228248 411166 228304
rect 411222 228248 564438 228304
rect 564494 228248 564499 228304
rect 411161 228246 564499 228248
rect 411161 228243 411227 228246
rect 564433 228243 564499 228246
rect 42057 227354 42123 227357
rect 42190 227354 42196 227356
rect 42057 227352 42196 227354
rect 42057 227296 42062 227352
rect 42118 227296 42196 227352
rect 42057 227294 42196 227296
rect 42057 227291 42123 227294
rect 42190 227292 42196 227294
rect 42260 227292 42266 227356
rect 380525 227354 380591 227357
rect 496905 227354 496971 227357
rect 380525 227352 496971 227354
rect 380525 227296 380530 227352
rect 380586 227296 496910 227352
rect 496966 227296 496971 227352
rect 380525 227294 496971 227296
rect 380525 227291 380591 227294
rect 496905 227291 496971 227294
rect 72969 227218 73035 227221
rect 201493 227218 201559 227221
rect 72969 227216 201559 227218
rect 72969 227160 72974 227216
rect 73030 227160 201498 227216
rect 201554 227160 201559 227216
rect 72969 227158 201559 227160
rect 72969 227155 73035 227158
rect 201493 227155 201559 227158
rect 383009 227218 383075 227221
rect 502517 227218 502583 227221
rect 383009 227216 502583 227218
rect 383009 227160 383014 227216
rect 383070 227160 502522 227216
rect 502578 227160 502583 227216
rect 383009 227158 502583 227160
rect 383009 227155 383075 227158
rect 502517 227155 502583 227158
rect 62757 227082 62823 227085
rect 197261 227082 197327 227085
rect 62757 227080 197327 227082
rect 62757 227024 62762 227080
rect 62818 227024 197266 227080
rect 197322 227024 197327 227080
rect 62757 227022 197327 227024
rect 62757 227019 62823 227022
rect 197261 227019 197327 227022
rect 388345 227082 388411 227085
rect 515489 227082 515555 227085
rect 388345 227080 515555 227082
rect 388345 227024 388350 227080
rect 388406 227024 515494 227080
rect 515550 227024 515555 227080
rect 388345 227022 515555 227024
rect 388345 227019 388411 227022
rect 515489 227019 515555 227022
rect 59261 226946 59327 226949
rect 195789 226946 195855 226949
rect 59261 226944 195855 226946
rect 59261 226888 59266 226944
rect 59322 226888 195794 226944
rect 195850 226888 195855 226944
rect 59261 226886 195855 226888
rect 59261 226883 59327 226886
rect 195789 226883 195855 226886
rect 407941 226946 408007 226949
rect 561673 226946 561739 226949
rect 407941 226944 561739 226946
rect 407941 226888 407946 226944
rect 408002 226888 561678 226944
rect 561734 226888 561739 226944
rect 407941 226886 561739 226888
rect 407941 226883 408007 226886
rect 561673 226883 561739 226886
rect 40534 226068 40540 226132
rect 40604 226130 40610 226132
rect 41781 226130 41847 226133
rect 40604 226128 41847 226130
rect 40604 226072 41786 226128
rect 41842 226072 41847 226128
rect 40604 226070 41847 226072
rect 40604 226068 40610 226070
rect 41781 226067 41847 226070
rect 390829 225994 390895 225997
rect 521653 225994 521719 225997
rect 390829 225992 521719 225994
rect 390829 225936 390834 225992
rect 390890 225936 521658 225992
rect 521714 225936 521719 225992
rect 390829 225934 521719 225936
rect 390829 225931 390895 225934
rect 521653 225931 521719 225934
rect 394049 225858 394115 225861
rect 528921 225858 528987 225861
rect 394049 225856 528987 225858
rect 394049 225800 394054 225856
rect 394110 225800 528926 225856
rect 528982 225800 528987 225856
rect 394049 225798 528987 225800
rect 394049 225795 394115 225798
rect 528921 225795 528987 225798
rect 93025 225722 93091 225725
rect 210049 225722 210115 225725
rect 93025 225720 210115 225722
rect 93025 225664 93030 225720
rect 93086 225664 210054 225720
rect 210110 225664 210115 225720
rect 93025 225662 210115 225664
rect 93025 225659 93091 225662
rect 210049 225659 210115 225662
rect 396441 225722 396507 225725
rect 534073 225722 534139 225725
rect 396441 225720 534139 225722
rect 396441 225664 396446 225720
rect 396502 225664 534078 225720
rect 534134 225664 534139 225720
rect 396441 225662 534139 225664
rect 396441 225659 396507 225662
rect 534073 225659 534139 225662
rect 89529 225586 89595 225589
rect 208669 225586 208735 225589
rect 89529 225584 208735 225586
rect 89529 225528 89534 225584
rect 89590 225528 208674 225584
rect 208730 225528 208735 225584
rect 89529 225526 208735 225528
rect 89529 225523 89595 225526
rect 208669 225523 208735 225526
rect 400489 225586 400555 225589
rect 544009 225586 544075 225589
rect 400489 225584 544075 225586
rect 400489 225528 400494 225584
rect 400550 225528 544014 225584
rect 544070 225528 544075 225584
rect 400489 225526 544075 225528
rect 400489 225523 400555 225526
rect 544009 225523 544075 225526
rect 78489 224634 78555 224637
rect 202597 224634 202663 224637
rect 78489 224632 202663 224634
rect 78489 224576 78494 224632
rect 78550 224576 202602 224632
rect 202658 224576 202663 224632
rect 78489 224574 202663 224576
rect 78489 224571 78555 224574
rect 202597 224571 202663 224574
rect 377673 224634 377739 224637
rect 490189 224634 490255 224637
rect 377673 224632 490255 224634
rect 377673 224576 377678 224632
rect 377734 224576 490194 224632
rect 490250 224576 490255 224632
rect 377673 224574 490255 224576
rect 377673 224571 377739 224574
rect 490189 224571 490255 224574
rect 72049 224498 72115 224501
rect 199745 224498 199811 224501
rect 72049 224496 199811 224498
rect 72049 224440 72054 224496
rect 72110 224440 199750 224496
rect 199806 224440 199811 224496
rect 72049 224438 199811 224440
rect 72049 224435 72115 224438
rect 199745 224435 199811 224438
rect 381905 224498 381971 224501
rect 499573 224498 499639 224501
rect 381905 224496 499639 224498
rect 381905 224440 381910 224496
rect 381966 224440 499578 224496
rect 499634 224440 499639 224496
rect 381905 224438 499639 224440
rect 381905 224435 381971 224438
rect 499573 224435 499639 224438
rect 69473 224362 69539 224365
rect 200113 224362 200179 224365
rect 69473 224360 200179 224362
rect 69473 224304 69478 224360
rect 69534 224304 200118 224360
rect 200174 224304 200179 224360
rect 69473 224302 200179 224304
rect 69473 224299 69539 224302
rect 200113 224299 200179 224302
rect 384021 224362 384087 224365
rect 505369 224362 505435 224365
rect 384021 224360 505435 224362
rect 384021 224304 384026 224360
rect 384082 224304 505374 224360
rect 505430 224304 505435 224360
rect 384021 224302 505435 224304
rect 384021 224299 384087 224302
rect 505369 224299 505435 224302
rect 62021 224226 62087 224229
rect 195421 224226 195487 224229
rect 62021 224224 195487 224226
rect 62021 224168 62026 224224
rect 62082 224168 195426 224224
rect 195482 224168 195487 224224
rect 62021 224166 195487 224168
rect 62021 224163 62087 224166
rect 195421 224163 195487 224166
rect 409597 224226 409663 224229
rect 556705 224226 556771 224229
rect 409597 224224 556771 224226
rect 409597 224168 409602 224224
rect 409658 224168 556710 224224
rect 556766 224168 556771 224224
rect 409597 224166 556771 224168
rect 409597 224163 409663 224166
rect 556705 224163 556771 224166
rect 676029 223546 676095 223549
rect 676029 223544 676292 223546
rect 676029 223488 676034 223544
rect 676090 223488 676292 223544
rect 676029 223486 676292 223488
rect 676029 223483 676095 223486
rect 376201 223410 376267 223413
rect 487797 223410 487863 223413
rect 376201 223408 487863 223410
rect 376201 223352 376206 223408
rect 376262 223352 487802 223408
rect 487858 223352 487863 223408
rect 376201 223350 487863 223352
rect 376201 223347 376267 223350
rect 487797 223347 487863 223350
rect 99005 223274 99071 223277
rect 211153 223274 211219 223277
rect 99005 223272 211219 223274
rect 99005 223216 99010 223272
rect 99066 223216 211158 223272
rect 211214 223216 211219 223272
rect 99005 223214 211219 223216
rect 99005 223211 99071 223214
rect 211153 223211 211219 223214
rect 379053 223274 379119 223277
rect 494053 223274 494119 223277
rect 379053 223272 494119 223274
rect 379053 223216 379058 223272
rect 379114 223216 494058 223272
rect 494114 223216 494119 223272
rect 379053 223214 494119 223216
rect 379053 223211 379119 223214
rect 494053 223211 494119 223214
rect 92289 223138 92355 223141
rect 208025 223138 208091 223141
rect 92289 223136 208091 223138
rect 92289 223080 92294 223136
rect 92350 223080 208030 223136
rect 208086 223080 208091 223136
rect 92289 223078 208091 223080
rect 92289 223075 92355 223078
rect 208025 223075 208091 223078
rect 389357 223138 389423 223141
rect 518157 223138 518223 223141
rect 389357 223136 518223 223138
rect 389357 223080 389362 223136
rect 389418 223080 518162 223136
rect 518218 223080 518223 223136
rect 389357 223078 518223 223080
rect 389357 223075 389423 223078
rect 518157 223075 518223 223078
rect 675937 223138 676003 223141
rect 675937 223136 676292 223138
rect 675937 223080 675942 223136
rect 675998 223080 676292 223136
rect 675937 223078 676292 223080
rect 675937 223075 676003 223078
rect 58709 223002 58775 223005
rect 194041 223002 194107 223005
rect 58709 223000 194107 223002
rect 58709 222944 58714 223000
rect 58770 222944 194046 223000
rect 194102 222944 194107 223000
rect 58709 222942 194107 222944
rect 58709 222939 58775 222942
rect 194041 222939 194107 222942
rect 390461 223002 390527 223005
rect 520457 223002 520523 223005
rect 390461 223000 520523 223002
rect 390461 222944 390466 223000
rect 390522 222944 520462 223000
rect 520518 222944 520523 223000
rect 390461 222942 520523 222944
rect 390461 222939 390527 222942
rect 520457 222939 520523 222942
rect 55029 222866 55095 222869
rect 192385 222866 192451 222869
rect 55029 222864 192451 222866
rect 55029 222808 55034 222864
rect 55090 222808 192390 222864
rect 192446 222808 192451 222864
rect 55029 222806 192451 222808
rect 55029 222803 55095 222806
rect 192385 222803 192451 222806
rect 410977 222866 411043 222869
rect 569309 222866 569375 222869
rect 410977 222864 569375 222866
rect 410977 222808 410982 222864
rect 411038 222808 569314 222864
rect 569370 222808 569375 222864
rect 410977 222806 569375 222808
rect 410977 222803 411043 222806
rect 569309 222803 569375 222806
rect 675937 222730 676003 222733
rect 675937 222728 676292 222730
rect 675937 222672 675942 222728
rect 675998 222672 676292 222728
rect 675937 222670 676292 222672
rect 675937 222667 676003 222670
rect 674741 222322 674807 222325
rect 674741 222320 676292 222322
rect 674741 222264 674746 222320
rect 674802 222264 676292 222320
rect 674741 222262 676292 222264
rect 674741 222259 674807 222262
rect 73705 221914 73771 221917
rect 200573 221914 200639 221917
rect 73705 221912 200639 221914
rect 73705 221856 73710 221912
rect 73766 221856 200578 221912
rect 200634 221856 200639 221912
rect 73705 221854 200639 221856
rect 73705 221851 73771 221854
rect 200573 221851 200639 221854
rect 400949 221914 401015 221917
rect 528093 221914 528159 221917
rect 400949 221912 528159 221914
rect 400949 221856 400954 221912
rect 401010 221856 528098 221912
rect 528154 221856 528159 221912
rect 400949 221854 528159 221856
rect 400949 221851 401015 221854
rect 528093 221851 528159 221854
rect 676029 221914 676095 221917
rect 676029 221912 676292 221914
rect 676029 221856 676034 221912
rect 676090 221856 676292 221912
rect 676029 221854 676292 221856
rect 676029 221851 676095 221854
rect 70209 221778 70275 221781
rect 199101 221778 199167 221781
rect 70209 221776 199167 221778
rect 70209 221720 70214 221776
rect 70270 221720 199106 221776
rect 199162 221720 199167 221776
rect 70209 221718 199167 221720
rect 70209 221715 70275 221718
rect 199101 221715 199167 221718
rect 392853 221778 392919 221781
rect 525885 221778 525951 221781
rect 392853 221776 525951 221778
rect 392853 221720 392858 221776
rect 392914 221720 525890 221776
rect 525946 221720 525951 221776
rect 392853 221718 525951 221720
rect 392853 221715 392919 221718
rect 525885 221715 525951 221718
rect 66989 221642 67055 221645
rect 197721 221642 197787 221645
rect 66989 221640 197787 221642
rect 66989 221584 66994 221640
rect 67050 221584 197726 221640
rect 197782 221584 197787 221640
rect 66989 221582 197787 221584
rect 66989 221579 67055 221582
rect 197721 221579 197787 221582
rect 397177 221642 397243 221645
rect 536005 221642 536071 221645
rect 397177 221640 536071 221642
rect 397177 221584 397182 221640
rect 397238 221584 536010 221640
rect 536066 221584 536071 221640
rect 397177 221582 536071 221584
rect 397177 221579 397243 221582
rect 536005 221579 536071 221582
rect 56869 221506 56935 221509
rect 193397 221506 193463 221509
rect 56869 221504 193463 221506
rect 56869 221448 56874 221504
rect 56930 221448 193402 221504
rect 193458 221448 193463 221504
rect 56869 221446 193463 221448
rect 56869 221443 56935 221446
rect 193397 221443 193463 221446
rect 404997 221506 405063 221509
rect 546677 221506 546743 221509
rect 404997 221504 546743 221506
rect 404997 221448 405002 221504
rect 405058 221448 546682 221504
rect 546738 221448 546743 221504
rect 404997 221446 546743 221448
rect 404997 221443 405063 221446
rect 546677 221443 546743 221446
rect 676029 221506 676095 221509
rect 676029 221504 676292 221506
rect 676029 221448 676034 221504
rect 676090 221448 676292 221504
rect 676029 221446 676292 221448
rect 676029 221443 676095 221446
rect 6022 221353 55460 221382
rect 6022 220209 6150 221353
rect 6854 221349 55460 221353
rect 6854 220245 54235 221349
rect 55339 220245 55460 221349
rect 676029 221098 676095 221101
rect 676029 221096 676292 221098
rect 676029 221040 676034 221096
rect 676090 221040 676292 221096
rect 676029 221038 676292 221040
rect 676029 221035 676095 221038
rect 676029 220690 676095 220693
rect 676029 220688 676292 220690
rect 676029 220632 676034 220688
rect 676090 220632 676292 220688
rect 676029 220630 676292 220632
rect 676029 220627 676095 220630
rect 389173 220554 389239 220557
rect 495617 220554 495683 220557
rect 389173 220552 495683 220554
rect 389173 220496 389178 220552
rect 389234 220496 495622 220552
rect 495678 220496 495683 220552
rect 389173 220494 495683 220496
rect 389173 220491 389239 220494
rect 495617 220491 495683 220494
rect 382181 220418 382247 220421
rect 498653 220418 498719 220421
rect 382181 220416 498719 220418
rect 382181 220360 382186 220416
rect 382242 220360 498658 220416
rect 498714 220360 498719 220416
rect 382181 220358 498719 220360
rect 382181 220355 382247 220358
rect 498653 220355 498719 220358
rect 6854 220209 55460 220245
rect 74441 220282 74507 220285
rect 201585 220282 201651 220285
rect 74441 220280 201651 220282
rect 74441 220224 74446 220280
rect 74502 220224 201590 220280
rect 201646 220224 201651 220280
rect 74441 220222 201651 220224
rect 74441 220219 74507 220222
rect 201585 220219 201651 220222
rect 381905 220282 381971 220285
rect 499665 220282 499731 220285
rect 381905 220280 499731 220282
rect 381905 220224 381910 220280
rect 381966 220224 499670 220280
rect 499726 220224 499731 220280
rect 381905 220222 499731 220224
rect 381905 220219 381971 220222
rect 499665 220219 499731 220222
rect 676029 220282 676095 220285
rect 676029 220280 676292 220282
rect 676029 220224 676034 220280
rect 676090 220224 676292 220280
rect 676029 220222 676292 220224
rect 676029 220219 676095 220222
rect 6022 220182 55460 220209
rect 67541 220146 67607 220149
rect 196617 220146 196683 220149
rect 67541 220144 196683 220146
rect 67541 220088 67546 220144
rect 67602 220088 196622 220144
rect 196678 220088 196683 220144
rect 67541 220086 196683 220088
rect 67541 220083 67607 220086
rect 196617 220083 196683 220086
rect 384849 220146 384915 220149
rect 507209 220146 507275 220149
rect 384849 220144 507275 220146
rect 384849 220088 384854 220144
rect 384910 220088 507214 220144
rect 507270 220088 507275 220144
rect 384849 220086 507275 220088
rect 384849 220083 384915 220086
rect 507209 220083 507275 220086
rect 676029 219874 676095 219877
rect 676029 219872 676292 219874
rect 676029 219816 676034 219872
rect 676090 219816 676292 219872
rect 676029 219814 676292 219816
rect 676029 219811 676095 219814
rect 7236 219757 53816 219782
rect 7236 218613 7348 219757
rect 8052 219731 53816 219757
rect 8052 218627 52641 219731
rect 53745 218627 53816 219731
rect 507209 219466 507275 219469
rect 623957 219466 624023 219469
rect 507209 219464 624023 219466
rect 507209 219408 507214 219464
rect 507270 219408 623962 219464
rect 624018 219408 624023 219464
rect 507209 219406 624023 219408
rect 507209 219403 507275 219406
rect 623957 219403 624023 219406
rect 674741 219466 674807 219469
rect 674741 219464 676292 219466
rect 674741 219408 674746 219464
rect 674802 219408 676292 219464
rect 674741 219406 676292 219408
rect 674741 219403 674807 219406
rect 676029 219058 676095 219061
rect 676029 219056 676292 219058
rect 676029 219000 676034 219056
rect 676090 219000 676292 219056
rect 676029 218998 676292 219000
rect 676029 218995 676095 218998
rect 8052 218613 53816 218627
rect 7236 218582 53816 218613
rect 676024 218588 676030 218652
rect 676094 218650 676100 218652
rect 676094 218590 676292 218650
rect 676094 218588 676100 218590
rect 654133 218514 654199 218517
rect 55170 218512 654199 218514
rect 55170 218456 654138 218512
rect 654194 218456 654199 218512
rect 55170 218454 654199 218456
rect 53097 218378 53163 218381
rect 55170 218378 55230 218454
rect 654133 218451 654199 218454
rect 53097 218376 55230 218378
rect 53097 218320 53102 218376
rect 53158 218320 55230 218376
rect 53097 218318 55230 218320
rect 53097 218315 53163 218318
rect 675334 218180 675340 218244
rect 675404 218242 675410 218244
rect 675404 218182 676292 218242
rect 675404 218180 675410 218182
rect 675886 217772 675892 217836
rect 675956 217834 675962 217836
rect 675956 217774 676292 217834
rect 675956 217772 675962 217774
rect 679617 217426 679683 217429
rect 679604 217424 679683 217426
rect 679604 217368 679622 217424
rect 679678 217368 679683 217424
rect 679604 217366 679683 217368
rect 679617 217363 679683 217366
rect 676078 216958 676292 217018
rect 489085 216882 489151 216885
rect 610341 216882 610407 216885
rect 676078 216884 676138 216958
rect 489085 216880 610407 216882
rect 489085 216824 489090 216880
rect 489146 216824 610346 216880
rect 610402 216824 610407 216880
rect 489085 216822 610407 216824
rect 489085 216819 489151 216822
rect 610341 216819 610407 216822
rect 676070 216820 676076 216884
rect 676140 216820 676146 216884
rect 495985 216746 496051 216749
rect 622485 216746 622551 216749
rect 495985 216744 622551 216746
rect 495985 216688 495990 216744
rect 496046 216688 622490 216744
rect 622546 216688 622551 216744
rect 495985 216686 622551 216688
rect 495985 216683 496051 216686
rect 622485 216683 622551 216686
rect 676029 216610 676095 216613
rect 676029 216608 676292 216610
rect 676029 216552 676034 216608
rect 676090 216552 676292 216608
rect 676029 216550 676292 216552
rect 676029 216547 676095 216550
rect 578877 216202 578943 216205
rect 576380 216200 578943 216202
rect 576380 216144 578882 216200
rect 578938 216144 578943 216200
rect 576380 216142 578943 216144
rect 578877 216139 578943 216142
rect 676029 216202 676095 216205
rect 676029 216200 676292 216202
rect 676029 216144 676034 216200
rect 676090 216144 676292 216200
rect 676029 216142 676292 216144
rect 676029 216139 676095 216142
rect 676029 215794 676095 215797
rect 676029 215792 676292 215794
rect 676029 215736 676034 215792
rect 676090 215736 676292 215792
rect 676029 215734 676292 215736
rect 676029 215731 676095 215734
rect 675937 215386 676003 215389
rect 675937 215384 676292 215386
rect 675937 215328 675942 215384
rect 675998 215328 676292 215384
rect 675937 215326 676292 215328
rect 675937 215323 676003 215326
rect 675845 214978 675911 214981
rect 675845 214976 676292 214978
rect 35758 214709 35818 214948
rect 675845 214920 675850 214976
rect 675906 214920 676292 214976
rect 675845 214918 676292 214920
rect 675845 214915 675911 214918
rect 35617 214706 35683 214709
rect 35574 214704 35683 214706
rect 35574 214648 35622 214704
rect 35678 214648 35683 214704
rect 35574 214643 35683 214648
rect 35758 214704 35867 214709
rect 579061 214706 579127 214709
rect 35758 214648 35806 214704
rect 35862 214648 35867 214704
rect 35758 214646 35867 214648
rect 576380 214704 579127 214706
rect 576380 214648 579066 214704
rect 579122 214648 579127 214704
rect 576380 214646 579127 214648
rect 35801 214643 35867 214646
rect 579061 214643 579127 214646
rect 35574 214540 35634 214643
rect 676998 214334 677058 214540
rect 35709 214298 35775 214301
rect 35709 214296 35818 214298
rect 35709 214240 35714 214296
rect 35770 214240 35818 214296
rect 676990 214270 676996 214334
rect 677060 214270 677066 214334
rect 35709 214235 35818 214240
rect 35758 214132 35818 214235
rect 676029 214162 676095 214165
rect 676029 214160 676292 214162
rect 676029 214104 676034 214160
rect 676090 214104 676292 214160
rect 676029 214102 676292 214104
rect 676029 214099 676095 214102
rect 675702 213964 675708 214028
rect 675772 214026 675778 214028
rect 676029 214026 676095 214029
rect 675772 214024 676095 214026
rect 675772 213968 676034 214024
rect 676090 213968 676095 214024
rect 675772 213966 676095 213968
rect 675772 213964 675778 213966
rect 676029 213963 676095 213966
rect 42885 213754 42951 213757
rect 41492 213752 42951 213754
rect 41492 213696 42890 213752
rect 42946 213696 42951 213752
rect 41492 213694 42951 213696
rect 42885 213691 42951 213694
rect 676029 213754 676095 213757
rect 676029 213752 676292 213754
rect 676029 213696 676034 213752
rect 676090 213696 676292 213752
rect 676029 213694 676292 213696
rect 676029 213691 676095 213694
rect 46565 213346 46631 213349
rect 41492 213344 46631 213346
rect 41492 213288 46570 213344
rect 46626 213288 46631 213344
rect 41492 213286 46631 213288
rect 46565 213283 46631 213286
rect 676029 213346 676095 213349
rect 676029 213344 676292 213346
rect 676029 213288 676034 213344
rect 676090 213288 676292 213344
rect 676029 213286 676292 213288
rect 676029 213283 676095 213286
rect 578969 213210 579035 213213
rect 576380 213208 579035 213210
rect 576380 213152 578974 213208
rect 579030 213152 579035 213208
rect 576380 213150 579035 213152
rect 578969 213147 579035 213150
rect 647734 213012 647740 213076
rect 647804 213074 647810 213076
rect 648521 213074 648587 213077
rect 647804 213072 648587 213074
rect 647804 213016 648526 213072
rect 648582 213016 648587 213072
rect 647804 213014 648587 213016
rect 647804 213012 647810 213014
rect 648521 213011 648587 213014
rect 43069 212938 43135 212941
rect 41492 212936 43135 212938
rect 41492 212880 43074 212936
rect 43130 212880 43135 212936
rect 41492 212878 43135 212880
rect 43069 212875 43135 212878
rect 42793 212530 42859 212533
rect 41492 212528 42859 212530
rect 41492 212472 42798 212528
rect 42854 212472 42859 212528
rect 676262 212500 676322 212908
rect 41492 212470 42859 212472
rect 42793 212467 42859 212470
rect 44633 212122 44699 212125
rect 41492 212120 44699 212122
rect 41492 212064 44638 212120
rect 44694 212064 44699 212120
rect 41492 212062 44699 212064
rect 44633 212059 44699 212062
rect 676029 212122 676095 212125
rect 676029 212120 676292 212122
rect 676029 212064 676034 212120
rect 676090 212064 676292 212120
rect 676029 212062 676292 212064
rect 676029 212059 676095 212062
rect 41781 211714 41847 211717
rect 578417 211714 578483 211717
rect 41492 211712 41847 211714
rect 41492 211656 41786 211712
rect 41842 211656 41847 211712
rect 41492 211654 41847 211656
rect 576380 211712 578483 211714
rect 576380 211656 578422 211712
rect 578478 211656 578483 211712
rect 576380 211654 578483 211656
rect 41781 211651 41847 211654
rect 578417 211651 578483 211654
rect 675937 211442 676003 211445
rect 676622 211442 676628 211444
rect 675937 211440 676628 211442
rect 675937 211384 675942 211440
rect 675998 211384 676628 211440
rect 675937 211382 676628 211384
rect 675937 211379 676003 211382
rect 676622 211380 676628 211382
rect 676692 211380 676698 211444
rect 44265 211306 44331 211309
rect 41492 211304 44331 211306
rect 41492 211248 44270 211304
rect 44326 211248 44331 211304
rect 41492 211246 44331 211248
rect 44265 211243 44331 211246
rect 675845 211306 675911 211309
rect 676806 211306 676812 211308
rect 675845 211304 676812 211306
rect 675845 211248 675850 211304
rect 675906 211248 676812 211304
rect 675845 211246 676812 211248
rect 675845 211243 675911 211246
rect 676806 211244 676812 211246
rect 676876 211244 676882 211308
rect 41321 211034 41387 211037
rect 41278 211032 41387 211034
rect 41278 210976 41326 211032
rect 41382 210976 41387 211032
rect 41278 210971 41387 210976
rect 41278 210868 41338 210971
rect 31158 210221 31218 210460
rect 31158 210216 31267 210221
rect 578509 210218 578575 210221
rect 31158 210160 31206 210216
rect 31262 210160 31267 210216
rect 31158 210158 31267 210160
rect 576380 210216 578575 210218
rect 576380 210160 578514 210216
rect 578570 210160 578575 210216
rect 576380 210158 578575 210160
rect 31201 210155 31267 210158
rect 578509 210155 578575 210158
rect 30974 209813 31034 210052
rect 30974 209808 31083 209813
rect 30974 209752 31022 209808
rect 31078 209752 31083 209808
rect 30974 209750 31083 209752
rect 31017 209747 31083 209750
rect 40542 209404 40602 209644
rect 603073 209538 603139 209541
rect 603073 209536 606556 209538
rect 603073 209480 603078 209536
rect 603134 209480 606556 209536
rect 603073 209478 606556 209480
rect 603073 209475 603139 209478
rect 40534 209340 40540 209404
rect 40604 209340 40610 209404
rect 42793 209266 42859 209269
rect 666921 209266 666987 209269
rect 667933 209266 667999 209269
rect 41492 209264 42859 209266
rect 41492 209208 42798 209264
rect 42854 209208 42859 209264
rect 41492 209206 42859 209208
rect 666356 209264 667999 209266
rect 666356 209208 666926 209264
rect 666982 209208 667938 209264
rect 667994 209208 667999 209264
rect 666356 209206 667999 209208
rect 42793 209203 42859 209206
rect 666921 209203 666987 209206
rect 667933 209203 667999 209206
rect 39297 208586 39363 208589
rect 41462 208588 41522 208828
rect 579521 208722 579587 208725
rect 576380 208720 579587 208722
rect 576380 208664 579526 208720
rect 579582 208664 579587 208720
rect 576380 208662 579587 208664
rect 579521 208659 579587 208662
rect 39254 208584 39363 208586
rect 39254 208528 39302 208584
rect 39358 208528 39363 208584
rect 39254 208523 39363 208528
rect 41454 208524 41460 208588
rect 41524 208524 41530 208588
rect 603165 208586 603231 208589
rect 603165 208584 606556 208586
rect 603165 208528 603170 208584
rect 603226 208528 606556 208584
rect 603165 208526 606556 208528
rect 603165 208523 603231 208526
rect 39254 208420 39314 208523
rect 676070 208252 676076 208316
rect 676140 208314 676146 208316
rect 676857 208314 676923 208317
rect 676140 208312 676923 208314
rect 676140 208256 676862 208312
rect 676918 208256 676923 208312
rect 676140 208254 676923 208256
rect 676140 208252 676146 208254
rect 676857 208251 676923 208254
rect 44173 208042 44239 208045
rect 41492 208040 44239 208042
rect 41492 207984 44178 208040
rect 44234 207984 44239 208040
rect 41492 207982 44239 207984
rect 44173 207979 44239 207982
rect 42885 207634 42951 207637
rect 41492 207632 42951 207634
rect 41492 207576 42890 207632
rect 42946 207576 42951 207632
rect 41492 207574 42951 207576
rect 42885 207571 42951 207574
rect 603073 207498 603139 207501
rect 603073 207496 606556 207498
rect 603073 207440 603078 207496
rect 603134 207440 606556 207496
rect 603073 207438 606556 207440
rect 603073 207435 603139 207438
rect 578785 207226 578851 207229
rect 576380 207224 578851 207226
rect 40726 206956 40786 207196
rect 576380 207168 578790 207224
rect 578846 207168 578851 207224
rect 576380 207166 578851 207168
rect 578785 207163 578851 207166
rect 675518 207164 675524 207228
rect 675588 207226 675594 207228
rect 679617 207226 679683 207229
rect 675588 207224 679683 207226
rect 675588 207168 679622 207224
rect 679678 207168 679683 207224
rect 675588 207166 679683 207168
rect 675588 207164 675594 207166
rect 679617 207163 679683 207166
rect 40718 206892 40724 206956
rect 40788 206892 40794 206956
rect 44449 206818 44515 206821
rect 41492 206816 44515 206818
rect 41492 206760 44454 206816
rect 44510 206760 44515 206816
rect 41492 206758 44515 206760
rect 44449 206755 44515 206758
rect 603073 206546 603139 206549
rect 603073 206544 606556 206546
rect 603073 206488 603078 206544
rect 603134 206488 606556 206544
rect 603073 206486 606556 206488
rect 603073 206483 603139 206486
rect 42977 206410 43043 206413
rect 41492 206408 43043 206410
rect 41492 206352 42982 206408
rect 43038 206352 43043 206408
rect 41492 206350 43043 206352
rect 42977 206347 43043 206350
rect 44265 206002 44331 206005
rect 41492 206000 44331 206002
rect 41492 205944 44270 206000
rect 44326 205944 44331 206000
rect 41492 205942 44331 205944
rect 44265 205939 44331 205942
rect 667933 205866 667999 205869
rect 666356 205864 667999 205866
rect 666356 205808 667938 205864
rect 667994 205808 667999 205864
rect 666356 205806 667999 205808
rect 667933 205803 667999 205806
rect 579429 205730 579495 205733
rect 576380 205728 579495 205730
rect 576380 205672 579434 205728
rect 579490 205672 579495 205728
rect 576380 205670 579495 205672
rect 579429 205667 579495 205670
rect 43069 205594 43135 205597
rect 675385 205596 675451 205597
rect 675334 205594 675340 205596
rect 41492 205592 43135 205594
rect 41492 205536 43074 205592
rect 43130 205536 43135 205592
rect 41492 205534 43135 205536
rect 675294 205534 675340 205594
rect 675404 205592 675451 205596
rect 675446 205536 675451 205592
rect 43069 205531 43135 205534
rect 675334 205532 675340 205534
rect 675404 205532 675451 205536
rect 675385 205531 675451 205532
rect 603073 205458 603139 205461
rect 603073 205456 606556 205458
rect 603073 205400 603078 205456
rect 603134 205400 606556 205456
rect 603073 205398 606556 205400
rect 603073 205395 603139 205398
rect 44357 205186 44423 205189
rect 41492 205184 44423 205186
rect 41492 205128 44362 205184
rect 44418 205128 44423 205184
rect 41492 205126 44423 205128
rect 44357 205123 44423 205126
rect 675753 205050 675819 205053
rect 676070 205050 676076 205052
rect 675753 205048 676076 205050
rect 675753 204992 675758 205048
rect 675814 204992 676076 205048
rect 675753 204990 676076 204992
rect 675753 204987 675819 204990
rect 676070 204988 676076 204990
rect 676140 204988 676146 205052
rect 40861 204914 40927 204917
rect 40861 204912 40970 204914
rect 40861 204856 40866 204912
rect 40922 204856 40970 204912
rect 40861 204851 40970 204856
rect 40910 204748 40970 204851
rect 40677 204506 40743 204509
rect 603165 204506 603231 204509
rect 40677 204504 40786 204506
rect 40677 204448 40682 204504
rect 40738 204448 40786 204504
rect 40677 204443 40786 204448
rect 603165 204504 606556 204506
rect 603165 204448 603170 204504
rect 603226 204448 606556 204504
rect 603165 204446 606556 204448
rect 603165 204443 603231 204446
rect 40726 204340 40786 204443
rect 578877 204234 578943 204237
rect 666829 204234 666895 204237
rect 675753 204236 675819 204237
rect 675702 204234 675708 204236
rect 576380 204232 578943 204234
rect 576380 204176 578882 204232
rect 578938 204176 578943 204232
rect 576380 204174 578943 204176
rect 666356 204232 666895 204234
rect 666356 204176 666834 204232
rect 666890 204176 666895 204232
rect 666356 204174 666895 204176
rect 675662 204174 675708 204234
rect 675772 204232 675819 204236
rect 675814 204176 675819 204232
rect 578877 204171 578943 204174
rect 666829 204171 666895 204174
rect 675702 204172 675708 204174
rect 675772 204172 675819 204176
rect 675753 204171 675819 204172
rect 35758 203285 35818 203524
rect 603073 203418 603139 203421
rect 603073 203416 606556 203418
rect 603073 203360 603078 203416
rect 603134 203360 606556 203416
rect 603073 203358 606556 203360
rect 603073 203355 603139 203358
rect 35758 203280 35867 203285
rect 35758 203224 35806 203280
rect 35862 203224 35867 203280
rect 35758 203222 35867 203224
rect 35801 203219 35867 203222
rect 675109 202874 675175 202877
rect 676990 202874 676996 202876
rect 675109 202872 676996 202874
rect 675109 202816 675114 202872
rect 675170 202816 676996 202872
rect 675109 202814 676996 202816
rect 675109 202811 675175 202814
rect 676990 202812 676996 202814
rect 677060 202812 677066 202876
rect 579245 202738 579311 202741
rect 576380 202736 579311 202738
rect 576380 202680 579250 202736
rect 579306 202680 579311 202736
rect 576380 202678 579311 202680
rect 579245 202675 579311 202678
rect 675753 202738 675819 202741
rect 675886 202738 675892 202740
rect 675753 202736 675892 202738
rect 675753 202680 675758 202736
rect 675814 202680 675892 202736
rect 675753 202678 675892 202680
rect 675753 202675 675819 202678
rect 675886 202676 675892 202678
rect 675956 202676 675962 202740
rect 603073 202466 603139 202469
rect 603073 202464 606556 202466
rect 603073 202408 603078 202464
rect 603134 202408 606556 202464
rect 603073 202406 606556 202408
rect 603073 202403 603139 202406
rect 603073 201378 603139 201381
rect 674833 201378 674899 201381
rect 676806 201378 676812 201380
rect 603073 201376 606556 201378
rect 603073 201320 603078 201376
rect 603134 201320 606556 201376
rect 603073 201318 606556 201320
rect 674833 201376 676812 201378
rect 674833 201320 674838 201376
rect 674894 201320 676812 201376
rect 674833 201318 676812 201320
rect 603073 201315 603139 201318
rect 674833 201315 674899 201318
rect 676806 201316 676812 201318
rect 676876 201316 676882 201380
rect 578233 201242 578299 201245
rect 576380 201240 578299 201242
rect 576380 201184 578238 201240
rect 578294 201184 578299 201240
rect 576380 201182 578299 201184
rect 578233 201179 578299 201182
rect 666829 200834 666895 200837
rect 666356 200832 666895 200834
rect 666356 200776 666834 200832
rect 666890 200776 666895 200832
rect 666356 200774 666895 200776
rect 666829 200771 666895 200774
rect 603165 200426 603231 200429
rect 603165 200424 606556 200426
rect 603165 200368 603170 200424
rect 603226 200368 606556 200424
rect 603165 200366 606556 200368
rect 603165 200363 603231 200366
rect 578417 199746 578483 199749
rect 576380 199744 578483 199746
rect 576380 199688 578422 199744
rect 578478 199688 578483 199744
rect 576380 199686 578483 199688
rect 578417 199683 578483 199686
rect 31017 199474 31083 199477
rect 41638 199474 41644 199476
rect 31017 199472 41644 199474
rect 31017 199416 31022 199472
rect 31078 199416 41644 199472
rect 31017 199414 41644 199416
rect 31017 199411 31083 199414
rect 41638 199412 41644 199414
rect 41708 199412 41714 199476
rect 31201 199338 31267 199341
rect 41822 199338 41828 199340
rect 31201 199336 41828 199338
rect 31201 199280 31206 199336
rect 31262 199280 41828 199336
rect 31201 199278 41828 199280
rect 31201 199275 31267 199278
rect 41822 199276 41828 199278
rect 41892 199276 41898 199340
rect 603073 199338 603139 199341
rect 603073 199336 606556 199338
rect 603073 199280 603078 199336
rect 603134 199280 606556 199336
rect 603073 199278 606556 199280
rect 603073 199275 603139 199278
rect 666737 199066 666803 199069
rect 667933 199066 667999 199069
rect 666356 199064 667999 199066
rect 666356 199008 666742 199064
rect 666798 199008 667938 199064
rect 667994 199008 667999 199064
rect 666356 199006 667999 199008
rect 666737 199003 666803 199006
rect 667933 199003 667999 199006
rect 603073 198386 603139 198389
rect 675477 198388 675543 198389
rect 603073 198384 606556 198386
rect 603073 198328 603078 198384
rect 603134 198328 606556 198384
rect 603073 198326 606556 198328
rect 675477 198384 675524 198388
rect 675588 198386 675594 198388
rect 675477 198328 675482 198384
rect 603073 198323 603139 198326
rect 675477 198324 675524 198328
rect 675588 198326 675634 198386
rect 675588 198324 675594 198326
rect 675477 198323 675543 198324
rect 579061 198250 579127 198253
rect 576380 198248 579127 198250
rect 576380 198192 579066 198248
rect 579122 198192 579127 198248
rect 576380 198190 579127 198192
rect 579061 198187 579127 198190
rect 39297 197706 39363 197709
rect 39297 197704 41890 197706
rect 39297 197648 39302 197704
rect 39358 197648 41890 197704
rect 39297 197646 41890 197648
rect 39297 197643 39363 197646
rect 41830 197165 41890 197646
rect 603073 197298 603139 197301
rect 603073 197296 606556 197298
rect 603073 197240 603078 197296
rect 603134 197240 606556 197296
rect 603073 197238 606556 197240
rect 603073 197235 603139 197238
rect 41830 197160 41939 197165
rect 41830 197104 41878 197160
rect 41934 197104 41939 197160
rect 41830 197102 41939 197104
rect 41873 197099 41939 197102
rect 579521 196754 579587 196757
rect 576380 196752 579587 196754
rect 576380 196696 579526 196752
rect 579582 196696 579587 196752
rect 576380 196694 579587 196696
rect 579521 196691 579587 196694
rect 603165 196346 603231 196349
rect 603165 196344 606556 196346
rect 603165 196288 603170 196344
rect 603226 196288 606556 196344
rect 603165 196286 606556 196288
rect 603165 196283 603231 196286
rect 667933 195666 667999 195669
rect 666356 195664 667999 195666
rect 666356 195608 667938 195664
rect 667994 195608 667999 195664
rect 666356 195606 667999 195608
rect 667933 195603 667999 195606
rect 675753 195394 675819 195397
rect 676622 195394 676628 195396
rect 675753 195392 676628 195394
rect 675753 195336 675758 195392
rect 675814 195336 676628 195392
rect 675753 195334 676628 195336
rect 675753 195331 675819 195334
rect 676622 195332 676628 195334
rect 676692 195332 676698 195396
rect 41638 195196 41644 195260
rect 41708 195258 41714 195260
rect 41781 195258 41847 195261
rect 579521 195258 579587 195261
rect 41708 195256 41847 195258
rect 41708 195200 41786 195256
rect 41842 195200 41847 195256
rect 41708 195198 41847 195200
rect 576380 195256 579587 195258
rect 576380 195200 579526 195256
rect 579582 195200 579587 195256
rect 576380 195198 579587 195200
rect 41708 195196 41714 195198
rect 41781 195195 41847 195198
rect 579521 195195 579587 195198
rect 603073 195258 603139 195261
rect 603073 195256 606556 195258
rect 603073 195200 603078 195256
rect 603134 195200 606556 195256
rect 603073 195198 606556 195200
rect 603073 195195 603139 195198
rect 40718 194652 40724 194716
rect 40788 194714 40794 194716
rect 41822 194714 41828 194716
rect 40788 194654 41828 194714
rect 40788 194652 40794 194654
rect 41822 194652 41828 194654
rect 41892 194652 41898 194716
rect 603073 194306 603139 194309
rect 603073 194304 606556 194306
rect 603073 194248 603078 194304
rect 603134 194248 606556 194304
rect 603073 194246 606556 194248
rect 603073 194243 603139 194246
rect 666645 194034 666711 194037
rect 666356 194032 666711 194034
rect 666356 193976 666650 194032
rect 666706 193976 666711 194032
rect 666356 193974 666711 193976
rect 666645 193971 666711 193974
rect 579521 193626 579587 193629
rect 576380 193624 579587 193626
rect 576380 193568 579526 193624
rect 579582 193568 579587 193624
rect 576380 193566 579587 193568
rect 579521 193563 579587 193566
rect 603073 193218 603139 193221
rect 603073 193216 606556 193218
rect 603073 193160 603078 193216
rect 603134 193160 606556 193216
rect 603073 193158 606556 193160
rect 603073 193155 603139 193158
rect 603073 192266 603139 192269
rect 603073 192264 606556 192266
rect 603073 192208 603078 192264
rect 603134 192208 606556 192264
rect 603073 192206 606556 192208
rect 603073 192203 603139 192206
rect 579521 192130 579587 192133
rect 576380 192128 579587 192130
rect 576380 192072 579526 192128
rect 579582 192072 579587 192128
rect 576380 192070 579587 192072
rect 579521 192067 579587 192070
rect 603073 191178 603139 191181
rect 603073 191176 606556 191178
rect 603073 191120 603078 191176
rect 603134 191120 606556 191176
rect 603073 191118 606556 191120
rect 603073 191115 603139 191118
rect 579245 190634 579311 190637
rect 666645 190634 666711 190637
rect 576380 190632 579311 190634
rect 576380 190576 579250 190632
rect 579306 190576 579311 190632
rect 576380 190574 579311 190576
rect 666356 190632 666711 190634
rect 666356 190576 666650 190632
rect 666706 190576 666711 190632
rect 666356 190574 666711 190576
rect 579245 190571 579311 190574
rect 666645 190571 666711 190574
rect 675753 190362 675819 190365
rect 676254 190362 676260 190364
rect 675753 190360 676260 190362
rect 675753 190304 675758 190360
rect 675814 190304 676260 190360
rect 675753 190302 676260 190304
rect 675753 190299 675819 190302
rect 676254 190300 676260 190302
rect 676324 190300 676330 190364
rect 41454 190164 41460 190228
rect 41524 190226 41530 190228
rect 41781 190226 41847 190229
rect 41524 190224 41847 190226
rect 41524 190168 41786 190224
rect 41842 190168 41847 190224
rect 41524 190166 41847 190168
rect 41524 190164 41530 190166
rect 41781 190163 41847 190166
rect 603165 190226 603231 190229
rect 674833 190226 674899 190229
rect 676438 190226 676444 190228
rect 603165 190224 606556 190226
rect 603165 190168 603170 190224
rect 603226 190168 606556 190224
rect 603165 190166 606556 190168
rect 674833 190224 676444 190226
rect 674833 190168 674838 190224
rect 674894 190168 676444 190224
rect 674833 190166 676444 190168
rect 603165 190163 603231 190166
rect 674833 190163 674899 190166
rect 676438 190164 676444 190166
rect 676508 190164 676514 190228
rect 578233 189138 578299 189141
rect 576380 189136 578299 189138
rect 576380 189080 578238 189136
rect 578294 189080 578299 189136
rect 576380 189078 578299 189080
rect 578233 189075 578299 189078
rect 603073 189138 603139 189141
rect 603073 189136 606556 189138
rect 603073 189080 603078 189136
rect 603134 189080 606556 189136
rect 603073 189078 606556 189080
rect 603073 189075 603139 189078
rect 666553 189002 666619 189005
rect 666356 189000 666619 189002
rect 666356 188944 666558 189000
rect 666614 188944 666619 189000
rect 666356 188942 666619 188944
rect 666553 188939 666619 188942
rect 603073 188186 603139 188189
rect 603073 188184 606556 188186
rect 603073 188128 603078 188184
rect 603134 188128 606556 188184
rect 603073 188126 606556 188128
rect 603073 188123 603139 188126
rect 579245 187642 579311 187645
rect 576380 187640 579311 187642
rect 576380 187584 579250 187640
rect 579306 187584 579311 187640
rect 576380 187582 579311 187584
rect 579245 187579 579311 187582
rect 41781 187372 41847 187373
rect 41781 187368 41828 187372
rect 41892 187370 41898 187372
rect 41781 187312 41786 187368
rect 41781 187308 41828 187312
rect 41892 187310 41938 187370
rect 41892 187308 41898 187310
rect 41781 187307 41847 187308
rect 603073 187098 603139 187101
rect 603073 187096 606556 187098
rect 603073 187040 603078 187096
rect 603134 187040 606556 187096
rect 603073 187038 606556 187040
rect 603073 187035 603139 187038
rect 579521 186146 579587 186149
rect 576380 186144 579587 186146
rect 576380 186088 579526 186144
rect 579582 186088 579587 186144
rect 576380 186086 579587 186088
rect 579521 186083 579587 186086
rect 603165 186146 603231 186149
rect 603165 186144 606556 186146
rect 603165 186088 603170 186144
rect 603226 186088 606556 186144
rect 603165 186086 606556 186088
rect 603165 186083 603231 186086
rect 666553 185602 666619 185605
rect 666356 185600 666619 185602
rect 666356 185544 666558 185600
rect 666614 185544 666619 185600
rect 666356 185542 666619 185544
rect 666553 185539 666619 185542
rect 603073 185058 603139 185061
rect 603073 185056 606556 185058
rect 603073 185000 603078 185056
rect 603134 185000 606556 185056
rect 603073 184998 606556 185000
rect 603073 184995 603139 184998
rect 578785 184650 578851 184653
rect 576380 184648 578851 184650
rect 576380 184592 578790 184648
rect 578846 184592 578851 184648
rect 576380 184590 578851 184592
rect 578785 184587 578851 184590
rect 41638 184044 41644 184108
rect 41708 184106 41714 184108
rect 41781 184106 41847 184109
rect 41708 184104 41847 184106
rect 41708 184048 41786 184104
rect 41842 184048 41847 184104
rect 41708 184046 41847 184048
rect 41708 184044 41714 184046
rect 41781 184043 41847 184046
rect 603073 184106 603139 184109
rect 603073 184104 606556 184106
rect 603073 184048 603078 184104
rect 603134 184048 606556 184104
rect 603073 184046 606556 184048
rect 603073 184043 603139 184046
rect 668025 183834 668091 183837
rect 668301 183834 668367 183837
rect 666356 183832 668367 183834
rect 666356 183776 668030 183832
rect 668086 183776 668306 183832
rect 668362 183776 668367 183832
rect 666356 183774 668367 183776
rect 668025 183771 668091 183774
rect 668301 183771 668367 183774
rect 579337 183154 579403 183157
rect 576380 183152 579403 183154
rect 576380 183096 579342 183152
rect 579398 183096 579403 183152
rect 576380 183094 579403 183096
rect 579337 183091 579403 183094
rect 40534 182956 40540 183020
rect 40604 183018 40610 183020
rect 41781 183018 41847 183021
rect 40604 183016 41847 183018
rect 40604 182960 41786 183016
rect 41842 182960 41847 183016
rect 40604 182958 41847 182960
rect 40604 182956 40610 182958
rect 41781 182955 41847 182958
rect 603073 183018 603139 183021
rect 603073 183016 606556 183018
rect 603073 182960 603078 183016
rect 603134 182960 606556 183016
rect 603073 182958 606556 182960
rect 603073 182955 603139 182958
rect 603165 182066 603231 182069
rect 603165 182064 606556 182066
rect 603165 182008 603170 182064
rect 603226 182008 606556 182064
rect 603165 182006 606556 182008
rect 603165 182003 603231 182006
rect 579061 181658 579127 181661
rect 576380 181656 579127 181658
rect 576380 181600 579066 181656
rect 579122 181600 579127 181656
rect 576380 181598 579127 181600
rect 579061 181595 579127 181598
rect 603073 180978 603139 180981
rect 603073 180976 606556 180978
rect 603073 180920 603078 180976
rect 603134 180920 606556 180976
rect 603073 180918 606556 180920
rect 603073 180915 603139 180918
rect 668025 180434 668091 180437
rect 666356 180432 668091 180434
rect 666356 180376 668030 180432
rect 668086 180376 668091 180432
rect 666356 180374 668091 180376
rect 668025 180371 668091 180374
rect 578969 180162 579035 180165
rect 576380 180160 579035 180162
rect 576380 180104 578974 180160
rect 579030 180104 579035 180160
rect 576380 180102 579035 180104
rect 578969 180099 579035 180102
rect 603073 180026 603139 180029
rect 603073 180024 606556 180026
rect 603073 179968 603078 180024
rect 603134 179968 606556 180024
rect 603073 179966 606556 179968
rect 603073 179963 603139 179966
rect 603073 178938 603139 178941
rect 603073 178936 606556 178938
rect 603073 178880 603078 178936
rect 603134 178880 606556 178936
rect 603073 178878 606556 178880
rect 603073 178875 603139 178878
rect 667933 178802 667999 178805
rect 666356 178800 667999 178802
rect 666356 178744 667938 178800
rect 667994 178744 667999 178800
rect 666356 178742 667999 178744
rect 667933 178739 667999 178742
rect 579245 178666 579311 178669
rect 576380 178664 579311 178666
rect 576380 178608 579250 178664
rect 579306 178608 579311 178664
rect 576380 178606 579311 178608
rect 579245 178603 579311 178606
rect 676029 178530 676095 178533
rect 676029 178528 676292 178530
rect 676029 178472 676034 178528
rect 676090 178472 676292 178528
rect 676029 178470 676292 178472
rect 676029 178467 676095 178470
rect 676029 178122 676095 178125
rect 676029 178120 676292 178122
rect 676029 178064 676034 178120
rect 676090 178064 676292 178120
rect 676029 178062 676292 178064
rect 676029 178059 676095 178062
rect 603165 177986 603231 177989
rect 603165 177984 606556 177986
rect 603165 177928 603170 177984
rect 603226 177928 606556 177984
rect 603165 177926 606556 177928
rect 603165 177923 603231 177926
rect 675937 177714 676003 177717
rect 675937 177712 676292 177714
rect 675937 177656 675942 177712
rect 675998 177656 676292 177712
rect 675937 177654 676292 177656
rect 675937 177651 676003 177654
rect 676029 177306 676095 177309
rect 676029 177304 676292 177306
rect 676029 177248 676034 177304
rect 676090 177248 676292 177304
rect 676029 177246 676292 177248
rect 676029 177243 676095 177246
rect 578233 177170 578299 177173
rect 576380 177168 578299 177170
rect 576380 177112 578238 177168
rect 578294 177112 578299 177168
rect 576380 177110 578299 177112
rect 578233 177107 578299 177110
rect 603073 176898 603139 176901
rect 676029 176898 676095 176901
rect 603073 176896 606556 176898
rect 603073 176840 603078 176896
rect 603134 176840 606556 176896
rect 603073 176838 606556 176840
rect 676029 176896 676292 176898
rect 676029 176840 676034 176896
rect 676090 176840 676292 176896
rect 676029 176838 676292 176840
rect 603073 176835 603139 176838
rect 676029 176835 676095 176838
rect 676029 176490 676095 176493
rect 676029 176488 676292 176490
rect 676029 176432 676034 176488
rect 676090 176432 676292 176488
rect 676029 176430 676292 176432
rect 676029 176427 676095 176430
rect 676029 176082 676095 176085
rect 676029 176080 676292 176082
rect 676029 176024 676034 176080
rect 676090 176024 676292 176080
rect 676029 176022 676292 176024
rect 676029 176019 676095 176022
rect 603073 175946 603139 175949
rect 603073 175944 606556 175946
rect 603073 175888 603078 175944
rect 603134 175888 606556 175944
rect 603073 175886 606556 175888
rect 603073 175883 603139 175886
rect 578325 175674 578391 175677
rect 576380 175672 578391 175674
rect 576380 175616 578330 175672
rect 578386 175616 578391 175672
rect 576380 175614 578391 175616
rect 578325 175611 578391 175614
rect 676029 175674 676095 175677
rect 676029 175672 676292 175674
rect 676029 175616 676034 175672
rect 676090 175616 676292 175672
rect 676029 175614 676292 175616
rect 676029 175611 676095 175614
rect 667933 175402 667999 175405
rect 666356 175400 667999 175402
rect 666356 175344 667938 175400
rect 667994 175344 667999 175400
rect 666356 175342 667999 175344
rect 667933 175339 667999 175342
rect 676029 175266 676095 175269
rect 676029 175264 676292 175266
rect 676029 175208 676034 175264
rect 676090 175208 676292 175264
rect 676029 175206 676292 175208
rect 676029 175203 676095 175206
rect 603073 174858 603139 174861
rect 674741 174858 674807 174861
rect 603073 174856 606556 174858
rect 603073 174800 603078 174856
rect 603134 174800 606556 174856
rect 603073 174798 606556 174800
rect 674741 174856 676292 174858
rect 674741 174800 674746 174856
rect 674802 174800 676292 174856
rect 674741 174798 676292 174800
rect 603073 174795 603139 174798
rect 674741 174795 674807 174798
rect 676029 174450 676095 174453
rect 676029 174448 676292 174450
rect 676029 174392 676034 174448
rect 676090 174392 676292 174448
rect 676029 174390 676292 174392
rect 676029 174387 676095 174390
rect 578417 174178 578483 174181
rect 576380 174176 578483 174178
rect 576380 174120 578422 174176
rect 578478 174120 578483 174176
rect 576380 174118 578483 174120
rect 578417 174115 578483 174118
rect 678237 174042 678303 174045
rect 678237 174040 678316 174042
rect 678237 173984 678242 174040
rect 678298 173984 678316 174040
rect 678237 173982 678316 173984
rect 678237 173979 678303 173982
rect 603717 173906 603783 173909
rect 603717 173904 606556 173906
rect 603717 173848 603722 173904
rect 603778 173848 606556 173904
rect 603717 173846 606556 173848
rect 603717 173843 603783 173846
rect 667933 173634 667999 173637
rect 666356 173632 667999 173634
rect 666356 173576 667938 173632
rect 667994 173576 667999 173632
rect 666356 173574 667999 173576
rect 667933 173571 667999 173574
rect 676078 173574 676292 173634
rect 676078 173500 676138 173574
rect 676070 173436 676076 173500
rect 676140 173436 676146 173500
rect 676029 173226 676095 173229
rect 676029 173224 676292 173226
rect 676029 173168 676034 173224
rect 676090 173168 676292 173224
rect 676029 173166 676292 173168
rect 676029 173163 676095 173166
rect 603073 172818 603139 172821
rect 603073 172816 606556 172818
rect 603073 172760 603078 172816
rect 603134 172760 606556 172816
rect 603073 172758 606556 172760
rect 603073 172755 603139 172758
rect 675886 172756 675892 172820
rect 675956 172818 675962 172820
rect 675956 172758 676292 172818
rect 675956 172756 675962 172758
rect 578785 172682 578851 172685
rect 576380 172680 578851 172682
rect 576380 172624 578790 172680
rect 578846 172624 578851 172680
rect 576380 172622 578851 172624
rect 578785 172619 578851 172622
rect 680997 172410 681063 172413
rect 680997 172408 681076 172410
rect 680997 172352 681002 172408
rect 681058 172352 681076 172408
rect 680997 172350 681076 172352
rect 680997 172347 681063 172350
rect 676078 171942 676292 172002
rect 603073 171866 603139 171869
rect 676078 171868 676138 171942
rect 603073 171864 606556 171866
rect 603073 171808 603078 171864
rect 603134 171808 606556 171864
rect 603073 171806 606556 171808
rect 603073 171803 603139 171806
rect 676070 171804 676076 171868
rect 676140 171804 676146 171868
rect 676857 171594 676923 171597
rect 676844 171592 676923 171594
rect 676844 171536 676862 171592
rect 676918 171536 676923 171592
rect 676844 171534 676923 171536
rect 676857 171531 676923 171534
rect 578693 171186 578759 171189
rect 667933 171186 667999 171189
rect 576380 171184 578759 171186
rect 576380 171128 578698 171184
rect 578754 171128 578759 171184
rect 576380 171126 578759 171128
rect 578693 171123 578759 171126
rect 666510 171184 667999 171186
rect 666510 171128 667938 171184
rect 667994 171128 667999 171184
rect 666510 171126 667999 171128
rect 603165 170778 603231 170781
rect 603165 170776 606556 170778
rect 603165 170720 603170 170776
rect 603226 170720 606556 170776
rect 603165 170718 606556 170720
rect 603165 170715 603231 170718
rect 666510 170506 666570 171126
rect 667933 171123 667999 171126
rect 678421 171186 678487 171189
rect 678421 171184 678500 171186
rect 678421 171128 678426 171184
rect 678482 171128 678500 171184
rect 678421 171126 678500 171128
rect 678421 171123 678487 171126
rect 676029 170778 676095 170781
rect 676029 170776 676292 170778
rect 676029 170720 676034 170776
rect 676090 170720 676292 170776
rect 676029 170718 676292 170720
rect 676029 170715 676095 170718
rect 666510 170446 666754 170506
rect 666694 170234 666754 170446
rect 676029 170370 676095 170373
rect 676029 170368 676292 170370
rect 676029 170312 676034 170368
rect 676090 170312 676292 170368
rect 676029 170310 676292 170312
rect 676029 170307 676095 170310
rect 666356 170174 666754 170234
rect 676581 169962 676647 169965
rect 676581 169960 676660 169962
rect 676581 169904 676586 169960
rect 676642 169904 676660 169960
rect 676581 169902 676660 169904
rect 676581 169899 676647 169902
rect 603073 169826 603139 169829
rect 603073 169824 606556 169826
rect 603073 169768 603078 169824
rect 603134 169768 606556 169824
rect 603073 169766 606556 169768
rect 603073 169763 603139 169766
rect 579429 169554 579495 169557
rect 576380 169552 579495 169554
rect 576380 169496 579434 169552
rect 579490 169496 579495 169552
rect 576380 169494 579495 169496
rect 579429 169491 579495 169494
rect 676029 169554 676095 169557
rect 676029 169552 676292 169554
rect 676029 169496 676034 169552
rect 676090 169496 676292 169552
rect 676029 169494 676292 169496
rect 676029 169491 676095 169494
rect 676029 169146 676095 169149
rect 676029 169144 676292 169146
rect 676029 169088 676034 169144
rect 676090 169088 676292 169144
rect 676029 169086 676292 169088
rect 676029 169083 676095 169086
rect 603073 168738 603139 168741
rect 676029 168738 676095 168741
rect 603073 168736 606556 168738
rect 603073 168680 603078 168736
rect 603134 168680 606556 168736
rect 603073 168678 606556 168680
rect 676029 168736 676292 168738
rect 676029 168680 676034 168736
rect 676090 168680 676292 168736
rect 676029 168678 676292 168680
rect 603073 168675 603139 168678
rect 676029 168675 676095 168678
rect 667933 168602 667999 168605
rect 673862 168602 673868 168604
rect 666356 168600 673868 168602
rect 666356 168544 667938 168600
rect 667994 168544 673868 168600
rect 666356 168542 673868 168544
rect 667933 168539 667999 168542
rect 673862 168540 673868 168542
rect 673932 168540 673938 168604
rect 676029 168330 676095 168333
rect 676029 168328 676292 168330
rect 676029 168272 676034 168328
rect 676090 168272 676292 168328
rect 676029 168270 676292 168272
rect 676029 168267 676095 168270
rect 579245 168058 579311 168061
rect 576380 168056 579311 168058
rect 576380 168000 579250 168056
rect 579306 168000 579311 168056
rect 576380 167998 579311 168000
rect 579245 167995 579311 167998
rect 676029 167922 676095 167925
rect 676029 167920 676292 167922
rect 676029 167864 676034 167920
rect 676090 167864 676292 167920
rect 676029 167862 676292 167864
rect 676029 167859 676095 167862
rect 603073 167786 603139 167789
rect 603073 167784 606556 167786
rect 603073 167728 603078 167784
rect 603134 167728 606556 167784
rect 603073 167726 606556 167728
rect 603073 167723 603139 167726
rect 676029 167106 676095 167109
rect 676029 167104 676292 167106
rect 676029 167048 676034 167104
rect 676090 167048 676292 167104
rect 676029 167046 676292 167048
rect 676029 167043 676095 167046
rect 603073 166698 603139 166701
rect 603073 166696 606556 166698
rect 603073 166640 603078 166696
rect 603134 166640 606556 166696
rect 603073 166638 606556 166640
rect 603073 166635 603139 166638
rect 578693 166562 578759 166565
rect 576380 166560 578759 166562
rect 576380 166504 578698 166560
rect 578754 166504 578759 166560
rect 576380 166502 578759 166504
rect 578693 166499 578759 166502
rect 676581 166428 676647 166429
rect 676857 166428 676923 166429
rect 676581 166424 676628 166428
rect 676692 166426 676698 166428
rect 676581 166368 676586 166424
rect 676581 166364 676628 166368
rect 676692 166366 676738 166426
rect 676692 166364 676698 166366
rect 676806 166364 676812 166428
rect 676876 166426 676923 166428
rect 676876 166424 676968 166426
rect 676918 166368 676968 166424
rect 676876 166366 676968 166368
rect 676876 166364 676923 166366
rect 676581 166363 676647 166364
rect 676857 166363 676923 166364
rect 603809 165746 603875 165749
rect 603809 165744 606556 165746
rect 603809 165688 603814 165744
rect 603870 165688 606556 165744
rect 603809 165686 606556 165688
rect 603809 165683 603875 165686
rect 667933 165202 667999 165205
rect 666356 165200 667999 165202
rect 666356 165144 667938 165200
rect 667994 165144 667999 165200
rect 666356 165142 667999 165144
rect 667933 165139 667999 165142
rect 576350 164386 576410 165036
rect 603073 164658 603139 164661
rect 603073 164656 606556 164658
rect 603073 164600 603078 164656
rect 603134 164600 606556 164656
rect 603073 164598 606556 164600
rect 603073 164595 603139 164598
rect 578233 164386 578299 164389
rect 576350 164384 578299 164386
rect 576350 164328 578238 164384
rect 578294 164328 578299 164384
rect 576350 164326 578299 164328
rect 578233 164323 578299 164326
rect 603073 163706 603139 163709
rect 603073 163704 606556 163706
rect 603073 163648 603078 163704
rect 603134 163648 606556 163704
rect 603073 163646 606556 163648
rect 603073 163643 603139 163646
rect 579521 163570 579587 163573
rect 666553 163570 666619 163573
rect 668393 163570 668459 163573
rect 576380 163568 579587 163570
rect 576380 163512 579526 163568
rect 579582 163512 579587 163568
rect 576380 163510 579587 163512
rect 666356 163568 668459 163570
rect 666356 163512 666558 163568
rect 666614 163512 668398 163568
rect 668454 163512 668459 163568
rect 666356 163510 668459 163512
rect 579521 163507 579587 163510
rect 666553 163507 666619 163510
rect 668393 163507 668459 163510
rect 675518 162692 675524 162756
rect 675588 162754 675594 162756
rect 676213 162754 676279 162757
rect 675588 162752 676279 162754
rect 675588 162696 676218 162752
rect 676274 162696 676279 162752
rect 675588 162694 676279 162696
rect 675588 162692 675594 162694
rect 676213 162691 676279 162694
rect 603073 162618 603139 162621
rect 603073 162616 606556 162618
rect 603073 162560 603078 162616
rect 603134 162560 606556 162616
rect 603073 162558 606556 162560
rect 603073 162555 603139 162558
rect 675886 162556 675892 162620
rect 675956 162618 675962 162620
rect 678237 162618 678303 162621
rect 675956 162616 678303 162618
rect 675956 162560 678242 162616
rect 678298 162560 678303 162616
rect 675956 162558 678303 162560
rect 675956 162556 675962 162558
rect 678237 162555 678303 162558
rect 675702 162420 675708 162484
rect 675772 162482 675778 162484
rect 678421 162482 678487 162485
rect 675772 162480 678487 162482
rect 675772 162424 678426 162480
rect 678482 162424 678487 162480
rect 675772 162422 678487 162424
rect 675772 162420 675778 162422
rect 678421 162419 678487 162422
rect 675334 162284 675340 162348
rect 675404 162346 675410 162348
rect 680997 162346 681063 162349
rect 675404 162344 681063 162346
rect 675404 162288 681002 162344
rect 681058 162288 681063 162344
rect 675404 162286 681063 162288
rect 675404 162284 675410 162286
rect 680997 162283 681063 162286
rect 579153 162074 579219 162077
rect 576380 162072 579219 162074
rect 576380 162016 579158 162072
rect 579214 162016 579219 162072
rect 576380 162014 579219 162016
rect 579153 162011 579219 162014
rect 603717 161666 603783 161669
rect 603717 161664 606556 161666
rect 603717 161608 603722 161664
rect 603778 161608 606556 161664
rect 603717 161606 606556 161608
rect 603717 161603 603783 161606
rect 666553 161530 666619 161533
rect 666510 161528 666619 161530
rect 666510 161472 666558 161528
rect 666614 161472 666619 161528
rect 666510 161467 666619 161472
rect 579337 160578 579403 160581
rect 576380 160576 579403 160578
rect 576380 160520 579342 160576
rect 579398 160520 579403 160576
rect 576380 160518 579403 160520
rect 579337 160515 579403 160518
rect 603073 160578 603139 160581
rect 603073 160576 606556 160578
rect 603073 160520 603078 160576
rect 603134 160520 606556 160576
rect 603073 160518 606556 160520
rect 603073 160515 603139 160518
rect 666510 160442 666570 161467
rect 666510 160382 666754 160442
rect 666694 160170 666754 160382
rect 666356 160110 666754 160170
rect 675753 160034 675819 160037
rect 676806 160034 676812 160036
rect 675753 160032 676812 160034
rect 675753 159976 675758 160032
rect 675814 159976 676812 160032
rect 675753 159974 676812 159976
rect 675753 159971 675819 159974
rect 676806 159972 676812 159974
rect 676876 159972 676882 160036
rect 603073 159626 603139 159629
rect 603073 159624 606556 159626
rect 603073 159568 603078 159624
rect 603134 159568 606556 159624
rect 603073 159566 606556 159568
rect 603073 159563 603139 159566
rect 675753 159490 675819 159493
rect 675886 159490 675892 159492
rect 675753 159488 675892 159490
rect 675753 159432 675758 159488
rect 675814 159432 675892 159488
rect 675753 159430 675892 159432
rect 675753 159427 675819 159430
rect 675886 159428 675892 159430
rect 675956 159428 675962 159492
rect 579061 159082 579127 159085
rect 576380 159080 579127 159082
rect 576380 159024 579066 159080
rect 579122 159024 579127 159080
rect 576380 159022 579127 159024
rect 579061 159019 579127 159022
rect 603165 158538 603231 158541
rect 603165 158536 606556 158538
rect 603165 158480 603170 158536
rect 603226 158480 606556 158536
rect 603165 158478 606556 158480
rect 603165 158475 603231 158478
rect 667933 158402 667999 158405
rect 668577 158402 668643 158405
rect 666356 158400 668643 158402
rect 666356 158344 667938 158400
rect 667994 158344 668582 158400
rect 668638 158344 668643 158400
rect 666356 158342 668643 158344
rect 667933 158339 667999 158342
rect 668577 158339 668643 158342
rect 578969 157586 579035 157589
rect 576380 157584 579035 157586
rect 576380 157528 578974 157584
rect 579030 157528 579035 157584
rect 576380 157526 579035 157528
rect 578969 157523 579035 157526
rect 603073 157586 603139 157589
rect 603073 157584 606556 157586
rect 603073 157528 603078 157584
rect 603134 157528 606556 157584
rect 603073 157526 606556 157528
rect 603073 157523 603139 157526
rect 675753 157450 675819 157453
rect 676070 157450 676076 157452
rect 675753 157448 676076 157450
rect 675753 157392 675758 157448
rect 675814 157392 676076 157448
rect 675753 157390 676076 157392
rect 675753 157387 675819 157390
rect 676070 157388 676076 157390
rect 676140 157388 676146 157452
rect 675661 157044 675727 157045
rect 675661 157040 675708 157044
rect 675772 157042 675778 157044
rect 675661 156984 675666 157040
rect 675661 156980 675708 156984
rect 675772 156982 675818 157042
rect 675772 156980 675778 156982
rect 675661 156979 675727 156980
rect 603073 156498 603139 156501
rect 675569 156500 675635 156501
rect 675518 156498 675524 156500
rect 603073 156496 606556 156498
rect 603073 156440 603078 156496
rect 603134 156440 606556 156496
rect 603073 156438 606556 156440
rect 675478 156438 675524 156498
rect 675588 156496 675635 156500
rect 675630 156440 675635 156496
rect 603073 156435 603139 156438
rect 675518 156436 675524 156438
rect 675588 156436 675635 156440
rect 675569 156435 675635 156436
rect 578877 156090 578943 156093
rect 576380 156088 578943 156090
rect 576380 156032 578882 156088
rect 578938 156032 578943 156088
rect 576380 156030 578943 156032
rect 578877 156027 578943 156030
rect 603073 155546 603139 155549
rect 603073 155544 606556 155546
rect 603073 155488 603078 155544
rect 603134 155488 606556 155544
rect 603073 155486 606556 155488
rect 603073 155483 603139 155486
rect 667933 155002 667999 155005
rect 666356 155000 667999 155002
rect 666356 154944 667938 155000
rect 667994 154944 667999 155000
rect 666356 154942 667999 154944
rect 667933 154939 667999 154942
rect 578509 154594 578575 154597
rect 576380 154592 578575 154594
rect 576380 154536 578514 154592
rect 578570 154536 578575 154592
rect 576380 154534 578575 154536
rect 578509 154531 578575 154534
rect 603165 154458 603231 154461
rect 603165 154456 606556 154458
rect 603165 154400 603170 154456
rect 603226 154400 606556 154456
rect 603165 154398 606556 154400
rect 603165 154395 603231 154398
rect 603073 153506 603139 153509
rect 603073 153504 606556 153506
rect 603073 153448 603078 153504
rect 603134 153448 606556 153504
rect 603073 153446 606556 153448
rect 603073 153443 603139 153446
rect 666553 153370 666619 153373
rect 668669 153370 668735 153373
rect 666356 153368 668735 153370
rect 666356 153312 666558 153368
rect 666614 153312 668674 153368
rect 668730 153312 668735 153368
rect 666356 153310 668735 153312
rect 666553 153307 666619 153310
rect 668669 153307 668735 153310
rect 579245 153098 579311 153101
rect 675385 153100 675451 153101
rect 675334 153098 675340 153100
rect 576380 153096 579311 153098
rect 576380 153040 579250 153096
rect 579306 153040 579311 153096
rect 576380 153038 579311 153040
rect 675294 153038 675340 153098
rect 675404 153096 675451 153100
rect 675446 153040 675451 153096
rect 579245 153035 579311 153038
rect 675334 153036 675340 153038
rect 675404 153036 675451 153040
rect 675385 153035 675451 153036
rect 603073 152418 603139 152421
rect 603073 152416 606556 152418
rect 603073 152360 603078 152416
rect 603134 152360 606556 152416
rect 603073 152358 606556 152360
rect 603073 152355 603139 152358
rect 666553 151874 666619 151877
rect 666510 151872 666619 151874
rect 666510 151816 666558 151872
rect 666614 151816 666619 151872
rect 666510 151811 666619 151816
rect 666510 151770 666616 151811
rect 666556 151605 666616 151770
rect 579521 151602 579587 151605
rect 576380 151600 579587 151602
rect 576380 151544 579526 151600
rect 579582 151544 579587 151600
rect 576380 151542 579587 151544
rect 579521 151539 579587 151542
rect 666553 151600 666619 151605
rect 666553 151544 666558 151600
rect 666614 151544 666619 151600
rect 666553 151539 666619 151544
rect 675753 151602 675819 151605
rect 676622 151602 676628 151604
rect 675753 151600 676628 151602
rect 675753 151544 675758 151600
rect 675814 151544 676628 151600
rect 675753 151542 676628 151544
rect 675753 151539 675819 151542
rect 676622 151540 676628 151542
rect 676692 151540 676698 151604
rect 603073 151466 603139 151469
rect 603073 151464 606556 151466
rect 603073 151408 603078 151464
rect 603134 151408 606556 151464
rect 603073 151406 606556 151408
rect 603073 151403 603139 151406
rect 603165 150378 603231 150381
rect 603165 150376 606556 150378
rect 603165 150320 603170 150376
rect 603226 150320 606556 150376
rect 603165 150318 606556 150320
rect 603165 150315 603231 150318
rect 579429 150106 579495 150109
rect 576380 150104 579495 150106
rect 576380 150048 579434 150104
rect 579490 150048 579495 150104
rect 576380 150046 579495 150048
rect 579429 150043 579495 150046
rect 666553 149970 666619 149973
rect 666356 149968 666619 149970
rect 666356 149912 666558 149968
rect 666614 149912 666619 149968
rect 666356 149910 666619 149912
rect 666553 149907 666619 149910
rect 603073 149426 603139 149429
rect 603073 149424 606556 149426
rect 603073 149368 603078 149424
rect 603134 149368 606556 149424
rect 603073 149366 606556 149368
rect 603073 149363 603139 149366
rect 578509 148610 578575 148613
rect 576380 148608 578575 148610
rect 576380 148552 578514 148608
rect 578570 148552 578575 148608
rect 576380 148550 578575 148552
rect 578509 148547 578575 148550
rect 675753 148474 675819 148477
rect 676438 148474 676444 148476
rect 675753 148472 676444 148474
rect 675753 148416 675758 148472
rect 675814 148416 676444 148472
rect 675753 148414 676444 148416
rect 675753 148411 675819 148414
rect 676438 148412 676444 148414
rect 676508 148412 676514 148476
rect 603073 148338 603139 148341
rect 603073 148336 606556 148338
rect 603073 148280 603078 148336
rect 603134 148280 606556 148336
rect 603073 148278 606556 148280
rect 603073 148275 603139 148278
rect 668301 148202 668367 148205
rect 666356 148200 668367 148202
rect 666356 148144 668306 148200
rect 668362 148144 668367 148200
rect 666356 148142 668367 148144
rect 668301 148139 668367 148142
rect 603073 147386 603139 147389
rect 603073 147384 606556 147386
rect 603073 147328 603078 147384
rect 603134 147328 606556 147384
rect 603073 147326 606556 147328
rect 603073 147323 603139 147326
rect 578509 146978 578575 146981
rect 576380 146976 578575 146978
rect 576380 146920 578514 146976
rect 578570 146920 578575 146976
rect 576380 146918 578575 146920
rect 578509 146915 578575 146918
rect 603165 146298 603231 146301
rect 675753 146298 675819 146301
rect 676254 146298 676260 146300
rect 603165 146296 606556 146298
rect 603165 146240 603170 146296
rect 603226 146240 606556 146296
rect 603165 146238 606556 146240
rect 675753 146296 676260 146298
rect 675753 146240 675758 146296
rect 675814 146240 676260 146296
rect 675753 146238 676260 146240
rect 603165 146235 603231 146238
rect 675753 146235 675819 146238
rect 676254 146236 676260 146238
rect 676324 146236 676330 146300
rect 579521 145482 579587 145485
rect 576380 145480 579587 145482
rect 576380 145424 579526 145480
rect 579582 145424 579587 145480
rect 576380 145422 579587 145424
rect 579521 145419 579587 145422
rect 603901 145346 603967 145349
rect 603901 145344 606556 145346
rect 603901 145288 603906 145344
rect 603962 145288 606556 145344
rect 603901 145286 606556 145288
rect 603901 145283 603967 145286
rect 668301 144938 668367 144941
rect 666356 144936 668367 144938
rect 666356 144880 668306 144936
rect 668362 144880 668367 144936
rect 666356 144878 668367 144880
rect 668301 144875 668367 144878
rect 603073 144258 603139 144261
rect 603073 144256 606556 144258
rect 603073 144200 603078 144256
rect 603134 144200 606556 144256
rect 603073 144198 606556 144200
rect 603073 144195 603139 144198
rect 578601 143986 578667 143989
rect 576380 143984 578667 143986
rect 576380 143928 578606 143984
rect 578662 143928 578667 143984
rect 576380 143926 578667 143928
rect 578601 143923 578667 143926
rect 603717 143306 603783 143309
rect 603717 143304 606556 143306
rect 603717 143248 603722 143304
rect 603778 143248 606556 143304
rect 603717 143246 606556 143248
rect 603717 143243 603783 143246
rect 667933 143170 667999 143173
rect 666356 143168 667999 143170
rect 666356 143112 667938 143168
rect 667994 143112 667999 143168
rect 666356 143110 667999 143112
rect 579521 142490 579587 142493
rect 576380 142488 579587 142490
rect 576380 142432 579526 142488
rect 579582 142432 579587 142488
rect 576380 142430 579587 142432
rect 579521 142427 579587 142430
rect 603073 142218 603139 142221
rect 603073 142216 606556 142218
rect 603073 142160 603078 142216
rect 603134 142160 606556 142216
rect 603073 142158 606556 142160
rect 603073 142155 603139 142158
rect 666510 142085 666570 143110
rect 667933 143107 667999 143110
rect 666510 142080 666619 142085
rect 666510 142024 666558 142080
rect 666614 142024 666619 142080
rect 666510 142022 666619 142024
rect 666553 142019 666619 142022
rect 603073 141266 603139 141269
rect 603073 141264 606556 141266
rect 603073 141208 603078 141264
rect 603134 141208 606556 141264
rect 603073 141206 606556 141208
rect 603073 141203 603139 141206
rect 579337 140994 579403 140997
rect 576380 140992 579403 140994
rect 576380 140936 579342 140992
rect 579398 140936 579403 140992
rect 576380 140934 579403 140936
rect 579337 140931 579403 140934
rect 603073 140178 603139 140181
rect 603073 140176 606556 140178
rect 603073 140120 603078 140176
rect 603134 140120 606556 140176
rect 603073 140118 606556 140120
rect 603073 140115 603139 140118
rect 666553 139770 666619 139773
rect 666356 139768 666619 139770
rect 666356 139712 666558 139768
rect 666614 139712 666619 139768
rect 666356 139710 666619 139712
rect 666553 139707 666619 139710
rect 579245 139498 579311 139501
rect 576380 139496 579311 139498
rect 576380 139440 579250 139496
rect 579306 139440 579311 139496
rect 576380 139438 579311 139440
rect 579245 139435 579311 139438
rect 603165 139226 603231 139229
rect 603165 139224 606556 139226
rect 603165 139168 603170 139224
rect 603226 139168 606556 139224
rect 603165 139166 606556 139168
rect 603165 139163 603231 139166
rect 603073 138138 603139 138141
rect 668025 138138 668091 138141
rect 603073 138136 606556 138138
rect 603073 138080 603078 138136
rect 603134 138080 606556 138136
rect 603073 138078 606556 138080
rect 666356 138136 668091 138138
rect 666356 138080 668030 138136
rect 668086 138080 668091 138136
rect 666356 138078 668091 138080
rect 603073 138075 603139 138078
rect 668025 138075 668091 138078
rect 579521 138002 579587 138005
rect 576380 138000 579587 138002
rect 576380 137944 579526 138000
rect 579582 137944 579587 138000
rect 576380 137942 579587 137944
rect 579521 137939 579587 137942
rect 603073 137186 603139 137189
rect 603073 137184 606556 137186
rect 603073 137128 603078 137184
rect 603134 137128 606556 137184
rect 603073 137126 606556 137128
rect 603073 137123 603139 137126
rect 579521 136506 579587 136509
rect 576380 136504 579587 136506
rect 576380 136448 579526 136504
rect 579582 136448 579587 136504
rect 576380 136446 579587 136448
rect 579521 136443 579587 136446
rect 603073 136098 603139 136101
rect 603073 136096 606556 136098
rect 603073 136040 603078 136096
rect 603134 136040 606556 136096
rect 603073 136038 606556 136040
rect 603073 136035 603139 136038
rect 603165 135146 603231 135149
rect 603165 135144 606556 135146
rect 603165 135088 603170 135144
rect 603226 135088 606556 135144
rect 603165 135086 606556 135088
rect 603165 135083 603231 135086
rect 579153 135010 579219 135013
rect 576380 135008 579219 135010
rect 576380 134952 579158 135008
rect 579214 134952 579219 135008
rect 576380 134950 579219 134952
rect 579153 134947 579219 134950
rect 668025 134738 668091 134741
rect 666356 134736 668091 134738
rect 666356 134680 668030 134736
rect 668086 134680 668091 134736
rect 666356 134678 668091 134680
rect 668025 134675 668091 134678
rect 603073 134058 603139 134061
rect 603073 134056 606556 134058
rect 603073 134000 603078 134056
rect 603134 134000 606556 134056
rect 603073 133998 606556 134000
rect 603073 133995 603139 133998
rect 579061 133514 579127 133517
rect 576380 133512 579127 133514
rect 576380 133456 579066 133512
rect 579122 133456 579127 133512
rect 576380 133454 579127 133456
rect 579061 133451 579127 133454
rect 603073 133106 603139 133109
rect 676121 133106 676187 133109
rect 676262 133106 676322 133348
rect 603073 133104 606556 133106
rect 603073 133048 603078 133104
rect 603134 133048 606556 133104
rect 603073 133046 606556 133048
rect 676121 133104 676322 133106
rect 676121 133048 676126 133104
rect 676182 133048 676322 133104
rect 676121 133046 676322 133048
rect 603073 133043 603139 133046
rect 676121 133043 676187 133046
rect 668577 132970 668643 132973
rect 666356 132968 668643 132970
rect 666356 132912 668582 132968
rect 668638 132912 668643 132968
rect 666356 132910 668643 132912
rect 666510 132429 666570 132910
rect 668577 132907 668643 132910
rect 676029 132970 676095 132973
rect 676029 132968 676292 132970
rect 676029 132912 676034 132968
rect 676090 132912 676292 132968
rect 676029 132910 676292 132912
rect 676029 132907 676095 132910
rect 676213 132698 676279 132701
rect 676213 132696 676322 132698
rect 676213 132640 676218 132696
rect 676274 132640 676322 132696
rect 676213 132635 676322 132640
rect 676262 132532 676322 132635
rect 666510 132424 666619 132429
rect 666510 132368 666558 132424
rect 666614 132368 666619 132424
rect 666510 132366 666619 132368
rect 666553 132363 666619 132366
rect 676213 132290 676279 132293
rect 676213 132288 676322 132290
rect 676213 132232 676218 132288
rect 676274 132232 676322 132288
rect 676213 132227 676322 132232
rect 676262 132124 676322 132227
rect 578969 132018 579035 132021
rect 576380 132016 579035 132018
rect 576380 131960 578974 132016
rect 579030 131960 579035 132016
rect 576380 131958 579035 131960
rect 578969 131955 579035 131958
rect 603073 132018 603139 132021
rect 603073 132016 606556 132018
rect 603073 131960 603078 132016
rect 603134 131960 606556 132016
rect 603073 131958 606556 131960
rect 603073 131955 603139 131958
rect 676262 131477 676322 131716
rect 676213 131472 676322 131477
rect 676213 131416 676218 131472
rect 676274 131416 676322 131472
rect 676213 131414 676322 131416
rect 676213 131411 676279 131414
rect 676029 131338 676095 131341
rect 676029 131336 676292 131338
rect 676029 131280 676034 131336
rect 676090 131280 676292 131336
rect 676029 131278 676292 131280
rect 676029 131275 676095 131278
rect 603073 131066 603139 131069
rect 603073 131064 606556 131066
rect 603073 131008 603078 131064
rect 603134 131008 606556 131064
rect 603073 131006 606556 131008
rect 603073 131003 603139 131006
rect 676262 130661 676322 130900
rect 676213 130656 676322 130661
rect 676213 130600 676218 130656
rect 676274 130600 676322 130656
rect 676213 130598 676322 130600
rect 676213 130595 676279 130598
rect 579245 130522 579311 130525
rect 576380 130520 579311 130522
rect 576380 130464 579250 130520
rect 579306 130464 579311 130520
rect 576380 130462 579311 130464
rect 579245 130459 579311 130462
rect 676029 130522 676095 130525
rect 676029 130520 676292 130522
rect 676029 130464 676034 130520
rect 676090 130464 676292 130520
rect 676029 130462 676292 130464
rect 676029 130459 676095 130462
rect 603809 129978 603875 129981
rect 603809 129976 606556 129978
rect 603809 129920 603814 129976
rect 603870 129920 606556 129976
rect 603809 129918 606556 129920
rect 603809 129915 603875 129918
rect 676262 129845 676322 130084
rect 676213 129840 676322 129845
rect 676213 129784 676218 129840
rect 676274 129784 676322 129840
rect 676213 129782 676322 129784
rect 676213 129779 676279 129782
rect 666553 129570 666619 129573
rect 666356 129568 666619 129570
rect 666356 129512 666558 129568
rect 666614 129512 666619 129568
rect 666356 129510 666619 129512
rect 666553 129507 666619 129510
rect 676121 129434 676187 129437
rect 676262 129434 676322 129676
rect 676121 129432 676322 129434
rect 676121 129376 676126 129432
rect 676182 129376 676322 129432
rect 676121 129374 676322 129376
rect 676121 129371 676187 129374
rect 676262 129029 676322 129268
rect 578877 129026 578943 129029
rect 576380 129024 578943 129026
rect 576380 128968 578882 129024
rect 578938 128968 578943 129024
rect 576380 128966 578943 128968
rect 578877 128963 578943 128966
rect 603073 129026 603139 129029
rect 603073 129024 606556 129026
rect 603073 128968 603078 129024
rect 603134 128968 606556 129024
rect 603073 128966 606556 128968
rect 676213 129024 676322 129029
rect 676213 128968 676218 129024
rect 676274 128968 676322 129024
rect 676213 128966 676322 128968
rect 603073 128963 603139 128966
rect 676213 128963 676279 128966
rect 676070 128556 676076 128620
rect 676140 128618 676146 128620
rect 676262 128618 676322 128860
rect 676140 128558 676322 128618
rect 676140 128556 676146 128558
rect 683622 128213 683682 128452
rect 683622 128208 683731 128213
rect 683622 128152 683670 128208
rect 683726 128152 683731 128208
rect 683622 128150 683731 128152
rect 683665 128147 683731 128150
rect 676029 128074 676095 128077
rect 676029 128072 676292 128074
rect 676029 128016 676034 128072
rect 676090 128016 676292 128072
rect 676029 128014 676292 128016
rect 676029 128011 676095 128014
rect 603073 127938 603139 127941
rect 668025 127938 668091 127941
rect 603073 127936 606556 127938
rect 603073 127880 603078 127936
rect 603134 127880 606556 127936
rect 603073 127878 606556 127880
rect 666356 127936 668091 127938
rect 666356 127880 668030 127936
rect 668086 127880 668091 127936
rect 666356 127878 668091 127880
rect 603073 127875 603139 127878
rect 668025 127875 668091 127878
rect 578877 127530 578943 127533
rect 576380 127528 578943 127530
rect 576380 127472 578882 127528
rect 578938 127472 578943 127528
rect 576380 127470 578943 127472
rect 578877 127467 578943 127470
rect 683070 127397 683130 127636
rect 683070 127392 683179 127397
rect 683070 127336 683118 127392
rect 683174 127336 683179 127392
rect 683070 127334 683179 127336
rect 683113 127331 683179 127334
rect 676814 126989 676874 127228
rect 603165 126986 603231 126989
rect 603165 126984 606556 126986
rect 603165 126928 603170 126984
rect 603226 126928 606556 126984
rect 603165 126926 606556 126928
rect 676814 126984 676923 126989
rect 676814 126928 676862 126984
rect 676918 126928 676923 126984
rect 676814 126926 676923 126928
rect 603165 126923 603231 126926
rect 676857 126923 676923 126926
rect 676262 126580 676322 126820
rect 676254 126516 676260 126580
rect 676324 126516 676330 126580
rect 683254 126173 683314 126412
rect 683254 126168 683363 126173
rect 683254 126112 683302 126168
rect 683358 126112 683363 126168
rect 683254 126110 683363 126112
rect 683297 126107 683363 126110
rect 579061 126034 579127 126037
rect 576380 126032 579127 126034
rect 576380 125976 579066 126032
rect 579122 125976 579127 126032
rect 576380 125974 579127 125976
rect 579061 125971 579127 125974
rect 603073 125898 603139 125901
rect 603073 125896 606556 125898
rect 603073 125840 603078 125896
rect 603134 125840 606556 125896
rect 603073 125838 606556 125840
rect 603073 125835 603139 125838
rect 679574 125765 679634 126004
rect 679574 125760 679683 125765
rect 679574 125704 679622 125760
rect 679678 125704 679683 125760
rect 679574 125702 679683 125704
rect 679617 125699 679683 125702
rect 678286 125357 678346 125596
rect 676397 125354 676463 125357
rect 676397 125352 676506 125354
rect 676397 125296 676402 125352
rect 676458 125296 676506 125352
rect 676397 125291 676506 125296
rect 678237 125352 678346 125357
rect 678237 125296 678242 125352
rect 678298 125296 678346 125352
rect 678237 125294 678346 125296
rect 678237 125291 678303 125294
rect 676446 125188 676506 125291
rect 603073 124946 603139 124949
rect 603073 124944 606556 124946
rect 603073 124888 603078 124944
rect 603134 124888 606556 124944
rect 603073 124886 606556 124888
rect 603073 124883 603139 124886
rect 675886 124884 675892 124948
rect 675956 124946 675962 124948
rect 683113 124946 683179 124949
rect 675956 124944 683179 124946
rect 675956 124888 683118 124944
rect 683174 124888 683179 124944
rect 675956 124886 683179 124888
rect 675956 124884 675962 124886
rect 683113 124883 683179 124886
rect 578417 124538 578483 124541
rect 668025 124538 668091 124541
rect 676446 124540 676506 124780
rect 576380 124536 578483 124538
rect 576380 124480 578422 124536
rect 578478 124480 578483 124536
rect 576380 124478 578483 124480
rect 666356 124536 668091 124538
rect 666356 124480 668030 124536
rect 668086 124480 668091 124536
rect 666356 124478 668091 124480
rect 578417 124475 578483 124478
rect 668025 124475 668091 124478
rect 676438 124476 676444 124540
rect 676508 124476 676514 124540
rect 677550 124133 677610 124372
rect 677550 124128 677659 124133
rect 677550 124072 677598 124128
rect 677654 124072 677659 124128
rect 677550 124070 677659 124072
rect 677593 124067 677659 124070
rect 602429 123858 602495 123861
rect 602429 123856 606556 123858
rect 602429 123800 602434 123856
rect 602490 123800 606556 123856
rect 602429 123798 606556 123800
rect 602429 123795 602495 123798
rect 676262 123725 676322 123964
rect 676213 123720 676322 123725
rect 676213 123664 676218 123720
rect 676274 123664 676322 123720
rect 676213 123662 676322 123664
rect 676213 123659 676279 123662
rect 674741 123586 674807 123589
rect 674741 123584 676292 123586
rect 674741 123528 674746 123584
rect 674802 123528 676292 123584
rect 674741 123526 676292 123528
rect 674741 123523 674807 123526
rect 676262 122909 676322 123148
rect 579245 122906 579311 122909
rect 576380 122904 579311 122906
rect 576380 122848 579250 122904
rect 579306 122848 579311 122904
rect 576380 122846 579311 122848
rect 579245 122843 579311 122846
rect 603073 122906 603139 122909
rect 667933 122906 667999 122909
rect 603073 122904 606556 122906
rect 603073 122848 603078 122904
rect 603134 122848 606556 122904
rect 603073 122846 606556 122848
rect 666356 122904 667999 122906
rect 666356 122848 667938 122904
rect 667994 122848 667999 122904
rect 666356 122846 667999 122848
rect 603073 122843 603139 122846
rect 666510 122773 666570 122846
rect 667933 122843 667999 122846
rect 676213 122904 676322 122909
rect 676213 122848 676218 122904
rect 676274 122848 676322 122904
rect 676213 122846 676322 122848
rect 676213 122843 676279 122846
rect 666510 122768 666619 122773
rect 666510 122712 666558 122768
rect 666614 122712 666619 122768
rect 666510 122710 666619 122712
rect 666553 122707 666619 122710
rect 676121 122498 676187 122501
rect 676262 122498 676322 122740
rect 676121 122496 676322 122498
rect 676121 122440 676126 122496
rect 676182 122440 676322 122496
rect 676121 122438 676322 122440
rect 676121 122435 676187 122438
rect 603073 121818 603139 121821
rect 603073 121816 606556 121818
rect 603073 121760 603078 121816
rect 603134 121760 606556 121816
rect 603073 121758 606556 121760
rect 603073 121755 603139 121758
rect 676262 121685 676322 121924
rect 676213 121680 676322 121685
rect 676213 121624 676218 121680
rect 676274 121624 676322 121680
rect 676213 121622 676322 121624
rect 676213 121619 676279 121622
rect 676806 121620 676812 121684
rect 676876 121682 676882 121684
rect 683665 121682 683731 121685
rect 676876 121680 683731 121682
rect 676876 121624 683670 121680
rect 683726 121624 683731 121680
rect 676876 121622 683731 121624
rect 676876 121620 676882 121622
rect 683665 121619 683731 121622
rect 579521 121410 579587 121413
rect 576380 121408 579587 121410
rect 576380 121352 579526 121408
rect 579582 121352 579587 121408
rect 576380 121350 579587 121352
rect 579521 121347 579587 121350
rect 603073 120866 603139 120869
rect 603073 120864 606556 120866
rect 603073 120808 603078 120864
rect 603134 120808 606556 120864
rect 603073 120806 606556 120808
rect 603073 120803 603139 120806
rect 579245 119914 579311 119917
rect 576380 119912 579311 119914
rect 576380 119856 579250 119912
rect 579306 119856 579311 119912
rect 576380 119854 579311 119856
rect 579245 119851 579311 119854
rect 603073 119778 603139 119781
rect 603073 119776 606556 119778
rect 603073 119720 603078 119776
rect 603134 119720 606556 119776
rect 603073 119718 606556 119720
rect 603073 119715 603139 119718
rect 666553 119506 666619 119509
rect 666356 119504 666619 119506
rect 666356 119448 666558 119504
rect 666614 119448 666619 119504
rect 666356 119446 666619 119448
rect 666553 119443 666619 119446
rect 602337 118826 602403 118829
rect 602337 118824 606556 118826
rect 602337 118768 602342 118824
rect 602398 118768 606556 118824
rect 602337 118766 606556 118768
rect 602337 118763 602403 118766
rect 578601 118418 578667 118421
rect 576380 118416 578667 118418
rect 576380 118360 578606 118416
rect 578662 118360 578667 118416
rect 576380 118358 578667 118360
rect 578601 118355 578667 118358
rect 675702 117948 675708 118012
rect 675772 118010 675778 118012
rect 676857 118010 676923 118013
rect 675772 118008 676923 118010
rect 675772 117952 676862 118008
rect 676918 117952 676923 118008
rect 675772 117950 676923 117952
rect 675772 117948 675778 117950
rect 676857 117947 676923 117950
rect 603073 117738 603139 117741
rect 669221 117738 669287 117741
rect 603073 117736 606556 117738
rect 603073 117680 603078 117736
rect 603134 117680 606556 117736
rect 603073 117678 606556 117680
rect 666356 117736 669287 117738
rect 666356 117680 669226 117736
rect 669282 117680 669287 117736
rect 666356 117678 669287 117680
rect 603073 117675 603139 117678
rect 669221 117675 669287 117678
rect 675334 117268 675340 117332
rect 675404 117330 675410 117332
rect 676397 117330 676463 117333
rect 675404 117328 676463 117330
rect 675404 117272 676402 117328
rect 676458 117272 676463 117328
rect 675404 117270 676463 117272
rect 675404 117268 675410 117270
rect 676397 117267 676463 117270
rect 675518 117132 675524 117196
rect 675588 117194 675594 117196
rect 679617 117194 679683 117197
rect 675588 117192 679683 117194
rect 675588 117136 679622 117192
rect 679678 117136 679683 117192
rect 675588 117134 679683 117136
rect 675588 117132 675594 117134
rect 679617 117131 679683 117134
rect 579521 116922 579587 116925
rect 576380 116920 579587 116922
rect 576380 116864 579526 116920
rect 579582 116864 579587 116920
rect 576380 116862 579587 116864
rect 579521 116859 579587 116862
rect 603441 116786 603507 116789
rect 603441 116784 606556 116786
rect 603441 116728 603446 116784
rect 603502 116728 606556 116784
rect 603441 116726 606556 116728
rect 603441 116723 603507 116726
rect 668485 116106 668551 116109
rect 666356 116104 668551 116106
rect 666356 116048 668490 116104
rect 668546 116048 668551 116104
rect 666356 116046 668551 116048
rect 668485 116043 668551 116046
rect 603073 115698 603139 115701
rect 603073 115696 606556 115698
rect 603073 115640 603078 115696
rect 603134 115640 606556 115696
rect 603073 115638 606556 115640
rect 603073 115635 603139 115638
rect 579521 115426 579587 115429
rect 576380 115424 579587 115426
rect 576380 115368 579526 115424
rect 579582 115368 579587 115424
rect 576380 115366 579587 115368
rect 579521 115363 579587 115366
rect 603165 114746 603231 114749
rect 603165 114744 606556 114746
rect 603165 114688 603170 114744
rect 603226 114688 606556 114744
rect 603165 114686 606556 114688
rect 603165 114683 603231 114686
rect 668485 114338 668551 114341
rect 666356 114336 668551 114338
rect 666356 114280 668490 114336
rect 668546 114280 668551 114336
rect 666356 114278 668551 114280
rect 668485 114275 668551 114278
rect 675753 114202 675819 114205
rect 676070 114202 676076 114204
rect 675753 114200 676076 114202
rect 675753 114144 675758 114200
rect 675814 114144 676076 114200
rect 675753 114142 676076 114144
rect 675753 114139 675819 114142
rect 676070 114140 676076 114142
rect 676140 114140 676146 114204
rect 579245 113930 579311 113933
rect 576380 113928 579311 113930
rect 576380 113872 579250 113928
rect 579306 113872 579311 113928
rect 576380 113870 579311 113872
rect 579245 113867 579311 113870
rect 603073 113658 603139 113661
rect 603073 113656 606556 113658
rect 603073 113600 603078 113656
rect 603134 113600 606556 113656
rect 603073 113598 606556 113600
rect 603073 113595 603139 113598
rect 603073 112706 603139 112709
rect 668853 112706 668919 112709
rect 603073 112704 606556 112706
rect 603073 112648 603078 112704
rect 603134 112648 606556 112704
rect 603073 112646 606556 112648
rect 666356 112704 668919 112706
rect 666356 112648 668858 112704
rect 668914 112648 668919 112704
rect 666356 112646 668919 112648
rect 603073 112643 603139 112646
rect 668853 112643 668919 112646
rect 675753 112570 675819 112573
rect 675886 112570 675892 112572
rect 675753 112568 675892 112570
rect 675753 112512 675758 112568
rect 675814 112512 675892 112568
rect 675753 112510 675892 112512
rect 675753 112507 675819 112510
rect 675886 112508 675892 112510
rect 675956 112508 675962 112572
rect 578417 112434 578483 112437
rect 576380 112432 578483 112434
rect 576380 112376 578422 112432
rect 578478 112376 578483 112432
rect 576380 112374 578483 112376
rect 578417 112371 578483 112374
rect 675477 111756 675543 111757
rect 675477 111752 675524 111756
rect 675588 111754 675594 111756
rect 675477 111696 675482 111752
rect 675477 111692 675524 111696
rect 675588 111694 675634 111754
rect 675588 111692 675594 111694
rect 675477 111691 675543 111692
rect 603073 111618 603139 111621
rect 603073 111616 606556 111618
rect 603073 111560 603078 111616
rect 603134 111560 606556 111616
rect 603073 111558 606556 111560
rect 603073 111555 603139 111558
rect 578693 110938 578759 110941
rect 667933 110938 667999 110941
rect 576380 110936 578759 110938
rect 576380 110880 578698 110936
rect 578754 110880 578759 110936
rect 576380 110878 578759 110880
rect 666356 110936 667999 110938
rect 666356 110880 667938 110936
rect 667994 110880 667999 110936
rect 666356 110878 667999 110880
rect 578693 110875 578759 110878
rect 667933 110875 667999 110878
rect 603809 110666 603875 110669
rect 603809 110664 606556 110666
rect 603809 110608 603814 110664
rect 603870 110608 606556 110664
rect 603809 110606 606556 110608
rect 603809 110603 603875 110606
rect 603073 109578 603139 109581
rect 603073 109576 606556 109578
rect 603073 109520 603078 109576
rect 603134 109520 606556 109576
rect 603073 109518 606556 109520
rect 603073 109515 603139 109518
rect 579429 109442 579495 109445
rect 576380 109440 579495 109442
rect 576380 109384 579434 109440
rect 579490 109384 579495 109440
rect 576380 109382 579495 109384
rect 579429 109379 579495 109382
rect 667933 109306 667999 109309
rect 666356 109304 667999 109306
rect 666356 109248 667938 109304
rect 667994 109248 667999 109304
rect 666356 109246 667999 109248
rect 667933 109243 667999 109246
rect 675109 109034 675175 109037
rect 676438 109034 676444 109036
rect 675109 109032 676444 109034
rect 675109 108976 675114 109032
rect 675170 108976 676444 109032
rect 675109 108974 676444 108976
rect 675109 108971 675175 108974
rect 676438 108972 676444 108974
rect 676508 108972 676514 109036
rect 603073 108626 603139 108629
rect 603073 108624 606556 108626
rect 603073 108568 603078 108624
rect 603134 108568 606556 108624
rect 603073 108566 606556 108568
rect 603073 108563 603139 108566
rect 675753 108220 675819 108221
rect 675702 108218 675708 108220
rect 675662 108158 675708 108218
rect 675772 108216 675819 108220
rect 675814 108160 675819 108216
rect 675702 108156 675708 108158
rect 675772 108156 675819 108160
rect 675753 108155 675819 108156
rect 579245 107946 579311 107949
rect 576380 107944 579311 107946
rect 576380 107888 579250 107944
rect 579306 107888 579311 107944
rect 576380 107886 579311 107888
rect 579245 107883 579311 107886
rect 603073 107538 603139 107541
rect 668117 107538 668183 107541
rect 603073 107536 606556 107538
rect 603073 107480 603078 107536
rect 603134 107480 606556 107536
rect 603073 107478 606556 107480
rect 666356 107536 668183 107538
rect 666356 107480 668122 107536
rect 668178 107480 668183 107536
rect 666356 107478 668183 107480
rect 603073 107475 603139 107478
rect 668117 107475 668183 107478
rect 603165 106586 603231 106589
rect 603165 106584 606556 106586
rect 603165 106528 603170 106584
rect 603226 106528 606556 106584
rect 603165 106526 606556 106528
rect 603165 106523 603231 106526
rect 579521 106450 579587 106453
rect 576380 106448 579587 106450
rect 576380 106392 579526 106448
rect 579582 106392 579587 106448
rect 576380 106390 579587 106392
rect 579521 106387 579587 106390
rect 669221 105906 669287 105909
rect 666356 105904 669287 105906
rect 666356 105848 669226 105904
rect 669282 105848 669287 105904
rect 666356 105846 669287 105848
rect 669221 105843 669287 105846
rect 603073 105498 603139 105501
rect 603073 105496 606556 105498
rect 603073 105440 603078 105496
rect 603134 105440 606556 105496
rect 603073 105438 606556 105440
rect 603073 105435 603139 105438
rect 579521 104954 579587 104957
rect 576380 104952 579587 104954
rect 576380 104896 579526 104952
rect 579582 104896 579587 104952
rect 576380 104894 579587 104896
rect 579521 104891 579587 104894
rect 675334 104756 675340 104820
rect 675404 104818 675410 104820
rect 675477 104818 675543 104821
rect 675404 104816 675543 104818
rect 675404 104760 675482 104816
rect 675538 104760 675543 104816
rect 675404 104758 675543 104760
rect 675404 104756 675410 104758
rect 675477 104755 675543 104758
rect 603717 104546 603783 104549
rect 603717 104544 606556 104546
rect 603717 104488 603722 104544
rect 603778 104488 606556 104544
rect 603717 104486 606556 104488
rect 603717 104483 603783 104486
rect 668669 104138 668735 104141
rect 666356 104136 668735 104138
rect 666356 104080 668674 104136
rect 668730 104080 668735 104136
rect 666356 104078 668735 104080
rect 668669 104075 668735 104078
rect 578509 103458 578575 103461
rect 576380 103456 578575 103458
rect 576380 103400 578514 103456
rect 578570 103400 578575 103456
rect 576380 103398 578575 103400
rect 578509 103395 578575 103398
rect 603165 103458 603231 103461
rect 603165 103456 606556 103458
rect 603165 103400 603170 103456
rect 603226 103400 606556 103456
rect 603165 103398 606556 103400
rect 603165 103395 603231 103398
rect 675753 103186 675819 103189
rect 676806 103186 676812 103188
rect 675753 103184 676812 103186
rect 675753 103128 675758 103184
rect 675814 103128 676812 103184
rect 675753 103126 676812 103128
rect 675753 103123 675819 103126
rect 676806 103124 676812 103126
rect 676876 103124 676882 103188
rect 603073 102506 603139 102509
rect 668761 102506 668827 102509
rect 603073 102504 606556 102506
rect 603073 102448 603078 102504
rect 603134 102448 606556 102504
rect 603073 102446 606556 102448
rect 666356 102504 668827 102506
rect 666356 102448 668766 102504
rect 668822 102448 668827 102504
rect 666356 102446 668827 102448
rect 603073 102443 603139 102446
rect 668761 102443 668827 102446
rect 578325 101962 578391 101965
rect 576380 101960 578391 101962
rect 576380 101904 578330 101960
rect 578386 101904 578391 101960
rect 576380 101902 578391 101904
rect 578325 101899 578391 101902
rect 603073 101418 603139 101421
rect 675753 101418 675819 101421
rect 676254 101418 676260 101420
rect 603073 101416 606556 101418
rect 603073 101360 603078 101416
rect 603134 101360 606556 101416
rect 603073 101358 606556 101360
rect 675753 101416 676260 101418
rect 675753 101360 675758 101416
rect 675814 101360 676260 101416
rect 675753 101358 676260 101360
rect 603073 101355 603139 101358
rect 675753 101355 675819 101358
rect 676254 101356 676260 101358
rect 676324 101356 676330 101420
rect 668577 100874 668643 100877
rect 666356 100872 668643 100874
rect 666356 100816 668582 100872
rect 668638 100816 668643 100872
rect 666356 100814 668643 100816
rect 668577 100811 668643 100814
rect 603073 100466 603139 100469
rect 603073 100464 606556 100466
rect 603073 100408 603078 100464
rect 603134 100408 606556 100464
rect 603073 100406 606556 100408
rect 603073 100403 603139 100406
rect 578693 100330 578759 100333
rect 576380 100328 578759 100330
rect 576380 100272 578698 100328
rect 578754 100272 578759 100328
rect 576380 100270 578759 100272
rect 578693 100267 578759 100270
rect 579521 98834 579587 98837
rect 576380 98832 579587 98834
rect 576380 98776 579526 98832
rect 579582 98776 579587 98832
rect 576380 98774 579587 98776
rect 579521 98771 579587 98774
rect 579521 97338 579587 97341
rect 576380 97336 579587 97338
rect 576380 97280 579526 97336
rect 579582 97280 579587 97336
rect 576380 97278 579587 97280
rect 579521 97275 579587 97278
rect 641713 96660 641779 96661
rect 641662 96658 641668 96660
rect 641622 96598 641668 96658
rect 641732 96656 641779 96660
rect 641774 96600 641779 96656
rect 641662 96596 641668 96598
rect 641732 96596 641779 96600
rect 641713 96595 641779 96596
rect 639822 96460 639828 96524
rect 639892 96522 639898 96524
rect 642265 96522 642331 96525
rect 639892 96520 642331 96522
rect 639892 96464 642270 96520
rect 642326 96464 642331 96520
rect 639892 96462 642331 96464
rect 639892 96460 639898 96462
rect 642265 96459 642331 96462
rect 628281 95978 628347 95981
rect 628238 95976 628347 95978
rect 628238 95920 628286 95976
rect 628342 95920 628347 95976
rect 628238 95915 628347 95920
rect 578601 95842 578667 95845
rect 576380 95840 578667 95842
rect 576380 95784 578606 95840
rect 578662 95784 578667 95840
rect 576380 95782 578667 95784
rect 578601 95779 578667 95782
rect 628238 95404 628298 95915
rect 657353 94754 657419 94757
rect 657310 94752 657419 94754
rect 657310 94696 657358 94752
rect 657414 94696 657419 94752
rect 657310 94691 657419 94696
rect 644565 94618 644631 94621
rect 642988 94616 644631 94618
rect 642988 94560 644570 94616
rect 644626 94560 644631 94616
rect 642988 94558 644631 94560
rect 644565 94555 644631 94558
rect 627821 94482 627887 94485
rect 627821 94480 628268 94482
rect 627821 94424 627826 94480
rect 627882 94424 628268 94480
rect 627821 94422 628268 94424
rect 627821 94419 627887 94422
rect 578693 94346 578759 94349
rect 576380 94344 578759 94346
rect 576380 94288 578698 94344
rect 578754 94288 578759 94344
rect 576380 94286 578759 94288
rect 578693 94283 578759 94286
rect 657310 94180 657370 94691
rect 626533 93530 626599 93533
rect 626533 93528 628268 93530
rect 626533 93472 626538 93528
rect 626594 93472 628268 93528
rect 626533 93470 628268 93472
rect 626533 93467 626599 93470
rect 655329 93394 655395 93397
rect 665357 93394 665423 93397
rect 655329 93392 656788 93394
rect 655329 93336 655334 93392
rect 655390 93336 656788 93392
rect 655329 93334 656788 93336
rect 663596 93392 665423 93394
rect 663596 93336 665362 93392
rect 665418 93336 665423 93392
rect 663596 93334 665423 93336
rect 655329 93331 655395 93334
rect 665357 93331 665423 93334
rect 579521 92850 579587 92853
rect 576380 92848 579587 92850
rect 576380 92792 579526 92848
rect 579582 92792 579587 92848
rect 576380 92790 579587 92792
rect 579521 92787 579587 92790
rect 626349 92578 626415 92581
rect 654777 92578 654843 92581
rect 663793 92578 663859 92581
rect 626349 92576 628268 92578
rect 626349 92520 626354 92576
rect 626410 92520 628268 92576
rect 626349 92518 628268 92520
rect 654777 92576 656788 92578
rect 654777 92520 654782 92576
rect 654838 92520 656788 92576
rect 654777 92518 656788 92520
rect 663596 92576 663859 92578
rect 663596 92520 663798 92576
rect 663854 92520 663859 92576
rect 663596 92518 663859 92520
rect 626349 92515 626415 92518
rect 654777 92515 654843 92518
rect 663793 92515 663859 92518
rect 644657 92170 644723 92173
rect 642988 92168 644723 92170
rect 642988 92112 644662 92168
rect 644718 92112 644723 92168
rect 642988 92110 644723 92112
rect 644657 92107 644723 92110
rect 665173 91762 665239 91765
rect 663596 91760 665239 91762
rect 663596 91704 665178 91760
rect 665234 91704 665239 91760
rect 663596 91702 665239 91704
rect 665173 91699 665239 91702
rect 626441 91626 626507 91629
rect 626441 91624 628268 91626
rect 626441 91568 626446 91624
rect 626502 91568 628268 91624
rect 626441 91566 628268 91568
rect 626441 91563 626507 91566
rect 654317 91490 654383 91493
rect 654317 91488 656788 91490
rect 654317 91432 654322 91488
rect 654378 91432 656788 91488
rect 654317 91430 656788 91432
rect 654317 91427 654383 91430
rect 579521 91354 579587 91357
rect 576380 91352 579587 91354
rect 576380 91296 579526 91352
rect 579582 91296 579587 91352
rect 576380 91294 579587 91296
rect 579521 91291 579587 91294
rect 625981 90674 626047 90677
rect 654869 90674 654935 90677
rect 663885 90674 663951 90677
rect 625981 90672 628268 90674
rect 625981 90616 625986 90672
rect 626042 90616 628268 90672
rect 625981 90614 628268 90616
rect 654869 90672 656788 90674
rect 654869 90616 654874 90672
rect 654930 90616 656788 90672
rect 654869 90614 656788 90616
rect 663596 90672 663951 90674
rect 663596 90616 663890 90672
rect 663946 90616 663951 90672
rect 663596 90614 663951 90616
rect 625981 90611 626047 90614
rect 654869 90611 654935 90614
rect 663885 90611 663951 90614
rect 579521 89858 579587 89861
rect 576380 89856 579587 89858
rect 576380 89800 579526 89856
rect 579582 89800 579587 89856
rect 576380 89798 579587 89800
rect 579521 89795 579587 89798
rect 655421 89858 655487 89861
rect 665265 89858 665331 89861
rect 655421 89856 656788 89858
rect 655421 89800 655426 89856
rect 655482 89800 656788 89856
rect 655421 89798 656788 89800
rect 663596 89856 665331 89858
rect 663596 89800 665270 89856
rect 665326 89800 665331 89856
rect 663596 89798 665331 89800
rect 655421 89795 655487 89798
rect 665265 89795 665331 89798
rect 625797 89722 625863 89725
rect 625797 89720 628268 89722
rect 625797 89664 625802 89720
rect 625858 89664 628268 89720
rect 625797 89662 628268 89664
rect 625797 89659 625863 89662
rect 642958 89586 643018 89692
rect 643093 89586 643159 89589
rect 642958 89584 643159 89586
rect 642958 89528 643098 89584
rect 643154 89528 643159 89584
rect 642958 89526 643159 89528
rect 643093 89523 643159 89526
rect 664069 89042 664135 89045
rect 663596 89040 664135 89042
rect 663596 88984 664074 89040
rect 664130 88984 664135 89040
rect 663596 88982 664135 88984
rect 664069 88979 664135 88982
rect 626441 88906 626507 88909
rect 626441 88904 628268 88906
rect 626441 88848 626446 88904
rect 626502 88848 628268 88904
rect 626441 88846 628268 88848
rect 626441 88843 626507 88846
rect 579521 88362 579587 88365
rect 576380 88360 579587 88362
rect 576380 88304 579526 88360
rect 579582 88304 579587 88360
rect 576380 88302 579587 88304
rect 579521 88299 579587 88302
rect 626441 87954 626507 87957
rect 626441 87952 628268 87954
rect 626441 87896 626446 87952
rect 626502 87896 628268 87952
rect 626441 87894 628268 87896
rect 626441 87891 626507 87894
rect 644473 87138 644539 87141
rect 642988 87136 644539 87138
rect 642988 87080 644478 87136
rect 644534 87080 644539 87136
rect 642988 87078 644539 87080
rect 644473 87075 644539 87078
rect 626349 87002 626415 87005
rect 626349 87000 628268 87002
rect 626349 86944 626354 87000
rect 626410 86944 628268 87000
rect 626349 86942 628268 86944
rect 626349 86939 626415 86942
rect 579521 86866 579587 86869
rect 576380 86864 579587 86866
rect 576380 86808 579526 86864
rect 579582 86808 579587 86864
rect 576380 86806 579587 86808
rect 579521 86803 579587 86806
rect 626441 86050 626507 86053
rect 626441 86048 628268 86050
rect 626441 85992 626446 86048
rect 626502 85992 628268 86048
rect 626441 85990 628268 85992
rect 626441 85987 626507 85990
rect 579521 85370 579587 85373
rect 576380 85368 579587 85370
rect 576380 85312 579526 85368
rect 579582 85312 579587 85368
rect 576380 85310 579587 85312
rect 579521 85307 579587 85310
rect 643185 85234 643251 85237
rect 642958 85232 643251 85234
rect 642958 85176 643190 85232
rect 643246 85176 643251 85232
rect 642958 85174 643251 85176
rect 626441 85098 626507 85101
rect 626441 85096 628268 85098
rect 626441 85040 626446 85096
rect 626502 85040 628268 85096
rect 626441 85038 628268 85040
rect 626441 85035 626507 85038
rect 642958 84660 643018 85174
rect 643185 85171 643251 85174
rect 625613 84146 625679 84149
rect 625613 84144 628268 84146
rect 625613 84088 625618 84144
rect 625674 84088 628268 84144
rect 625613 84086 628268 84088
rect 625613 84083 625679 84086
rect 579521 83874 579587 83877
rect 576380 83872 579587 83874
rect 576380 83816 579526 83872
rect 579582 83816 579587 83872
rect 576380 83814 579587 83816
rect 579521 83811 579587 83814
rect 626441 83194 626507 83197
rect 626441 83192 628268 83194
rect 626441 83136 626446 83192
rect 626502 83136 628268 83192
rect 626441 83134 628268 83136
rect 626441 83131 626507 83134
rect 39456 82706 45844 82744
rect 39456 78242 41937 82706
rect 45681 78242 45844 82706
rect 579153 82378 579219 82381
rect 576380 82376 579219 82378
rect 576380 82320 579158 82376
rect 579214 82320 579219 82376
rect 576380 82318 579219 82320
rect 579153 82315 579219 82318
rect 626441 82242 626507 82245
rect 643277 82242 643343 82245
rect 626441 82240 628268 82242
rect 626441 82184 626446 82240
rect 626502 82184 628268 82240
rect 626441 82182 628268 82184
rect 642988 82240 643343 82242
rect 642988 82184 643282 82240
rect 643338 82184 643343 82240
rect 642988 82182 643343 82184
rect 626441 82179 626507 82182
rect 643277 82179 643343 82182
rect 578509 80882 578575 80885
rect 576380 80880 578575 80882
rect 576380 80824 578514 80880
rect 578570 80824 578575 80880
rect 576380 80822 578575 80824
rect 628790 80882 628850 81396
rect 629201 80882 629267 80885
rect 628790 80880 629267 80882
rect 628790 80824 629206 80880
rect 629262 80824 629267 80880
rect 628790 80822 629267 80824
rect 578509 80819 578575 80822
rect 629201 80819 629267 80822
rect 579061 79386 579127 79389
rect 576380 79384 579127 79386
rect 576380 79328 579066 79384
rect 579122 79328 579127 79384
rect 576380 79326 579127 79328
rect 579061 79323 579127 79326
rect 39456 78151 45844 78242
rect 579521 77890 579587 77893
rect 576380 77888 579587 77890
rect 576380 77832 579526 77888
rect 579582 77832 579587 77888
rect 576380 77830 579587 77832
rect 579521 77827 579587 77830
rect 633893 77890 633959 77893
rect 634670 77890 634676 77892
rect 633893 77888 634676 77890
rect 633893 77832 633898 77888
rect 633954 77832 634676 77888
rect 633893 77830 634676 77832
rect 633893 77827 633959 77830
rect 634670 77828 634676 77830
rect 634740 77828 634746 77892
rect 639597 77754 639663 77757
rect 639822 77754 639828 77756
rect 639597 77752 639828 77754
rect 639597 77696 639602 77752
rect 639658 77696 639828 77752
rect 639597 77694 639828 77696
rect 639597 77691 639663 77694
rect 639822 77692 639828 77694
rect 639892 77692 639898 77756
rect 578969 76258 579035 76261
rect 576380 76256 579035 76258
rect 576380 76200 578974 76256
rect 579030 76200 579035 76256
rect 576380 76198 579035 76200
rect 578969 76195 579035 76198
rect 638902 75108 638908 75172
rect 638972 75170 638978 75172
rect 639229 75170 639295 75173
rect 638972 75168 639295 75170
rect 638972 75112 639234 75168
rect 639290 75112 639295 75168
rect 638972 75110 639295 75112
rect 638972 75108 638978 75110
rect 639229 75107 639295 75110
rect 579521 74762 579587 74765
rect 576380 74760 579587 74762
rect 576380 74704 579526 74760
rect 579582 74704 579587 74760
rect 576380 74702 579587 74704
rect 579521 74699 579587 74702
rect 623773 74762 623839 74765
rect 633525 74762 633591 74765
rect 623773 74760 633591 74762
rect 623773 74704 623778 74760
rect 623834 74704 633530 74760
rect 633586 74704 633591 74760
rect 623773 74702 633591 74704
rect 623773 74699 623839 74702
rect 633525 74699 633591 74702
rect 646865 74490 646931 74493
rect 646668 74488 646931 74490
rect 646668 74432 646870 74488
rect 646926 74432 646931 74488
rect 646668 74430 646931 74432
rect 646865 74427 646931 74430
rect 578877 73266 578943 73269
rect 576380 73264 578943 73266
rect 576380 73208 578882 73264
rect 578938 73208 578943 73264
rect 576380 73206 578943 73208
rect 578877 73203 578943 73206
rect 646957 72994 647023 72997
rect 646668 72992 647023 72994
rect 646668 72936 646962 72992
rect 647018 72936 647023 72992
rect 646668 72934 647023 72936
rect 646957 72931 647023 72934
rect 39456 72802 45844 72900
rect 39456 68338 41913 72802
rect 45657 68338 45844 72802
rect 579521 71770 579587 71773
rect 646129 71770 646195 71773
rect 576380 71768 579587 71770
rect 576380 71712 579526 71768
rect 579582 71712 579587 71768
rect 576380 71710 579587 71712
rect 579521 71707 579587 71710
rect 646086 71768 646195 71770
rect 646086 71712 646134 71768
rect 646190 71712 646195 71768
rect 646086 71707 646195 71712
rect 646086 71468 646146 71707
rect 579521 70274 579587 70277
rect 576380 70272 579587 70274
rect 576380 70216 579526 70272
rect 579582 70216 579587 70272
rect 576380 70214 579587 70216
rect 579521 70211 579587 70214
rect 647233 70002 647299 70005
rect 646668 70000 647299 70002
rect 646668 69944 647238 70000
rect 647294 69944 647299 70000
rect 646668 69942 647299 69944
rect 647233 69939 647299 69942
rect 578325 68778 578391 68781
rect 576380 68776 578391 68778
rect 576380 68720 578330 68776
rect 578386 68720 578391 68776
rect 576380 68718 578391 68720
rect 578325 68715 578391 68718
rect 648797 68506 648863 68509
rect 646668 68504 648863 68506
rect 646668 68448 648802 68504
rect 648858 68448 648863 68504
rect 646668 68446 648863 68448
rect 648797 68443 648863 68446
rect 39456 68256 45844 68338
rect 579521 67282 579587 67285
rect 576380 67280 579587 67282
rect 576380 67224 579526 67280
rect 579582 67224 579587 67280
rect 576380 67222 579587 67224
rect 579521 67219 579587 67222
rect 647417 67010 647483 67013
rect 646668 67008 647483 67010
rect 646668 66952 647422 67008
rect 647478 66952 647483 67008
rect 646668 66950 647483 66952
rect 647417 66947 647483 66950
rect 646129 66058 646195 66061
rect 646086 66056 646195 66058
rect 646086 66000 646134 66056
rect 646190 66000 646195 66056
rect 646086 65995 646195 66000
rect 579245 65786 579311 65789
rect 576380 65784 579311 65786
rect 576380 65728 579250 65784
rect 579306 65728 579311 65784
rect 576380 65726 579311 65728
rect 579245 65723 579311 65726
rect 646086 65484 646146 65995
rect 646129 64426 646195 64429
rect 646086 64424 646195 64426
rect 646086 64368 646134 64424
rect 646190 64368 646195 64424
rect 646086 64363 646195 64368
rect 579521 64290 579587 64293
rect 576380 64288 579587 64290
rect 576380 64232 579526 64288
rect 579582 64232 579587 64288
rect 576380 64230 579587 64232
rect 579521 64227 579587 64230
rect 646086 63988 646146 64363
rect 579521 62794 579587 62797
rect 576380 62792 579587 62794
rect 576380 62736 579526 62792
rect 579582 62736 579587 62792
rect 576380 62734 579587 62736
rect 579521 62731 579587 62734
rect 578693 61298 578759 61301
rect 576380 61296 578759 61298
rect 576380 61240 578698 61296
rect 578754 61240 578759 61296
rect 576380 61238 578759 61240
rect 578693 61235 578759 61238
rect 578969 59802 579035 59805
rect 576380 59800 579035 59802
rect 576380 59744 578974 59800
rect 579030 59744 579035 59800
rect 576380 59742 579035 59744
rect 578969 59739 579035 59742
rect 578877 58306 578943 58309
rect 576380 58304 578943 58306
rect 576380 58248 578882 58304
rect 578938 58248 578943 58304
rect 576380 58246 578943 58248
rect 578877 58243 578943 58246
rect 578877 56810 578943 56813
rect 576380 56808 578943 56810
rect 576380 56752 578882 56808
rect 578938 56752 578943 56808
rect 576380 56750 578943 56752
rect 578877 56747 578943 56750
rect 578233 55314 578299 55317
rect 576380 55312 578299 55314
rect 576380 55256 578238 55312
rect 578294 55256 578299 55312
rect 576380 55254 578299 55256
rect 578233 55251 578299 55254
rect 578325 53818 578391 53821
rect 576380 53816 578391 53818
rect 576380 53760 578330 53816
rect 578386 53760 578391 53816
rect 576380 53758 578391 53760
rect 578325 53755 578391 53758
rect 189073 51778 189139 51781
rect 638902 51778 638908 51780
rect 189073 51776 638908 51778
rect 189073 51720 189078 51776
rect 189134 51720 638908 51776
rect 189073 51718 638908 51720
rect 189073 51715 189139 51718
rect 638902 51716 638908 51718
rect 638972 51716 638978 51780
rect 281441 50554 281507 50557
rect 520222 50554 520228 50556
rect 281441 50552 520228 50554
rect 281441 50496 281446 50552
rect 281502 50496 520228 50552
rect 281441 50494 520228 50496
rect 281441 50491 281507 50494
rect 520222 50492 520228 50494
rect 520292 50492 520298 50556
rect 216121 50418 216187 50421
rect 521694 50418 521700 50420
rect 216121 50416 521700 50418
rect 216121 50360 216126 50416
rect 216182 50360 521700 50416
rect 216121 50358 521700 50360
rect 216121 50355 216187 50358
rect 521694 50356 521700 50358
rect 521764 50356 521770 50420
rect 85113 50282 85179 50285
rect 514702 50282 514708 50284
rect 85113 50280 514708 50282
rect 85113 50224 85118 50280
rect 85174 50224 514708 50280
rect 85113 50222 514708 50224
rect 85113 50219 85179 50222
rect 514702 50220 514708 50222
rect 514772 50220 514778 50284
rect 529790 50220 529796 50284
rect 529860 50282 529866 50284
rect 542997 50282 543063 50285
rect 529860 50280 543063 50282
rect 529860 50224 543002 50280
rect 543058 50224 543063 50280
rect 529860 50222 543063 50224
rect 529860 50220 529866 50222
rect 542997 50219 543063 50222
rect 664437 48514 664503 48517
rect 662094 48512 664503 48514
rect 661480 48456 664442 48512
rect 664498 48456 664503 48512
rect 661480 48454 664503 48456
rect 661480 48452 662154 48454
rect 664437 48451 664503 48454
rect 661174 47565 661234 47761
rect 661125 47560 661234 47565
rect 661125 47504 661130 47560
rect 661186 47504 661234 47560
rect 661125 47502 661234 47504
rect 661125 47499 661191 47502
rect 662413 47426 662479 47429
rect 661388 47424 662479 47426
rect 661388 47368 662418 47424
rect 662474 47368 662479 47424
rect 661388 47366 662479 47368
rect 662413 47363 662479 47366
rect 648104 47124 649670 47188
rect 241690 46621 246049 46686
rect 187550 44916 187556 44980
rect 187620 44978 187626 44980
rect 241513 44978 241579 44981
rect 187620 44976 241579 44978
rect 187620 44920 241518 44976
rect 241574 44920 241579 44976
rect 187620 44918 241579 44920
rect 187620 44916 187626 44918
rect 241513 44915 241579 44918
rect 194358 44780 194364 44844
rect 194428 44842 194434 44844
rect 241513 44842 241579 44845
rect 194428 44840 241579 44842
rect 194428 44784 241518 44840
rect 241574 44784 241579 44840
rect 194428 44782 241579 44784
rect 194428 44780 194434 44782
rect 241513 44779 241579 44782
rect 142337 44298 142403 44301
rect 142110 44296 142403 44298
rect 142110 44240 142342 44296
rect 142398 44240 142403 44296
rect 142110 44238 142403 44240
rect 141918 43964 141924 44028
rect 141988 44026 141994 44028
rect 142110 44026 142170 44238
rect 142337 44235 142403 44238
rect 141988 43966 142170 44026
rect 141988 43964 141994 43966
rect 241690 42837 241731 46621
rect 245995 42837 246049 46621
rect 251300 46635 255702 46686
rect 246113 44978 246179 44981
rect 251081 44978 251147 44981
rect 246113 44976 251147 44978
rect 246113 44920 246118 44976
rect 246174 44920 251086 44976
rect 251142 44920 251147 44976
rect 246113 44918 251147 44920
rect 246113 44915 246179 44918
rect 251081 44915 251147 44918
rect 246113 44842 246179 44845
rect 251081 44842 251147 44845
rect 246113 44840 251147 44842
rect 246113 44784 246118 44840
rect 246174 44784 251086 44840
rect 251142 44784 251147 44840
rect 246113 44782 251147 44784
rect 246113 44779 246179 44782
rect 251081 44779 251147 44782
rect 187509 42124 187575 42125
rect 194317 42124 194383 42125
rect 187509 42122 187556 42124
rect 187464 42120 187556 42122
rect 187464 42064 187514 42120
rect 187464 42062 187556 42064
rect 187509 42060 187556 42062
rect 187620 42060 187626 42124
rect 194317 42122 194364 42124
rect 194272 42120 194364 42122
rect 194272 42064 194322 42120
rect 194272 42062 194364 42064
rect 194317 42060 194364 42062
rect 194428 42060 194434 42124
rect 187509 42059 187575 42060
rect 194317 42059 194383 42060
rect 141693 40354 141759 40357
rect 141918 40354 141924 40356
rect 141693 40352 141924 40354
rect 141693 40296 141698 40352
rect 141754 40296 141924 40352
rect 141693 40294 141924 40296
rect 141693 40291 141759 40294
rect 141918 40292 141924 40294
rect 141988 40292 141994 40356
rect 241690 39426 246049 42837
rect 251300 42851 251383 46635
rect 255647 42851 255702 46635
rect 648104 46660 648155 47124
rect 649619 46660 649670 47124
rect 412449 46610 412515 46613
rect 518566 46610 518572 46612
rect 412449 46608 518572 46610
rect 412449 46552 412454 46608
rect 412510 46552 518572 46608
rect 412449 46550 518572 46552
rect 412449 46547 412515 46550
rect 518566 46548 518572 46550
rect 518636 46548 518642 46612
rect 648104 46590 649670 46660
rect 471646 46412 471652 46476
rect 471716 46474 471722 46476
rect 611445 46474 611511 46477
rect 471716 46472 611511 46474
rect 471716 46416 611450 46472
rect 611506 46416 611511 46472
rect 471716 46414 611511 46416
rect 471716 46412 471722 46414
rect 611445 46411 611511 46414
rect 473169 46338 473235 46341
rect 612825 46338 612891 46341
rect 473169 46336 612891 46338
rect 473169 46280 473174 46336
rect 473230 46280 612830 46336
rect 612886 46280 612891 46336
rect 473169 46278 612891 46280
rect 473169 46275 473235 46278
rect 612825 46275 612891 46278
rect 470133 46202 470199 46205
rect 612733 46202 612799 46205
rect 470133 46200 612799 46202
rect 470133 46144 470138 46200
rect 470194 46144 612738 46200
rect 612794 46144 612799 46200
rect 470133 46142 612799 46144
rect 470133 46139 470199 46142
rect 612733 46139 612799 46142
rect 419717 45522 419783 45525
rect 610065 45522 610131 45525
rect 419717 45520 610131 45522
rect 419717 45464 419722 45520
rect 419778 45464 610070 45520
rect 610126 45464 610131 45520
rect 419717 45462 610131 45464
rect 419717 45459 419783 45462
rect 610065 45459 610131 45462
rect 415393 45386 415459 45389
rect 610157 45386 610223 45389
rect 415393 45384 610223 45386
rect 415393 45328 415398 45384
rect 415454 45328 610162 45384
rect 610218 45328 610223 45384
rect 415393 45326 610223 45328
rect 415393 45323 415459 45326
rect 610157 45323 610223 45326
rect 365110 45188 365116 45252
rect 365180 45250 365186 45252
rect 607305 45250 607371 45253
rect 365180 45248 607371 45250
rect 365180 45192 607310 45248
rect 607366 45192 607371 45248
rect 365180 45190 607371 45192
rect 365180 45188 365186 45190
rect 607305 45187 607371 45190
rect 310094 45052 310100 45116
rect 310164 45114 310170 45116
rect 608593 45114 608659 45117
rect 310164 45112 608659 45114
rect 310164 45056 608598 45112
rect 608654 45056 608659 45112
rect 310164 45054 608659 45056
rect 310164 45052 310170 45054
rect 608593 45051 608659 45054
rect 255865 44978 255931 44981
rect 576117 44978 576183 44981
rect 255865 44976 576183 44978
rect 255865 44920 255870 44976
rect 255926 44920 576122 44976
rect 576178 44920 576183 44976
rect 255865 44918 576183 44920
rect 255865 44915 255931 44918
rect 576117 44915 576183 44918
rect 255865 44842 255931 44845
rect 661125 44842 661191 44845
rect 255865 44840 661191 44842
rect 255865 44784 255870 44840
rect 255926 44784 661130 44840
rect 661186 44784 661191 44840
rect 255865 44782 661191 44784
rect 255865 44779 255931 44782
rect 661125 44779 661191 44782
rect 478781 44706 478847 44709
rect 525926 44706 525932 44708
rect 478781 44704 525932 44706
rect 478781 44648 478786 44704
rect 478842 44648 525932 44704
rect 478781 44646 525932 44648
rect 478781 44643 478847 44646
rect 525926 44644 525932 44646
rect 525996 44644 526002 44708
rect 361757 43618 361823 43621
rect 605833 43618 605899 43621
rect 361757 43616 605899 43618
rect 361757 43560 361762 43616
rect 361818 43560 605838 43616
rect 605894 43560 605899 43616
rect 361757 43558 605899 43560
rect 361757 43555 361823 43558
rect 605833 43555 605899 43558
rect 307293 43482 307359 43485
rect 607213 43482 607279 43485
rect 307293 43480 607279 43482
rect 307293 43424 307298 43480
rect 307354 43424 607218 43480
rect 607274 43424 607279 43480
rect 307293 43422 607279 43424
rect 307293 43419 307359 43422
rect 607213 43419 607279 43422
rect 251300 39426 255702 42851
rect 310099 42396 310165 42397
rect 518617 42396 518683 42397
rect 310094 42394 310100 42396
rect 310008 42334 310100 42394
rect 310094 42332 310100 42334
rect 310164 42332 310170 42396
rect 518566 42332 518572 42396
rect 518636 42394 518683 42396
rect 518636 42392 518728 42394
rect 518678 42336 518728 42392
rect 518636 42334 518728 42336
rect 518636 42332 518683 42334
rect 310099 42331 310165 42332
rect 518617 42331 518683 42332
rect 365069 42124 365135 42125
rect 471605 42124 471671 42125
rect 365069 42122 365116 42124
rect 365024 42120 365116 42122
rect 365024 42064 365074 42120
rect 365024 42062 365116 42064
rect 365069 42060 365116 42062
rect 365180 42060 365186 42124
rect 471605 42122 471652 42124
rect 471560 42120 471652 42122
rect 471560 42064 471610 42120
rect 471560 42062 471652 42064
rect 471605 42060 471652 42062
rect 471716 42060 471722 42124
rect 514702 42060 514708 42124
rect 514772 42122 514778 42124
rect 514845 42122 514911 42125
rect 514772 42120 514911 42122
rect 514772 42064 514850 42120
rect 514906 42064 514911 42120
rect 514772 42062 514911 42064
rect 514772 42060 514778 42062
rect 365069 42059 365135 42060
rect 471605 42059 471671 42060
rect 514845 42059 514911 42062
rect 520222 42060 520228 42124
rect 520292 42122 520298 42124
rect 520365 42122 520431 42125
rect 521745 42124 521811 42125
rect 525977 42124 526043 42125
rect 520292 42120 520431 42122
rect 520292 42064 520370 42120
rect 520426 42064 520431 42120
rect 520292 42062 520431 42064
rect 520292 42060 520298 42062
rect 520365 42059 520431 42062
rect 521694 42060 521700 42124
rect 521764 42122 521811 42124
rect 521764 42120 521856 42122
rect 521806 42064 521856 42120
rect 521764 42062 521856 42064
rect 521764 42060 521811 42062
rect 525926 42060 525932 42124
rect 525996 42122 526043 42124
rect 529657 42122 529723 42125
rect 529790 42122 529796 42124
rect 525996 42120 526088 42122
rect 526038 42064 526088 42120
rect 525996 42062 526088 42064
rect 529657 42120 529796 42122
rect 529657 42064 529662 42120
rect 529718 42064 529796 42120
rect 529657 42062 529796 42064
rect 525996 42060 526043 42062
rect 521745 42059 521811 42060
rect 525977 42059 526043 42060
rect 529657 42059 529723 42062
rect 529790 42060 529796 42062
rect 529860 42060 529866 42124
rect 416681 41850 416747 41853
rect 460565 41850 460631 41853
rect 416681 41848 422310 41850
rect 416681 41792 416686 41848
rect 416742 41792 422310 41848
rect 416681 41790 422310 41792
rect 416681 41787 416747 41790
rect 422250 41442 422310 41790
rect 460565 41848 460950 41850
rect 460565 41792 460570 41848
rect 460626 41792 460950 41848
rect 460565 41790 460950 41792
rect 460565 41787 460631 41790
rect 460890 41578 460950 41790
rect 611353 41578 611419 41581
rect 460890 41576 611419 41578
rect 460890 41520 611358 41576
rect 611414 41520 611419 41576
rect 460890 41518 611419 41520
rect 611353 41515 611419 41518
rect 609973 41442 610039 41445
rect 422250 41440 610039 41442
rect 422250 41384 609978 41440
rect 610034 41384 610039 41440
rect 422250 41382 610039 41384
rect 609973 41379 610039 41382
<< via3 >>
rect 114809 1030864 115953 1031568
rect 113213 1029666 114357 1030370
rect 85252 997188 85316 997252
rect 84700 996916 84764 996980
rect 84700 995616 84764 995620
rect 84700 995560 84714 995616
rect 84714 995560 84764 995616
rect 84700 995556 84764 995560
rect 85252 995616 85316 995620
rect 85252 995560 85266 995616
rect 85266 995560 85316 995616
rect 85252 995556 85316 995560
rect 113227 995573 114331 996677
rect 88932 995480 88996 995484
rect 88932 995424 88946 995480
rect 88946 995424 88996 995480
rect 88932 995420 88996 995424
rect 166209 1030864 167353 1031568
rect 164613 1029666 165757 1030370
rect 136772 996100 136836 996164
rect 164627 995573 165731 996677
rect 114845 993979 115949 995083
rect 217609 1030864 218753 1031568
rect 216013 1029666 217157 1030370
rect 216027 995573 217131 996677
rect 136772 995012 136836 995076
rect 166245 993979 167349 995083
rect 269009 1030864 270153 1031568
rect 267413 1029666 268557 1030370
rect 243860 996372 243924 996436
rect 243860 995752 243924 995756
rect 243860 995696 243874 995752
rect 243874 995696 243924 995752
rect 243860 995692 243924 995696
rect 267427 995573 268531 996677
rect 217645 993979 218749 995083
rect 320609 1030864 321753 1031568
rect 319013 1029666 320157 1030370
rect 292436 997052 292500 997116
rect 292436 995480 292500 995484
rect 292436 995424 292450 995480
rect 292450 995424 292500 995480
rect 292436 995420 292500 995424
rect 269045 993979 270149 995083
rect 319027 995573 320131 996677
rect 371009 1030864 372153 1031568
rect 369413 1029666 370557 1030370
rect 369427 995573 370531 996677
rect 320645 993979 321749 995083
rect 438409 1030864 439553 1031568
rect 436813 1029666 437957 1030370
rect 383700 997732 383764 997796
rect 387564 996236 387628 996300
rect 390324 996100 390388 996164
rect 383700 995964 383764 996028
rect 389036 995828 389100 995892
rect 389404 995828 389468 995892
rect 390324 995692 390388 995756
rect 436827 995573 437931 996677
rect 371045 993979 372149 995083
rect 515409 1030864 516553 1031568
rect 513813 1029666 514957 1030370
rect 485636 995752 485700 995756
rect 485636 995696 485650 995752
rect 485650 995696 485700 995752
rect 485636 995692 485700 995696
rect 506428 995828 506492 995892
rect 513827 995573 514931 996677
rect 387564 995012 387628 995076
rect 438445 993979 439549 995083
rect 566809 1030864 567953 1031568
rect 565213 1029666 566357 1030370
rect 565227 995573 566331 996677
rect 515445 993979 516549 995083
rect 566845 993979 567949 995083
rect 575774 995123 580398 997067
rect 585744 995129 590368 997073
rect 114508 990932 114572 990996
rect 40540 968764 40604 968828
rect 40724 967268 40788 967332
rect 676444 966452 676508 966516
rect 676260 966180 676324 966244
rect 41644 965092 41708 965156
rect 676628 964956 676692 965020
rect 40908 963460 40972 963524
rect 676076 963324 676140 963388
rect 675708 962840 675772 962844
rect 675708 962784 675722 962840
rect 675722 962784 675772 962840
rect 675708 962780 675772 962784
rect 41828 962160 41892 962164
rect 41828 962104 41842 962160
rect 41842 962104 41892 962160
rect 41828 962100 41892 962104
rect 675524 961888 675588 961892
rect 675524 961832 675538 961888
rect 675538 961832 675588 961888
rect 675524 961828 675588 961832
rect 675892 959108 675956 959172
rect 42012 958488 42076 958492
rect 42012 958432 42062 958488
rect 42062 958432 42076 958488
rect 42012 958428 42076 958432
rect 676812 957884 676876 957948
rect 41460 957748 41524 957812
rect 676996 957612 677060 957676
rect 675340 954000 675404 954004
rect 675340 953944 675390 954000
rect 675390 953944 675404 954000
rect 675340 953940 675404 953944
rect 41828 952852 41892 952916
rect 42012 952308 42076 952372
rect 41644 952172 41708 952236
rect 6150 948809 6854 949953
rect 54235 948845 55339 949949
rect 675708 949724 675772 949788
rect 63339 948525 63883 949629
rect 675524 949588 675588 949652
rect 675340 949452 675404 949516
rect 7348 947213 8052 948357
rect 52641 947227 53745 948331
rect 62371 947017 62915 948121
rect 40724 943740 40788 943804
rect 42012 937756 42076 937820
rect 41828 936804 41892 936868
rect 676628 935580 676692 935644
rect 42012 934900 42076 934964
rect 676444 934764 676508 934828
rect 676076 933948 676140 934012
rect 675892 933812 675956 933876
rect 676628 933132 676692 933196
rect 676996 931500 677060 931564
rect 676812 931092 676876 931156
rect 675156 877236 675220 877300
rect 676260 876556 676324 876620
rect 676076 875876 676140 875940
rect 675892 873972 675956 874036
rect 676444 866764 676508 866828
rect 675708 864784 675772 864788
rect 675708 864728 675758 864784
rect 675758 864728 675772 864784
rect 675708 864724 675772 864728
rect 47909 837790 49693 842334
rect 47909 827858 49693 832402
rect 667276 828626 669740 833210
rect 6150 823009 6854 824153
rect 54235 823045 55339 824149
rect 63339 823025 63883 824129
rect 7348 821413 8052 822557
rect 52641 821427 53745 822531
rect 62371 821417 62915 822521
rect 667262 818632 669726 823216
rect 42012 816036 42076 816100
rect 41828 814404 41892 814468
rect 42196 811956 42260 812020
rect 41828 807876 41892 807940
rect 41644 802572 41708 802636
rect 42012 802436 42076 802500
rect 41828 801620 41892 801684
rect 41460 800940 41524 801004
rect 40540 796724 40604 796788
rect 42012 791964 42076 792028
rect 42196 791828 42260 791892
rect 41460 788156 41524 788220
rect 41828 788020 41892 788084
rect 41644 786116 41708 786180
rect 675708 785164 675772 785228
rect 675892 784892 675956 784956
rect 675524 784816 675588 784820
rect 675524 784760 675538 784816
rect 675538 784760 675588 784816
rect 675524 784756 675588 784760
rect 675156 784212 675220 784276
rect 675708 784212 675772 784276
rect 676628 784076 676692 784140
rect 63339 781025 63883 782129
rect 6150 779809 6854 780953
rect 54235 779845 55339 780949
rect 677180 779860 677244 779924
rect 7348 778213 8052 779357
rect 52641 778227 53745 779331
rect 62371 778217 62915 779321
rect 675156 775644 675220 775708
rect 675340 774828 675404 774892
rect 676812 774828 676876 774892
rect 40172 773468 40236 773532
rect 675708 773392 675772 773396
rect 675708 773336 675758 773392
rect 675758 773336 675772 773392
rect 675708 773332 675772 773336
rect 675892 772652 675956 772716
rect 39988 771836 40052 771900
rect 39988 771020 40052 771084
rect 40908 766124 40972 766188
rect 40540 764900 40604 764964
rect 40724 764492 40788 764556
rect 672764 759052 672828 759116
rect 41644 758236 41708 758300
rect 672764 757828 672828 757892
rect 41460 757692 41524 757756
rect 676076 757148 676140 757212
rect 42748 756528 42812 756532
rect 42748 756472 42762 756528
rect 42762 756472 42812 756528
rect 42748 756468 42812 756472
rect 676812 755924 676876 755988
rect 40908 755244 40972 755308
rect 41828 755244 41892 755308
rect 676260 754700 676324 754764
rect 676444 753476 676508 753540
rect 41828 753128 41892 753132
rect 41828 753072 41842 753128
rect 41842 753072 41892 753128
rect 41828 753068 41892 753072
rect 40724 751708 40788 751772
rect 40540 750348 40604 750412
rect 42748 749320 42812 749324
rect 42748 749264 42762 749320
rect 42762 749264 42812 749320
rect 42748 749260 42812 749264
rect 41644 746540 41708 746604
rect 41460 742324 41524 742388
rect 675340 741644 675404 741708
rect 675892 739876 675956 739940
rect 675708 739256 675772 739260
rect 675708 739200 675722 739256
rect 675722 739200 675772 739256
rect 675708 739196 675772 739200
rect 6150 736609 6854 737753
rect 54235 736645 55339 737749
rect 63339 736625 63883 737729
rect 7348 735013 8052 736157
rect 52641 735027 53745 736131
rect 62371 735017 62915 736121
rect 676812 734300 676876 734364
rect 676996 732940 677060 733004
rect 40172 729404 40236 729468
rect 39988 728588 40052 728652
rect 39988 727772 40052 727836
rect 675156 727228 675220 727292
rect 41460 726140 41524 726204
rect 40540 721244 40604 721308
rect 41828 715532 41892 715596
rect 41644 715396 41708 715460
rect 40908 714036 40972 714100
rect 42012 713824 42076 713828
rect 42012 713768 42062 713824
rect 42062 713768 42076 713824
rect 42012 713764 42076 713768
rect 677364 713488 677428 713492
rect 677364 713432 677378 713488
rect 677378 713432 677428 713488
rect 677364 713428 677428 713432
rect 42196 713220 42260 713284
rect 42380 712268 42444 712332
rect 42196 711784 42260 711788
rect 42196 711728 42210 711784
rect 42210 711728 42260 711784
rect 42196 711724 42260 711728
rect 676076 711044 676140 711108
rect 40540 710772 40604 710836
rect 675524 710772 675588 710836
rect 40908 709820 40972 709884
rect 676076 708868 676140 708932
rect 42380 708460 42444 708524
rect 42012 706556 42076 706620
rect 41828 704924 41892 704988
rect 676260 704380 676324 704444
rect 41644 702884 41708 702948
rect 41460 699348 41524 699412
rect 674604 697308 674668 697372
rect 675708 696960 675772 696964
rect 675708 696904 675722 696960
rect 675722 696904 675772 696960
rect 675708 696900 675772 696904
rect 676076 694996 676140 695060
rect 6150 693409 6854 694553
rect 54235 693445 55339 694549
rect 63339 693425 63883 694529
rect 676444 694180 676508 694244
rect 7348 691813 8052 692957
rect 52641 691827 53745 692931
rect 62371 691817 62915 692921
rect 40172 687108 40236 687172
rect 39988 685476 40052 685540
rect 39988 684660 40052 684724
rect 41460 682212 41524 682276
rect 40540 679356 40604 679420
rect 675340 678948 675404 679012
rect 40724 678132 40788 678196
rect 30604 677724 30668 677788
rect 30604 676500 30668 676564
rect 41644 671332 41708 671396
rect 41828 670924 41892 670988
rect 42012 670712 42076 670716
rect 42012 670656 42062 670712
rect 42062 670656 42076 670712
rect 42012 670652 42076 670656
rect 42196 670108 42260 670172
rect 675892 665620 675956 665684
rect 40724 665348 40788 665412
rect 40540 664532 40604 664596
rect 42012 663368 42076 663372
rect 42012 663312 42062 663368
rect 42062 663312 42076 663368
rect 42012 663308 42076 663312
rect 676260 663308 676324 663372
rect 676996 663308 677060 663372
rect 676812 662900 676876 662964
rect 41460 661268 41524 661332
rect 42196 660512 42260 660516
rect 42196 660456 42210 660512
rect 42210 660456 42260 660512
rect 42196 660452 42260 660456
rect 41828 660316 41892 660380
rect 673868 659908 673932 659972
rect 41644 658276 41708 658340
rect 674420 652156 674484 652220
rect 675892 651476 675956 651540
rect 6150 650209 6854 651353
rect 54235 650245 55339 651349
rect 63339 650225 63883 651329
rect 7348 648613 8052 649757
rect 52641 648627 53745 649731
rect 62371 648617 62915 649721
rect 673316 649164 673380 649228
rect 676260 648620 676324 648684
rect 676628 644676 676692 644740
rect 676996 644540 677060 644604
rect 39988 642228 40052 642292
rect 39988 641412 40052 641476
rect 41460 640596 41524 640660
rect 675524 640384 675588 640388
rect 675524 640328 675538 640384
rect 675538 640328 675588 640384
rect 675524 640324 675588 640328
rect 675524 638148 675588 638212
rect 40908 636516 40972 636580
rect 40540 636108 40604 636172
rect 40724 634884 40788 634948
rect 675708 633388 675772 633452
rect 41828 629852 41892 629916
rect 42012 629172 42076 629236
rect 41644 629036 41708 629100
rect 42196 628900 42260 628964
rect 40908 625228 40972 625292
rect 40724 623732 40788 623796
rect 40540 621420 40604 621484
rect 676076 620740 676140 620804
rect 674604 619380 674668 619444
rect 42012 618972 42076 619036
rect 676444 618700 676508 618764
rect 41828 616796 41892 616860
rect 42196 616040 42260 616044
rect 42196 615984 42246 616040
rect 42246 615984 42260 616040
rect 42196 615980 42260 615984
rect 41460 614076 41524 614140
rect 41644 612716 41708 612780
rect 6150 607009 6854 608153
rect 54235 607045 55339 608149
rect 63339 607025 63883 608129
rect 675524 607880 675588 607884
rect 675524 607824 675538 607880
rect 675538 607824 675588 607880
rect 675524 607820 675588 607824
rect 7348 605413 8052 606557
rect 52641 605427 53745 606531
rect 62371 605417 62915 606521
rect 675340 606520 675404 606524
rect 675340 606464 675390 606520
rect 675390 606464 675404 606520
rect 675340 606460 675404 606464
rect 675340 605780 675404 605844
rect 675708 605780 675772 605844
rect 675708 600884 675772 600948
rect 675524 600264 675588 600268
rect 675524 600208 675574 600264
rect 675574 600208 675588 600264
rect 675524 600204 675588 600208
rect 39988 598980 40052 599044
rect 676444 598980 676508 599044
rect 39988 598164 40052 598228
rect 676812 597756 676876 597820
rect 41460 596532 41524 596596
rect 41644 594900 41708 594964
rect 675524 593192 675588 593196
rect 675524 593136 675538 593192
rect 675538 593136 675588 593192
rect 675524 593132 675588 593136
rect 675708 593192 675772 593196
rect 675708 593136 675722 593192
rect 675722 593136 675772 593192
rect 675708 593132 675772 593136
rect 40540 592044 40604 592108
rect 40724 591636 40788 591700
rect 676076 589188 676140 589252
rect 42380 585108 42444 585172
rect 41828 584216 41892 584220
rect 41828 584160 41842 584216
rect 41842 584160 41892 584216
rect 41828 584156 41892 584160
rect 42012 584216 42076 584220
rect 42012 584160 42026 584216
rect 42026 584160 42076 584216
rect 42012 584156 42076 584160
rect 42564 583612 42628 583676
rect 42012 582176 42076 582180
rect 42012 582120 42026 582176
rect 42026 582120 42076 582176
rect 42012 582116 42076 582120
rect 41828 580272 41892 580276
rect 41828 580216 41842 580272
rect 41842 580216 41892 580272
rect 41828 580212 41892 580216
rect 40724 578988 40788 579052
rect 40540 577492 40604 577556
rect 42196 576812 42260 576876
rect 42196 575860 42260 575924
rect 674420 574092 674484 574156
rect 41828 573684 41892 573748
rect 42012 572792 42076 572796
rect 42012 572736 42026 572792
rect 42026 572736 42076 572792
rect 42012 572732 42076 572736
rect 673316 572732 673380 572796
rect 676260 573140 676324 573204
rect 676996 573140 677060 573204
rect 676628 572732 676692 572796
rect 41460 571508 41524 571572
rect 41644 570420 41708 570484
rect 676996 568516 677060 568580
rect 6150 563809 6854 564953
rect 54235 563845 55339 564949
rect 63339 563825 63883 564929
rect 7348 562213 8052 563357
rect 52641 562227 53745 563331
rect 62371 562217 62915 563321
rect 675892 562668 675956 562732
rect 676076 561172 676140 561236
rect 675340 559540 675404 559604
rect 676260 558316 676324 558380
rect 39988 555868 40052 555932
rect 676628 551924 676692 551988
rect 40540 550564 40604 550628
rect 40724 549340 40788 549404
rect 40908 548932 40972 548996
rect 675524 546484 675588 546548
rect 41460 545124 41524 545188
rect 675708 543764 675772 543828
rect 41644 542948 41708 543012
rect 41828 542812 41892 542876
rect 42012 542268 42076 542332
rect 42012 535876 42076 535940
rect 40908 534516 40972 534580
rect 40724 533836 40788 533900
rect 41828 532612 41892 532676
rect 40540 530708 40604 530772
rect 676996 530164 677060 530228
rect 41460 529892 41524 529956
rect 41644 529348 41708 529412
rect 676812 528124 676876 528188
rect 676444 527716 676508 527780
rect 667329 514047 669713 518591
rect 667343 504057 669727 508601
rect 675892 503644 675956 503708
rect 675340 503508 675404 503572
rect 50356 493239 52100 497743
rect 50344 483249 52088 487753
rect 676076 487732 676140 487796
rect 676260 484570 676324 484634
rect 676076 483788 676140 483852
rect 6150 436209 6854 437353
rect 54235 436245 55339 437349
rect 63339 436225 63883 437329
rect 7348 434613 8052 435757
rect 52641 434627 53745 435731
rect 62371 434617 62915 435721
rect 42196 425988 42260 426052
rect 664125 425685 666549 430389
rect 41828 425580 41892 425644
rect 40724 425068 40788 425072
rect 40724 425012 40774 425068
rect 40774 425012 40788 425068
rect 40724 425008 40788 425012
rect 41828 423948 41892 424012
rect 42012 423540 42076 423604
rect 41828 422724 41892 422788
rect 30604 420868 30668 420932
rect 30604 418780 30668 418844
rect 41644 417964 41708 418028
rect 664108 415847 666532 420471
rect 41828 414564 41892 414628
rect 42380 411164 42444 411228
rect 41092 409396 41156 409460
rect 41644 406268 41708 406332
rect 41460 402460 41524 402524
rect 42012 401840 42076 401844
rect 42012 401784 42026 401840
rect 42026 401784 42076 401840
rect 42012 401780 42076 401784
rect 40724 400012 40788 400076
rect 40908 399604 40972 399668
rect 675708 399332 675772 399396
rect 40540 398788 40604 398852
rect 676260 398788 676324 398852
rect 676444 397156 676508 397220
rect 676076 395524 676140 395588
rect 675892 395252 675956 395316
rect 6150 393009 6854 394153
rect 54235 393045 55339 394149
rect 63339 393025 63883 394129
rect 7348 391413 8052 392557
rect 52641 391427 53745 392531
rect 62371 391417 62915 392521
rect 675524 388452 675588 388516
rect 675340 388180 675404 388244
rect 675708 384976 675772 384980
rect 675708 384920 675758 384976
rect 675758 384920 675772 384976
rect 675708 384916 675772 384920
rect 40724 383012 40788 383076
rect 40540 382196 40604 382260
rect 675340 382256 675404 382260
rect 675340 382200 675390 382256
rect 675390 382200 675404 382256
rect 675340 382196 675404 382200
rect 41460 381788 41524 381852
rect 40908 379748 40972 379812
rect 675524 378720 675588 378724
rect 675524 378664 675538 378720
rect 675538 378664 675588 378720
rect 675524 378660 675588 378664
rect 675892 377300 675956 377364
rect 676076 374988 676140 375052
rect 676260 373628 676324 373692
rect 676444 371996 676508 372060
rect 42012 371860 42076 371924
rect 41644 371316 41708 371380
rect 41828 370288 41892 370292
rect 41828 370232 41842 370288
rect 41842 370232 41892 370288
rect 41828 370228 41892 370232
rect 41828 366344 41892 366348
rect 41828 366288 41878 366344
rect 41878 366288 41892 366344
rect 41828 366284 41892 366288
rect 42012 363760 42076 363764
rect 42012 363704 42026 363760
rect 42026 363704 42076 363760
rect 42012 363700 42076 363704
rect 41644 362884 41708 362948
rect 40908 360164 40972 360228
rect 41460 358668 41524 358732
rect 40724 356900 40788 356964
rect 40540 355676 40604 355740
rect 675892 354180 675956 354244
rect 676076 353636 676140 353700
rect 675708 353364 675772 353428
rect 675340 352956 675404 353020
rect 676076 352004 676140 352068
rect 6150 349809 6854 350953
rect 54235 349845 55339 350949
rect 63339 350625 63883 351729
rect 7348 348213 8052 349357
rect 52641 348227 53745 349331
rect 62371 348217 62915 349321
rect 676996 346564 677060 346628
rect 676628 346428 676692 346492
rect 676812 346488 676876 346492
rect 676812 346432 676826 346488
rect 676826 346432 676876 346488
rect 676812 346428 676876 346432
rect 676076 342348 676140 342412
rect 675708 340776 675772 340780
rect 675708 340720 675722 340776
rect 675722 340720 675772 340776
rect 675708 340716 675772 340720
rect 40724 339764 40788 339828
rect 675892 339356 675956 339420
rect 40540 338948 40604 339012
rect 41460 338540 41524 338604
rect 675340 337860 675404 337924
rect 40908 337316 40972 337380
rect 41644 336908 41708 336972
rect 676996 335820 677060 335884
rect 41276 335684 41340 335748
rect 41092 335276 41156 335340
rect 676812 335276 676876 335340
rect 41828 334052 41892 334116
rect 676076 333508 676140 333572
rect 676628 332556 676692 332620
rect 42012 328340 42076 328404
rect 676444 325620 676508 325684
rect 676260 325484 676324 325548
rect 41828 324864 41892 324868
rect 41828 324808 41842 324864
rect 41842 324808 41892 324864
rect 41828 324804 41892 324808
rect 41276 321132 41340 321196
rect 42012 319968 42076 319972
rect 42012 319912 42026 319968
rect 42026 319912 42076 319968
rect 42012 319908 42076 319912
rect 41092 317324 41156 317388
rect 41644 315828 41708 315892
rect 41460 315420 41524 315484
rect 40724 313788 40788 313852
rect 40908 313108 40972 313172
rect 40540 312292 40604 312356
rect 676444 308620 676508 308684
rect 6150 306609 6854 307753
rect 54235 306645 55339 307749
rect 63339 306625 63883 307729
rect 676076 307396 676140 307460
rect 676260 306988 676324 307052
rect 7348 305013 8052 306157
rect 52641 305027 53745 306131
rect 62371 305017 62915 306121
rect 676628 304948 676692 305012
rect 675892 299372 675956 299436
rect 675708 297740 675772 297804
rect 675340 297468 675404 297532
rect 675524 297332 675588 297396
rect 42380 296788 42444 296852
rect 41828 295972 41892 296036
rect 42196 295564 42260 295628
rect 42012 295156 42076 295220
rect 675892 294748 675956 294812
rect 41828 294340 41892 294404
rect 41828 293932 41892 293996
rect 675708 292632 675772 292636
rect 41460 292528 41524 292592
rect 675708 292576 675722 292632
rect 675722 292576 675772 292632
rect 675708 292572 675772 292576
rect 675524 292088 675588 292092
rect 675524 292032 675538 292088
rect 675538 292032 675588 292088
rect 675524 292028 675588 292032
rect 676076 288356 676140 288420
rect 41828 288084 41892 288148
rect 41828 287812 41892 287876
rect 676628 287268 676692 287332
rect 675340 285500 675404 285564
rect 41644 284956 41708 285020
rect 42012 284956 42076 285020
rect 41460 284820 41524 284884
rect 676444 283596 676508 283660
rect 41460 281420 41524 281484
rect 676260 281420 676324 281484
rect 40908 278700 40972 278764
rect 40908 277340 40972 277404
rect 41828 276720 41892 276724
rect 41828 276664 41842 276720
rect 41842 276664 41892 276720
rect 41828 276660 41892 276664
rect 41644 272308 41708 272372
rect 42012 270464 42076 270468
rect 42012 270408 42026 270464
rect 42026 270408 42076 270464
rect 42012 270404 42076 270408
rect 40724 269724 40788 269788
rect 40540 269044 40604 269108
rect 6150 263409 6854 264553
rect 54235 263445 55339 264549
rect 675892 264148 675956 264212
rect 676996 263570 677060 263634
rect 7348 261813 8052 262957
rect 52641 261827 53745 262931
rect 675708 262924 675772 262988
rect 677180 261972 677244 262036
rect 677364 261564 677428 261628
rect 676076 260340 676140 260404
rect 42196 253540 42260 253604
rect 41828 253132 41892 253196
rect 40540 252588 40604 252652
rect 674788 252588 674852 252652
rect 41644 252180 41708 252244
rect 676444 251500 676508 251564
rect 677364 251500 677428 251564
rect 676444 250276 676508 250340
rect 40172 249732 40236 249796
rect 674788 249732 674852 249796
rect 675892 249732 675956 249796
rect 673868 249656 673932 249660
rect 673868 249600 673882 249656
rect 673882 249600 673932 249656
rect 673868 249596 673932 249600
rect 675708 249596 675772 249660
rect 676076 249596 676140 249660
rect 40356 249324 40420 249388
rect 39988 248916 40052 248980
rect 674972 246196 675036 246260
rect 675340 246196 675404 246260
rect 673868 246120 673932 246124
rect 673868 246064 673882 246120
rect 673882 246064 673932 246120
rect 673868 246060 673932 246064
rect 42196 245788 42260 245852
rect 41828 245652 41892 245716
rect 39988 244624 40052 244628
rect 39988 244568 40038 244624
rect 40038 244568 40052 244624
rect 39988 244564 40052 244568
rect 40172 244156 40236 244220
rect 674972 241844 675036 241908
rect 675340 240272 675404 240276
rect 675340 240216 675390 240272
rect 675390 240216 675404 240272
rect 675340 240212 675404 240216
rect 40724 238988 40788 239052
rect 40356 238444 40420 238508
rect 40540 238172 40604 238236
rect 676996 238444 677060 238508
rect 41092 238036 41156 238100
rect 41276 238036 41340 238100
rect 41460 238036 41524 238100
rect 41644 238036 41708 238100
rect 42196 238036 42260 238100
rect 42564 237900 42628 237964
rect 677180 236812 677244 236876
rect 40540 236676 40604 236740
rect 41276 234772 41340 234836
rect 41460 233276 41524 233340
rect 40724 230420 40788 230484
rect 647740 230420 647804 230484
rect 42564 229876 42628 229940
rect 41644 228924 41708 228988
rect 42196 227292 42260 227356
rect 40540 226068 40604 226132
rect 6150 220209 6854 221353
rect 54235 220245 55339 221349
rect 7348 218613 8052 219757
rect 52641 218627 53745 219731
rect 676030 218588 676094 218652
rect 675340 218180 675404 218244
rect 675892 217772 675956 217836
rect 676076 216820 676140 216884
rect 676996 214270 677060 214334
rect 675708 213964 675772 214028
rect 647740 213012 647804 213076
rect 676628 211380 676692 211444
rect 676812 211244 676876 211308
rect 40540 209340 40604 209404
rect 41460 208524 41524 208588
rect 676076 208252 676140 208316
rect 675524 207164 675588 207228
rect 40724 206892 40788 206956
rect 675340 205592 675404 205596
rect 675340 205536 675390 205592
rect 675390 205536 675404 205592
rect 675340 205532 675404 205536
rect 676076 204988 676140 205052
rect 675708 204232 675772 204236
rect 675708 204176 675758 204232
rect 675758 204176 675772 204232
rect 675708 204172 675772 204176
rect 676996 202812 677060 202876
rect 675892 202676 675956 202740
rect 676812 201316 676876 201380
rect 41644 199412 41708 199476
rect 41828 199276 41892 199340
rect 675524 198384 675588 198388
rect 675524 198328 675538 198384
rect 675538 198328 675588 198384
rect 675524 198324 675588 198328
rect 676628 195332 676692 195396
rect 41644 195196 41708 195260
rect 40724 194652 40788 194716
rect 41828 194652 41892 194716
rect 676260 190300 676324 190364
rect 41460 190164 41524 190228
rect 676444 190164 676508 190228
rect 41828 187368 41892 187372
rect 41828 187312 41842 187368
rect 41842 187312 41892 187368
rect 41828 187308 41892 187312
rect 41644 184044 41708 184108
rect 40540 182956 40604 183020
rect 676076 173436 676140 173500
rect 675892 172756 675956 172820
rect 676076 171804 676140 171868
rect 673868 168540 673932 168604
rect 676628 166424 676692 166428
rect 676628 166368 676642 166424
rect 676642 166368 676692 166424
rect 676628 166364 676692 166368
rect 676812 166424 676876 166428
rect 676812 166368 676862 166424
rect 676862 166368 676876 166424
rect 676812 166364 676876 166368
rect 675524 162692 675588 162756
rect 675892 162556 675956 162620
rect 675708 162420 675772 162484
rect 675340 162284 675404 162348
rect 676812 159972 676876 160036
rect 675892 159428 675956 159492
rect 676076 157388 676140 157452
rect 675708 157040 675772 157044
rect 675708 156984 675722 157040
rect 675722 156984 675772 157040
rect 675708 156980 675772 156984
rect 675524 156496 675588 156500
rect 675524 156440 675574 156496
rect 675574 156440 675588 156496
rect 675524 156436 675588 156440
rect 675340 153096 675404 153100
rect 675340 153040 675390 153096
rect 675390 153040 675404 153096
rect 675340 153036 675404 153040
rect 676628 151540 676692 151604
rect 676444 148412 676508 148476
rect 676260 146236 676324 146300
rect 676076 128556 676140 128620
rect 676260 126516 676324 126580
rect 675892 124884 675956 124948
rect 676444 124476 676508 124540
rect 676812 121620 676876 121684
rect 675708 117948 675772 118012
rect 675340 117268 675404 117332
rect 675524 117132 675588 117196
rect 676076 114140 676140 114204
rect 675892 112508 675956 112572
rect 675524 111752 675588 111756
rect 675524 111696 675538 111752
rect 675538 111696 675588 111752
rect 675524 111692 675588 111696
rect 676444 108972 676508 109036
rect 675708 108216 675772 108220
rect 675708 108160 675758 108216
rect 675758 108160 675772 108216
rect 675708 108156 675772 108160
rect 675340 104756 675404 104820
rect 676812 103124 676876 103188
rect 676260 101356 676324 101420
rect 641668 96656 641732 96660
rect 641668 96600 641718 96656
rect 641718 96600 641732 96656
rect 641668 96596 641732 96600
rect 639828 96460 639892 96524
rect 41937 78242 45681 82706
rect 634676 77828 634740 77892
rect 639828 77692 639892 77756
rect 638908 75108 638972 75172
rect 41913 68338 45657 72802
rect 638908 51716 638972 51780
rect 520228 50492 520292 50556
rect 521700 50356 521764 50420
rect 514708 50220 514772 50284
rect 529796 50220 529860 50284
rect 187556 44916 187620 44980
rect 194364 44780 194428 44844
rect 141924 43964 141988 44028
rect 241731 42837 245995 46621
rect 187556 42120 187620 42124
rect 187556 42064 187570 42120
rect 187570 42064 187620 42120
rect 187556 42060 187620 42064
rect 194364 42120 194428 42124
rect 194364 42064 194378 42120
rect 194378 42064 194428 42120
rect 194364 42060 194428 42064
rect 141924 40292 141988 40356
rect 251383 42851 255647 46635
rect 648155 47120 649619 47124
rect 648155 46664 648159 47120
rect 648159 46664 649615 47120
rect 649615 46664 649619 47120
rect 648155 46660 649619 46664
rect 518572 46548 518636 46612
rect 471652 46412 471716 46476
rect 365116 45188 365180 45252
rect 310100 45052 310164 45116
rect 525932 44644 525996 44708
rect 310100 42392 310164 42396
rect 310100 42336 310104 42392
rect 310104 42336 310160 42392
rect 310160 42336 310164 42392
rect 310100 42332 310164 42336
rect 518572 42392 518636 42396
rect 518572 42336 518622 42392
rect 518622 42336 518636 42392
rect 518572 42332 518636 42336
rect 365116 42120 365180 42124
rect 365116 42064 365130 42120
rect 365130 42064 365180 42120
rect 365116 42060 365180 42064
rect 471652 42120 471716 42124
rect 471652 42064 471666 42120
rect 471666 42064 471716 42120
rect 471652 42060 471716 42064
rect 514708 42060 514772 42124
rect 520228 42060 520292 42124
rect 521700 42120 521764 42124
rect 521700 42064 521750 42120
rect 521750 42064 521764 42120
rect 521700 42060 521764 42064
rect 525932 42120 525996 42124
rect 525932 42064 525982 42120
rect 525982 42064 525996 42120
rect 525932 42060 525996 42064
rect 529796 42060 529860 42124
<< metal4 >>
rect 99346 1030812 99391 1031612
rect 99787 1030812 102778 1031612
rect 103174 1030812 106148 1031612
rect 106544 1031568 116070 1031612
rect 106544 1030864 114809 1031568
rect 115953 1030864 116070 1031568
rect 106544 1030812 116070 1030864
rect 150746 1030812 150791 1031612
rect 151187 1030812 154178 1031612
rect 154574 1030812 157548 1031612
rect 157944 1031568 167470 1031612
rect 157944 1030864 166209 1031568
rect 167353 1030864 167470 1031568
rect 157944 1030812 167470 1030864
rect 202146 1030812 202191 1031612
rect 202587 1030812 205578 1031612
rect 205974 1030812 208948 1031612
rect 209344 1031568 218870 1031612
rect 209344 1030864 217609 1031568
rect 218753 1030864 218870 1031568
rect 209344 1030812 218870 1030864
rect 253546 1030812 253591 1031612
rect 253987 1030812 256978 1031612
rect 257374 1030812 260348 1031612
rect 260744 1031568 270270 1031612
rect 260744 1030864 269009 1031568
rect 270153 1030864 270270 1031568
rect 260744 1030812 270270 1030864
rect 305146 1030812 305191 1031612
rect 305587 1030812 308578 1031612
rect 308974 1030812 311948 1031612
rect 312344 1031568 321870 1031612
rect 312344 1030864 320609 1031568
rect 321753 1030864 321870 1031568
rect 312344 1030812 321870 1030864
rect 355546 1030812 355591 1031612
rect 355987 1030812 358978 1031612
rect 359374 1030812 362348 1031612
rect 362744 1031568 372270 1031612
rect 362744 1030864 371009 1031568
rect 372153 1030864 372270 1031568
rect 362744 1030812 372270 1030864
rect 422946 1030812 422991 1031612
rect 423387 1030812 426378 1031612
rect 426774 1030812 429748 1031612
rect 430144 1031568 439670 1031612
rect 430144 1030864 438409 1031568
rect 439553 1030864 439670 1031568
rect 430144 1030812 439670 1030864
rect 499946 1030812 499991 1031612
rect 500387 1030812 503378 1031612
rect 503774 1030812 506748 1031612
rect 507144 1031568 516670 1031612
rect 507144 1030864 515409 1031568
rect 516553 1030864 516670 1031568
rect 507144 1030812 516670 1030864
rect 551346 1030812 551391 1031612
rect 551787 1030812 554778 1031612
rect 555174 1030812 558148 1031612
rect 558544 1031568 568070 1031612
rect 558544 1030864 566809 1031568
rect 567953 1030864 568070 1031568
rect 558544 1030812 568070 1030864
rect 101076 1029612 101079 1030412
rect 101475 1029612 104462 1030412
rect 104858 1029612 107838 1030412
rect 108234 1030370 114442 1030412
rect 108234 1029666 113213 1030370
rect 114357 1029666 114442 1030370
rect 108234 1029612 114442 1029666
rect 152476 1029612 152479 1030412
rect 152875 1029612 155862 1030412
rect 156258 1029612 159238 1030412
rect 159634 1030370 165842 1030412
rect 159634 1029666 164613 1030370
rect 165757 1029666 165842 1030370
rect 159634 1029612 165842 1029666
rect 203876 1029612 203879 1030412
rect 204275 1029612 207262 1030412
rect 207658 1029612 210638 1030412
rect 211034 1030370 217242 1030412
rect 211034 1029666 216013 1030370
rect 217157 1029666 217242 1030370
rect 211034 1029612 217242 1029666
rect 255276 1029612 255279 1030412
rect 255675 1029612 258662 1030412
rect 259058 1029612 262038 1030412
rect 262434 1030370 268642 1030412
rect 262434 1029666 267413 1030370
rect 268557 1029666 268642 1030370
rect 262434 1029612 268642 1029666
rect 306876 1029612 306879 1030412
rect 307275 1029612 310262 1030412
rect 310658 1029612 313638 1030412
rect 314034 1030370 320242 1030412
rect 314034 1029666 319013 1030370
rect 320157 1029666 320242 1030370
rect 314034 1029612 320242 1029666
rect 357276 1029612 357279 1030412
rect 357675 1029612 360662 1030412
rect 361058 1029612 364038 1030412
rect 364434 1030370 370642 1030412
rect 364434 1029666 369413 1030370
rect 370557 1029666 370642 1030370
rect 364434 1029612 370642 1029666
rect 424676 1029612 424679 1030412
rect 425075 1029612 428062 1030412
rect 428458 1029612 431438 1030412
rect 431834 1030370 438042 1030412
rect 431834 1029666 436813 1030370
rect 437957 1029666 438042 1030370
rect 431834 1029612 438042 1029666
rect 501676 1029612 501679 1030412
rect 502075 1029612 505062 1030412
rect 505458 1029612 508438 1030412
rect 508834 1030370 515042 1030412
rect 508834 1029666 513813 1030370
rect 514957 1029666 515042 1030370
rect 508834 1029612 515042 1029666
rect 553076 1029612 553079 1030412
rect 553475 1029612 556462 1030412
rect 556858 1029612 559838 1030412
rect 560234 1030370 566442 1030412
rect 560234 1029666 565213 1030370
rect 566357 1029666 566442 1030370
rect 560234 1029612 566442 1029666
rect 383699 997796 383765 997797
rect 383699 997732 383700 997796
rect 383764 997732 383765 997796
rect 383699 997731 383765 997732
rect 85251 997252 85317 997253
rect 85251 997188 85252 997252
rect 85316 997188 85317 997252
rect 85251 997187 85317 997188
rect 84699 996980 84765 996981
rect 84699 996916 84700 996980
rect 84764 996916 84765 996980
rect 84699 996915 84765 996916
rect 84702 995621 84762 996915
rect 85254 995621 85314 997187
rect 292435 997116 292501 997117
rect 84699 995620 84765 995621
rect 84699 995556 84700 995620
rect 84764 995556 84765 995620
rect 84699 995555 84765 995556
rect 85251 995620 85317 995621
rect 85251 995556 85252 995620
rect 85316 995556 85317 995620
rect 85251 995555 85317 995556
rect 88934 995485 88994 997102
rect 113174 996723 114388 996738
rect 113174 995532 113181 996723
rect 114377 995532 114388 996723
rect 88931 995484 88997 995485
rect 88931 995420 88932 995484
rect 88996 995420 88997 995484
rect 88931 995419 88997 995420
rect 114510 990997 114570 997102
rect 292435 997052 292436 997116
rect 292500 997052 292501 997116
rect 292435 997051 292501 997052
rect 164574 996723 165788 996738
rect 136771 996164 136837 996165
rect 136771 996100 136772 996164
rect 136836 996100 136837 996164
rect 136771 996099 136837 996100
rect 114774 995129 115988 995134
rect 114774 993933 114799 995129
rect 136774 995077 136834 996099
rect 164574 995532 164581 996723
rect 165777 995532 165788 996723
rect 215974 996723 217188 996738
rect 215974 995532 215981 996723
rect 217177 995532 217188 996723
rect 267374 996723 268588 996738
rect 243859 996436 243925 996437
rect 243859 996372 243860 996436
rect 243924 996372 243925 996436
rect 243859 996371 243925 996372
rect 243862 995757 243922 996371
rect 243859 995756 243925 995757
rect 243859 995692 243860 995756
rect 243924 995692 243925 995756
rect 243859 995691 243925 995692
rect 267374 995532 267381 996723
rect 268577 995532 268588 996723
rect 292438 995485 292498 997051
rect 318974 996723 320188 996738
rect 318974 995532 318981 996723
rect 320177 995532 320188 996723
rect 369374 996723 370588 996738
rect 369374 995532 369381 996723
rect 370577 995532 370588 996723
rect 383702 996029 383762 997731
rect 436774 996723 437988 996738
rect 387563 996300 387629 996301
rect 387563 996236 387564 996300
rect 387628 996236 387629 996300
rect 387563 996235 387629 996236
rect 383699 996028 383765 996029
rect 383699 995964 383700 996028
rect 383764 995964 383765 996028
rect 383699 995963 383765 995964
rect 292435 995484 292501 995485
rect 292435 995420 292436 995484
rect 292500 995420 292501 995484
rect 292435 995419 292501 995420
rect 166174 995129 167388 995134
rect 217574 995129 218788 995134
rect 268974 995129 270188 995134
rect 320574 995129 321788 995134
rect 370974 995129 372188 995134
rect 136771 995076 136837 995077
rect 136771 995012 136772 995076
rect 136836 995012 136837 995076
rect 136771 995011 136837 995012
rect 166174 993933 166199 995129
rect 217574 993933 217599 995129
rect 268974 993933 268999 995129
rect 320574 993933 320599 995129
rect 370974 993933 370999 995129
rect 387566 995077 387626 996235
rect 390323 996164 390389 996165
rect 390323 996100 390324 996164
rect 390388 996100 390389 996164
rect 390323 996099 390389 996100
rect 389035 995892 389101 995893
rect 389035 995828 389036 995892
rect 389100 995890 389101 995892
rect 389403 995892 389469 995893
rect 389403 995890 389404 995892
rect 389100 995830 389404 995890
rect 389100 995828 389101 995830
rect 389035 995827 389101 995828
rect 389403 995828 389404 995830
rect 389468 995828 389469 995892
rect 389403 995827 389469 995828
rect 390326 995757 390386 996099
rect 390323 995756 390389 995757
rect 390323 995692 390324 995756
rect 390388 995692 390389 995756
rect 390323 995691 390389 995692
rect 436774 995532 436781 996723
rect 437977 995532 437988 996723
rect 485638 995757 485698 997102
rect 506430 995893 506490 997102
rect 575680 997067 580478 997130
rect 513774 996723 514988 996738
rect 506427 995892 506493 995893
rect 506427 995828 506428 995892
rect 506492 995828 506493 995892
rect 506427 995827 506493 995828
rect 485635 995756 485701 995757
rect 485635 995692 485636 995756
rect 485700 995692 485701 995756
rect 485635 995691 485701 995692
rect 513774 995532 513781 996723
rect 514977 995532 514988 996723
rect 565174 996723 566388 996738
rect 565174 995532 565181 996723
rect 566377 995532 566388 996723
rect 438374 995129 439588 995134
rect 515374 995129 516588 995134
rect 566774 995129 567988 995134
rect 387563 995076 387629 995077
rect 387563 995012 387564 995076
rect 387628 995012 387629 995076
rect 387563 995011 387629 995012
rect 438374 993933 438399 995129
rect 515374 993933 515399 995129
rect 566774 993933 566799 995129
rect 575680 995123 575774 997067
rect 580398 995123 580478 997067
rect 114774 993928 115988 993933
rect 166174 993928 167388 993933
rect 217574 993928 218788 993933
rect 268974 993928 270188 993933
rect 320574 993928 321788 993933
rect 370974 993928 372188 993933
rect 438374 993928 439588 993933
rect 515374 993928 516588 993933
rect 566774 993928 567988 993933
rect 575680 993337 580478 995123
rect 114507 990996 114573 990997
rect 114507 990932 114508 990996
rect 114572 990932 114573 990996
rect 114507 990931 114573 990932
rect 575680 990861 575715 993337
rect 580431 990861 580478 993337
rect 575680 990788 580478 990861
rect 585670 997073 590468 997144
rect 585670 995129 585744 997073
rect 590368 995129 590468 997073
rect 670816 996692 673426 996696
rect 670808 996624 676654 996692
rect 670808 995588 670876 996624
rect 676552 995588 676654 996624
rect 670808 995492 676654 995588
rect 585670 993351 590468 995129
rect 585670 990875 585711 993351
rect 590427 990875 590468 993351
rect 585670 990802 590468 990875
rect 670816 992520 673426 995492
rect 670816 990364 670962 992520
rect 673278 990364 673426 992520
rect 47796 990286 56582 990310
rect 47796 990285 55829 990286
rect 49790 989730 55829 990285
rect 56385 989730 56582 990286
rect 670816 990200 673426 990364
rect 49790 989729 56582 989730
rect 47796 989692 56582 989729
rect 50194 989326 56434 989348
rect 50194 989321 55833 989326
rect 50194 988765 50200 989321
rect 52196 988770 55833 989321
rect 56389 988770 56434 989326
rect 52196 988765 56434 988770
rect 50194 988736 56434 988765
rect 658380 987407 669826 987436
rect 658380 987402 667281 987407
rect 658380 986846 658417 987402
rect 663133 986851 667281 987402
rect 669757 986851 669826 987407
rect 663133 986846 669826 986851
rect 658380 986812 669826 986846
rect 52596 984517 56404 984548
rect 52596 983961 52599 984517
rect 53795 983961 55811 984517
rect 56367 983961 56404 984517
rect 52596 983928 56404 983961
rect 40539 968828 40605 968829
rect 40539 968764 40540 968828
rect 40604 968764 40605 968828
rect 40539 968763 40605 968764
rect 6106 949953 6906 950070
rect 6106 948809 6150 949953
rect 6854 948809 6906 949953
rect 6106 940543 6906 948809
rect 7306 948357 8106 948442
rect 7306 947213 7348 948357
rect 8052 947213 8106 948357
rect 7306 942235 8106 947213
rect 6106 937177 6906 940147
rect 7306 938855 8106 941839
rect 6106 933787 6906 936781
rect 7306 935475 8106 938459
rect 40542 936050 40602 968763
rect 40723 967332 40789 967333
rect 40723 967268 40724 967332
rect 40788 967268 40789 967332
rect 40723 967267 40789 967268
rect 40726 943805 40786 967267
rect 676443 966516 676509 966517
rect 676443 966452 676444 966516
rect 676508 966452 676509 966516
rect 676443 966451 676509 966452
rect 676259 966244 676325 966245
rect 676259 966180 676260 966244
rect 676324 966180 676325 966244
rect 676259 966179 676325 966180
rect 41643 965156 41709 965157
rect 41643 965092 41644 965156
rect 41708 965092 41709 965156
rect 41643 965091 41709 965092
rect 40907 963524 40973 963525
rect 40907 963460 40908 963524
rect 40972 963460 40973 963524
rect 40907 963459 40973 963460
rect 40723 943804 40789 943805
rect 40723 943740 40724 943804
rect 40788 943740 40789 943804
rect 40723 943739 40789 943740
rect 40910 937050 40970 963459
rect 41459 957812 41525 957813
rect 41459 957748 41460 957812
rect 41524 957748 41525 957812
rect 41459 957747 41525 957748
rect 41462 943950 41522 957747
rect 41646 952237 41706 965091
rect 676075 963388 676141 963389
rect 676075 963324 676076 963388
rect 676140 963324 676141 963388
rect 676075 963323 676141 963324
rect 675707 962844 675773 962845
rect 675707 962780 675708 962844
rect 675772 962780 675773 962844
rect 675707 962779 675773 962780
rect 41827 962164 41893 962165
rect 41827 962100 41828 962164
rect 41892 962100 41893 962164
rect 41827 962099 41893 962100
rect 41830 952917 41890 962099
rect 675523 961892 675589 961893
rect 675523 961828 675524 961892
rect 675588 961828 675589 961892
rect 675523 961827 675589 961828
rect 42011 958492 42077 958493
rect 42011 958428 42012 958492
rect 42076 958428 42077 958492
rect 42011 958427 42077 958428
rect 41827 952916 41893 952917
rect 41827 952852 41828 952916
rect 41892 952852 41893 952916
rect 41827 952851 41893 952852
rect 42014 952373 42074 958427
rect 675339 954004 675405 954005
rect 675339 953940 675340 954004
rect 675404 953940 675405 954004
rect 675339 953939 675405 953940
rect 42011 952372 42077 952373
rect 42011 952308 42012 952372
rect 42076 952308 42077 952372
rect 42011 952307 42077 952308
rect 41643 952236 41709 952237
rect 41643 952172 41644 952236
rect 41708 952172 41709 952236
rect 41643 952171 41709 952172
rect 54184 948799 54189 949988
rect 55385 948799 55390 949988
rect 63350 949629 63872 949632
rect 54184 948774 55390 948799
rect 675342 949517 675402 953939
rect 675526 949653 675586 961827
rect 675710 949789 675770 962779
rect 675891 959172 675957 959173
rect 675891 959108 675892 959172
rect 675956 959108 675957 959172
rect 675891 959107 675957 959108
rect 675707 949788 675773 949789
rect 675707 949724 675708 949788
rect 675772 949724 675773 949788
rect 675707 949723 675773 949724
rect 675523 949652 675589 949653
rect 675523 949588 675524 949652
rect 675588 949588 675589 949652
rect 675523 949587 675589 949588
rect 675339 949516 675405 949517
rect 675339 949452 675340 949516
rect 675404 949452 675405 949516
rect 675339 949451 675405 949452
rect 63350 948522 63872 948525
rect 52580 948377 53786 948388
rect 52580 947181 52595 948377
rect 62382 948121 62904 948124
rect 52580 947174 53786 947181
rect 62382 947014 62904 947017
rect 41462 943890 42074 943950
rect 42014 937821 42074 943890
rect 42011 937820 42077 937821
rect 42011 937756 42012 937820
rect 42076 937756 42077 937820
rect 42011 937755 42077 937756
rect 40910 936990 42074 937050
rect 41827 936868 41893 936869
rect 41827 936866 41828 936868
rect 41462 936806 41828 936866
rect 41462 936050 41522 936806
rect 41827 936804 41828 936806
rect 41892 936804 41893 936868
rect 41827 936803 41893 936804
rect 40542 935990 41522 936050
rect 7306 935076 8106 935079
rect 42014 934965 42074 936990
rect 42011 934964 42077 934965
rect 42011 934900 42012 934964
rect 42076 934900 42077 934964
rect 42011 934899 42077 934900
rect 675894 933877 675954 959107
rect 676078 934013 676138 963323
rect 676262 934290 676322 966179
rect 676446 934829 676506 966451
rect 676627 965020 676693 965021
rect 676627 964956 676628 965020
rect 676692 964956 676693 965020
rect 676627 964955 676693 964956
rect 676630 935645 676690 964955
rect 676811 957948 676877 957949
rect 676811 957884 676812 957948
rect 676876 957884 676877 957948
rect 676811 957883 676877 957884
rect 676627 935644 676693 935645
rect 676627 935580 676628 935644
rect 676692 935580 676693 935644
rect 676627 935579 676693 935580
rect 676443 934828 676509 934829
rect 676443 934764 676444 934828
rect 676508 934764 676509 934828
rect 676443 934763 676509 934764
rect 676262 934230 676690 934290
rect 676075 934012 676141 934013
rect 676075 933948 676076 934012
rect 676140 933948 676141 934012
rect 676075 933947 676141 933948
rect 675891 933876 675957 933877
rect 675891 933812 675892 933876
rect 675956 933812 675957 933876
rect 675891 933811 675957 933812
rect 6106 933346 6906 933391
rect 676630 933197 676690 934230
rect 676627 933196 676693 933197
rect 676627 933132 676628 933196
rect 676692 933132 676693 933196
rect 676627 933131 676693 933132
rect 676814 931157 676874 957883
rect 676995 957676 677061 957677
rect 676995 957612 676996 957676
rect 677060 957612 677061 957676
rect 676995 957611 677061 957612
rect 676998 931565 677058 957611
rect 676995 931564 677061 931565
rect 676995 931500 676996 931564
rect 677060 931500 677061 931564
rect 676995 931499 677061 931500
rect 676811 931156 676877 931157
rect 676811 931092 676812 931156
rect 676876 931092 676877 931156
rect 676811 931091 676877 931092
rect 675155 877300 675221 877301
rect 675155 877236 675156 877300
rect 675220 877236 675221 877300
rect 675155 877235 675221 877236
rect 47792 842340 49822 842462
rect 47792 837784 47883 842340
rect 49719 837784 49822 842340
rect 47792 837658 49822 837784
rect 667202 833210 669802 833310
rect 667202 833196 667276 833210
rect 669740 833196 669802 833210
rect 47792 832408 49822 832506
rect 47792 827852 47883 832408
rect 49719 827852 49822 832408
rect 667202 828640 667270 833196
rect 669746 828640 669802 833196
rect 667202 828626 667276 828640
rect 669740 828626 669802 828640
rect 667202 828520 669802 828626
rect 47792 827702 49822 827852
rect 6106 824153 6906 824270
rect 6106 823009 6150 824153
rect 6854 823009 6906 824153
rect 6106 814743 6906 823009
rect 54184 822999 54189 824188
rect 55385 822999 55390 824188
rect 63350 824129 63872 824132
rect 667214 823216 669814 823336
rect 667214 823202 667262 823216
rect 669726 823202 669814 823216
rect 63350 823022 63872 823025
rect 54184 822974 55390 822999
rect 7306 822557 8106 822642
rect 7306 821413 7348 822557
rect 8052 821413 8106 822557
rect 7306 816435 8106 821413
rect 52580 822577 53786 822588
rect 52580 821381 52595 822577
rect 62382 822521 62904 822524
rect 62382 821414 62904 821417
rect 52580 821374 53786 821381
rect 667214 818646 667256 823202
rect 669732 818646 669814 823202
rect 667214 818632 667262 818646
rect 669726 818632 669814 818646
rect 667214 818546 669814 818632
rect 42011 816100 42077 816101
rect 6106 811377 6906 814347
rect 7306 813055 8106 816039
rect 42011 816036 42012 816100
rect 42076 816036 42077 816100
rect 42011 816035 42077 816036
rect 41827 814468 41893 814469
rect 41827 814404 41828 814468
rect 41892 814404 41893 814468
rect 41827 814403 41893 814404
rect 41830 813650 41890 814403
rect 39990 813590 41890 813650
rect 6106 807987 6906 810981
rect 7306 809675 8106 812659
rect 7306 809276 8106 809279
rect 6106 807546 6906 807591
rect 6106 780953 6906 781070
rect 6106 779809 6150 780953
rect 6854 779809 6906 780953
rect 6106 771543 6906 779809
rect 7306 779357 8106 779442
rect 7306 778213 7348 779357
rect 8052 778213 8106 779357
rect 7306 773235 8106 778213
rect 6106 768177 6906 771147
rect 7306 769855 8106 772839
rect 39990 771901 40050 813590
rect 42014 812290 42074 816035
rect 40174 812230 42074 812290
rect 40174 773533 40234 812230
rect 42195 812020 42261 812021
rect 42195 811956 42196 812020
rect 42260 811956 42261 812020
rect 42195 811955 42261 811956
rect 41827 807940 41893 807941
rect 41827 807876 41828 807940
rect 41892 807876 41893 807940
rect 41827 807875 41893 807876
rect 41830 807530 41890 807875
rect 40542 807470 41890 807530
rect 40542 796789 40602 807470
rect 41643 802636 41709 802637
rect 41643 802572 41644 802636
rect 41708 802572 41709 802636
rect 41643 802571 41709 802572
rect 41459 801004 41525 801005
rect 41459 800940 41460 801004
rect 41524 800940 41525 801004
rect 41459 800939 41525 800940
rect 40539 796788 40605 796789
rect 40539 796724 40540 796788
rect 40604 796724 40605 796788
rect 40539 796723 40605 796724
rect 41462 788221 41522 800939
rect 41459 788220 41525 788221
rect 41459 788156 41460 788220
rect 41524 788156 41525 788220
rect 41459 788155 41525 788156
rect 41646 786181 41706 802571
rect 42011 802500 42077 802501
rect 42011 802436 42012 802500
rect 42076 802436 42077 802500
rect 42011 802435 42077 802436
rect 41827 801684 41893 801685
rect 41827 801620 41828 801684
rect 41892 801620 41893 801684
rect 41827 801619 41893 801620
rect 41830 788085 41890 801619
rect 42014 792029 42074 802435
rect 42011 792028 42077 792029
rect 42011 791964 42012 792028
rect 42076 791964 42077 792028
rect 42011 791963 42077 791964
rect 42198 791893 42258 811955
rect 42195 791892 42261 791893
rect 42195 791828 42196 791892
rect 42260 791828 42261 791892
rect 42195 791827 42261 791828
rect 41827 788084 41893 788085
rect 41827 788020 41828 788084
rect 41892 788020 41893 788084
rect 41827 788019 41893 788020
rect 41643 786180 41709 786181
rect 41643 786116 41644 786180
rect 41708 786116 41709 786180
rect 41643 786115 41709 786116
rect 675158 784277 675218 877235
rect 676259 876620 676325 876621
rect 676259 876556 676260 876620
rect 676324 876556 676325 876620
rect 676259 876555 676325 876556
rect 676075 875940 676141 875941
rect 676075 875876 676076 875940
rect 676140 875876 676141 875940
rect 676075 875875 676141 875876
rect 675891 874036 675957 874037
rect 675891 873972 675892 874036
rect 675956 873972 675957 874036
rect 675891 873971 675957 873972
rect 675707 864788 675773 864789
rect 675707 864724 675708 864788
rect 675772 864724 675773 864788
rect 675707 864723 675773 864724
rect 675710 785229 675770 864723
rect 675707 785228 675773 785229
rect 675707 785164 675708 785228
rect 675772 785164 675773 785228
rect 675707 785163 675773 785164
rect 675894 785090 675954 873971
rect 675342 785030 675954 785090
rect 675155 784276 675221 784277
rect 675155 784212 675156 784276
rect 675220 784212 675221 784276
rect 675155 784211 675221 784212
rect 63350 782129 63872 782132
rect 63350 781022 63872 781025
rect 54184 779799 54189 780988
rect 55385 779799 55390 780988
rect 54184 779774 55390 779799
rect 52580 779377 53786 779388
rect 52580 778181 52595 779377
rect 62382 779321 62904 779324
rect 62382 778214 62904 778217
rect 52580 778174 53786 778181
rect 675155 775708 675221 775709
rect 675155 775644 675156 775708
rect 675220 775644 675221 775708
rect 675155 775643 675221 775644
rect 40171 773532 40237 773533
rect 40171 773468 40172 773532
rect 40236 773468 40237 773532
rect 40171 773467 40237 773468
rect 39987 771900 40053 771901
rect 39987 771836 39988 771900
rect 40052 771836 40053 771900
rect 39987 771835 40053 771836
rect 39987 771084 40053 771085
rect 39987 771020 39988 771084
rect 40052 771020 40053 771084
rect 39987 771019 40053 771020
rect 6106 764787 6906 767781
rect 7306 766475 8106 769459
rect 7306 766076 8106 766079
rect 6106 764346 6906 764391
rect 6106 737753 6906 737870
rect 6106 736609 6150 737753
rect 6854 736609 6906 737753
rect 6106 728343 6906 736609
rect 7306 736157 8106 736242
rect 7306 735013 7348 736157
rect 8052 735013 8106 736157
rect 7306 730035 8106 735013
rect 6106 724977 6906 727947
rect 7306 726655 8106 729639
rect 39990 728653 40050 771019
rect 40907 766188 40973 766189
rect 40907 766124 40908 766188
rect 40972 766124 40973 766188
rect 40907 766123 40973 766124
rect 40539 764964 40605 764965
rect 40539 764900 40540 764964
rect 40604 764900 40605 764964
rect 40539 764899 40605 764900
rect 40542 750413 40602 764899
rect 40723 764556 40789 764557
rect 40723 764492 40724 764556
rect 40788 764492 40789 764556
rect 40723 764491 40789 764492
rect 40726 751773 40786 764491
rect 40910 755309 40970 766123
rect 672763 759116 672829 759117
rect 672763 759052 672764 759116
rect 672828 759052 672829 759116
rect 672763 759051 672829 759052
rect 41643 758300 41709 758301
rect 41643 758236 41644 758300
rect 41708 758236 41709 758300
rect 41643 758235 41709 758236
rect 41459 757756 41525 757757
rect 41459 757692 41460 757756
rect 41524 757692 41525 757756
rect 41459 757691 41525 757692
rect 40907 755308 40973 755309
rect 40907 755244 40908 755308
rect 40972 755244 40973 755308
rect 40907 755243 40973 755244
rect 40723 751772 40789 751773
rect 40723 751708 40724 751772
rect 40788 751708 40789 751772
rect 40723 751707 40789 751708
rect 40539 750412 40605 750413
rect 40539 750348 40540 750412
rect 40604 750348 40605 750412
rect 40539 750347 40605 750348
rect 41462 742389 41522 757691
rect 41646 746605 41706 758235
rect 672766 757893 672826 759051
rect 672763 757892 672829 757893
rect 672763 757828 672764 757892
rect 672828 757828 672829 757892
rect 672763 757827 672829 757828
rect 42747 756532 42813 756533
rect 42747 756468 42748 756532
rect 42812 756468 42813 756532
rect 42747 756467 42813 756468
rect 41827 755308 41893 755309
rect 41827 755244 41828 755308
rect 41892 755244 41893 755308
rect 41827 755243 41893 755244
rect 41830 753133 41890 755243
rect 41827 753132 41893 753133
rect 41827 753068 41828 753132
rect 41892 753068 41893 753132
rect 41827 753067 41893 753068
rect 42750 749325 42810 756467
rect 42747 749324 42813 749325
rect 42747 749260 42748 749324
rect 42812 749260 42813 749324
rect 42747 749259 42813 749260
rect 41643 746604 41709 746605
rect 41643 746540 41644 746604
rect 41708 746540 41709 746604
rect 41643 746539 41709 746540
rect 41459 742388 41525 742389
rect 41459 742324 41460 742388
rect 41524 742324 41525 742388
rect 41459 742323 41525 742324
rect 54184 736599 54189 737788
rect 55385 736599 55390 737788
rect 63350 737729 63872 737732
rect 63350 736622 63872 736625
rect 54184 736574 55390 736599
rect 52580 736177 53786 736188
rect 52580 734981 52595 736177
rect 62382 736121 62904 736124
rect 62382 735014 62904 735017
rect 52580 734974 53786 734981
rect 40171 729468 40237 729469
rect 40171 729404 40172 729468
rect 40236 729404 40237 729468
rect 40171 729403 40237 729404
rect 39987 728652 40053 728653
rect 39987 728588 39988 728652
rect 40052 728588 40053 728652
rect 39987 728587 40053 728588
rect 39987 727836 40053 727837
rect 39987 727772 39988 727836
rect 40052 727772 40053 727836
rect 39987 727771 40053 727772
rect 6106 721587 6906 724581
rect 7306 723275 8106 726259
rect 7306 722876 8106 722879
rect 6106 721146 6906 721191
rect 6106 694553 6906 694670
rect 6106 693409 6150 694553
rect 6854 693409 6906 694553
rect 6106 685143 6906 693409
rect 7306 692957 8106 693042
rect 7306 691813 7348 692957
rect 8052 691813 8106 692957
rect 7306 686835 8106 691813
rect 6106 681777 6906 684747
rect 7306 683455 8106 686439
rect 39990 685541 40050 727771
rect 40174 687173 40234 729403
rect 675158 727293 675218 775643
rect 675342 774893 675402 785030
rect 675891 784956 675957 784957
rect 675891 784892 675892 784956
rect 675956 784892 675957 784956
rect 675891 784891 675957 784892
rect 675523 784820 675589 784821
rect 675523 784756 675524 784820
rect 675588 784756 675589 784820
rect 675523 784755 675589 784756
rect 675339 774892 675405 774893
rect 675339 774828 675340 774892
rect 675404 774828 675405 774892
rect 675339 774827 675405 774828
rect 675339 741708 675405 741709
rect 675339 741644 675340 741708
rect 675404 741644 675405 741708
rect 675339 741643 675405 741644
rect 675155 727292 675221 727293
rect 675155 727228 675156 727292
rect 675220 727228 675221 727292
rect 675155 727227 675221 727228
rect 41459 726204 41525 726205
rect 41459 726140 41460 726204
rect 41524 726140 41525 726204
rect 41459 726139 41525 726140
rect 40539 721308 40605 721309
rect 40539 721244 40540 721308
rect 40604 721244 40605 721308
rect 40539 721243 40605 721244
rect 40542 710837 40602 721243
rect 40907 714100 40973 714101
rect 40907 714036 40908 714100
rect 40972 714036 40973 714100
rect 40907 714035 40973 714036
rect 40539 710836 40605 710837
rect 40539 710772 40540 710836
rect 40604 710772 40605 710836
rect 40539 710771 40605 710772
rect 40910 709885 40970 714035
rect 40907 709884 40973 709885
rect 40907 709820 40908 709884
rect 40972 709820 40973 709884
rect 40907 709819 40973 709820
rect 41462 699413 41522 726139
rect 41827 715596 41893 715597
rect 41827 715532 41828 715596
rect 41892 715532 41893 715596
rect 41827 715531 41893 715532
rect 41643 715460 41709 715461
rect 41643 715396 41644 715460
rect 41708 715396 41709 715460
rect 41643 715395 41709 715396
rect 41646 702949 41706 715395
rect 41830 704989 41890 715531
rect 42011 713828 42077 713829
rect 42011 713764 42012 713828
rect 42076 713764 42077 713828
rect 42011 713763 42077 713764
rect 42014 706621 42074 713763
rect 42195 713284 42261 713285
rect 42195 713220 42196 713284
rect 42260 713220 42261 713284
rect 42195 713219 42261 713220
rect 42198 711789 42258 713219
rect 42379 712332 42445 712333
rect 42379 712268 42380 712332
rect 42444 712268 42445 712332
rect 42379 712267 42445 712268
rect 42195 711788 42261 711789
rect 42195 711724 42196 711788
rect 42260 711724 42261 711788
rect 42195 711723 42261 711724
rect 42382 708525 42442 712267
rect 42379 708524 42445 708525
rect 42379 708460 42380 708524
rect 42444 708460 42445 708524
rect 42379 708459 42445 708460
rect 42011 706620 42077 706621
rect 42011 706556 42012 706620
rect 42076 706556 42077 706620
rect 42011 706555 42077 706556
rect 41827 704988 41893 704989
rect 41827 704924 41828 704988
rect 41892 704924 41893 704988
rect 41827 704923 41893 704924
rect 41643 702948 41709 702949
rect 41643 702884 41644 702948
rect 41708 702884 41709 702948
rect 41643 702883 41709 702884
rect 41459 699412 41525 699413
rect 41459 699348 41460 699412
rect 41524 699348 41525 699412
rect 41459 699347 41525 699348
rect 674603 697372 674669 697373
rect 674603 697308 674604 697372
rect 674668 697308 674669 697372
rect 674603 697307 674669 697308
rect 54184 693399 54189 694588
rect 55385 693399 55390 694588
rect 63350 694529 63872 694532
rect 63350 693422 63872 693425
rect 54184 693374 55390 693399
rect 52580 692977 53786 692988
rect 52580 691781 52595 692977
rect 62382 692921 62904 692924
rect 62382 691814 62904 691817
rect 52580 691774 53786 691781
rect 40171 687172 40237 687173
rect 40171 687108 40172 687172
rect 40236 687108 40237 687172
rect 40171 687107 40237 687108
rect 39987 685540 40053 685541
rect 39987 685476 39988 685540
rect 40052 685476 40053 685540
rect 39987 685475 40053 685476
rect 39987 684724 40053 684725
rect 39987 684660 39988 684724
rect 40052 684660 40053 684724
rect 39987 684659 40053 684660
rect 6106 678387 6906 681381
rect 7306 680075 8106 683059
rect 7306 679676 8106 679679
rect 6106 677946 6906 677991
rect 30603 677788 30669 677789
rect 30603 677724 30604 677788
rect 30668 677724 30669 677788
rect 30603 677723 30669 677724
rect 30606 676565 30666 677723
rect 30603 676564 30669 676565
rect 30603 676500 30604 676564
rect 30668 676500 30669 676564
rect 30603 676499 30669 676500
rect 6106 651353 6906 651470
rect 6106 650209 6150 651353
rect 6854 650209 6906 651353
rect 6106 641943 6906 650209
rect 7306 649757 8106 649842
rect 7306 648613 7348 649757
rect 8052 648613 8106 649757
rect 7306 643635 8106 648613
rect 6106 638577 6906 641547
rect 7306 640255 8106 643239
rect 39990 642293 40050 684659
rect 41459 682276 41525 682277
rect 41459 682212 41460 682276
rect 41524 682212 41525 682276
rect 41459 682211 41525 682212
rect 40539 679420 40605 679421
rect 40539 679356 40540 679420
rect 40604 679356 40605 679420
rect 40539 679355 40605 679356
rect 40542 664597 40602 679355
rect 40723 678196 40789 678197
rect 40723 678132 40724 678196
rect 40788 678132 40789 678196
rect 40723 678131 40789 678132
rect 40726 665413 40786 678131
rect 40723 665412 40789 665413
rect 40723 665348 40724 665412
rect 40788 665348 40789 665412
rect 40723 665347 40789 665348
rect 40539 664596 40605 664597
rect 40539 664532 40540 664596
rect 40604 664532 40605 664596
rect 40539 664531 40605 664532
rect 41462 661333 41522 682211
rect 41643 671396 41709 671397
rect 41643 671332 41644 671396
rect 41708 671332 41709 671396
rect 41643 671331 41709 671332
rect 41459 661332 41525 661333
rect 41459 661268 41460 661332
rect 41524 661268 41525 661332
rect 41459 661267 41525 661268
rect 41646 658341 41706 671331
rect 41827 670988 41893 670989
rect 41827 670924 41828 670988
rect 41892 670924 41893 670988
rect 41827 670923 41893 670924
rect 41830 660381 41890 670923
rect 42011 670716 42077 670717
rect 42011 670652 42012 670716
rect 42076 670652 42077 670716
rect 42011 670651 42077 670652
rect 42014 663373 42074 670651
rect 42195 670172 42261 670173
rect 42195 670108 42196 670172
rect 42260 670108 42261 670172
rect 42195 670107 42261 670108
rect 42011 663372 42077 663373
rect 42011 663308 42012 663372
rect 42076 663308 42077 663372
rect 42011 663307 42077 663308
rect 42198 660517 42258 670107
rect 42195 660516 42261 660517
rect 42195 660452 42196 660516
rect 42260 660452 42261 660516
rect 42195 660451 42261 660452
rect 41827 660380 41893 660381
rect 41827 660316 41828 660380
rect 41892 660316 41893 660380
rect 41827 660315 41893 660316
rect 673867 659972 673933 659973
rect 673867 659908 673868 659972
rect 673932 659908 673933 659972
rect 673867 659907 673933 659908
rect 41643 658340 41709 658341
rect 41643 658276 41644 658340
rect 41708 658276 41709 658340
rect 41643 658275 41709 658276
rect 54184 650199 54189 651388
rect 55385 650199 55390 651388
rect 63350 651329 63872 651332
rect 63350 650222 63872 650225
rect 54184 650174 55390 650199
rect 52580 649777 53786 649788
rect 52580 648581 52595 649777
rect 62382 649721 62904 649724
rect 673315 649228 673381 649229
rect 673315 649164 673316 649228
rect 673380 649164 673381 649228
rect 673315 649163 673381 649164
rect 62382 648614 62904 648617
rect 52580 648574 53786 648581
rect 39987 642292 40053 642293
rect 39987 642228 39988 642292
rect 40052 642228 40053 642292
rect 39987 642227 40053 642228
rect 39987 641476 40053 641477
rect 39987 641412 39988 641476
rect 40052 641412 40053 641476
rect 39987 641411 40053 641412
rect 6106 635187 6906 638181
rect 7306 636875 8106 639859
rect 7306 636476 8106 636479
rect 6106 634746 6906 634791
rect 6106 608153 6906 608270
rect 6106 607009 6150 608153
rect 6854 607009 6906 608153
rect 6106 598743 6906 607009
rect 7306 606557 8106 606642
rect 7306 605413 7348 606557
rect 8052 605413 8106 606557
rect 7306 600435 8106 605413
rect 6106 595377 6906 598347
rect 7306 597055 8106 600039
rect 39990 599045 40050 641411
rect 41459 640660 41525 640661
rect 41459 640596 41460 640660
rect 41524 640596 41525 640660
rect 41459 640595 41525 640596
rect 40907 636580 40973 636581
rect 40907 636516 40908 636580
rect 40972 636516 40973 636580
rect 40907 636515 40973 636516
rect 40539 636172 40605 636173
rect 40539 636108 40540 636172
rect 40604 636108 40605 636172
rect 40539 636107 40605 636108
rect 40542 621485 40602 636107
rect 40723 634948 40789 634949
rect 40723 634884 40724 634948
rect 40788 634884 40789 634948
rect 40723 634883 40789 634884
rect 40726 623797 40786 634883
rect 40910 625293 40970 636515
rect 40907 625292 40973 625293
rect 40907 625228 40908 625292
rect 40972 625228 40973 625292
rect 40907 625227 40973 625228
rect 40723 623796 40789 623797
rect 40723 623732 40724 623796
rect 40788 623732 40789 623796
rect 40723 623731 40789 623732
rect 40539 621484 40605 621485
rect 40539 621420 40540 621484
rect 40604 621420 40605 621484
rect 40539 621419 40605 621420
rect 41462 614141 41522 640595
rect 41827 629916 41893 629917
rect 41827 629852 41828 629916
rect 41892 629852 41893 629916
rect 41827 629851 41893 629852
rect 41643 629100 41709 629101
rect 41643 629036 41644 629100
rect 41708 629036 41709 629100
rect 41643 629035 41709 629036
rect 41459 614140 41525 614141
rect 41459 614076 41460 614140
rect 41524 614076 41525 614140
rect 41459 614075 41525 614076
rect 41646 612781 41706 629035
rect 41830 616861 41890 629851
rect 42011 629236 42077 629237
rect 42011 629172 42012 629236
rect 42076 629172 42077 629236
rect 42011 629171 42077 629172
rect 42014 619037 42074 629171
rect 42195 628964 42261 628965
rect 42195 628900 42196 628964
rect 42260 628900 42261 628964
rect 42195 628899 42261 628900
rect 42011 619036 42077 619037
rect 42011 618972 42012 619036
rect 42076 618972 42077 619036
rect 42011 618971 42077 618972
rect 41827 616860 41893 616861
rect 41827 616796 41828 616860
rect 41892 616796 41893 616860
rect 41827 616795 41893 616796
rect 42198 616045 42258 628899
rect 42195 616044 42261 616045
rect 42195 615980 42196 616044
rect 42260 615980 42261 616044
rect 42195 615979 42261 615980
rect 41643 612780 41709 612781
rect 41643 612716 41644 612780
rect 41708 612716 41709 612780
rect 41643 612715 41709 612716
rect 54184 606999 54189 608188
rect 55385 606999 55390 608188
rect 63350 608129 63872 608132
rect 63350 607022 63872 607025
rect 54184 606974 55390 606999
rect 52580 606577 53786 606588
rect 52580 605381 52595 606577
rect 62382 606521 62904 606524
rect 62382 605414 62904 605417
rect 52580 605374 53786 605381
rect 39987 599044 40053 599045
rect 39987 598980 39988 599044
rect 40052 598980 40053 599044
rect 39987 598979 40053 598980
rect 39987 598228 40053 598229
rect 39987 598164 39988 598228
rect 40052 598164 40053 598228
rect 39987 598163 40053 598164
rect 6106 591987 6906 594981
rect 7306 593675 8106 596659
rect 7306 593276 8106 593279
rect 6106 591546 6906 591591
rect 6106 564953 6906 565070
rect 6106 563809 6150 564953
rect 6854 563809 6906 564953
rect 6106 555543 6906 563809
rect 7306 563357 8106 563442
rect 7306 562213 7348 563357
rect 8052 562213 8106 563357
rect 7306 557235 8106 562213
rect 6106 552177 6906 555147
rect 7306 553855 8106 556839
rect 39990 555933 40050 598163
rect 41459 596596 41525 596597
rect 41459 596532 41460 596596
rect 41524 596532 41525 596596
rect 41459 596531 41525 596532
rect 40539 592108 40605 592109
rect 40539 592044 40540 592108
rect 40604 592044 40605 592108
rect 40539 592043 40605 592044
rect 40542 577557 40602 592043
rect 40723 591700 40789 591701
rect 40723 591636 40724 591700
rect 40788 591636 40789 591700
rect 40723 591635 40789 591636
rect 40726 579053 40786 591635
rect 40723 579052 40789 579053
rect 40723 578988 40724 579052
rect 40788 578988 40789 579052
rect 40723 578987 40789 578988
rect 40539 577556 40605 577557
rect 40539 577492 40540 577556
rect 40604 577492 40605 577556
rect 40539 577491 40605 577492
rect 41462 571573 41522 596531
rect 41643 594964 41709 594965
rect 41643 594900 41644 594964
rect 41708 594900 41709 594964
rect 41643 594899 41709 594900
rect 41459 571572 41525 571573
rect 41459 571508 41460 571572
rect 41524 571508 41525 571572
rect 41459 571507 41525 571508
rect 41646 570485 41706 594899
rect 42379 585172 42445 585173
rect 42379 585108 42380 585172
rect 42444 585108 42445 585172
rect 42379 585107 42445 585108
rect 41827 584220 41893 584221
rect 41827 584156 41828 584220
rect 41892 584156 41893 584220
rect 41827 584155 41893 584156
rect 42011 584220 42077 584221
rect 42011 584156 42012 584220
rect 42076 584156 42077 584220
rect 42011 584155 42077 584156
rect 41830 580277 41890 584155
rect 42014 582181 42074 584155
rect 42011 582180 42077 582181
rect 42011 582116 42012 582180
rect 42076 582116 42077 582180
rect 42011 582115 42077 582116
rect 41827 580276 41893 580277
rect 41827 580212 41828 580276
rect 41892 580212 41893 580276
rect 41827 580211 41893 580212
rect 42382 579730 42442 585107
rect 42563 583676 42629 583677
rect 42563 583612 42564 583676
rect 42628 583612 42629 583676
rect 42563 583611 42629 583612
rect 41830 579670 42442 579730
rect 41830 573749 41890 579670
rect 42566 579050 42626 583611
rect 42014 578990 42626 579050
rect 41827 573748 41893 573749
rect 41827 573684 41828 573748
rect 41892 573684 41893 573748
rect 41827 573683 41893 573684
rect 42014 572797 42074 578990
rect 42195 576876 42261 576877
rect 42195 576812 42196 576876
rect 42260 576812 42261 576876
rect 42195 576811 42261 576812
rect 42198 575925 42258 576811
rect 42195 575924 42261 575925
rect 42195 575860 42196 575924
rect 42260 575860 42261 575924
rect 42195 575859 42261 575860
rect 673318 572797 673378 649163
rect 42011 572796 42077 572797
rect 42011 572732 42012 572796
rect 42076 572732 42077 572796
rect 42011 572731 42077 572732
rect 673315 572796 673381 572797
rect 673315 572732 673316 572796
rect 673380 572732 673381 572796
rect 673315 572731 673381 572732
rect 41643 570484 41709 570485
rect 41643 570420 41644 570484
rect 41708 570420 41709 570484
rect 41643 570419 41709 570420
rect 54184 563799 54189 564988
rect 55385 563799 55390 564988
rect 63350 564929 63872 564932
rect 63350 563822 63872 563825
rect 54184 563774 55390 563799
rect 52580 563377 53786 563388
rect 52580 562181 52595 563377
rect 62382 563321 62904 563324
rect 62382 562214 62904 562217
rect 52580 562174 53786 562181
rect 39987 555932 40053 555933
rect 39987 555868 39988 555932
rect 40052 555868 40053 555932
rect 39987 555867 40053 555868
rect 6106 548787 6906 551781
rect 7306 550475 8106 553459
rect 40539 550628 40605 550629
rect 40539 550564 40540 550628
rect 40604 550564 40605 550628
rect 40539 550563 40605 550564
rect 7306 550076 8106 550079
rect 6106 548346 6906 548391
rect 40542 530773 40602 550563
rect 40723 549404 40789 549405
rect 40723 549340 40724 549404
rect 40788 549340 40789 549404
rect 40723 549339 40789 549340
rect 40726 533901 40786 549339
rect 40907 548996 40973 548997
rect 40907 548932 40908 548996
rect 40972 548932 40973 548996
rect 40907 548931 40973 548932
rect 40910 534581 40970 548931
rect 41459 545188 41525 545189
rect 41459 545124 41460 545188
rect 41524 545124 41525 545188
rect 41459 545123 41525 545124
rect 40907 534580 40973 534581
rect 40907 534516 40908 534580
rect 40972 534516 40973 534580
rect 40907 534515 40973 534516
rect 40723 533900 40789 533901
rect 40723 533836 40724 533900
rect 40788 533836 40789 533900
rect 40723 533835 40789 533836
rect 40539 530772 40605 530773
rect 40539 530708 40540 530772
rect 40604 530708 40605 530772
rect 40539 530707 40605 530708
rect 41462 529957 41522 545123
rect 41643 543012 41709 543013
rect 41643 542948 41644 543012
rect 41708 542948 41709 543012
rect 41643 542947 41709 542948
rect 41459 529956 41525 529957
rect 41459 529892 41460 529956
rect 41524 529892 41525 529956
rect 41459 529891 41525 529892
rect 41646 529413 41706 542947
rect 41827 542876 41893 542877
rect 41827 542812 41828 542876
rect 41892 542812 41893 542876
rect 41827 542811 41893 542812
rect 41830 532677 41890 542811
rect 42011 542332 42077 542333
rect 42011 542268 42012 542332
rect 42076 542268 42077 542332
rect 42011 542267 42077 542268
rect 42014 535941 42074 542267
rect 42011 535940 42077 535941
rect 42011 535876 42012 535940
rect 42076 535876 42077 535940
rect 42011 535875 42077 535876
rect 41827 532676 41893 532677
rect 41827 532612 41828 532676
rect 41892 532612 41893 532676
rect 41827 532611 41893 532612
rect 41643 529412 41709 529413
rect 41643 529348 41644 529412
rect 41708 529348 41709 529412
rect 41643 529347 41709 529348
rect 667206 518597 669814 518696
rect 667206 514041 667283 518597
rect 669759 514041 669814 518597
rect 667206 513920 669814 514041
rect 667218 508607 669826 508726
rect 667218 504051 667297 508607
rect 669773 504051 669826 508607
rect 667218 503950 669826 504051
rect 50172 497769 52196 497874
rect 50172 493213 50310 497769
rect 52146 493213 52196 497769
rect 50172 493084 52196 493213
rect 50198 487779 52222 487884
rect 50198 483223 50298 487779
rect 52134 483223 52222 487779
rect 50198 483094 52222 483223
rect 6106 437353 6906 437470
rect 6106 436209 6150 437353
rect 6854 436209 6906 437353
rect 6106 427943 6906 436209
rect 54184 436199 54189 437388
rect 55385 436199 55390 437388
rect 63350 437329 63872 437332
rect 63350 436222 63872 436225
rect 54184 436174 55390 436199
rect 7306 435757 8106 435842
rect 7306 434613 7348 435757
rect 8052 434613 8106 435757
rect 7306 429635 8106 434613
rect 52580 435777 53786 435788
rect 52580 434581 52595 435777
rect 62382 435721 62904 435724
rect 62382 434614 62904 434617
rect 52580 434574 53786 434581
rect 664008 430395 666612 430490
rect 6106 424577 6906 427547
rect 7306 426255 8106 429239
rect 42195 426052 42261 426053
rect 42195 425988 42196 426052
rect 42260 425988 42261 426052
rect 42195 425987 42261 425988
rect 6106 421187 6906 424181
rect 7306 422875 8106 425859
rect 41827 425644 41893 425645
rect 41827 425580 41828 425644
rect 41892 425580 41893 425644
rect 41827 425579 41893 425580
rect 41830 425370 41890 425579
rect 40542 425310 41890 425370
rect 7306 422476 8106 422479
rect 30603 420932 30669 420933
rect 30603 420868 30604 420932
rect 30668 420868 30669 420932
rect 30603 420867 30669 420868
rect 6106 420746 6906 420791
rect 30606 418845 30666 420867
rect 30603 418844 30669 418845
rect 30603 418780 30604 418844
rect 30668 418780 30669 418844
rect 30603 418779 30669 418780
rect 40542 398853 40602 425310
rect 40723 425072 40789 425073
rect 40723 425008 40724 425072
rect 40788 425008 40789 425072
rect 42198 425070 42258 425987
rect 664008 425679 664099 430395
rect 666575 425679 666612 430395
rect 664008 425572 666612 425679
rect 42198 425010 42442 425070
rect 40723 425007 40789 425008
rect 40726 400077 40786 425007
rect 41827 424012 41893 424013
rect 41827 424010 41828 424012
rect 40910 423950 41828 424010
rect 40723 400076 40789 400077
rect 40723 400012 40724 400076
rect 40788 400012 40789 400076
rect 40723 400011 40789 400012
rect 40910 399669 40970 423950
rect 41827 423948 41828 423950
rect 41892 423948 41893 424012
rect 41827 423947 41893 423948
rect 42011 423604 42077 423605
rect 42011 423540 42012 423604
rect 42076 423540 42077 423604
rect 42011 423539 42077 423540
rect 41827 422788 41893 422789
rect 41827 422724 41828 422788
rect 41892 422724 41893 422788
rect 41827 422723 41893 422724
rect 41830 422650 41890 422723
rect 41094 422590 41890 422650
rect 41094 409461 41154 422590
rect 42014 421970 42074 423539
rect 41830 421910 42074 421970
rect 41830 418170 41890 421910
rect 41462 418110 41890 418170
rect 41091 409460 41157 409461
rect 41091 409396 41092 409460
rect 41156 409396 41157 409460
rect 41091 409395 41157 409396
rect 41462 402525 41522 418110
rect 41643 418028 41709 418029
rect 41643 417964 41644 418028
rect 41708 417964 41709 418028
rect 41643 417963 41709 417964
rect 41646 406333 41706 417963
rect 41827 414628 41893 414629
rect 41827 414564 41828 414628
rect 41892 414564 41893 414628
rect 41827 414563 41893 414564
rect 41830 408510 41890 414563
rect 42382 411229 42442 425010
rect 664018 420517 666634 420524
rect 664018 415801 664082 420517
rect 666558 415801 666634 420517
rect 664018 415760 666634 415801
rect 42379 411228 42445 411229
rect 42379 411164 42380 411228
rect 42444 411164 42445 411228
rect 42379 411163 42445 411164
rect 41830 408450 42074 408510
rect 41643 406332 41709 406333
rect 41643 406268 41644 406332
rect 41708 406268 41709 406332
rect 41643 406267 41709 406268
rect 41459 402524 41525 402525
rect 41459 402460 41460 402524
rect 41524 402460 41525 402524
rect 41459 402459 41525 402460
rect 42014 401845 42074 408450
rect 42011 401844 42077 401845
rect 42011 401780 42012 401844
rect 42076 401780 42077 401844
rect 42011 401779 42077 401780
rect 40907 399668 40973 399669
rect 40907 399604 40908 399668
rect 40972 399604 40973 399668
rect 40907 399603 40973 399604
rect 40539 398852 40605 398853
rect 40539 398788 40540 398852
rect 40604 398788 40605 398852
rect 40539 398787 40605 398788
rect 6106 394153 6906 394270
rect 6106 393009 6150 394153
rect 6854 393009 6906 394153
rect 6106 384743 6906 393009
rect 54184 392999 54189 394188
rect 55385 392999 55390 394188
rect 63350 394129 63872 394132
rect 63350 393022 63872 393025
rect 54184 392974 55390 392999
rect 7306 392557 8106 392642
rect 7306 391413 7348 392557
rect 8052 391413 8106 392557
rect 7306 386435 8106 391413
rect 52580 392577 53786 392588
rect 52580 391381 52595 392577
rect 62382 392521 62904 392524
rect 62382 391414 62904 391417
rect 52580 391374 53786 391381
rect 6106 381377 6906 384347
rect 7306 383055 8106 386039
rect 40723 383076 40789 383077
rect 40723 383012 40724 383076
rect 40788 383012 40789 383076
rect 40723 383011 40789 383012
rect 6106 377987 6906 380981
rect 7306 379675 8106 382659
rect 40539 382260 40605 382261
rect 40539 382196 40540 382260
rect 40604 382196 40605 382260
rect 40539 382195 40605 382196
rect 7306 379276 8106 379279
rect 6106 377546 6906 377591
rect 40542 355741 40602 382195
rect 40726 356965 40786 383011
rect 41459 381852 41525 381853
rect 41459 381788 41460 381852
rect 41524 381788 41525 381852
rect 41459 381787 41525 381788
rect 40907 379812 40973 379813
rect 40907 379748 40908 379812
rect 40972 379748 40973 379812
rect 40907 379747 40973 379748
rect 40910 360229 40970 379747
rect 40907 360228 40973 360229
rect 40907 360164 40908 360228
rect 40972 360164 40973 360228
rect 40907 360163 40973 360164
rect 41462 358733 41522 381787
rect 42011 371924 42077 371925
rect 42011 371860 42012 371924
rect 42076 371860 42077 371924
rect 42011 371859 42077 371860
rect 41643 371380 41709 371381
rect 41643 371316 41644 371380
rect 41708 371316 41709 371380
rect 41643 371315 41709 371316
rect 41646 362949 41706 371315
rect 41827 370292 41893 370293
rect 41827 370228 41828 370292
rect 41892 370228 41893 370292
rect 41827 370227 41893 370228
rect 41830 366349 41890 370227
rect 41827 366348 41893 366349
rect 41827 366284 41828 366348
rect 41892 366284 41893 366348
rect 41827 366283 41893 366284
rect 42014 363765 42074 371859
rect 42011 363764 42077 363765
rect 42011 363700 42012 363764
rect 42076 363700 42077 363764
rect 42011 363699 42077 363700
rect 41643 362948 41709 362949
rect 41643 362884 41644 362948
rect 41708 362884 41709 362948
rect 41643 362883 41709 362884
rect 41459 358732 41525 358733
rect 41459 358668 41460 358732
rect 41524 358668 41525 358732
rect 41459 358667 41525 358668
rect 40723 356964 40789 356965
rect 40723 356900 40724 356964
rect 40788 356900 40789 356964
rect 40723 356899 40789 356900
rect 40539 355740 40605 355741
rect 40539 355676 40540 355740
rect 40604 355676 40605 355740
rect 40539 355675 40605 355676
rect 63350 351729 63872 351732
rect 6106 350953 6906 351070
rect 6106 349809 6150 350953
rect 6854 349809 6906 350953
rect 6106 341543 6906 349809
rect 54184 349799 54189 350988
rect 55385 349799 55390 350988
rect 63350 350622 63872 350625
rect 54184 349774 55390 349799
rect 7306 349357 8106 349442
rect 7306 348213 7348 349357
rect 8052 348213 8106 349357
rect 7306 343235 8106 348213
rect 52580 349377 53786 349388
rect 52580 348181 52595 349377
rect 62382 349321 62904 349324
rect 62382 348214 62904 348217
rect 52580 348174 53786 348181
rect 6106 338177 6906 341147
rect 7306 339855 8106 342839
rect 40723 339828 40789 339829
rect 40723 339764 40724 339828
rect 40788 339764 40789 339828
rect 40723 339763 40789 339764
rect 6106 334787 6906 337781
rect 7306 336475 8106 339459
rect 40539 339012 40605 339013
rect 40539 338948 40540 339012
rect 40604 338948 40605 339012
rect 40539 338947 40605 338948
rect 7306 336076 8106 336079
rect 6106 334346 6906 334391
rect 40542 312357 40602 338947
rect 40726 313853 40786 339763
rect 41459 338604 41525 338605
rect 41459 338540 41460 338604
rect 41524 338540 41525 338604
rect 41459 338539 41525 338540
rect 40907 337380 40973 337381
rect 40907 337316 40908 337380
rect 40972 337316 40973 337380
rect 40907 337315 40973 337316
rect 40723 313852 40789 313853
rect 40723 313788 40724 313852
rect 40788 313788 40789 313852
rect 40723 313787 40789 313788
rect 40910 313173 40970 337315
rect 41275 335748 41341 335749
rect 41275 335684 41276 335748
rect 41340 335684 41341 335748
rect 41275 335683 41341 335684
rect 41091 335340 41157 335341
rect 41091 335276 41092 335340
rect 41156 335276 41157 335340
rect 41091 335275 41157 335276
rect 41094 317389 41154 335275
rect 41278 321197 41338 335683
rect 41275 321196 41341 321197
rect 41275 321132 41276 321196
rect 41340 321132 41341 321196
rect 41275 321131 41341 321132
rect 41091 317388 41157 317389
rect 41091 317324 41092 317388
rect 41156 317324 41157 317388
rect 41091 317323 41157 317324
rect 41462 315485 41522 338539
rect 41643 336972 41709 336973
rect 41643 336908 41644 336972
rect 41708 336908 41709 336972
rect 41643 336907 41709 336908
rect 41646 315893 41706 336907
rect 41827 334116 41893 334117
rect 41827 334052 41828 334116
rect 41892 334052 41893 334116
rect 41827 334051 41893 334052
rect 41830 324869 41890 334051
rect 42011 328404 42077 328405
rect 42011 328340 42012 328404
rect 42076 328340 42077 328404
rect 42011 328339 42077 328340
rect 41827 324868 41893 324869
rect 41827 324804 41828 324868
rect 41892 324804 41893 324868
rect 41827 324803 41893 324804
rect 42014 319973 42074 328339
rect 42011 319972 42077 319973
rect 42011 319908 42012 319972
rect 42076 319908 42077 319972
rect 42011 319907 42077 319908
rect 41643 315892 41709 315893
rect 41643 315828 41644 315892
rect 41708 315828 41709 315892
rect 41643 315827 41709 315828
rect 41459 315484 41525 315485
rect 41459 315420 41460 315484
rect 41524 315420 41525 315484
rect 41459 315419 41525 315420
rect 40907 313172 40973 313173
rect 40907 313108 40908 313172
rect 40972 313108 40973 313172
rect 40907 313107 40973 313108
rect 40539 312356 40605 312357
rect 40539 312292 40540 312356
rect 40604 312292 40605 312356
rect 40539 312291 40605 312292
rect 6106 307753 6906 307870
rect 6106 306609 6150 307753
rect 6854 306609 6906 307753
rect 6106 298343 6906 306609
rect 54184 306599 54189 307788
rect 55385 306599 55390 307788
rect 63350 307729 63872 307732
rect 63350 306622 63872 306625
rect 54184 306574 55390 306599
rect 7306 306157 8106 306242
rect 7306 305013 7348 306157
rect 8052 305013 8106 306157
rect 7306 300035 8106 305013
rect 52580 306177 53786 306188
rect 52580 304981 52595 306177
rect 62382 306121 62904 306124
rect 62382 305014 62904 305017
rect 52580 304974 53786 304981
rect 6106 294977 6906 297947
rect 7306 296655 8106 299639
rect 42379 296852 42445 296853
rect 42379 296788 42380 296852
rect 42444 296788 42445 296852
rect 42379 296787 42445 296788
rect 6106 291587 6906 294581
rect 7306 293275 8106 296259
rect 40542 296110 41890 296170
rect 7306 292876 8106 292879
rect 6106 291146 6906 291191
rect 40542 269109 40602 296110
rect 41830 296037 41890 296110
rect 41827 296036 41893 296037
rect 41827 295972 41828 296036
rect 41892 295972 41893 296036
rect 41827 295971 41893 295972
rect 42195 295628 42261 295629
rect 42195 295564 42196 295628
rect 42260 295564 42261 295628
rect 42195 295563 42261 295564
rect 42011 295220 42077 295221
rect 42011 295156 42012 295220
rect 42076 295156 42077 295220
rect 42011 295155 42077 295156
rect 41827 294404 41893 294405
rect 41827 294340 41828 294404
rect 41892 294340 41893 294404
rect 41827 294339 41893 294340
rect 41830 294130 41890 294339
rect 40726 294070 41890 294130
rect 40726 269789 40786 294070
rect 41827 293996 41893 293997
rect 41827 293932 41828 293996
rect 41892 293932 41893 293996
rect 41827 293931 41893 293932
rect 41830 293450 41890 293931
rect 41094 293390 41890 293450
rect 41094 287070 41154 293390
rect 42014 292770 42074 295155
rect 40910 287010 41154 287070
rect 41278 292710 41522 292770
rect 40910 278765 40970 287010
rect 40907 278764 40973 278765
rect 40907 278700 40908 278764
rect 40972 278700 40973 278764
rect 40907 278699 40973 278700
rect 41278 278490 41338 292710
rect 41462 292593 41522 292710
rect 41830 292710 42074 292770
rect 41459 292592 41525 292593
rect 41459 292528 41460 292592
rect 41524 292528 41525 292592
rect 41459 292527 41525 292528
rect 41830 288149 41890 292710
rect 42198 292590 42258 295563
rect 42014 292530 42258 292590
rect 41827 288148 41893 288149
rect 41827 288084 41828 288148
rect 41892 288084 41893 288148
rect 41827 288083 41893 288084
rect 41827 287876 41893 287877
rect 41827 287812 41828 287876
rect 41892 287812 41893 287876
rect 41827 287811 41893 287812
rect 41643 285020 41709 285021
rect 41643 284956 41644 285020
rect 41708 284956 41709 285020
rect 41643 284955 41709 284956
rect 41459 284884 41525 284885
rect 41459 284820 41460 284884
rect 41524 284820 41525 284884
rect 41459 284819 41525 284820
rect 41462 281485 41522 284819
rect 41459 281484 41525 281485
rect 41459 281420 41460 281484
rect 41524 281420 41525 281484
rect 41459 281419 41525 281420
rect 40910 278430 41338 278490
rect 40910 277405 40970 278430
rect 40907 277404 40973 277405
rect 40907 277340 40908 277404
rect 40972 277340 40973 277404
rect 40907 277339 40973 277340
rect 41646 272373 41706 284955
rect 41830 276725 41890 287811
rect 42014 285021 42074 292530
rect 42011 285020 42077 285021
rect 42011 284956 42012 285020
rect 42076 284956 42077 285020
rect 42011 284955 42077 284956
rect 42382 277410 42442 296787
rect 42014 277350 42442 277410
rect 41827 276724 41893 276725
rect 41827 276660 41828 276724
rect 41892 276660 41893 276724
rect 41827 276659 41893 276660
rect 41643 272372 41709 272373
rect 41643 272308 41644 272372
rect 41708 272308 41709 272372
rect 41643 272307 41709 272308
rect 42014 270469 42074 277350
rect 52582 276850 52593 278046
rect 53789 277446 53800 278046
rect 53789 277415 56416 277446
rect 53789 276859 55806 277415
rect 56362 276859 56416 277415
rect 53789 276850 56416 276859
rect 52582 276822 56416 276850
rect 50186 273412 52198 273438
rect 50186 272056 50193 273412
rect 52189 272638 52198 273412
rect 52189 272613 56406 272638
rect 52189 272057 55802 272613
rect 56358 272057 56406 272613
rect 52189 272056 56406 272057
rect 50186 272026 56406 272056
rect 47792 271659 56616 271688
rect 42011 270468 42077 270469
rect 42011 270404 42012 270468
rect 42076 270404 42077 270468
rect 42011 270403 42077 270404
rect 47792 270303 47799 271659
rect 49795 271650 56616 271659
rect 49795 271094 55776 271650
rect 56492 271094 56616 271650
rect 49795 271082 56616 271094
rect 49795 271058 57202 271082
rect 49795 270303 49802 271058
rect 47792 270258 49802 270303
rect 40723 269788 40789 269789
rect 40723 269724 40724 269788
rect 40788 269724 40789 269788
rect 40723 269723 40789 269724
rect 40539 269108 40605 269109
rect 40539 269044 40540 269108
rect 40604 269044 40605 269108
rect 40539 269043 40605 269044
rect 6106 264553 6906 264670
rect 6106 263409 6150 264553
rect 6854 263409 6906 264553
rect 6106 255143 6906 263409
rect 54184 263399 54189 264588
rect 55385 263399 55390 264588
rect 54184 263374 55390 263399
rect 7306 262957 8106 263042
rect 7306 261813 7348 262957
rect 8052 261813 8106 262957
rect 7306 256835 8106 261813
rect 52580 262977 53786 262988
rect 52580 261781 52595 262977
rect 52580 261774 53786 261781
rect 56572 261466 57202 271058
rect 57542 264698 58162 272042
rect 58502 269444 59122 272992
rect 58502 266488 58529 269444
rect 59085 266488 59122 269444
rect 58502 266408 59122 266488
rect 59462 266618 60082 273952
rect 60422 267578 61042 274922
rect 61382 268538 62002 275876
rect 62342 269498 62962 276834
rect 63302 270458 63922 277792
rect 63302 269838 67172 270458
rect 62342 268878 66212 269498
rect 61382 267918 65252 268538
rect 60422 266958 64292 267578
rect 59462 265998 63332 266618
rect 62712 265440 63332 265998
rect 57542 264078 61412 264698
rect 47770 261325 59470 261466
rect 47770 258689 47991 261325
rect 49667 261264 59470 261325
rect 49667 258689 56555 261264
rect 47770 258628 56555 258689
rect 59351 258628 59470 261264
rect 47770 258466 59470 258628
rect 60792 257466 61412 264078
rect 62712 262484 62737 265440
rect 63293 262484 63332 265440
rect 62712 262402 63332 262484
rect 50170 257442 61412 257466
rect 50170 257325 60820 257442
rect 6106 251777 6906 254747
rect 7306 253455 8106 256439
rect 50170 254689 50391 257325
rect 52067 257264 60820 257325
rect 52067 254689 56564 257264
rect 50170 254628 56564 254689
rect 60320 254628 60820 257264
rect 50170 254486 60820 254628
rect 61376 254486 61412 257442
rect 50170 254466 61412 254486
rect 60792 254422 61412 254466
rect 42195 253604 42261 253605
rect 42195 253540 42196 253604
rect 42260 253540 42261 253604
rect 42195 253539 42261 253540
rect 41827 253196 41893 253197
rect 41827 253132 41828 253196
rect 41892 253132 41893 253196
rect 41827 253131 41893 253132
rect 6106 248387 6906 251381
rect 7306 250075 8106 253059
rect 40539 252652 40605 252653
rect 40539 252588 40540 252652
rect 40604 252588 40605 252652
rect 40539 252587 40605 252588
rect 40171 249796 40237 249797
rect 40171 249732 40172 249796
rect 40236 249732 40237 249796
rect 40171 249731 40237 249732
rect 7306 249676 8106 249679
rect 39987 248980 40053 248981
rect 39987 248916 39988 248980
rect 40052 248916 40053 248980
rect 39987 248915 40053 248916
rect 6106 247946 6906 247991
rect 39990 244629 40050 248915
rect 39987 244628 40053 244629
rect 39987 244564 39988 244628
rect 40052 244564 40053 244628
rect 39987 244563 40053 244564
rect 40174 244490 40234 249731
rect 40355 249388 40421 249389
rect 40355 249324 40356 249388
rect 40420 249324 40421 249388
rect 40355 249323 40421 249324
rect 39990 244430 40234 244490
rect 39990 238098 40050 244430
rect 40171 244220 40237 244221
rect 40171 244156 40172 244220
rect 40236 244156 40237 244220
rect 40171 244155 40237 244156
rect 40174 238370 40234 244155
rect 40358 238509 40418 249323
rect 40355 238508 40421 238509
rect 40355 238444 40356 238508
rect 40420 238444 40421 238508
rect 40542 238506 40602 252587
rect 41643 252244 41709 252245
rect 41643 252180 41644 252244
rect 41708 252180 41709 252244
rect 41643 252179 41709 252180
rect 41646 248430 41706 252179
rect 41462 248370 41706 248430
rect 41462 245850 41522 248370
rect 40726 245790 41522 245850
rect 40726 239053 40786 245790
rect 41830 245717 41890 253131
rect 42198 245853 42258 253539
rect 52578 253450 63292 253466
rect 52578 253448 56152 253450
rect 52578 250492 52602 253448
rect 53798 250494 56152 253448
rect 63268 250494 63292 253450
rect 53798 250492 63292 250494
rect 52578 250466 63292 250492
rect 42195 245852 42261 245853
rect 42195 245788 42196 245852
rect 42260 245788 42261 245852
rect 42195 245787 42261 245788
rect 41827 245716 41893 245717
rect 41827 245652 41828 245716
rect 41892 245652 41893 245716
rect 41827 245651 41893 245652
rect 63672 245466 64292 266958
rect 40984 245450 64292 245466
rect 40984 245433 63703 245450
rect 40723 239052 40789 239053
rect 40723 238988 40724 239052
rect 40788 238988 40789 239052
rect 40723 238987 40789 238988
rect 40542 238446 40786 238506
rect 40355 238443 40421 238444
rect 40174 238310 40602 238370
rect 40542 238237 40602 238310
rect 40539 238236 40605 238237
rect 40539 238172 40540 238236
rect 40604 238172 40605 238236
rect 40539 238171 40605 238172
rect 39990 238038 40602 238098
rect 40542 236741 40602 238038
rect 40539 236740 40605 236741
rect 40539 236676 40540 236740
rect 40604 236676 40605 236740
rect 40539 236675 40605 236676
rect 40726 234562 40786 238446
rect 40984 238317 41060 245433
rect 43536 245341 63703 245433
rect 43536 242545 56391 245341
rect 63347 242545 63703 245341
rect 43536 242494 63703 242545
rect 64259 242494 64292 245450
rect 43536 242466 64292 242494
rect 43536 238317 43612 242466
rect 63672 242358 64292 242466
rect 64632 241466 65252 267918
rect 65592 253438 66212 268878
rect 65592 250482 65615 253438
rect 66171 250482 66212 253438
rect 65592 250386 66212 250482
rect 66552 249450 67172 269838
rect 393442 269361 394228 269470
rect 393442 266565 393481 269361
rect 394197 266565 394228 269361
rect 393442 266474 394228 266565
rect 394044 262208 394224 266474
rect 409094 265462 409274 265476
rect 408466 265368 409274 265462
rect 408466 262892 408507 265368
rect 409223 262892 409274 265368
rect 408466 262854 409274 262892
rect 409094 262244 409274 262854
rect 394504 261349 395406 261450
rect 394504 258553 394597 261349
rect 395313 258553 395406 261349
rect 394504 258468 395406 258553
rect 409686 257366 410808 257470
rect 409686 254570 409735 257366
rect 410771 254570 410808 257366
rect 409686 254452 410808 254570
rect 211712 253376 212610 253472
rect 211712 250580 211801 253376
rect 212517 250580 212610 253376
rect 211712 250470 212610 250580
rect 241812 253376 242710 253472
rect 272232 253376 272620 253472
rect 302162 253376 302714 253472
rect 332112 253376 333010 253472
rect 241812 250580 241901 253376
rect 242617 250580 242710 253376
rect 332112 250580 332201 253376
rect 332917 250580 333010 253376
rect 241812 250470 242710 250580
rect 272232 250470 272620 250580
rect 302162 250470 302714 250580
rect 332112 250470 333010 250580
rect 362212 253376 363110 253472
rect 392572 253376 393110 253472
rect 362212 250580 362301 253376
rect 363017 250580 363110 253376
rect 393073 250580 393110 253376
rect 362212 250470 363110 250580
rect 392572 250470 393110 250580
rect 66552 246494 66579 249450
rect 67135 246494 67172 249450
rect 66552 246348 67172 246494
rect 196676 249367 197618 249464
rect 196676 246571 196785 249367
rect 197501 246571 197618 249367
rect 196676 246468 197618 246571
rect 226776 249367 227718 249464
rect 226776 246571 226885 249367
rect 227601 246571 227718 249367
rect 226776 246468 227718 246571
rect 256876 249367 257818 249464
rect 287156 249405 287658 249464
rect 256876 246571 256985 249367
rect 257701 246571 257818 249367
rect 347176 249367 348118 249464
rect 256876 246468 257818 246571
rect 347176 246571 347285 249367
rect 348001 246571 348118 249367
rect 317354 246468 317802 246541
rect 347176 246468 348118 246571
rect 377176 249367 378118 249464
rect 377176 246571 377285 249367
rect 378001 246571 378118 249367
rect 377176 246468 378118 246571
rect 407176 249367 408118 249464
rect 407176 246571 407285 249367
rect 408001 246571 408118 249367
rect 407176 246468 408118 246571
rect 650618 249455 651238 277798
rect 651578 253437 652198 276844
rect 651578 250481 651614 253437
rect 652170 250481 652198 253437
rect 651578 250392 652198 250481
rect 650618 246499 650648 249455
rect 651204 246499 651238 249455
rect 650618 246296 651238 246499
rect 212568 245451 213540 245462
rect 212568 242495 212605 245451
rect 213481 242495 213540 245451
rect 212568 242464 213540 242495
rect 242668 245451 243640 245462
rect 272982 245451 273314 245462
rect 303168 245451 303460 245462
rect 332968 245451 333940 245462
rect 242668 242495 242705 245451
rect 243581 242495 243640 245451
rect 332968 242495 333005 245451
rect 333881 242495 333940 245451
rect 242668 242464 243640 242495
rect 272982 242464 273314 242495
rect 303168 242464 303460 242495
rect 332968 242464 333940 242495
rect 363068 245451 364040 245462
rect 363068 242495 363105 245451
rect 363981 242495 364040 245451
rect 363068 242464 364040 242495
rect 393210 245451 393800 245462
rect 393210 242495 393227 245451
rect 393783 242495 393800 245451
rect 393210 242464 393800 242495
rect 40984 238266 43612 238317
rect 44196 241446 65252 241466
rect 44196 241375 64653 241446
rect 44196 241343 56406 241375
rect 41091 238100 41157 238101
rect 41091 238036 41092 238100
rect 41156 238036 41157 238100
rect 41091 238035 41157 238036
rect 41275 238100 41341 238101
rect 41275 238036 41276 238100
rect 41340 238036 41341 238100
rect 41275 238035 41341 238036
rect 41459 238100 41525 238101
rect 41459 238036 41460 238100
rect 41524 238036 41525 238100
rect 41459 238035 41525 238036
rect 41643 238100 41709 238101
rect 41643 238036 41644 238100
rect 41708 238036 41709 238100
rect 41643 238035 41709 238036
rect 42195 238100 42261 238101
rect 42195 238036 42196 238100
rect 42260 238036 42261 238100
rect 42195 238035 42261 238036
rect 40542 234502 40786 234562
rect 40542 226133 40602 234502
rect 41094 231870 41154 238035
rect 41278 234837 41338 238035
rect 41275 234836 41341 234837
rect 41275 234772 41276 234836
rect 41340 234772 41341 234836
rect 41275 234771 41341 234772
rect 41462 233341 41522 238035
rect 41459 233340 41525 233341
rect 41459 233276 41460 233340
rect 41524 233276 41525 233340
rect 41459 233275 41525 233276
rect 40726 231810 41154 231870
rect 40726 230485 40786 231810
rect 40723 230484 40789 230485
rect 40723 230420 40724 230484
rect 40788 230420 40789 230484
rect 40723 230419 40789 230420
rect 41646 228989 41706 238035
rect 41643 228988 41709 228989
rect 41643 228924 41644 228988
rect 41708 228924 41709 228988
rect 41643 228923 41709 228924
rect 42198 227357 42258 238035
rect 42563 237964 42629 237965
rect 42563 237900 42564 237964
rect 42628 237900 42629 237964
rect 42563 237899 42629 237900
rect 42566 229941 42626 237899
rect 44196 234547 44248 241343
rect 46724 238579 56406 241343
rect 63362 238579 64653 241375
rect 46724 238490 64653 238579
rect 65209 238490 65252 241446
rect 46724 238466 65252 238490
rect 197542 241446 198398 241470
rect 197542 238490 197619 241446
rect 198335 238490 198398 241446
rect 197542 238480 198398 238490
rect 227642 241446 228498 241470
rect 227642 238490 227719 241446
rect 228435 238490 228498 241446
rect 227642 238480 228498 238490
rect 257742 241446 258598 241470
rect 288068 241446 288566 241470
rect 318226 241446 318574 241470
rect 348042 241446 348898 241470
rect 257742 238490 257819 241446
rect 258535 238490 258598 241446
rect 348042 238490 348119 241446
rect 348835 238490 348898 241446
rect 257742 238480 258598 238490
rect 288068 238480 288566 238490
rect 318226 238480 318574 238490
rect 348042 238480 348898 238490
rect 378042 241446 378898 241470
rect 408410 241446 408734 241470
rect 652538 241451 653158 275876
rect 653498 245453 654118 274916
rect 658950 274532 669812 274574
rect 658950 274525 667288 274532
rect 658950 273969 659025 274525
rect 663101 273969 667288 274525
rect 654458 265439 655078 273956
rect 658950 273938 667288 273969
rect 667216 273176 667288 273938
rect 669764 273176 669812 274532
rect 667216 273138 669812 273176
rect 655418 269441 656038 273004
rect 655418 266485 655447 269441
rect 656003 266485 656038 269441
rect 655418 266386 656038 266485
rect 654458 262483 654489 265439
rect 655045 262483 655078 265439
rect 654458 262362 655078 262483
rect 656378 257435 656998 272036
rect 657338 261453 657958 271082
rect 657338 258497 657363 261453
rect 657919 258497 657958 261453
rect 657338 258390 657958 258497
rect 656378 254479 656401 257435
rect 656957 254479 656998 257435
rect 656378 254386 656998 254479
rect 673870 249661 673930 659907
rect 674419 652220 674485 652221
rect 674419 652156 674420 652220
rect 674484 652156 674485 652220
rect 674419 652155 674485 652156
rect 674422 574157 674482 652155
rect 674606 619445 674666 697307
rect 675342 679013 675402 741643
rect 675526 710837 675586 784755
rect 675707 784276 675773 784277
rect 675707 784212 675708 784276
rect 675772 784212 675773 784276
rect 675707 784211 675773 784212
rect 675710 773397 675770 784211
rect 675707 773396 675773 773397
rect 675707 773332 675708 773396
rect 675772 773332 675773 773396
rect 675707 773331 675773 773332
rect 675894 772717 675954 784891
rect 675891 772716 675957 772717
rect 675891 772652 675892 772716
rect 675956 772652 675957 772716
rect 675891 772651 675957 772652
rect 676078 757213 676138 875875
rect 676075 757212 676141 757213
rect 676075 757148 676076 757212
rect 676140 757148 676141 757212
rect 676075 757147 676141 757148
rect 676262 754765 676322 876555
rect 676443 866828 676509 866829
rect 676443 866764 676444 866828
rect 676508 866764 676509 866828
rect 676443 866763 676509 866764
rect 676259 754764 676325 754765
rect 676259 754700 676260 754764
rect 676324 754700 676325 754764
rect 676259 754699 676325 754700
rect 676446 753541 676506 866763
rect 676627 784140 676693 784141
rect 676627 784076 676628 784140
rect 676692 784076 676693 784140
rect 676627 784075 676693 784076
rect 676443 753540 676509 753541
rect 676443 753476 676444 753540
rect 676508 753476 676509 753540
rect 676443 753475 676509 753476
rect 675710 741030 676322 741090
rect 675710 739261 675770 741030
rect 675891 739940 675957 739941
rect 675891 739876 675892 739940
rect 675956 739876 675957 739940
rect 675891 739875 675957 739876
rect 675707 739260 675773 739261
rect 675707 739196 675708 739260
rect 675772 739196 675773 739260
rect 675707 739195 675773 739196
rect 675523 710836 675589 710837
rect 675523 710772 675524 710836
rect 675588 710772 675589 710836
rect 675523 710771 675589 710772
rect 675707 696964 675773 696965
rect 675707 696900 675708 696964
rect 675772 696900 675773 696964
rect 675707 696899 675773 696900
rect 675339 679012 675405 679013
rect 675339 678948 675340 679012
rect 675404 678948 675405 679012
rect 675339 678947 675405 678948
rect 675523 640388 675589 640389
rect 675523 640324 675524 640388
rect 675588 640324 675589 640388
rect 675523 640323 675589 640324
rect 675526 638213 675586 640323
rect 675523 638212 675589 638213
rect 675523 638148 675524 638212
rect 675588 638148 675589 638212
rect 675523 638147 675589 638148
rect 675710 633453 675770 696899
rect 675894 665685 675954 739875
rect 676262 713490 676322 741030
rect 676078 713430 676322 713490
rect 676078 711109 676138 713430
rect 676075 711108 676141 711109
rect 676075 711044 676076 711108
rect 676140 711044 676141 711108
rect 676075 711043 676141 711044
rect 676630 710970 676690 784075
rect 677179 779924 677245 779925
rect 677179 779860 677180 779924
rect 677244 779860 677245 779924
rect 677179 779859 677245 779860
rect 676811 774892 676877 774893
rect 676811 774828 676812 774892
rect 676876 774828 676877 774892
rect 676811 774827 676877 774828
rect 676814 755989 676874 774827
rect 676811 755988 676877 755989
rect 676811 755924 676812 755988
rect 676876 755924 676877 755988
rect 676811 755923 676877 755924
rect 676811 734364 676877 734365
rect 676811 734300 676812 734364
rect 676876 734300 676877 734364
rect 676811 734299 676877 734300
rect 676078 710910 676690 710970
rect 676078 708933 676138 710910
rect 676075 708932 676141 708933
rect 676075 708868 676076 708932
rect 676140 708868 676141 708932
rect 676075 708867 676141 708868
rect 676259 704444 676325 704445
rect 676259 704380 676260 704444
rect 676324 704380 676325 704444
rect 676259 704379 676325 704380
rect 676075 695060 676141 695061
rect 676075 694996 676076 695060
rect 676140 694996 676141 695060
rect 676075 694995 676141 694996
rect 675891 665684 675957 665685
rect 675891 665620 675892 665684
rect 675956 665620 675957 665684
rect 675891 665619 675957 665620
rect 675891 651540 675957 651541
rect 675891 651476 675892 651540
rect 675956 651476 675957 651540
rect 675891 651475 675957 651476
rect 675707 633452 675773 633453
rect 675707 633388 675708 633452
rect 675772 633388 675773 633452
rect 675707 633387 675773 633388
rect 674603 619444 674669 619445
rect 674603 619380 674604 619444
rect 674668 619380 674669 619444
rect 674603 619379 674669 619380
rect 675894 615510 675954 651475
rect 676078 620805 676138 694995
rect 676262 663373 676322 704379
rect 676443 694244 676509 694245
rect 676443 694180 676444 694244
rect 676508 694180 676509 694244
rect 676443 694179 676509 694180
rect 676259 663372 676325 663373
rect 676259 663308 676260 663372
rect 676324 663308 676325 663372
rect 676259 663307 676325 663308
rect 676259 648684 676325 648685
rect 676259 648620 676260 648684
rect 676324 648620 676325 648684
rect 676259 648619 676325 648620
rect 676075 620804 676141 620805
rect 676075 620740 676076 620804
rect 676140 620740 676141 620804
rect 676075 620739 676141 620740
rect 675894 615450 676138 615510
rect 675523 607884 675589 607885
rect 675523 607820 675524 607884
rect 675588 607820 675589 607884
rect 675523 607819 675589 607820
rect 675339 606524 675405 606525
rect 675339 606460 675340 606524
rect 675404 606460 675405 606524
rect 675339 606459 675405 606460
rect 675342 605845 675402 606459
rect 675339 605844 675405 605845
rect 675339 605780 675340 605844
rect 675404 605780 675405 605844
rect 675339 605779 675405 605780
rect 675526 602850 675586 607819
rect 675707 605844 675773 605845
rect 675707 605780 675708 605844
rect 675772 605780 675773 605844
rect 675707 605779 675773 605780
rect 675710 605570 675770 605779
rect 675710 605510 675954 605570
rect 675158 602790 675586 602850
rect 675158 586530 675218 602790
rect 675707 600948 675773 600949
rect 675707 600884 675708 600948
rect 675772 600884 675773 600948
rect 675707 600883 675773 600884
rect 675523 600268 675589 600269
rect 675523 600204 675524 600268
rect 675588 600204 675589 600268
rect 675523 600203 675589 600204
rect 675526 593197 675586 600203
rect 675710 593197 675770 600883
rect 675523 593196 675589 593197
rect 675523 593132 675524 593196
rect 675588 593132 675589 593196
rect 675523 593131 675589 593132
rect 675707 593196 675773 593197
rect 675707 593132 675708 593196
rect 675772 593132 675773 593196
rect 675707 593131 675773 593132
rect 675894 586530 675954 605510
rect 676078 589253 676138 615450
rect 676075 589252 676141 589253
rect 676075 589188 676076 589252
rect 676140 589188 676141 589252
rect 676075 589187 676141 589188
rect 675158 586470 675586 586530
rect 674419 574156 674485 574157
rect 674419 574092 674420 574156
rect 674484 574092 674485 574156
rect 674419 574091 674485 574092
rect 675339 559604 675405 559605
rect 675339 559540 675340 559604
rect 675404 559540 675405 559604
rect 675339 559539 675405 559540
rect 675342 503573 675402 559539
rect 675526 546549 675586 586470
rect 675710 586470 675954 586530
rect 675523 546548 675589 546549
rect 675523 546484 675524 546548
rect 675588 546484 675589 546548
rect 675523 546483 675589 546484
rect 675710 543829 675770 586470
rect 676262 573205 676322 648619
rect 676446 618765 676506 694179
rect 676814 662965 676874 734299
rect 676995 733004 677061 733005
rect 676995 732940 676996 733004
rect 677060 732940 677061 733004
rect 676995 732939 677061 732940
rect 676998 663373 677058 732939
rect 677182 717630 677242 779859
rect 677182 717570 677426 717630
rect 677366 713493 677426 717570
rect 677363 713492 677429 713493
rect 677363 713428 677364 713492
rect 677428 713428 677429 713492
rect 677363 713427 677429 713428
rect 676995 663372 677061 663373
rect 676995 663308 676996 663372
rect 677060 663308 677061 663372
rect 676995 663307 677061 663308
rect 676811 662964 676877 662965
rect 676811 662900 676812 662964
rect 676876 662900 676877 662964
rect 676811 662899 676877 662900
rect 676627 644740 676693 644741
rect 676627 644676 676628 644740
rect 676692 644676 676693 644740
rect 676627 644675 676693 644676
rect 676443 618764 676509 618765
rect 676443 618700 676444 618764
rect 676508 618700 676509 618764
rect 676443 618699 676509 618700
rect 676443 599044 676509 599045
rect 676443 598980 676444 599044
rect 676508 598980 676509 599044
rect 676443 598979 676509 598980
rect 676259 573204 676325 573205
rect 676259 573140 676260 573204
rect 676324 573140 676325 573204
rect 676259 573139 676325 573140
rect 675891 562732 675957 562733
rect 675891 562668 675892 562732
rect 675956 562668 675957 562732
rect 675891 562667 675957 562668
rect 675707 543828 675773 543829
rect 675707 543764 675708 543828
rect 675772 543764 675773 543828
rect 675707 543763 675773 543764
rect 675894 503709 675954 562667
rect 676075 561236 676141 561237
rect 676075 561172 676076 561236
rect 676140 561172 676141 561236
rect 676075 561171 676141 561172
rect 675891 503708 675957 503709
rect 675891 503644 675892 503708
rect 675956 503644 675957 503708
rect 675891 503643 675957 503644
rect 675339 503572 675405 503573
rect 675339 503508 675340 503572
rect 675404 503508 675405 503572
rect 675339 503507 675405 503508
rect 676078 487797 676138 561171
rect 676259 558380 676325 558381
rect 676259 558316 676260 558380
rect 676324 558316 676325 558380
rect 676259 558315 676325 558316
rect 676075 487796 676141 487797
rect 676075 487732 676076 487796
rect 676140 487732 676141 487796
rect 676075 487731 676141 487732
rect 676262 484635 676322 558315
rect 676446 527781 676506 598979
rect 676630 572797 676690 644675
rect 676995 644604 677061 644605
rect 676995 644540 676996 644604
rect 677060 644540 677061 644604
rect 676995 644539 677061 644540
rect 676811 597820 676877 597821
rect 676811 597756 676812 597820
rect 676876 597756 676877 597820
rect 676811 597755 676877 597756
rect 676627 572796 676693 572797
rect 676627 572732 676628 572796
rect 676692 572732 676693 572796
rect 676627 572731 676693 572732
rect 676627 551988 676693 551989
rect 676627 551924 676628 551988
rect 676692 551924 676693 551988
rect 676627 551923 676693 551924
rect 676443 527780 676509 527781
rect 676443 527716 676444 527780
rect 676508 527716 676509 527780
rect 676443 527715 676509 527716
rect 676259 484634 676325 484635
rect 676259 484570 676260 484634
rect 676324 484570 676325 484634
rect 676259 484569 676325 484570
rect 676075 483852 676141 483853
rect 676075 483788 676076 483852
rect 676140 483850 676141 483852
rect 676630 483850 676690 551923
rect 676814 528189 676874 597755
rect 676998 573205 677058 644539
rect 676995 573204 677061 573205
rect 676995 573140 676996 573204
rect 677060 573140 677061 573204
rect 676995 573139 677061 573140
rect 676995 568580 677061 568581
rect 676995 568516 676996 568580
rect 677060 568516 677061 568580
rect 676995 568515 677061 568516
rect 676998 530229 677058 568515
rect 676995 530228 677061 530229
rect 676995 530164 676996 530228
rect 677060 530164 677061 530228
rect 676995 530163 677061 530164
rect 676811 528188 676877 528189
rect 676811 528124 676812 528188
rect 676876 528124 676877 528188
rect 676811 528123 676877 528124
rect 676140 483790 676690 483850
rect 676140 483788 676141 483790
rect 676075 483787 676141 483788
rect 675707 399396 675773 399397
rect 675707 399332 675708 399396
rect 675772 399332 675773 399396
rect 675707 399331 675773 399332
rect 675523 388516 675589 388517
rect 675523 388452 675524 388516
rect 675588 388452 675589 388516
rect 675523 388451 675589 388452
rect 675339 388244 675405 388245
rect 675339 388180 675340 388244
rect 675404 388180 675405 388244
rect 675339 388179 675405 388180
rect 675342 382261 675402 388179
rect 675339 382260 675405 382261
rect 675339 382196 675340 382260
rect 675404 382196 675405 382260
rect 675339 382195 675405 382196
rect 675526 378725 675586 388451
rect 675710 384981 675770 399331
rect 676259 398852 676325 398853
rect 676259 398788 676260 398852
rect 676324 398788 676325 398852
rect 676259 398787 676325 398788
rect 676075 395588 676141 395589
rect 676075 395524 676076 395588
rect 676140 395524 676141 395588
rect 676075 395523 676141 395524
rect 675891 395316 675957 395317
rect 675891 395252 675892 395316
rect 675956 395252 675957 395316
rect 675891 395251 675957 395252
rect 675707 384980 675773 384981
rect 675707 384916 675708 384980
rect 675772 384916 675773 384980
rect 675707 384915 675773 384916
rect 675523 378724 675589 378725
rect 675523 378660 675524 378724
rect 675588 378660 675589 378724
rect 675523 378659 675589 378660
rect 675894 377365 675954 395251
rect 675891 377364 675957 377365
rect 675891 377300 675892 377364
rect 675956 377300 675957 377364
rect 675891 377299 675957 377300
rect 676078 375053 676138 395523
rect 676075 375052 676141 375053
rect 676075 374988 676076 375052
rect 676140 374988 676141 375052
rect 676075 374987 676141 374988
rect 676262 373693 676322 398787
rect 676443 397220 676509 397221
rect 676443 397156 676444 397220
rect 676508 397156 676509 397220
rect 676443 397155 676509 397156
rect 676259 373692 676325 373693
rect 676259 373628 676260 373692
rect 676324 373628 676325 373692
rect 676259 373627 676325 373628
rect 676446 372061 676506 397155
rect 676443 372060 676509 372061
rect 676443 371996 676444 372060
rect 676508 371996 676509 372060
rect 676443 371995 676509 371996
rect 675891 354244 675957 354245
rect 675891 354180 675892 354244
rect 675956 354180 675957 354244
rect 675891 354179 675957 354180
rect 675707 353428 675773 353429
rect 675707 353364 675708 353428
rect 675772 353364 675773 353428
rect 675707 353363 675773 353364
rect 675339 353020 675405 353021
rect 675339 352956 675340 353020
rect 675404 352956 675405 353020
rect 675339 352955 675405 352956
rect 675342 337925 675402 352955
rect 675710 340781 675770 353363
rect 675707 340780 675773 340781
rect 675707 340716 675708 340780
rect 675772 340716 675773 340780
rect 675707 340715 675773 340716
rect 675894 339421 675954 354179
rect 676075 353700 676141 353701
rect 676075 353636 676076 353700
rect 676140 353698 676141 353700
rect 676140 353638 676506 353698
rect 676140 353636 676141 353638
rect 676075 353635 676141 353636
rect 676075 352068 676141 352069
rect 676075 352004 676076 352068
rect 676140 352004 676141 352068
rect 676075 352003 676141 352004
rect 676078 351930 676138 352003
rect 676078 351870 676322 351930
rect 676075 342412 676141 342413
rect 676075 342348 676076 342412
rect 676140 342348 676141 342412
rect 676075 342347 676141 342348
rect 675891 339420 675957 339421
rect 675891 339356 675892 339420
rect 675956 339356 675957 339420
rect 675891 339355 675957 339356
rect 675339 337924 675405 337925
rect 675339 337860 675340 337924
rect 675404 337860 675405 337924
rect 675339 337859 675405 337860
rect 676078 333573 676138 342347
rect 676075 333572 676141 333573
rect 676075 333508 676076 333572
rect 676140 333508 676141 333572
rect 676075 333507 676141 333508
rect 676262 325549 676322 351870
rect 676446 325685 676506 353638
rect 676995 346628 677061 346629
rect 676995 346564 676996 346628
rect 677060 346564 677061 346628
rect 676995 346563 677061 346564
rect 676627 346492 676693 346493
rect 676627 346428 676628 346492
rect 676692 346428 676693 346492
rect 676627 346427 676693 346428
rect 676811 346492 676877 346493
rect 676811 346428 676812 346492
rect 676876 346428 676877 346492
rect 676811 346427 676877 346428
rect 676630 332621 676690 346427
rect 676814 335341 676874 346427
rect 676998 335885 677058 346563
rect 676995 335884 677061 335885
rect 676995 335820 676996 335884
rect 677060 335820 677061 335884
rect 676995 335819 677061 335820
rect 676811 335340 676877 335341
rect 676811 335276 676812 335340
rect 676876 335276 676877 335340
rect 676811 335275 676877 335276
rect 676627 332620 676693 332621
rect 676627 332556 676628 332620
rect 676692 332556 676693 332620
rect 676627 332555 676693 332556
rect 676443 325684 676509 325685
rect 676443 325620 676444 325684
rect 676508 325620 676509 325684
rect 676443 325619 676509 325620
rect 676259 325548 676325 325549
rect 676259 325484 676260 325548
rect 676324 325484 676325 325548
rect 676259 325483 676325 325484
rect 676443 308684 676509 308685
rect 676443 308620 676444 308684
rect 676508 308620 676509 308684
rect 676443 308619 676509 308620
rect 676075 307460 676141 307461
rect 676075 307396 676076 307460
rect 676140 307396 676141 307460
rect 676075 307395 676141 307396
rect 675891 299436 675957 299437
rect 675891 299372 675892 299436
rect 675956 299372 675957 299436
rect 675891 299371 675957 299372
rect 675707 297804 675773 297805
rect 675707 297740 675708 297804
rect 675772 297740 675773 297804
rect 675707 297739 675773 297740
rect 675339 297532 675405 297533
rect 675339 297468 675340 297532
rect 675404 297468 675405 297532
rect 675339 297467 675405 297468
rect 675342 285565 675402 297467
rect 675523 297396 675589 297397
rect 675523 297332 675524 297396
rect 675588 297332 675589 297396
rect 675523 297331 675589 297332
rect 675526 292093 675586 297331
rect 675710 292637 675770 297739
rect 675894 294813 675954 299371
rect 675891 294812 675957 294813
rect 675891 294748 675892 294812
rect 675956 294748 675957 294812
rect 675891 294747 675957 294748
rect 675707 292636 675773 292637
rect 675707 292572 675708 292636
rect 675772 292572 675773 292636
rect 675707 292571 675773 292572
rect 675523 292092 675589 292093
rect 675523 292028 675524 292092
rect 675588 292028 675589 292092
rect 675523 292027 675589 292028
rect 676078 288421 676138 307395
rect 676259 307052 676325 307053
rect 676259 306988 676260 307052
rect 676324 306988 676325 307052
rect 676259 306987 676325 306988
rect 676075 288420 676141 288421
rect 676075 288356 676076 288420
rect 676140 288356 676141 288420
rect 676075 288355 676141 288356
rect 675339 285564 675405 285565
rect 675339 285500 675340 285564
rect 675404 285500 675405 285564
rect 675339 285499 675405 285500
rect 676262 281485 676322 306987
rect 676446 283661 676506 308619
rect 676627 305012 676693 305013
rect 676627 304948 676628 305012
rect 676692 304948 676693 305012
rect 676627 304947 676693 304948
rect 676630 287333 676690 304947
rect 676627 287332 676693 287333
rect 676627 287268 676628 287332
rect 676692 287268 676693 287332
rect 676627 287267 676693 287268
rect 676443 283660 676509 283661
rect 676443 283596 676444 283660
rect 676508 283596 676509 283660
rect 676443 283595 676509 283596
rect 676259 281484 676325 281485
rect 676259 281420 676260 281484
rect 676324 281420 676325 281484
rect 676259 281419 676325 281420
rect 675891 264212 675957 264213
rect 675891 264148 675892 264212
rect 675956 264148 675957 264212
rect 675891 264147 675957 264148
rect 675707 262988 675773 262989
rect 675707 262924 675708 262988
rect 675772 262924 675773 262988
rect 675707 262923 675773 262924
rect 674787 252652 674853 252653
rect 674787 252588 674788 252652
rect 674852 252588 674853 252652
rect 674787 252587 674853 252588
rect 674790 249797 674850 252587
rect 674787 249796 674853 249797
rect 674787 249732 674788 249796
rect 674852 249732 674853 249796
rect 674787 249731 674853 249732
rect 675710 249661 675770 262923
rect 675894 249797 675954 264147
rect 676995 263634 677061 263635
rect 676995 263570 676996 263634
rect 677060 263570 677061 263634
rect 676995 263569 677061 263570
rect 676075 260404 676141 260405
rect 676075 260340 676076 260404
rect 676140 260340 676141 260404
rect 676075 260339 676141 260340
rect 675891 249796 675957 249797
rect 675891 249732 675892 249796
rect 675956 249732 675957 249796
rect 675891 249731 675957 249732
rect 676078 249661 676138 260339
rect 676443 251564 676509 251565
rect 676443 251500 676444 251564
rect 676508 251500 676509 251564
rect 676443 251499 676509 251500
rect 676446 250341 676506 251499
rect 676443 250340 676509 250341
rect 676443 250276 676444 250340
rect 676508 250276 676509 250340
rect 676443 250275 676509 250276
rect 673867 249660 673933 249661
rect 673867 249596 673868 249660
rect 673932 249596 673933 249660
rect 673867 249595 673933 249596
rect 675707 249660 675773 249661
rect 675707 249596 675708 249660
rect 675772 249596 675773 249660
rect 675707 249595 675773 249596
rect 676075 249660 676141 249661
rect 676075 249596 676076 249660
rect 676140 249596 676141 249660
rect 676075 249595 676141 249596
rect 666890 249354 676670 249476
rect 666890 249293 674146 249354
rect 666890 246657 667032 249293
rect 669668 246657 674146 249293
rect 666890 246558 674146 246657
rect 676462 246558 676670 249354
rect 666890 246466 676670 246558
rect 674971 246260 675037 246261
rect 674971 246196 674972 246260
rect 675036 246196 675037 246260
rect 674971 246195 675037 246196
rect 675339 246260 675405 246261
rect 675339 246196 675340 246260
rect 675404 246196 675405 246260
rect 675339 246195 675405 246196
rect 673867 246124 673933 246125
rect 673867 246060 673868 246124
rect 673932 246060 673933 246124
rect 673867 246059 673933 246060
rect 653498 242497 653519 245453
rect 654075 242497 654118 245453
rect 653498 242362 654118 242497
rect 378042 238490 378119 241446
rect 378835 238490 378898 241446
rect 652538 238495 652561 241451
rect 653117 238495 653158 241451
rect 378042 238480 378898 238490
rect 408410 238480 408734 238490
rect 46724 234547 46802 238466
rect 64632 238400 65252 238466
rect 652538 238266 653158 238495
rect 44196 234466 46802 234547
rect 47786 237381 63250 237466
rect 47786 237375 56375 237381
rect 47786 234579 47931 237375
rect 50727 234585 56375 237375
rect 63171 234585 63250 237381
rect 50727 234579 63250 234585
rect 47786 234466 63250 234579
rect 210866 237441 211814 237474
rect 210866 234485 210902 237441
rect 211778 234485 211814 237441
rect 210866 234448 211814 234485
rect 240966 237441 241914 237474
rect 240966 234485 241002 237441
rect 241878 234485 241914 237441
rect 240966 234448 241914 234485
rect 271344 237441 272014 237474
rect 331414 237441 332214 237474
rect 271344 234485 271355 237441
rect 271911 234485 272014 237441
rect 302046 234517 302114 237290
rect 271344 234448 272014 234485
rect 301514 234448 302114 234517
rect 332126 234485 332214 237441
rect 331414 234448 332214 234485
rect 361366 237441 362314 237474
rect 391834 237441 392314 237474
rect 361366 234485 361402 237441
rect 362278 234485 362314 237441
rect 392226 234485 392314 237441
rect 361366 234448 362314 234485
rect 391834 234448 392314 234485
rect 44186 233371 63160 233466
rect 44186 230575 56394 233371
rect 63030 230575 63160 233371
rect 89776 232124 90096 233636
rect 93776 232124 94096 233606
rect 89776 232086 94096 232124
rect 89776 231370 89903 232086
rect 93979 231370 94096 232086
rect 89776 231308 94096 231370
rect 169776 232162 170096 233642
rect 173776 232162 174096 233642
rect 169776 232108 174096 232162
rect 169776 231392 169887 232108
rect 173963 231392 174096 232108
rect 169776 231346 174096 231392
rect 195988 233442 196616 233464
rect 44186 230466 63160 230575
rect 195988 230486 196029 233442
rect 196585 230486 196616 233442
rect 195988 230466 196616 230486
rect 226088 233442 226716 233464
rect 226088 230486 226129 233442
rect 226685 230486 226716 233442
rect 226088 230466 226716 230486
rect 256188 233442 256816 233464
rect 256188 230486 256229 233442
rect 256785 230486 256816 233442
rect 256188 230466 256816 230486
rect 286288 233442 286916 233464
rect 286288 230486 286329 233442
rect 286885 230486 286916 233442
rect 286288 230466 286916 230486
rect 316388 233442 317016 233464
rect 316388 230486 316429 233442
rect 316985 230486 317016 233442
rect 316388 230466 317016 230486
rect 346488 233442 347116 233464
rect 346488 230486 346529 233442
rect 347085 230486 347116 233442
rect 346488 230466 347116 230486
rect 376488 233442 377116 233464
rect 376488 230486 376529 233442
rect 377085 230486 377116 233442
rect 376488 230466 377116 230486
rect 406660 233442 407116 233464
rect 407056 230486 407116 233442
rect 429776 232184 430096 233640
rect 433776 232184 434096 233610
rect 429776 232120 434096 232184
rect 429776 231404 429905 232120
rect 433981 231404 434096 232120
rect 429776 231368 434096 231404
rect 406660 230466 407116 230486
rect 647739 230484 647805 230485
rect 42563 229940 42629 229941
rect 42563 229876 42564 229940
rect 42628 229876 42629 229940
rect 42563 229875 42629 229876
rect 42195 227356 42261 227357
rect 42195 227292 42196 227356
rect 42260 227292 42261 227356
rect 42195 227291 42261 227292
rect 40539 226132 40605 226133
rect 40539 226068 40540 226132
rect 40604 226068 40605 226132
rect 40539 226067 40605 226068
rect 6106 221353 6906 221470
rect 6106 220209 6150 221353
rect 6854 220209 6906 221353
rect 6106 211943 6906 220209
rect 7306 219757 8106 219842
rect 7306 218613 7348 219757
rect 8052 218613 8106 219757
rect 7306 213635 8106 218613
rect 6106 208577 6906 211547
rect 7306 210255 8106 213239
rect 6106 205187 6906 208181
rect 7306 206875 8106 209859
rect 40539 209404 40605 209405
rect 40539 209340 40540 209404
rect 40604 209340 40605 209404
rect 40539 209339 40605 209340
rect 7306 206476 8106 206479
rect 6106 204746 6906 204791
rect 40542 183021 40602 209339
rect 41459 208588 41525 208589
rect 41459 208524 41460 208588
rect 41524 208524 41525 208588
rect 41459 208523 41525 208524
rect 40723 206956 40789 206957
rect 40723 206892 40724 206956
rect 40788 206892 40789 206956
rect 40723 206891 40789 206892
rect 40726 194717 40786 206891
rect 40723 194716 40789 194717
rect 40723 194652 40724 194716
rect 40788 194652 40789 194716
rect 40723 194651 40789 194652
rect 41462 190229 41522 208523
rect 41643 199476 41709 199477
rect 41643 199412 41644 199476
rect 41708 199412 41709 199476
rect 41643 199411 41709 199412
rect 41646 195261 41706 199411
rect 41827 199340 41893 199341
rect 41827 199276 41828 199340
rect 41892 199276 41893 199340
rect 41827 199275 41893 199276
rect 41643 195260 41709 195261
rect 41643 195196 41644 195260
rect 41708 195196 41709 195260
rect 41643 195195 41709 195196
rect 41830 194850 41890 199275
rect 41646 194790 41890 194850
rect 44198 197498 46798 230466
rect 647739 230420 647740 230484
rect 647804 230420 647805 230484
rect 647739 230419 647805 230420
rect 54184 220199 54189 221388
rect 55385 220199 55390 221388
rect 54184 220174 55390 220199
rect 52580 219777 53786 219788
rect 52580 218581 52595 219777
rect 52580 218574 53786 218581
rect 647742 213077 647802 230419
rect 647739 213076 647805 213077
rect 647739 213012 647740 213076
rect 647804 213012 647805 213076
rect 647739 213011 647805 213012
rect 598368 212351 610962 212504
rect 598368 209715 598610 212351
rect 601086 209715 607464 212351
rect 609940 209715 610962 212351
rect 598368 209504 610962 209715
rect 641044 212394 642108 212460
rect 641044 209598 641143 212394
rect 642019 209598 642108 212394
rect 641044 209528 642108 209598
rect 596262 208462 605388 208502
rect 596262 207906 596320 208462
rect 597676 207906 602413 208462
rect 605369 207906 605388 208462
rect 596262 207862 605388 207906
rect 610642 207692 610962 209504
rect 641362 207684 641682 209528
rect 598496 197801 601174 197876
rect 44198 197472 52344 197498
rect 44198 196916 51413 197472
rect 52289 196916 52344 197472
rect 598496 197085 598703 197801
rect 601019 197528 601174 197801
rect 601019 197483 606976 197528
rect 601019 197247 605958 197483
rect 601019 197208 606976 197247
rect 601019 197085 601174 197208
rect 598496 196992 601174 197085
rect 44198 196858 52344 196916
rect 41459 190228 41525 190229
rect 41459 190164 41460 190228
rect 41524 190164 41525 190228
rect 41459 190163 41525 190164
rect 41646 184109 41706 194790
rect 41827 194716 41893 194717
rect 41827 194652 41828 194716
rect 41892 194652 41893 194716
rect 41827 194651 41893 194652
rect 41830 187373 41890 194651
rect 41827 187372 41893 187373
rect 41827 187308 41828 187372
rect 41892 187308 41893 187372
rect 41827 187307 41893 187308
rect 41643 184108 41709 184109
rect 41643 184044 41644 184108
rect 41708 184044 41709 184108
rect 41643 184043 41709 184044
rect 40539 183020 40605 183021
rect 40539 182956 40540 183020
rect 40604 182956 40605 183020
rect 40539 182955 40605 182956
rect 44198 176742 46798 196858
rect 596072 184450 605388 184502
rect 596072 183894 596124 184450
rect 596840 184446 605388 184450
rect 596840 183894 602413 184446
rect 596072 183890 602413 183894
rect 605369 183890 605388 184446
rect 596072 183862 605388 183890
rect 41864 176665 46798 176742
rect 41864 173229 42007 176665
rect 45603 173229 46798 176665
rect 41864 173126 46798 173229
rect 42646 171458 52246 171498
rect 42646 171454 51305 171458
rect 42646 170898 42777 171454
rect 45733 170902 51305 171454
rect 52181 170902 52246 171458
rect 45733 170898 52246 170902
rect 42646 170858 52246 170898
rect 673870 168605 673930 246059
rect 674974 241909 675034 246195
rect 674971 241908 675037 241909
rect 674971 241844 674972 241908
rect 675036 241844 675037 241908
rect 674971 241843 675037 241844
rect 675342 240277 675402 246195
rect 675339 240276 675405 240277
rect 675339 240212 675340 240276
rect 675404 240212 675405 240276
rect 675339 240211 675405 240212
rect 676998 238509 677058 263569
rect 677179 262036 677245 262037
rect 677179 261972 677180 262036
rect 677244 261972 677245 262036
rect 677179 261971 677245 261972
rect 676995 238508 677061 238509
rect 676995 238444 676996 238508
rect 677060 238444 677061 238508
rect 676995 238443 677061 238444
rect 677182 236877 677242 261971
rect 677363 261628 677429 261629
rect 677363 261564 677364 261628
rect 677428 261564 677429 261628
rect 677363 261563 677429 261564
rect 677366 251565 677426 261563
rect 677363 251564 677429 251565
rect 677363 251500 677364 251564
rect 677428 251500 677429 251564
rect 677363 251499 677429 251500
rect 677179 236876 677245 236877
rect 677179 236812 677180 236876
rect 677244 236812 677245 236876
rect 677179 236811 677245 236812
rect 676029 218652 676095 218653
rect 676029 218588 676030 218652
rect 676094 218650 676095 218652
rect 676094 218590 676506 218650
rect 676094 218588 676095 218590
rect 676029 218587 676095 218588
rect 675339 218244 675405 218245
rect 675339 218180 675340 218244
rect 675404 218180 675405 218244
rect 675339 218179 675405 218180
rect 675342 205597 675402 218179
rect 675891 217836 675957 217837
rect 675891 217772 675892 217836
rect 675956 217772 675957 217836
rect 675891 217771 675957 217772
rect 675707 214028 675773 214029
rect 675707 213964 675708 214028
rect 675772 213964 675773 214028
rect 675707 213963 675773 213964
rect 675523 207228 675589 207229
rect 675523 207164 675524 207228
rect 675588 207164 675589 207228
rect 675523 207163 675589 207164
rect 675339 205596 675405 205597
rect 675339 205532 675340 205596
rect 675404 205532 675405 205596
rect 675339 205531 675405 205532
rect 675526 198389 675586 207163
rect 675710 204237 675770 213963
rect 675707 204236 675773 204237
rect 675707 204172 675708 204236
rect 675772 204172 675773 204236
rect 675707 204171 675773 204172
rect 675894 202741 675954 217771
rect 676075 216884 676141 216885
rect 676075 216820 676076 216884
rect 676140 216820 676141 216884
rect 676075 216819 676141 216820
rect 676078 216610 676138 216819
rect 676078 216550 676322 216610
rect 676075 208316 676141 208317
rect 676075 208252 676076 208316
rect 676140 208252 676141 208316
rect 676075 208251 676141 208252
rect 676078 205053 676138 208251
rect 676075 205052 676141 205053
rect 676075 204988 676076 205052
rect 676140 204988 676141 205052
rect 676075 204987 676141 204988
rect 675891 202740 675957 202741
rect 675891 202676 675892 202740
rect 675956 202676 675957 202740
rect 675891 202675 675957 202676
rect 675523 198388 675589 198389
rect 675523 198324 675524 198388
rect 675588 198324 675589 198388
rect 675523 198323 675589 198324
rect 676262 190365 676322 216550
rect 676259 190364 676325 190365
rect 676259 190300 676260 190364
rect 676324 190300 676325 190364
rect 676259 190299 676325 190300
rect 676446 190229 676506 218590
rect 676995 214334 677061 214335
rect 676995 214270 676996 214334
rect 677060 214270 677061 214334
rect 676995 214269 677061 214270
rect 676627 211444 676693 211445
rect 676627 211380 676628 211444
rect 676692 211380 676693 211444
rect 676627 211379 676693 211380
rect 676630 195397 676690 211379
rect 676811 211308 676877 211309
rect 676811 211244 676812 211308
rect 676876 211244 676877 211308
rect 676811 211243 676877 211244
rect 676814 201381 676874 211243
rect 676998 202877 677058 214269
rect 676995 202876 677061 202877
rect 676995 202812 676996 202876
rect 677060 202812 677061 202876
rect 676995 202811 677061 202812
rect 676811 201380 676877 201381
rect 676811 201316 676812 201380
rect 676876 201316 676877 201380
rect 676811 201315 676877 201316
rect 676627 195396 676693 195397
rect 676627 195332 676628 195396
rect 676692 195332 676693 195396
rect 676627 195331 676693 195332
rect 676443 190228 676509 190229
rect 676443 190164 676444 190228
rect 676508 190164 676509 190228
rect 676443 190163 676509 190164
rect 676078 173710 676322 173770
rect 676078 173501 676138 173710
rect 676075 173500 676141 173501
rect 676075 173436 676076 173500
rect 676140 173436 676141 173500
rect 676075 173435 676141 173436
rect 676262 173090 676322 173710
rect 676262 173030 676506 173090
rect 675891 172820 675957 172821
rect 675891 172756 675892 172820
rect 675956 172756 675957 172820
rect 675891 172755 675957 172756
rect 673867 168604 673933 168605
rect 673867 168540 673868 168604
rect 673932 168540 673933 168604
rect 673867 168539 673933 168540
rect 598496 167161 601174 167236
rect 598496 166445 598703 167161
rect 601019 166892 601174 167161
rect 675894 167010 675954 172755
rect 676075 171868 676141 171869
rect 676075 171804 676076 171868
rect 676140 171804 676141 171868
rect 676075 171803 676141 171804
rect 676078 171730 676138 171803
rect 676078 171670 676322 171730
rect 675894 166950 676138 167010
rect 601019 166855 606976 166892
rect 601019 166619 605941 166855
rect 601019 166572 606976 166619
rect 601019 166445 601174 166572
rect 598496 166352 601174 166445
rect 675523 162756 675589 162757
rect 675523 162692 675524 162756
rect 675588 162692 675589 162756
rect 675523 162691 675589 162692
rect 675339 162348 675405 162349
rect 675339 162284 675340 162348
rect 675404 162284 675405 162348
rect 675339 162283 675405 162284
rect 594072 158458 605388 158502
rect 594072 158454 602387 158458
rect 594072 157898 594082 158454
rect 596878 157902 602387 158454
rect 605343 157902 605388 158458
rect 596878 157898 605388 157902
rect 594072 157862 605388 157898
rect 675342 153101 675402 162283
rect 675526 156501 675586 162691
rect 675891 162620 675957 162621
rect 675891 162556 675892 162620
rect 675956 162556 675957 162620
rect 675891 162555 675957 162556
rect 675707 162484 675773 162485
rect 675707 162420 675708 162484
rect 675772 162420 675773 162484
rect 675707 162419 675773 162420
rect 675710 157045 675770 162419
rect 675894 159493 675954 162555
rect 675891 159492 675957 159493
rect 675891 159428 675892 159492
rect 675956 159428 675957 159492
rect 675891 159427 675957 159428
rect 676078 157453 676138 166950
rect 676075 157452 676141 157453
rect 676075 157388 676076 157452
rect 676140 157388 676141 157452
rect 676075 157387 676141 157388
rect 675707 157044 675773 157045
rect 675707 156980 675708 157044
rect 675772 156980 675773 157044
rect 675707 156979 675773 156980
rect 675523 156500 675589 156501
rect 675523 156436 675524 156500
rect 675588 156436 675589 156500
rect 675523 156435 675589 156436
rect 675339 153100 675405 153101
rect 675339 153036 675340 153100
rect 675404 153036 675405 153100
rect 675339 153035 675405 153036
rect 676262 146301 676322 171670
rect 676446 148477 676506 173030
rect 676627 166428 676693 166429
rect 676627 166364 676628 166428
rect 676692 166364 676693 166428
rect 676627 166363 676693 166364
rect 676811 166428 676877 166429
rect 676811 166364 676812 166428
rect 676876 166364 676877 166428
rect 676811 166363 676877 166364
rect 676630 151605 676690 166363
rect 676814 160037 676874 166363
rect 676811 160036 676877 160037
rect 676811 159972 676812 160036
rect 676876 159972 676877 160036
rect 676811 159971 676877 159972
rect 676627 151604 676693 151605
rect 676627 151540 676628 151604
rect 676692 151540 676693 151604
rect 676627 151539 676693 151540
rect 676443 148476 676509 148477
rect 676443 148412 676444 148476
rect 676508 148412 676509 148476
rect 676443 148411 676509 148412
rect 676259 146300 676325 146301
rect 676259 146236 676260 146300
rect 676324 146236 676325 146300
rect 676259 146235 676325 146236
rect 42578 145460 52178 145498
rect 42578 144904 42791 145460
rect 45747 145450 52178 145460
rect 45747 144904 51239 145450
rect 42578 144894 51239 144904
rect 52115 144894 52178 145450
rect 42578 144858 52178 144894
rect 598496 136521 601174 136596
rect 598496 135805 598703 136521
rect 601019 136256 601174 136521
rect 601019 136215 606976 136256
rect 601019 135979 605931 136215
rect 606967 135979 606976 136215
rect 601019 135936 606976 135979
rect 601019 135805 601174 135936
rect 598496 135712 601174 135805
rect 594072 132448 605388 132502
rect 594072 131892 594092 132448
rect 596888 132442 605388 132448
rect 596888 131892 602413 132442
rect 594072 131886 602413 131892
rect 605369 131886 605388 132442
rect 594072 131862 605388 131886
rect 676075 128620 676141 128621
rect 676075 128556 676076 128620
rect 676140 128556 676141 128620
rect 676075 128555 676141 128556
rect 675891 124948 675957 124949
rect 675891 124884 675892 124948
rect 675956 124884 675957 124948
rect 675891 124883 675957 124884
rect 42578 119456 52178 119498
rect 42578 118900 42781 119456
rect 45737 118900 51235 119456
rect 52111 118900 52178 119456
rect 42578 118858 52178 118900
rect 675707 118012 675773 118013
rect 675707 117948 675708 118012
rect 675772 117948 675773 118012
rect 675707 117947 675773 117948
rect 675339 117332 675405 117333
rect 675339 117268 675340 117332
rect 675404 117268 675405 117332
rect 675339 117267 675405 117268
rect 594072 106454 605388 106502
rect 594072 105898 594094 106454
rect 596890 105898 602417 106454
rect 605373 105898 605388 106454
rect 594072 105862 605388 105898
rect 598496 105620 601174 105676
rect 598496 105601 606976 105620
rect 598496 104885 598703 105601
rect 601019 105578 606976 105601
rect 601019 105342 605943 105578
rect 601019 105300 606976 105342
rect 601019 104885 601174 105300
rect 598496 104792 601174 104885
rect 675342 104821 675402 117267
rect 675523 117196 675589 117197
rect 675523 117132 675524 117196
rect 675588 117132 675589 117196
rect 675523 117131 675589 117132
rect 675526 111757 675586 117131
rect 675523 111756 675589 111757
rect 675523 111692 675524 111756
rect 675588 111692 675589 111756
rect 675523 111691 675589 111692
rect 675710 108221 675770 117947
rect 675894 112573 675954 124883
rect 676078 114205 676138 128555
rect 676259 126580 676325 126581
rect 676259 126516 676260 126580
rect 676324 126516 676325 126580
rect 676259 126515 676325 126516
rect 676075 114204 676141 114205
rect 676075 114140 676076 114204
rect 676140 114140 676141 114204
rect 676075 114139 676141 114140
rect 675891 112572 675957 112573
rect 675891 112508 675892 112572
rect 675956 112508 675957 112572
rect 675891 112507 675957 112508
rect 675707 108220 675773 108221
rect 675707 108156 675708 108220
rect 675772 108156 675773 108220
rect 675707 108155 675773 108156
rect 675339 104820 675405 104821
rect 675339 104756 675340 104820
rect 675404 104756 675405 104820
rect 675339 104755 675405 104756
rect 626002 98760 626322 102316
rect 656722 98804 657042 102238
rect 676262 101421 676322 126515
rect 676443 124540 676509 124541
rect 676443 124476 676444 124540
rect 676508 124476 676509 124540
rect 676443 124475 676509 124476
rect 676446 109037 676506 124475
rect 676811 121684 676877 121685
rect 676811 121620 676812 121684
rect 676876 121620 676877 121684
rect 676811 121619 676877 121620
rect 676443 109036 676509 109037
rect 676443 108972 676444 109036
rect 676508 108972 676509 109036
rect 676443 108971 676509 108972
rect 676814 103189 676874 121619
rect 676811 103188 676877 103189
rect 676811 103124 676812 103188
rect 676876 103124 676877 103188
rect 676811 103123 676877 103124
rect 676259 101420 676325 101421
rect 676259 101356 676260 101420
rect 676324 101356 676325 101420
rect 676259 101355 676325 101356
rect 625442 98683 626852 98760
rect 625442 96047 625552 98683
rect 626748 96047 626852 98683
rect 636080 98681 636994 98758
rect 636080 96525 636179 98681
rect 636895 96525 636994 98681
rect 656284 98745 657602 98804
rect 641667 96660 641733 96661
rect 641667 96596 641668 96660
rect 641732 96596 641733 96660
rect 641667 96595 641733 96596
rect 636080 96434 636994 96525
rect 639827 96524 639893 96525
rect 639827 96460 639828 96524
rect 639892 96460 639893 96524
rect 639827 96459 639893 96460
rect 625442 95956 626852 96047
rect 636354 94448 636674 96434
rect 42578 93454 52178 93498
rect 42578 92898 42777 93454
rect 45733 93452 52178 93454
rect 45733 92898 51239 93452
rect 42578 92896 51239 92898
rect 52115 92896 52178 93452
rect 42578 92858 52178 92896
rect 41864 82752 45778 82794
rect 41864 78196 41931 82752
rect 45687 78196 45778 82752
rect 632354 80924 632674 82062
rect 632072 80789 633010 80924
rect 594072 80466 605388 80502
rect 594072 80464 602411 80466
rect 594072 79908 594088 80464
rect 596884 79910 602411 80464
rect 605367 79910 605388 80466
rect 596884 79908 605388 79910
rect 594072 79862 605388 79908
rect 632072 78313 632174 80789
rect 632890 78313 633010 80789
rect 632072 78198 633010 78313
rect 41864 78154 45778 78196
rect 634678 77893 634738 94062
rect 634675 77892 634741 77893
rect 634675 77828 634676 77892
rect 634740 77828 634741 77892
rect 634675 77827 634741 77828
rect 639830 77757 639890 96459
rect 641670 94298 641730 96595
rect 656284 96109 656363 98745
rect 657559 96109 657602 98745
rect 656284 96050 657602 96109
rect 640354 81016 640674 82000
rect 640098 80896 640922 81016
rect 640098 78260 640152 80896
rect 640868 78260 640922 80896
rect 640098 78134 640922 78260
rect 639827 77756 639893 77757
rect 639827 77692 639828 77756
rect 639892 77692 639893 77756
rect 639827 77691 639893 77692
rect 629888 77193 630208 77374
rect 629888 76317 629919 77193
rect 630155 76317 630208 77193
rect 629888 74104 630208 76317
rect 631438 75791 631758 77374
rect 631438 74915 631471 75791
rect 631707 74915 631758 75791
rect 631438 74104 631758 74915
rect 632988 77207 633308 77374
rect 632988 76331 633031 77207
rect 633267 76331 633308 77207
rect 632988 74104 633308 76331
rect 634538 75795 634858 77374
rect 634538 74919 634565 75795
rect 634801 74919 634858 75795
rect 634538 74104 634858 74919
rect 636088 77203 636408 77374
rect 636088 76327 636121 77203
rect 636357 76327 636408 77203
rect 636088 74104 636408 76327
rect 637638 75799 637958 77374
rect 637638 74923 637673 75799
rect 637909 74923 637958 75799
rect 639188 77203 639508 77374
rect 639188 76327 639215 77203
rect 639451 76327 639508 77203
rect 638907 75172 638973 75173
rect 638907 75108 638908 75172
rect 638972 75108 638973 75172
rect 638907 75107 638973 75108
rect 637638 74104 637958 74923
rect 41858 72848 45772 72890
rect 41858 68292 41907 72848
rect 45663 68292 45772 72848
rect 41858 68250 45772 68292
rect 41862 67454 52362 67498
rect 41862 67448 51437 67454
rect 41862 66892 41935 67448
rect 45691 66898 51437 67448
rect 52313 66898 52362 67454
rect 45691 66892 52362 66898
rect 41862 66858 52362 66892
rect 41874 51994 58536 52122
rect 41874 48398 42000 51994
rect 45596 51960 58536 51994
rect 45596 48398 54490 51960
rect 41874 48364 54490 48398
rect 58246 48364 58536 51960
rect 638910 51781 638970 75107
rect 639188 74104 639508 76327
rect 640738 75791 641058 77374
rect 640738 74915 640777 75791
rect 641013 74915 641058 75791
rect 640738 74104 641058 74915
rect 642288 77215 642608 77374
rect 642288 76339 642323 77215
rect 642559 76339 642608 77215
rect 642288 74104 642608 76339
rect 643838 75817 644158 77374
rect 643838 74941 643879 75817
rect 644115 74941 644158 75817
rect 643838 74104 644158 74941
rect 638907 51780 638973 51781
rect 638907 51716 638908 51780
rect 638972 51716 638973 51780
rect 638907 51715 638973 51716
rect 143324 50672 144738 50688
rect 143324 49956 143343 50672
rect 144699 49956 144738 50672
rect 520227 50556 520293 50557
rect 520227 50492 520228 50556
rect 520292 50492 520293 50556
rect 520227 50491 520293 50492
rect 514707 50284 514773 50285
rect 514707 50220 514708 50284
rect 514772 50220 514773 50284
rect 514707 50219 514773 50220
rect 143324 49936 144738 49956
rect 143860 49638 144040 49936
rect 41874 48222 58536 48364
rect 142560 45396 142740 47256
rect 241680 46621 246056 46692
rect 141776 45394 142866 45396
rect 141376 45354 142866 45394
rect 141376 44158 141448 45354
rect 142804 44158 142866 45354
rect 187555 44980 187621 44981
rect 187555 44916 187556 44980
rect 187620 44916 187621 44980
rect 187555 44915 187621 44916
rect 141376 44130 142866 44158
rect 141923 44028 141989 44029
rect 141923 43964 141924 44028
rect 141988 43964 141989 44028
rect 141923 43963 141989 43964
rect 141926 40357 141986 43963
rect 187558 42125 187618 44915
rect 194363 44844 194429 44845
rect 194363 44780 194364 44844
rect 194428 44780 194429 44844
rect 194363 44779 194429 44780
rect 194366 42125 194426 44779
rect 241680 42837 241731 46621
rect 245995 42837 246056 46621
rect 241680 42784 246056 42837
rect 251302 46635 255700 46684
rect 251302 42851 251383 46635
rect 255647 42851 255700 46635
rect 471651 46476 471717 46477
rect 471651 46412 471652 46476
rect 471716 46412 471717 46476
rect 471651 46411 471717 46412
rect 365115 45252 365181 45253
rect 365115 45188 365116 45252
rect 365180 45188 365181 45252
rect 365115 45187 365181 45188
rect 310099 45116 310165 45117
rect 310099 45052 310100 45116
rect 310164 45052 310165 45116
rect 310099 45051 310165 45052
rect 251302 42788 255700 42851
rect 310102 42397 310162 45051
rect 310099 42396 310165 42397
rect 310099 42332 310100 42396
rect 310164 42332 310165 42396
rect 310099 42331 310165 42332
rect 365118 42125 365178 45187
rect 471654 42125 471714 46411
rect 514710 42125 514770 50219
rect 518571 46612 518637 46613
rect 518571 46548 518572 46612
rect 518636 46548 518637 46612
rect 518571 46547 518637 46548
rect 518574 42397 518634 46547
rect 518571 42396 518637 42397
rect 518571 42332 518572 42396
rect 518636 42332 518637 42396
rect 518571 42331 518637 42332
rect 520230 42125 520290 50491
rect 521699 50420 521765 50421
rect 521699 50356 521700 50420
rect 521764 50356 521765 50420
rect 521699 50355 521765 50356
rect 521702 42125 521762 50355
rect 529795 50284 529861 50285
rect 529795 50220 529796 50284
rect 529860 50220 529861 50284
rect 529795 50219 529861 50220
rect 525931 44708 525997 44709
rect 525931 44644 525932 44708
rect 525996 44644 525997 44708
rect 525931 44643 525997 44644
rect 525934 42125 525994 44643
rect 529798 42125 529858 50219
rect 661270 47274 669426 47320
rect 648104 47170 649670 47188
rect 648104 46614 648129 47170
rect 649645 46614 649670 47170
rect 661270 47038 666442 47274
rect 669398 47038 669426 47274
rect 661270 46991 669426 47038
rect 648104 46590 649670 46614
rect 187555 42124 187621 42125
rect 187555 42060 187556 42124
rect 187620 42060 187621 42124
rect 187555 42059 187621 42060
rect 194363 42124 194429 42125
rect 194363 42060 194364 42124
rect 194428 42060 194429 42124
rect 194363 42059 194429 42060
rect 365115 42124 365181 42125
rect 365115 42060 365116 42124
rect 365180 42060 365181 42124
rect 365115 42059 365181 42060
rect 471651 42124 471717 42125
rect 471651 42060 471652 42124
rect 471716 42060 471717 42124
rect 471651 42059 471717 42060
rect 514707 42124 514773 42125
rect 514707 42060 514708 42124
rect 514772 42060 514773 42124
rect 514707 42059 514773 42060
rect 520227 42124 520293 42125
rect 520227 42060 520228 42124
rect 520292 42060 520293 42124
rect 520227 42059 520293 42060
rect 521699 42124 521765 42125
rect 521699 42060 521700 42124
rect 521764 42060 521765 42124
rect 521699 42059 521765 42060
rect 525931 42124 525997 42125
rect 525931 42060 525932 42124
rect 525996 42060 525997 42124
rect 525931 42059 525997 42060
rect 529795 42124 529861 42125
rect 529795 42060 529796 42124
rect 529860 42060 529861 42124
rect 529795 42059 529861 42060
rect 141923 40356 141989 40357
rect 141923 40292 141924 40356
rect 141988 40292 141989 40356
rect 141923 40291 141989 40292
<< via4 >>
rect 99391 1030771 99787 1031647
rect 102778 1030775 103174 1031651
rect 106148 1030773 106544 1031649
rect 150791 1030771 151187 1031647
rect 154178 1030775 154574 1031651
rect 157548 1030773 157944 1031649
rect 202191 1030771 202587 1031647
rect 205578 1030775 205974 1031651
rect 208948 1030773 209344 1031649
rect 253591 1030771 253987 1031647
rect 256978 1030775 257374 1031651
rect 260348 1030773 260744 1031649
rect 305191 1030771 305587 1031647
rect 308578 1030775 308974 1031651
rect 311948 1030773 312344 1031649
rect 355591 1030771 355987 1031647
rect 358978 1030775 359374 1031651
rect 362348 1030773 362744 1031649
rect 422991 1030771 423387 1031647
rect 426378 1030775 426774 1031651
rect 429748 1030773 430144 1031649
rect 499991 1030771 500387 1031647
rect 503378 1030775 503774 1031651
rect 506748 1030773 507144 1031649
rect 551391 1030771 551787 1031647
rect 554778 1030775 555174 1031651
rect 558148 1030773 558544 1031649
rect 101079 1029577 101475 1030453
rect 104462 1029577 104858 1030453
rect 107838 1029575 108234 1030451
rect 152479 1029577 152875 1030453
rect 155862 1029577 156258 1030453
rect 159238 1029575 159634 1030451
rect 203879 1029577 204275 1030453
rect 207262 1029577 207658 1030453
rect 210638 1029575 211034 1030451
rect 255279 1029577 255675 1030453
rect 258662 1029577 259058 1030453
rect 262038 1029575 262434 1030451
rect 306879 1029577 307275 1030453
rect 310262 1029577 310658 1030453
rect 313638 1029575 314034 1030451
rect 357279 1029577 357675 1030453
rect 360662 1029577 361058 1030453
rect 364038 1029575 364434 1030451
rect 424679 1029577 425075 1030453
rect 428062 1029577 428458 1030453
rect 431438 1029575 431834 1030451
rect 501679 1029577 502075 1030453
rect 505062 1029577 505458 1030453
rect 508438 1029575 508834 1030451
rect 553079 1029577 553475 1030453
rect 556462 1029577 556858 1030453
rect 559838 1029575 560234 1030451
rect 88846 997102 89082 997338
rect 114422 997102 114658 997338
rect 113181 996677 114377 996723
rect 113181 995573 113227 996677
rect 113227 995573 114331 996677
rect 114331 995573 114377 996677
rect 113181 995527 114377 995573
rect 114799 995083 115995 995129
rect 114799 993979 114845 995083
rect 114845 993979 115949 995083
rect 115949 993979 115995 995083
rect 164581 996677 165777 996723
rect 164581 995573 164627 996677
rect 164627 995573 165731 996677
rect 165731 995573 165777 996677
rect 164581 995527 165777 995573
rect 215981 996677 217177 996723
rect 215981 995573 216027 996677
rect 216027 995573 217131 996677
rect 217131 995573 217177 996677
rect 215981 995527 217177 995573
rect 267381 996677 268577 996723
rect 267381 995573 267427 996677
rect 267427 995573 268531 996677
rect 268531 995573 268577 996677
rect 267381 995527 268577 995573
rect 318981 996677 320177 996723
rect 318981 995573 319027 996677
rect 319027 995573 320131 996677
rect 320131 995573 320177 996677
rect 318981 995527 320177 995573
rect 369381 996677 370577 996723
rect 369381 995573 369427 996677
rect 369427 995573 370531 996677
rect 370531 995573 370577 996677
rect 369381 995527 370577 995573
rect 485550 997102 485786 997338
rect 506342 997102 506578 997338
rect 114799 993933 115995 993979
rect 166199 995083 167395 995129
rect 166199 993979 166245 995083
rect 166245 993979 167349 995083
rect 167349 993979 167395 995083
rect 166199 993933 167395 993979
rect 217599 995083 218795 995129
rect 217599 993979 217645 995083
rect 217645 993979 218749 995083
rect 218749 993979 218795 995083
rect 217599 993933 218795 993979
rect 268999 995083 270195 995129
rect 268999 993979 269045 995083
rect 269045 993979 270149 995083
rect 270149 993979 270195 995083
rect 268999 993933 270195 993979
rect 320599 995083 321795 995129
rect 320599 993979 320645 995083
rect 320645 993979 321749 995083
rect 321749 993979 321795 995083
rect 320599 993933 321795 993979
rect 370999 995083 372195 995129
rect 370999 993979 371045 995083
rect 371045 993979 372149 995083
rect 372149 993979 372195 995083
rect 436781 996677 437977 996723
rect 436781 995573 436827 996677
rect 436827 995573 437931 996677
rect 437931 995573 437977 996677
rect 436781 995527 437977 995573
rect 513781 996677 514977 996723
rect 513781 995573 513827 996677
rect 513827 995573 514931 996677
rect 514931 995573 514977 996677
rect 513781 995527 514977 995573
rect 565181 996677 566377 996723
rect 565181 995573 565227 996677
rect 565227 995573 566331 996677
rect 566331 995573 566377 996677
rect 565181 995527 566377 995573
rect 370999 993933 372195 993979
rect 438399 995083 439595 995129
rect 438399 993979 438445 995083
rect 438445 993979 439549 995083
rect 439549 993979 439595 995083
rect 438399 993933 439595 993979
rect 515399 995083 516595 995129
rect 515399 993979 515445 995083
rect 515445 993979 516549 995083
rect 516549 993979 516595 995083
rect 515399 993933 516595 993979
rect 566799 995083 567995 995129
rect 566799 993979 566845 995083
rect 566845 993979 567949 995083
rect 567949 993979 567995 995083
rect 566799 993933 567995 993979
rect 575715 990861 580431 993337
rect 670876 995588 676552 996624
rect 585711 990875 590427 993351
rect 670962 990364 673278 992520
rect 47794 989729 49790 990285
rect 55829 989730 56385 990286
rect 50200 988765 52196 989321
rect 55833 988770 56389 989326
rect 658417 986846 663133 987402
rect 667281 986851 669757 987407
rect 52599 983961 53795 984517
rect 55811 983961 56367 984517
rect 7267 941839 8143 942235
rect 6064 940147 6940 940543
rect 7268 938459 8144 938855
rect 6070 936781 6946 937177
rect 54189 949949 55385 949995
rect 54189 948845 54235 949949
rect 54235 948845 55339 949949
rect 55339 948845 55385 949949
rect 54189 948799 55385 948845
rect 52595 948331 53791 948377
rect 52595 947227 52641 948331
rect 52641 947227 53745 948331
rect 53745 947227 53791 948331
rect 52595 947181 53791 947227
rect 7265 935079 8141 935475
rect 6071 933391 6947 933787
rect 47883 842334 49719 842340
rect 47883 837790 47909 842334
rect 47909 837790 49693 842334
rect 49693 837790 49719 842334
rect 47883 837784 49719 837790
rect 47883 832402 49719 832408
rect 47883 827858 47909 832402
rect 47909 827858 49693 832402
rect 49693 827858 49719 832402
rect 47883 827852 49719 827858
rect 667270 828640 667276 833196
rect 667276 828640 669740 833196
rect 669740 828640 669746 833196
rect 54189 824149 55385 824195
rect 54189 823045 54235 824149
rect 54235 823045 55339 824149
rect 55339 823045 55385 824149
rect 54189 822999 55385 823045
rect 52595 822531 53791 822577
rect 52595 821427 52641 822531
rect 52641 821427 53745 822531
rect 53745 821427 53791 822531
rect 52595 821381 53791 821427
rect 667256 818646 667262 823202
rect 667262 818646 669726 823202
rect 669726 818646 669732 823202
rect 7267 816039 8143 816435
rect 6064 814347 6940 814743
rect 7268 812659 8144 813055
rect 6070 810981 6946 811377
rect 7265 809279 8141 809675
rect 6071 807591 6947 807987
rect 7267 772839 8143 773235
rect 6064 771147 6940 771543
rect 54189 780949 55385 780995
rect 54189 779845 54235 780949
rect 54235 779845 55339 780949
rect 55339 779845 55385 780949
rect 54189 779799 55385 779845
rect 52595 779331 53791 779377
rect 52595 778227 52641 779331
rect 52641 778227 53745 779331
rect 53745 778227 53791 779331
rect 52595 778181 53791 778227
rect 7268 769459 8144 769855
rect 6070 767781 6946 768177
rect 7265 766079 8141 766475
rect 6071 764391 6947 764787
rect 7267 729639 8143 730035
rect 6064 727947 6940 728343
rect 54189 737749 55385 737795
rect 54189 736645 54235 737749
rect 54235 736645 55339 737749
rect 55339 736645 55385 737749
rect 54189 736599 55385 736645
rect 52595 736131 53791 736177
rect 52595 735027 52641 736131
rect 52641 735027 53745 736131
rect 53745 735027 53791 736131
rect 52595 734981 53791 735027
rect 7268 726259 8144 726655
rect 6070 724581 6946 724977
rect 7265 722879 8141 723275
rect 6071 721191 6947 721587
rect 7267 686439 8143 686835
rect 6064 684747 6940 685143
rect 54189 694549 55385 694595
rect 54189 693445 54235 694549
rect 54235 693445 55339 694549
rect 55339 693445 55385 694549
rect 54189 693399 55385 693445
rect 52595 692931 53791 692977
rect 52595 691827 52641 692931
rect 52641 691827 53745 692931
rect 53745 691827 53791 692931
rect 52595 691781 53791 691827
rect 7268 683059 8144 683455
rect 6070 681381 6946 681777
rect 7265 679679 8141 680075
rect 6071 677991 6947 678387
rect 7267 643239 8143 643635
rect 6064 641547 6940 641943
rect 54189 651349 55385 651395
rect 54189 650245 54235 651349
rect 54235 650245 55339 651349
rect 55339 650245 55385 651349
rect 54189 650199 55385 650245
rect 52595 649731 53791 649777
rect 52595 648627 52641 649731
rect 52641 648627 53745 649731
rect 53745 648627 53791 649731
rect 52595 648581 53791 648627
rect 7268 639859 8144 640255
rect 6070 638181 6946 638577
rect 7265 636479 8141 636875
rect 6071 634791 6947 635187
rect 7267 600039 8143 600435
rect 6064 598347 6940 598743
rect 54189 608149 55385 608195
rect 54189 607045 54235 608149
rect 54235 607045 55339 608149
rect 55339 607045 55385 608149
rect 54189 606999 55385 607045
rect 52595 606531 53791 606577
rect 52595 605427 52641 606531
rect 52641 605427 53745 606531
rect 53745 605427 53791 606531
rect 52595 605381 53791 605427
rect 7268 596659 8144 597055
rect 6070 594981 6946 595377
rect 7265 593279 8141 593675
rect 6071 591591 6947 591987
rect 7267 556839 8143 557235
rect 6064 555147 6940 555543
rect 54189 564949 55385 564995
rect 54189 563845 54235 564949
rect 54235 563845 55339 564949
rect 55339 563845 55385 564949
rect 54189 563799 55385 563845
rect 52595 563331 53791 563377
rect 52595 562227 52641 563331
rect 52641 562227 53745 563331
rect 53745 562227 53791 563331
rect 52595 562181 53791 562227
rect 7268 553459 8144 553855
rect 6070 551781 6946 552177
rect 7265 550079 8141 550475
rect 6071 548391 6947 548787
rect 667283 518591 669759 518597
rect 667283 514047 667329 518591
rect 667329 514047 669713 518591
rect 669713 514047 669759 518591
rect 667283 514041 669759 514047
rect 667297 508601 669773 508607
rect 667297 504057 667343 508601
rect 667343 504057 669727 508601
rect 669727 504057 669773 508601
rect 667297 504051 669773 504057
rect 50310 497743 52146 497769
rect 50310 493239 50356 497743
rect 50356 493239 52100 497743
rect 52100 493239 52146 497743
rect 50310 493213 52146 493239
rect 50298 487753 52134 487779
rect 50298 483249 50344 487753
rect 50344 483249 52088 487753
rect 52088 483249 52134 487753
rect 50298 483223 52134 483249
rect 54189 437349 55385 437395
rect 54189 436245 54235 437349
rect 54235 436245 55339 437349
rect 55339 436245 55385 437349
rect 54189 436199 55385 436245
rect 52595 435731 53791 435777
rect 52595 434627 52641 435731
rect 52641 434627 53745 435731
rect 53745 434627 53791 435731
rect 52595 434581 53791 434627
rect 7267 429239 8143 429635
rect 6064 427547 6940 427943
rect 7268 425859 8144 426255
rect 6070 424181 6946 424577
rect 7265 422479 8141 422875
rect 6071 420791 6947 421187
rect 664099 430389 666575 430395
rect 664099 425685 664125 430389
rect 664125 425685 666549 430389
rect 666549 425685 666575 430389
rect 664099 425679 666575 425685
rect 664082 420471 666558 420517
rect 664082 415847 664108 420471
rect 664108 415847 666532 420471
rect 666532 415847 666558 420471
rect 664082 415801 666558 415847
rect 54189 394149 55385 394195
rect 54189 393045 54235 394149
rect 54235 393045 55339 394149
rect 55339 393045 55385 394149
rect 54189 392999 55385 393045
rect 52595 392531 53791 392577
rect 52595 391427 52641 392531
rect 52641 391427 53745 392531
rect 53745 391427 53791 392531
rect 52595 391381 53791 391427
rect 7267 386039 8143 386435
rect 6064 384347 6940 384743
rect 7268 382659 8144 383055
rect 6070 380981 6946 381377
rect 7265 379279 8141 379675
rect 6071 377591 6947 377987
rect 54189 350949 55385 350995
rect 54189 349845 54235 350949
rect 54235 349845 55339 350949
rect 55339 349845 55385 350949
rect 54189 349799 55385 349845
rect 52595 349331 53791 349377
rect 52595 348227 52641 349331
rect 52641 348227 53745 349331
rect 53745 348227 53791 349331
rect 52595 348181 53791 348227
rect 7267 342839 8143 343235
rect 6064 341147 6940 341543
rect 7268 339459 8144 339855
rect 6070 337781 6946 338177
rect 7265 336079 8141 336475
rect 6071 334391 6947 334787
rect 54189 307749 55385 307795
rect 54189 306645 54235 307749
rect 54235 306645 55339 307749
rect 55339 306645 55385 307749
rect 54189 306599 55385 306645
rect 52595 306131 53791 306177
rect 52595 305027 52641 306131
rect 52641 305027 53745 306131
rect 53745 305027 53791 306131
rect 52595 304981 53791 305027
rect 7267 299639 8143 300035
rect 6064 297947 6940 298343
rect 7268 296259 8144 296655
rect 6070 294581 6946 294977
rect 7265 292879 8141 293275
rect 6071 291191 6947 291587
rect 52593 276850 53789 278046
rect 55806 276859 56362 277415
rect 50193 272056 52189 273412
rect 55802 272057 56358 272613
rect 47799 270303 49795 271659
rect 55776 271094 56492 271650
rect 54189 264549 55385 264595
rect 54189 263445 54235 264549
rect 54235 263445 55339 264549
rect 55339 263445 55385 264549
rect 54189 263399 55385 263445
rect 52595 262931 53791 262977
rect 52595 261827 52641 262931
rect 52641 261827 53745 262931
rect 53745 261827 53791 262931
rect 52595 261781 53791 261827
rect 58529 266488 59085 269444
rect 47991 258689 49667 261325
rect 56555 258628 59351 261264
rect 62737 262484 63293 265440
rect 7267 256439 8143 256835
rect 6064 254747 6940 255143
rect 50391 254689 52067 257325
rect 56564 254628 60320 257264
rect 60820 254486 61376 257442
rect 7268 253059 8144 253455
rect 6070 251381 6946 251777
rect 7265 249679 8141 250075
rect 6071 247991 6947 248387
rect 52602 250492 53798 253448
rect 56152 250494 63268 253450
rect 41060 238317 43536 245433
rect 56391 242545 63347 245341
rect 63703 242494 64259 245450
rect 65615 250482 66171 253438
rect 393481 266565 394197 269361
rect 408507 262892 409223 265368
rect 394597 258553 395313 261349
rect 409735 254570 410771 257366
rect 211801 250580 212517 253376
rect 241901 250580 242617 253376
rect 272228 250580 272624 253376
rect 302160 250580 302716 253376
rect 332201 250580 332917 253376
rect 362301 250580 363017 253376
rect 392517 250580 393073 253376
rect 66579 246494 67135 249450
rect 196785 246571 197501 249367
rect 226885 246571 227601 249367
rect 256985 246571 257701 249367
rect 287129 246769 287685 249405
rect 317300 246541 317856 249337
rect 347285 246571 348001 249367
rect 377285 246571 378001 249367
rect 407285 246571 408001 249367
rect 651614 250481 652170 253437
rect 650648 246499 651204 249455
rect 212605 242495 213481 245451
rect 242705 242495 243581 245451
rect 272950 242495 273346 245451
rect 303116 242495 303512 245451
rect 333005 242495 333881 245451
rect 363105 242495 363981 245451
rect 393227 242495 393783 245451
rect 44248 234547 46724 241343
rect 56406 238579 63362 241375
rect 64653 238490 65209 241446
rect 197619 238490 198335 241446
rect 227719 238490 228435 241446
rect 257819 238490 258535 241446
rect 288039 238490 288595 241446
rect 318202 238490 318598 241446
rect 348119 238490 348835 241446
rect 659025 273969 663101 274525
rect 667288 273176 669764 274532
rect 655447 266485 656003 269441
rect 654489 262483 655045 265439
rect 657363 258497 657919 261453
rect 656401 254479 656957 257435
rect 667032 246657 669668 249293
rect 674146 246558 676462 249354
rect 653519 242497 654075 245453
rect 378119 238490 378835 241446
rect 408374 238490 408770 241446
rect 652561 238495 653117 241451
rect 47931 234579 50727 237375
rect 56375 234585 63171 237381
rect 210902 234485 211778 237441
rect 241002 234485 241878 237441
rect 271355 234485 271911 237441
rect 301490 234517 302046 237313
rect 331410 234485 332126 237441
rect 361402 234485 362278 237441
rect 391830 234485 392226 237441
rect 56394 230575 63030 233371
rect 89903 231370 93979 232086
rect 169887 231392 173963 232108
rect 196029 230486 196585 233442
rect 226129 230486 226685 233442
rect 256229 230486 256785 233442
rect 286329 230486 286885 233442
rect 316429 230486 316985 233442
rect 346529 230486 347085 233442
rect 376529 230486 377085 233442
rect 406660 230486 407056 233442
rect 429905 231404 433981 232120
rect 7267 213239 8143 213635
rect 6064 211547 6940 211943
rect 7268 209859 8144 210255
rect 6070 208181 6946 208577
rect 7265 206479 8141 206875
rect 6071 204791 6947 205187
rect 54189 221349 55385 221395
rect 54189 220245 54235 221349
rect 54235 220245 55339 221349
rect 55339 220245 55385 221349
rect 54189 220199 55385 220245
rect 52595 219731 53791 219777
rect 52595 218627 52641 219731
rect 52641 218627 53745 219731
rect 53745 218627 53791 219731
rect 52595 218581 53791 218627
rect 598610 209715 601086 212351
rect 607464 209715 609940 212351
rect 641143 209598 642019 212394
rect 596320 207906 597676 208462
rect 602413 207906 605369 208462
rect 51413 196916 52289 197472
rect 598703 197085 601019 197801
rect 605958 197247 606994 197483
rect 596124 183894 596840 184450
rect 602413 183890 605369 184446
rect 42007 173229 45603 176665
rect 42777 170898 45733 171454
rect 51305 170902 52181 171458
rect 598703 166445 601019 167161
rect 605941 166619 606977 166855
rect 594082 157898 596878 158454
rect 602387 157902 605343 158458
rect 42791 144904 45747 145460
rect 51239 144894 52115 145450
rect 598703 135805 601019 136521
rect 605931 135979 606967 136215
rect 594092 131892 596888 132448
rect 602413 131886 605369 132442
rect 42781 118900 45737 119456
rect 51235 118900 52111 119456
rect 594094 105898 596890 106454
rect 602417 105898 605373 106454
rect 598703 104885 601019 105601
rect 605943 105342 606979 105578
rect 625552 96047 626748 98683
rect 636179 96525 636895 98681
rect 634590 94062 634826 94298
rect 42777 92898 45733 93454
rect 51239 92896 52115 93452
rect 41931 82706 45687 82752
rect 41931 78242 41937 82706
rect 41937 78242 45681 82706
rect 45681 78242 45687 82706
rect 41931 78196 45687 78242
rect 594088 79908 596884 80464
rect 602411 79910 605367 80466
rect 632174 78313 632890 80789
rect 656363 96109 657559 98745
rect 641582 94062 641818 94298
rect 640152 78260 640868 80896
rect 629919 76317 630155 77193
rect 631471 74915 631707 75791
rect 633031 76331 633267 77207
rect 634565 74919 634801 75795
rect 636121 76327 636357 77203
rect 637673 74923 637909 75799
rect 639215 76327 639451 77203
rect 41907 72802 45663 72848
rect 41907 68338 41913 72802
rect 41913 68338 45657 72802
rect 45657 68338 45663 72802
rect 41907 68292 45663 68338
rect 41935 66892 45691 67448
rect 51437 66898 52313 67454
rect 42000 48398 45596 51994
rect 54490 48364 58246 51960
rect 640777 74915 641013 75791
rect 642323 76339 642559 77215
rect 643879 74941 644115 75817
rect 143343 49956 144699 50672
rect 141448 44158 142804 45354
rect 241745 42851 245981 46607
rect 251397 42865 255633 46621
rect 648129 47124 649645 47170
rect 648129 46660 648155 47124
rect 648155 46660 649619 47124
rect 649619 46660 649645 47124
rect 648129 46614 649645 46660
rect 666442 47038 669398 47274
<< metal5 >>
rect 102802 1031651 103148 1031678
rect 78440 1018512 90960 1031002
rect 106166 1031649 106512 1031674
rect 154202 1031651 154548 1031678
rect 99428 1029104 99748 1030771
rect 101118 1029104 101438 1029577
rect 102808 1029136 103128 1030775
rect 104480 1030453 104826 1030464
rect 104498 1029136 104818 1029577
rect 106188 1029136 106508 1030773
rect 107868 1030451 108214 1030470
rect 107878 1029136 108198 1029575
rect 129840 1018512 142360 1031002
rect 157566 1031649 157912 1031674
rect 205602 1031651 205948 1031678
rect 150828 1029104 151148 1030771
rect 152518 1029104 152838 1029577
rect 154208 1029136 154528 1030775
rect 155880 1030453 156226 1030464
rect 155898 1029136 156218 1029577
rect 157588 1029136 157908 1030773
rect 159268 1030451 159614 1030470
rect 159278 1029136 159598 1029575
rect 181240 1018512 193760 1031002
rect 208966 1031649 209312 1031674
rect 257002 1031651 257348 1031678
rect 202228 1029104 202548 1030771
rect 203918 1029104 204238 1029577
rect 205608 1029136 205928 1030775
rect 207280 1030453 207626 1030464
rect 207298 1029136 207618 1029577
rect 208988 1029136 209308 1030773
rect 210668 1030451 211014 1030470
rect 210678 1029136 210998 1029575
rect 232640 1018512 245160 1031002
rect 260366 1031649 260712 1031674
rect 308602 1031651 308948 1031678
rect 253628 1029104 253948 1030771
rect 255318 1029104 255638 1029577
rect 257008 1029136 257328 1030775
rect 258680 1030453 259026 1030464
rect 258698 1029136 259018 1029577
rect 260388 1029136 260708 1030773
rect 262068 1030451 262414 1030470
rect 262078 1029136 262398 1029575
rect 284240 1018512 296760 1031002
rect 311966 1031649 312312 1031674
rect 359002 1031651 359348 1031678
rect 305228 1029104 305548 1030771
rect 306918 1029104 307238 1029577
rect 308608 1029136 308928 1030775
rect 310280 1030453 310626 1030464
rect 310298 1029136 310618 1029577
rect 311988 1029136 312308 1030773
rect 313668 1030451 314014 1030470
rect 313678 1029136 313998 1029575
rect 334810 1018624 346978 1030789
rect 362366 1031649 362712 1031674
rect 426402 1031651 426748 1031678
rect 355628 1029104 355948 1030771
rect 357318 1029104 357638 1029577
rect 359008 1029136 359328 1030775
rect 360680 1030453 361026 1030464
rect 360698 1029136 361018 1029577
rect 362388 1029136 362708 1030773
rect 364068 1030451 364414 1030470
rect 364078 1029136 364398 1029575
rect 386040 1018512 398560 1031002
rect 429766 1031649 430112 1031674
rect 503402 1031651 503748 1031678
rect 423028 1029104 423348 1030771
rect 424718 1029104 425038 1029577
rect 426408 1029136 426728 1030775
rect 428080 1030453 428426 1030464
rect 428098 1029136 428418 1029577
rect 429788 1029136 430108 1030773
rect 431468 1030451 431814 1030470
rect 431478 1029136 431798 1029575
rect 475040 1018512 487560 1031002
rect 506766 1031649 507112 1031674
rect 554802 1031651 555148 1031678
rect 500028 1029104 500348 1030771
rect 501718 1029104 502038 1029577
rect 503408 1029136 503728 1030775
rect 505080 1030453 505426 1030464
rect 505098 1029136 505418 1029577
rect 506788 1029136 507108 1030773
rect 508468 1030451 508814 1030470
rect 508478 1029136 508798 1029575
rect 526440 1018512 538960 1031002
rect 558166 1031649 558512 1031674
rect 551428 1029104 551748 1030771
rect 553118 1029104 553438 1029577
rect 554808 1029136 555128 1030775
rect 556480 1030453 556826 1030464
rect 556498 1029136 556818 1029577
rect 558188 1029136 558508 1030773
rect 559868 1030451 560214 1030470
rect 559878 1029136 560198 1029575
rect 577010 1018624 589178 1030789
rect 628240 1018512 640760 1031002
rect 88804 997338 114700 997380
rect 88804 997102 88846 997338
rect 89082 997102 114422 997338
rect 114658 997102 114700 997338
rect 88804 997060 114700 997102
rect 485508 997338 506620 997380
rect 485508 997102 485550 997338
rect 485786 997102 506342 997338
rect 506578 997102 506620 997338
rect 485508 997060 506620 997102
rect 52598 995527 113181 996702
rect 114377 995527 164581 996702
rect 165777 995527 215981 996702
rect 217177 995527 267381 996702
rect 268577 995527 318981 996702
rect 320177 995527 369381 996702
rect 370577 995527 436781 996702
rect 437977 995527 513781 996702
rect 514977 995527 565181 996702
rect 566377 996624 676660 996702
rect 566377 995588 670876 996624
rect 676552 995588 676660 996624
rect 566377 995527 676660 995588
rect 52598 995502 676660 995527
rect 47798 990285 49798 990466
rect 49790 989729 49798 990285
rect 6598 956440 19088 968960
rect 7260 941878 7267 942198
rect 8143 941878 8582 942198
rect 6048 940188 6064 940508
rect 6940 940188 8582 940508
rect 7266 938498 7268 938818
rect 8144 938498 8582 938818
rect 6034 936806 6070 937154
rect 6946 936808 8582 937128
rect 8141 935438 8172 935453
rect 8141 935118 8614 935438
rect 8141 935102 8172 935118
rect 6947 933748 6980 933770
rect 6947 933428 8614 933748
rect 6947 933408 6980 933428
rect 6167 914054 19620 924934
rect 6811 871210 18976 883378
rect 47798 842340 49798 989729
rect 6811 829010 18976 841178
rect 47798 837784 47883 842340
rect 49719 837784 49798 842340
rect 47798 832408 49798 837784
rect 47798 827852 47883 832408
rect 49719 827852 49798 832408
rect 7260 816078 7267 816398
rect 8143 816078 8582 816398
rect 6048 814388 6064 814708
rect 6940 814388 8582 814708
rect 7266 812698 7268 813018
rect 8144 812698 8582 813018
rect 6034 811006 6070 811354
rect 6946 811008 8582 811328
rect 8141 809638 8172 809653
rect 8141 809318 8614 809638
rect 8141 809302 8172 809318
rect 6947 807948 6980 807970
rect 6947 807628 8614 807948
rect 6947 807608 6980 807628
rect 6598 786640 19088 799160
rect 7260 772878 7267 773198
rect 8143 772878 8582 773198
rect 6048 771188 6064 771508
rect 6940 771188 8582 771508
rect 7266 769498 7268 769818
rect 8144 769498 8582 769818
rect 6034 767806 6070 768154
rect 6946 767808 8582 768128
rect 8141 766438 8172 766453
rect 8141 766118 8614 766438
rect 8141 766102 8172 766118
rect 6947 764748 6980 764770
rect 6947 764428 8614 764748
rect 6947 764408 6980 764428
rect 6598 743440 19088 755960
rect 7260 729678 7267 729998
rect 8143 729678 8582 729998
rect 6048 727988 6064 728308
rect 6940 727988 8582 728308
rect 7266 726298 7268 726618
rect 8144 726298 8582 726618
rect 6034 724606 6070 724954
rect 6946 724608 8582 724928
rect 8141 723238 8172 723253
rect 8141 722918 8614 723238
rect 8141 722902 8172 722918
rect 6947 721548 6980 721570
rect 6947 721228 8614 721548
rect 6947 721208 6980 721228
rect 6598 700240 19088 712760
rect 7260 686478 7267 686798
rect 8143 686478 8582 686798
rect 6048 684788 6064 685108
rect 6940 684788 8582 685108
rect 7266 683098 7268 683418
rect 8144 683098 8582 683418
rect 6034 681406 6070 681754
rect 6946 681408 8582 681728
rect 8141 680038 8172 680053
rect 8141 679718 8614 680038
rect 8141 679702 8172 679718
rect 6947 678348 6980 678370
rect 6947 678028 8614 678348
rect 6947 678008 6980 678028
rect 6598 657040 19088 669560
rect 7260 643278 7267 643598
rect 8143 643278 8582 643598
rect 6048 641588 6064 641908
rect 6940 641588 8582 641908
rect 7266 639898 7268 640218
rect 8144 639898 8582 640218
rect 6034 638206 6070 638554
rect 6946 638208 8582 638528
rect 8141 636838 8172 636853
rect 8141 636518 8614 636838
rect 8141 636502 8172 636518
rect 6947 635148 6980 635170
rect 6947 634828 8614 635148
rect 6947 634808 6980 634828
rect 6598 613840 19088 626360
rect 7260 600078 7267 600398
rect 8143 600078 8582 600398
rect 6048 598388 6064 598708
rect 6940 598388 8582 598708
rect 7266 596698 7268 597018
rect 8144 596698 8582 597018
rect 6034 595006 6070 595354
rect 6946 595008 8582 595328
rect 8141 593638 8172 593653
rect 8141 593318 8614 593638
rect 8141 593302 8172 593318
rect 6947 591948 6980 591970
rect 6947 591628 8614 591948
rect 6947 591608 6980 591628
rect 6598 570640 19088 583160
rect 7260 556878 7267 557198
rect 8143 556878 8582 557198
rect 6048 555188 6064 555508
rect 6940 555188 8582 555508
rect 7266 553498 7268 553818
rect 8144 553498 8582 553818
rect 6034 551806 6070 552154
rect 6946 551808 8582 552128
rect 8141 550438 8172 550453
rect 8141 550118 8614 550438
rect 8141 550102 8172 550118
rect 6947 548748 6980 548770
rect 6947 548428 8614 548748
rect 6947 548408 6980 548428
rect 6598 527440 19088 539960
rect 6811 484410 18976 496578
rect 6167 442854 19620 453734
rect 7260 429278 7267 429598
rect 8143 429278 8582 429598
rect 6048 427588 6064 427908
rect 6940 427588 8582 427908
rect 7266 425898 7268 426218
rect 8144 425898 8582 426218
rect 6034 424206 6070 424554
rect 6946 424208 8582 424528
rect 8141 422838 8172 422853
rect 8141 422518 8614 422838
rect 8141 422502 8172 422518
rect 6947 421148 6980 421170
rect 6947 420828 8614 421148
rect 6947 420808 6980 420828
rect 6598 399840 19088 412360
rect 7260 386078 7267 386398
rect 8143 386078 8582 386398
rect 6048 384388 6064 384708
rect 6940 384388 8582 384708
rect 7266 382698 7268 383018
rect 8144 382698 8582 383018
rect 6034 381006 6070 381354
rect 6946 381008 8582 381328
rect 8141 379638 8172 379653
rect 8141 379318 8614 379638
rect 8141 379302 8172 379318
rect 6947 377948 6980 377970
rect 6947 377628 8614 377948
rect 6947 377608 6980 377628
rect 6598 356640 19088 369160
rect 7260 342878 7267 343198
rect 8143 342878 8582 343198
rect 6048 341188 6064 341508
rect 6940 341188 8582 341508
rect 7266 339498 7268 339818
rect 8144 339498 8582 339818
rect 6034 337806 6070 338154
rect 6946 337808 8582 338128
rect 8141 336438 8172 336453
rect 8141 336118 8614 336438
rect 8141 336102 8172 336118
rect 6947 334748 6980 334770
rect 6947 334428 8614 334748
rect 6947 334408 6980 334428
rect 6598 313440 19088 325960
rect 7260 299678 7267 299998
rect 8143 299678 8582 299998
rect 6048 297988 6064 298308
rect 6940 297988 8582 298308
rect 7266 296298 7268 296618
rect 8144 296298 8582 296618
rect 6034 294606 6070 294954
rect 6946 294608 8582 294928
rect 8141 293238 8172 293253
rect 8141 292918 8614 293238
rect 8141 292902 8172 292918
rect 6947 291548 6980 291570
rect 6947 291228 8614 291548
rect 6947 291208 6980 291228
rect 6598 270240 19088 282760
rect 47798 271659 49798 827852
rect 50198 989321 52198 990466
rect 50198 988765 50200 989321
rect 52196 988765 52198 989321
rect 50198 497769 52198 988765
rect 52598 984517 53798 995502
rect 52598 983961 52599 984517
rect 53795 983961 53798 984517
rect 52598 948377 53798 983961
rect 54198 993933 114799 995102
rect 115995 993933 166199 995102
rect 167395 993933 217599 995102
rect 218795 993933 268999 995102
rect 270195 993933 320599 995102
rect 321795 993933 370999 995102
rect 372195 993933 438399 995102
rect 439595 993933 515399 995102
rect 516595 993933 566799 995102
rect 567995 993933 676620 995102
rect 54198 993902 676620 993933
rect 54198 983588 55398 993902
rect 575640 993351 666620 993396
rect 575640 993337 585711 993351
rect 575640 990861 575715 993337
rect 580431 990875 585711 993337
rect 590427 990875 666620 993351
rect 674020 992696 676620 993902
rect 670976 992520 673264 992530
rect 580431 990861 666620 990875
rect 575640 990796 666620 990861
rect 55776 990286 56596 990308
rect 55776 989730 55829 990286
rect 56385 989730 56596 990286
rect 55776 989688 56596 989730
rect 55776 989326 57552 989348
rect 55776 988770 55833 989326
rect 56389 988770 57552 989326
rect 55776 988728 57552 988770
rect 664020 988388 666620 990796
rect 670976 990354 673264 990364
rect 656038 987768 666620 988388
rect 655078 987402 663178 987428
rect 655078 986846 658417 987402
rect 663133 986846 663178 987402
rect 655078 986808 663178 986846
rect 55776 984517 62358 984548
rect 55776 983961 55811 984517
rect 56367 983961 62358 984517
rect 55776 983928 62358 983961
rect 54198 982968 63316 983588
rect 54198 949995 55398 982968
rect 55385 948799 55398 949995
rect 53791 947181 53798 948377
rect 52598 822577 53798 947181
rect 54198 824195 55398 948799
rect 55385 822999 55398 824195
rect 53791 821381 53798 822577
rect 52598 779377 53798 821381
rect 54198 780995 55398 822999
rect 55385 779799 55398 780995
rect 53791 778181 53798 779377
rect 52598 736177 53798 778181
rect 54198 737795 55398 779799
rect 55385 736599 55398 737795
rect 53791 734981 53798 736177
rect 52598 692977 53798 734981
rect 54198 694595 55398 736599
rect 55385 693399 55398 694595
rect 53791 691781 53798 692977
rect 52598 649777 53798 691781
rect 54198 651395 55398 693399
rect 55385 650199 55398 651395
rect 53791 648581 53798 649777
rect 52598 606577 53798 648581
rect 54198 608195 55398 650199
rect 55385 606999 55398 608195
rect 53791 605381 53798 606577
rect 52598 563377 53798 605381
rect 54198 564995 55398 606999
rect 55385 563799 55398 564995
rect 53791 562181 53798 563377
rect 50198 493213 50310 497769
rect 52146 493213 52198 497769
rect 50198 487779 52198 493213
rect 50198 483223 50298 487779
rect 52134 483223 52198 487779
rect 50198 273412 52198 483223
rect 52598 435777 53798 562181
rect 54198 437395 55398 563799
rect 55385 436199 55398 437395
rect 53791 434581 53798 435777
rect 52598 392577 53798 434581
rect 54198 394195 55398 436199
rect 55385 392999 55398 394195
rect 53791 391381 53798 392577
rect 52598 349377 53798 391381
rect 54198 350995 55398 392999
rect 55385 349799 55398 350995
rect 53791 348181 53798 349377
rect 52598 306177 53798 348181
rect 54198 307795 55398 349799
rect 55385 306599 55398 307795
rect 53791 304981 53798 306177
rect 52598 278046 53798 304981
rect 53789 276850 53798 278046
rect 52189 272056 52198 273412
rect 47798 270303 47799 271659
rect 49795 270303 49798 271659
rect 47798 261325 49798 270303
rect 47798 258689 47991 261325
rect 49667 258689 49798 261325
rect 47798 258484 49798 258689
rect 50198 257325 52198 272056
rect 52598 262977 53798 276850
rect 54198 278404 55398 306599
rect 664020 430395 666620 987768
rect 664020 425679 664099 430395
rect 666575 425679 666620 430395
rect 664020 420517 666620 425679
rect 664020 415801 664082 420517
rect 666558 415801 666620 420517
rect 54198 277784 63312 278404
rect 54198 264595 55398 277784
rect 55754 277415 62352 277444
rect 55754 276859 55806 277415
rect 56362 276859 62352 277415
rect 55754 276824 62352 276859
rect 655060 274525 663158 274564
rect 655060 273969 659025 274525
rect 663101 273969 663158 274525
rect 655060 273944 663158 273969
rect 664020 273604 666620 415801
rect 656026 272984 666620 273604
rect 55754 272613 57546 272644
rect 55754 272057 55802 272613
rect 56358 272057 57546 272613
rect 55754 272024 57546 272057
rect 55754 271650 56590 271684
rect 55754 271094 55776 271650
rect 56492 271094 56590 271650
rect 55754 271064 56590 271094
rect 664020 269466 666620 272984
rect 58388 269444 666620 269466
rect 58388 266488 58529 269444
rect 59085 269441 666620 269444
rect 59085 269361 655447 269441
rect 59085 266565 393481 269361
rect 394197 266565 655447 269361
rect 59085 266488 655447 266565
rect 58388 266485 655447 266488
rect 656003 266485 666620 269441
rect 58388 266466 666620 266485
rect 667220 987407 669820 987566
rect 667220 986851 667281 987407
rect 669757 986851 669820 987407
rect 667220 833196 669820 986851
rect 698512 952840 711002 965360
rect 697980 909666 711433 920546
rect 698512 863640 711002 876160
rect 667220 828640 667270 833196
rect 669746 828640 669820 833196
rect 667220 823202 669820 828640
rect 667220 818646 667256 823202
rect 669732 818646 669820 823202
rect 698624 819822 710789 831990
rect 667220 518597 669820 818646
rect 698512 774440 711002 786960
rect 698512 729440 711002 741960
rect 698512 684440 711002 696960
rect 698512 639240 711002 651760
rect 698512 594240 711002 606760
rect 698512 549040 711002 561560
rect 667220 514041 667283 518597
rect 669759 514041 669820 518597
rect 667220 508607 669820 514041
rect 667220 504051 667297 508607
rect 669773 504051 669820 508607
rect 698624 505222 710789 517390
rect 667220 274532 669820 504051
rect 697980 461866 711433 472746
rect 698624 417022 710789 429190
rect 698512 371840 711002 384360
rect 698512 326640 711002 339160
rect 698512 281640 711002 294160
rect 667220 273176 667288 274532
rect 669764 273176 669820 274532
rect 667220 265466 669820 273176
rect 55385 263399 55398 264595
rect 53791 261781 53798 262977
rect 7260 256478 7267 256798
rect 8143 256478 8582 256798
rect 6048 254788 6064 255108
rect 6940 254788 8582 255108
rect 50198 254689 50391 257325
rect 52067 254689 52198 257325
rect 50198 254498 52198 254689
rect 7266 253098 7268 253418
rect 52598 253448 53798 261781
rect 8144 253098 8582 253418
rect 6034 251406 6070 251754
rect 6946 251408 8582 251728
rect 52598 250492 52602 253448
rect 8141 250038 8172 250053
rect 8141 249718 8614 250038
rect 8141 249702 8172 249718
rect 6947 248348 6980 248370
rect 6947 248028 8614 248348
rect 6947 248008 6980 248028
rect 6598 227040 19088 239560
rect 44254 241343 46718 241358
rect 47836 237375 50836 237612
rect 47836 234579 47931 237375
rect 50727 234579 50836 237375
rect 44254 234532 46718 234547
rect 7260 213278 7267 213598
rect 8143 213278 8582 213598
rect 6048 211588 6064 211908
rect 6940 211588 8582 211908
rect 47836 210498 50836 234579
rect 52598 219777 53798 250492
rect 54198 249466 55398 263399
rect 62534 265440 669820 265466
rect 62534 262484 62737 265440
rect 63293 265439 669820 265440
rect 63293 265368 654489 265439
rect 63293 262892 408507 265368
rect 409223 262892 654489 265368
rect 63293 262484 654489 262892
rect 62534 262483 654489 262484
rect 655045 262483 669820 265439
rect 62534 262466 669820 262483
rect 56370 261453 658090 261466
rect 56370 261349 657363 261453
rect 56370 261264 394597 261349
rect 56370 258628 56555 261264
rect 59351 258628 394597 261264
rect 56370 258553 394597 258628
rect 395313 258553 657363 261349
rect 56370 258497 657363 258553
rect 657919 258497 658090 261453
rect 56370 258466 658090 258497
rect 56370 257442 657076 257466
rect 56370 257264 60820 257442
rect 56370 254628 56564 257264
rect 60320 254628 60820 257264
rect 56370 254486 60820 254628
rect 61376 257435 657076 257442
rect 61376 257366 656401 257435
rect 61376 254570 409735 257366
rect 410771 254570 656401 257366
rect 61376 254486 656401 254570
rect 56370 254479 656401 254486
rect 656957 254479 657076 257435
rect 56370 254466 657076 254479
rect 56126 253450 670986 253466
rect 56126 250494 56152 253450
rect 63268 253438 670986 253450
rect 63268 250494 65615 253438
rect 56126 250482 65615 250494
rect 66171 253437 670986 253438
rect 66171 253376 651614 253437
rect 66171 250580 211801 253376
rect 212517 250580 241901 253376
rect 242617 250580 272228 253376
rect 272624 250580 302160 253376
rect 302716 250580 332201 253376
rect 332917 250580 362301 253376
rect 363017 250580 392517 253376
rect 393073 250580 651614 253376
rect 66171 250482 651614 250580
rect 56126 250481 651614 250482
rect 652170 250481 670986 253437
rect 56126 250466 670986 250481
rect 54198 249455 669890 249466
rect 54198 249450 650648 249455
rect 54198 246494 66579 249450
rect 67135 249405 650648 249450
rect 67135 249367 287129 249405
rect 67135 246571 196785 249367
rect 197501 246571 226885 249367
rect 227601 246571 256985 249367
rect 257701 246769 287129 249367
rect 287685 249367 650648 249405
rect 287685 249337 347285 249367
rect 287685 246769 317300 249337
rect 257701 246571 317300 246769
rect 67135 246541 317300 246571
rect 317856 246571 347285 249337
rect 348001 246571 377285 249367
rect 378001 246571 407285 249367
rect 408001 246571 650648 249367
rect 317856 246541 650648 246571
rect 67135 246499 650648 246541
rect 651204 249293 669890 249455
rect 651204 246657 667032 249293
rect 669668 246657 669890 249293
rect 651204 246499 669890 246657
rect 67135 246494 669890 246499
rect 54198 246466 669890 246494
rect 54198 221395 55398 246466
rect 56278 245453 654222 245466
rect 56278 245451 653519 245453
rect 56278 245450 212605 245451
rect 56278 245341 63703 245450
rect 56278 242545 56391 245341
rect 63347 242545 63703 245341
rect 56278 242494 63703 242545
rect 64259 242495 212605 245450
rect 213481 242495 242705 245451
rect 243581 242495 272950 245451
rect 273346 242495 303116 245451
rect 303512 242495 333005 245451
rect 333881 242495 363105 245451
rect 363981 242495 393227 245451
rect 393783 242497 653519 245451
rect 654075 242497 654222 245453
rect 393783 242495 654222 242497
rect 64259 242494 654222 242495
rect 56278 242466 654222 242494
rect 56278 241451 653306 241466
rect 56278 241446 652561 241451
rect 56278 241375 64653 241446
rect 56278 238579 56406 241375
rect 63362 238579 64653 241375
rect 56278 238490 64653 238579
rect 65209 238490 197619 241446
rect 198335 238490 227719 241446
rect 228435 238490 257819 241446
rect 258535 238490 288039 241446
rect 288595 238490 318202 241446
rect 318598 238490 348119 241446
rect 348835 238490 378119 241446
rect 378835 238490 408374 241446
rect 408770 238495 652561 241446
rect 653117 238495 653306 241451
rect 408770 238490 653306 238495
rect 56278 238466 653306 238490
rect 56288 237441 605390 237466
rect 56288 237381 210902 237441
rect 56288 234585 56375 237381
rect 63171 234585 210902 237381
rect 56288 234485 210902 234585
rect 211778 234485 241002 237441
rect 241878 234485 271355 237441
rect 271911 237313 331410 237441
rect 271911 234517 301490 237313
rect 302046 234517 331410 237313
rect 271911 234485 331410 234517
rect 332126 234485 361402 237441
rect 362278 234485 391830 237441
rect 392226 234485 605390 237441
rect 698512 236640 711002 249160
rect 56288 234466 605390 234485
rect 56296 233442 601374 233466
rect 56296 233371 196029 233442
rect 56296 230575 56394 233371
rect 63030 232108 196029 233371
rect 63030 232086 169887 232108
rect 63030 231370 89903 232086
rect 93979 231392 169887 232086
rect 173963 231392 196029 232108
rect 93979 231370 196029 231392
rect 63030 230575 196029 231370
rect 56296 230486 196029 230575
rect 196585 230486 226129 233442
rect 226685 230486 256229 233442
rect 256785 230486 286329 233442
rect 286885 230486 316429 233442
rect 316985 230486 346529 233442
rect 347085 230486 376529 233442
rect 377085 230486 406660 233442
rect 407056 232120 601374 233442
rect 407056 231404 429905 232120
rect 433981 231404 601374 232120
rect 407056 230486 601374 231404
rect 56296 230466 601374 230486
rect 55385 220199 55398 221395
rect 53791 218581 53798 219777
rect 54198 219342 55398 220199
rect 52598 217742 53798 218581
rect 598374 212351 601374 230466
rect 7266 209898 7268 210218
rect 8144 209898 8582 210218
rect 47836 209858 53232 210498
rect 574646 209858 596910 210498
rect 6034 208206 6070 208554
rect 6946 208208 8582 208528
rect 8141 206838 8172 206853
rect 8141 206518 8614 206838
rect 8141 206502 8172 206518
rect 6947 205148 6980 205170
rect 6947 204828 8614 205148
rect 6947 204808 6980 204828
rect 6598 183840 19088 196360
rect 47836 184498 50836 209858
rect 596270 208502 596910 209858
rect 598374 209715 598610 212351
rect 601086 209715 601374 212351
rect 596270 208462 597742 208502
rect 596270 207906 596320 208462
rect 597676 207906 597742 208462
rect 596270 207862 597742 207906
rect 598374 197801 601374 209715
rect 598374 197498 598703 197801
rect 51344 197472 53216 197498
rect 51344 196916 51413 197472
rect 52289 196916 53216 197472
rect 51344 196858 53216 196916
rect 574646 197085 598703 197498
rect 601019 197085 601374 197801
rect 574646 196858 601374 197085
rect 47836 183858 53212 184498
rect 574646 184450 596910 184498
rect 574646 183894 596124 184450
rect 596840 183894 596910 184450
rect 574646 183858 596910 183894
rect 41768 176665 45768 176874
rect 41768 173229 42007 176665
rect 45603 173229 45768 176665
rect 41768 171454 45768 173229
rect 41768 170898 42777 171454
rect 45733 170898 45768 171454
rect 41768 145460 45768 170898
rect 47836 166788 50836 183858
rect 598374 171498 601374 196858
rect 51246 171458 53240 171498
rect 51246 170902 51305 171458
rect 52181 170902 53240 171458
rect 51246 170858 53240 170902
rect 574646 170858 601374 171498
rect 41768 144904 42791 145460
rect 45747 144904 45768 145460
rect 6811 111610 18976 123778
rect 41768 119456 45768 144904
rect 41768 118900 42781 119456
rect 45737 118900 45768 119456
rect 41768 93454 45768 118900
rect 41768 92898 42777 93454
rect 45733 92898 45768 93454
rect 41768 82752 45768 92898
rect 6167 70054 19620 80934
rect 41768 78196 41931 82752
rect 45687 78196 45768 82752
rect 41768 72848 45768 78196
rect 41768 68292 41907 72848
rect 45663 68292 45768 72848
rect 41768 67448 45768 68292
rect 41768 66892 41935 67448
rect 45691 66892 45768 67448
rect 41768 51994 45768 66892
rect 41768 48398 42000 51994
rect 45596 48398 45768 51994
rect 41768 48074 45768 48398
rect 46836 158498 50836 166788
rect 598374 167161 601374 170858
rect 598374 166445 598703 167161
rect 601019 166445 601374 167161
rect 46836 157858 53220 158498
rect 574646 158454 596910 158498
rect 574646 157898 594082 158454
rect 596878 157898 596910 158454
rect 574646 157858 596910 157898
rect 46836 132498 50836 157858
rect 598374 145498 601374 166445
rect 602390 226084 605390 234466
rect 602390 224192 640366 226084
rect 648608 225872 651358 226192
rect 602390 224082 641998 224192
rect 602390 208462 605390 224082
rect 639466 223872 641998 224082
rect 650224 222192 651358 225872
rect 648640 221872 651358 222192
rect 650224 212504 651358 221872
rect 607252 212394 669426 212504
rect 607252 212351 641143 212394
rect 607252 209715 607464 212351
rect 609940 209715 641143 212351
rect 607252 209598 641143 209715
rect 642019 209598 669426 212394
rect 607252 209504 669426 209598
rect 602390 207906 602413 208462
rect 605369 207906 605390 208462
rect 602390 184446 605390 207906
rect 666426 197528 669426 209504
rect 605976 197483 607594 197528
rect 606994 197247 607594 197483
rect 605976 197208 607594 197247
rect 665238 197208 669426 197528
rect 602390 183890 602413 184446
rect 605369 183890 605390 184446
rect 602390 182210 605390 183890
rect 602390 181890 607594 182210
rect 602390 158458 605390 181890
rect 666426 166892 669426 197208
rect 698512 191440 711002 203960
rect 605952 166855 607594 166892
rect 606977 166619 607594 166855
rect 605952 166572 607594 166619
rect 665206 166572 669426 166892
rect 605343 157902 605390 158458
rect 51178 145450 53266 145498
rect 51178 144894 51239 145450
rect 52115 144894 53266 145450
rect 51178 144858 53266 144894
rect 574646 144858 601374 145498
rect 598374 136521 601374 144858
rect 598374 135805 598703 136521
rect 601019 135805 601374 136521
rect 46836 131858 53206 132498
rect 574646 132448 596910 132498
rect 574646 131892 594092 132448
rect 596888 131892 596910 132448
rect 574646 131858 596910 131892
rect 46836 106498 50836 131858
rect 598374 119498 601374 135805
rect 51178 119456 53266 119498
rect 51178 118900 51235 119456
rect 52111 118900 53266 119456
rect 51178 118858 53266 118900
rect 574646 118858 601374 119498
rect 46836 105858 53222 106498
rect 574646 106454 596910 106498
rect 574646 105898 594094 106454
rect 596890 105898 596910 106454
rect 574646 105858 596910 105898
rect 46836 80498 50836 105858
rect 598374 105601 601374 118858
rect 598374 104885 598703 105601
rect 601019 104885 601374 105601
rect 598374 93498 601374 104885
rect 51178 93452 53266 93498
rect 51178 92896 51239 93452
rect 52115 92896 53266 93452
rect 51178 92858 53266 92896
rect 574646 92858 601374 93498
rect 46836 79858 53168 80498
rect 574646 80464 596910 80498
rect 574646 79908 594088 80464
rect 596884 79908 596910 80464
rect 574646 79858 596910 79908
rect 46836 46788 50836 79858
rect 598374 67498 601374 92858
rect 51362 67454 53172 67498
rect 51362 66898 51437 67454
rect 52313 66898 53172 67454
rect 51362 66858 53172 66898
rect 574754 66858 601374 67498
rect 598374 52222 601374 66858
rect 54374 51960 601374 52222
rect 54374 48364 54490 51960
rect 58246 50672 601374 51960
rect 58246 49956 143343 50672
rect 144699 49956 601374 50672
rect 58246 48364 601374 49956
rect 54374 48222 601374 48364
rect 602390 151574 605390 157902
rect 602390 151254 607594 151574
rect 602390 132442 605390 151254
rect 666426 136256 669426 166572
rect 698512 146440 711002 158960
rect 605940 136215 607594 136256
rect 606967 135979 607594 136215
rect 605940 135936 607594 135979
rect 665164 135936 669426 136256
rect 602390 131886 602413 132442
rect 605369 131886 605390 132442
rect 602390 120938 605390 131886
rect 602390 120618 607610 120938
rect 602390 106454 605390 120618
rect 602390 105898 602417 106454
rect 605373 105898 605390 106454
rect 602390 98956 605390 105898
rect 666426 105620 669426 135936
rect 605940 105578 607594 105620
rect 605940 105342 605943 105578
rect 606979 105342 607594 105578
rect 605940 105300 607594 105342
rect 665176 105300 669426 105620
rect 602390 98745 657728 98956
rect 602390 98683 656363 98745
rect 602390 96047 625552 98683
rect 626748 98681 656363 98683
rect 626748 96525 636179 98681
rect 636895 96525 656363 98681
rect 626748 96109 656363 96525
rect 657559 96109 657728 98745
rect 626748 96047 657728 96109
rect 602390 95956 657728 96047
rect 602390 80466 605390 95956
rect 624824 89474 627824 95956
rect 634548 94298 641860 94340
rect 634548 94062 634590 94298
rect 634826 94062 641582 94298
rect 641818 94062 641860 94298
rect 634548 94020 641860 94062
rect 643544 93474 646544 93588
rect 641906 93154 646544 93474
rect 624824 89154 629362 89474
rect 624824 89012 627824 89154
rect 602390 79910 602411 80466
rect 605367 79910 605390 80466
rect 602390 47188 605390 79910
rect 625618 75868 627034 89012
rect 643544 85474 646544 93154
rect 650994 92590 653994 95956
rect 666426 93406 669426 105300
rect 698512 101240 711002 113760
rect 662522 93086 669426 93406
rect 650994 92270 657754 92590
rect 650994 90958 653994 92270
rect 666426 91774 669426 93086
rect 662484 91454 669426 91774
rect 650994 90638 657784 90958
rect 650994 90522 653994 90638
rect 666426 90142 669426 91454
rect 662504 89822 669426 90142
rect 641968 85154 646544 85474
rect 643544 81082 646544 85154
rect 666426 81082 669426 89822
rect 632002 80896 669426 81082
rect 632002 80789 640152 80896
rect 632002 78313 632174 80789
rect 632890 78313 640152 80789
rect 632002 78260 640152 78313
rect 640868 78260 669426 80896
rect 632002 78082 669426 78260
rect 645256 77268 647084 78082
rect 629786 77215 647084 77268
rect 629786 77207 642323 77215
rect 629786 77193 633031 77207
rect 629786 76317 629919 77193
rect 630155 76331 633031 77193
rect 633267 77203 642323 77207
rect 633267 76331 636121 77203
rect 630155 76327 636121 76331
rect 636357 76327 639215 77203
rect 639451 76339 642323 77203
rect 642559 76339 647084 77215
rect 639451 76327 647084 76339
rect 630155 76317 647084 76327
rect 629786 76268 647084 76317
rect 625618 75817 644188 75868
rect 625618 75799 643879 75817
rect 625618 75795 637673 75799
rect 625618 75791 634565 75795
rect 625618 74915 631471 75791
rect 631707 74919 634565 75791
rect 634801 74923 637673 75795
rect 637909 75791 643879 75799
rect 637909 74923 640777 75791
rect 634801 74919 640777 74923
rect 631707 74915 640777 74919
rect 641013 74941 643879 75791
rect 644115 74941 644188 75817
rect 641013 74915 644188 74941
rect 625618 74868 644188 74915
rect 625618 71796 626418 74868
rect 646284 73486 647084 76268
rect 645536 73166 647084 73486
rect 625618 71476 626968 71796
rect 625618 68416 626418 71476
rect 646284 70106 647084 73166
rect 645502 69786 647084 70106
rect 625618 68096 626846 68416
rect 646284 66726 647084 69786
rect 645624 66406 647084 66726
rect 666426 47274 669426 78082
rect 602390 47170 649668 47188
rect 602390 46788 648129 47170
rect 46836 46621 648129 46788
rect 46836 46607 251397 46621
rect 46836 45354 241745 46607
rect 46836 44158 141448 45354
rect 142804 44158 241745 45354
rect 46836 42851 241745 44158
rect 245981 42865 251397 46607
rect 255633 46614 648129 46621
rect 649645 46614 649668 47170
rect 666426 47038 666442 47274
rect 669398 47038 669426 47274
rect 666426 46978 669426 47038
rect 255633 46588 649668 46614
rect 255633 45788 605390 46588
rect 255633 42865 605396 45788
rect 245981 42851 605396 42865
rect 46836 42788 605396 42851
rect 80222 6811 92390 18976
rect 136713 7143 144150 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19620
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18976
rect 624222 6811 636390 18976
use user_id_programming  user_id_value
timestamp 1648835380
transform 1 0 656624 0 1 88126
box 0 0 7109 7077
use mgmt_core_wrapper  soc
timestamp 1648835380
transform 1 0 52034 0 1 53002
box 382 -400 524400 164400
use xres_buf  rstb_level
timestamp 1648835380
transform -1 0 145710 0 -1 50488
box 414 -400 3522 3800
use simple_por  por
timestamp 1648835380
transform 1 0 650146 0 -1 55282
box 25 11 11344 8291
use digital_pll  pll
timestamp 1648835380
transform 1 0 628146 0 1 80944
box 0 0 15000 15000
use housekeeping  housekeeping
timestamp 1648835380
transform 1 0 606434 0 1 100002
box 0 0 60046 110190
use gpio_defaults_block  gpio_defaults_block_0\[0\]
timestamp 1648835380
transform -1 0 709467 0 1 134000
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_1\[0\]
timestamp 1648835380
transform -1 0 710203 0 1 121000
box 14 416 34000 13000
use caravel_clocking  clocking
timestamp 1648835380
transform 1 0 626764 0 1 63284
box -38 -48 20000 12000
use gpio_control_block  gpio_control_bidir_2\[2\]
timestamp 1648835380
transform 1 0 7631 0 1 202600
box 14 416 34000 13000
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1648835380
transform -1 0 710203 0 1 166200
box 14 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_0\[1\]
timestamp 1648835380
transform -1 0 709467 0 1 179200
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1648835380
transform 1 0 7631 0 1 245800
box 14 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_37
timestamp 1648835380
transform 1 0 8367 0 1 215600
box -38 0 6018 2224
use mgmt_protect  mgmt_buffers
timestamp 1648835380
transform 1 0 192180 0 1 232036
box -400 -400 220400 32400
use spare_logic_block  spare_logic\[0\]
timestamp 1648835380
transform 1 0 88632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[1\]
timestamp 1648835380
transform 1 0 168632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[3\]
timestamp 1648835380
transform 1 0 428632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[2\]
timestamp 1648835380
transform 1 0 640874 0 1 220592
box 0 0 9000 9000
use gpio_control_block  gpio_control_in_1a\[0\]
timestamp 1648835380
transform -1 0 710203 0 1 211200
box 14 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_2\[0\]
timestamp 1648835380
transform -1 0 709467 0 1 224200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_36
timestamp 1648835380
transform 1 0 8367 0 1 258800
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[1\]
timestamp 1648835380
transform -1 0 710203 0 1 256400
box 14 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_2\[1\]
timestamp 1648835380
transform -1 0 709467 0 1 269400
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1648835380
transform 1 0 7631 0 1 289000
box 14 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_35
timestamp 1648835380
transform 1 0 8367 0 1 302000
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[2\]
timestamp 1648835380
transform -1 0 710203 0 1 301400
box 14 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_2\[2\]
timestamp 1648835380
transform -1 0 709467 0 1 314400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[13\]
timestamp 1648835380
transform 1 0 7631 0 1 418600
box 14 416 34000 13000
use gpio_control_block  gpio_control_in_2\[14\]
timestamp 1648835380
transform 1 0 7631 0 1 375400
box 14 416 34000 13000
use gpio_control_block  gpio_control_in_2\[15\]
timestamp 1648835380
transform 1 0 7631 0 1 332200
box 14 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_32
timestamp 1648835380
transform 1 0 8367 0 1 431600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_33
timestamp 1648835380
transform 1 0 8367 0 1 388400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_34
timestamp 1648835380
transform 1 0 8367 0 1 345200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[3\]
timestamp 1648835380
transform -1 0 710203 0 1 346400
box 14 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[4\]
timestamp 1648835380
transform -1 0 710203 0 1 391600
box 14 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[5\]
timestamp 1648835380
transform -1 0 710203 0 1 479800
box 14 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_5
timestamp 1648835380
transform -1 0 709467 0 1 359400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_6
timestamp 1648835380
transform -1 0 709467 0 1 404600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_7
timestamp 1648835380
transform -1 0 709467 0 1 492800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_31
timestamp 1648835380
transform 1 0 8367 0 1 559200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_30
timestamp 1648835380
transform 1 0 8367 0 1 602400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[12\]
timestamp 1648835380
transform 1 0 7631 0 1 546200
box 14 416 34000 13000
use gpio_control_block  gpio_control_in_2\[11\]
timestamp 1648835380
transform 1 0 7631 0 1 589400
box 14 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_9
timestamp 1648835380
transform -1 0 709467 0 1 581800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_8
timestamp 1648835380
transform -1 0 709467 0 1 536800
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1648835380
transform -1 0 710203 0 1 568800
box 14 416 34000 13000
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1648835380
transform -1 0 710203 0 1 523800
box 14 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_29
timestamp 1648835380
transform 1 0 8367 0 1 645600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_28
timestamp 1648835380
transform 1 0 8367 0 1 688800
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1648835380
transform 1 0 7631 0 1 675800
box 14 416 34000 13000
use gpio_control_block  gpio_control_in_2\[10\]
timestamp 1648835380
transform 1 0 7631 0 1 632600
box 14 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_11
timestamp 1648835380
transform -1 0 709467 0 1 672000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_10
timestamp 1648835380
transform -1 0 709467 0 1 627000
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1648835380
transform -1 0 710203 0 1 659000
box 14 416 34000 13000
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1648835380
transform -1 0 710203 0 1 614000
box 14 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_27
timestamp 1648835380
transform 1 0 8367 0 1 732000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_26
timestamp 1648835380
transform 1 0 8367 0 1 775200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1648835380
transform 1 0 7631 0 1 719000
box 14 416 34000 13000
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1648835380
transform 1 0 7631 0 1 762200
box 14 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_13
timestamp 1648835380
transform -1 0 709467 0 1 762200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_12
timestamp 1648835380
transform -1 0 709467 0 1 717200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1648835380
transform -1 0 710203 0 1 749200
box 14 416 34000 13000
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1648835380
transform -1 0 710203 0 1 704200
box 14 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_25
timestamp 1648835380
transform 1 0 8367 0 1 818400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1648835380
transform 1 0 7631 0 1 805400
box 14 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_24
timestamp 1648835380
transform 1 0 8367 0 1 944200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1648835380
transform 1 0 7631 0 1 931200
box 14 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_14
timestamp 1648835380
transform -1 0 709467 0 1 940600
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[6\]
timestamp 1648835380
transform -1 0 710203 0 1 927600
box 14 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_23
timestamp 1648835380
transform 0 1 110194 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_22
timestamp 1648835380
transform 0 1 161594 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1648835380
transform 0 1 97200 -1 0 1030077
box 14 416 34000 13000
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1648835380
transform 0 1 148600 -1 0 1030077
box 14 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_21
timestamp 1648835380
transform 0 1 212994 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1648835380
transform 0 1 200000 -1 0 1030077
box 14 416 34000 13000
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1648835380
transform 0 1 251400 -1 0 1030077
box 14 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_20
timestamp 1648835380
transform 0 1 264394 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_19
timestamp 1648835380
transform 0 1 315994 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1648835380
transform 0 1 303000 -1 0 1030077
box 14 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_18
timestamp 1648835380
transform 0 1 366394 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_17
timestamp 1648835380
transform 0 1 433794 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[9\]
timestamp 1648835380
transform 0 1 420800 -1 0 1030077
box 14 416 34000 13000
use gpio_control_block  gpio_control_in_1\[10\]
timestamp 1648835380
transform 0 1 353400 -1 0 1030077
box 14 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_16
timestamp 1648835380
transform 0 1 510794 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[8\]
timestamp 1648835380
transform 0 1 497800 -1 0 1030077
box 14 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_15
timestamp 1648835380
transform 0 1 562194 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[7\]
timestamp 1648835380
transform 0 1 549200 -1 0 1030077
box 14 416 34000 13000
use user_project_wrapper  mprj
timestamp 1648835380
transform 1 0 65308 0 1 278718
box -8726 -7654 592650 711590
use chip_io  padframe
timestamp 1648835380
transform 1 0 0 0 1 0
box 0 0 717600 1037600
<< labels >>
rlabel metal5 s 187640 6598 200160 19088 6 clock
port 0 nsew signal input
rlabel metal5 s 351040 6598 363560 19088 6 flash_clk
port 1 nsew signal tristate
rlabel metal5 s 296240 6598 308760 19088 6 flash_csb
port 2 nsew signal tristate
rlabel metal5 s 405840 6598 418360 19088 6 flash_io0
port 3 nsew signal tristate
rlabel metal5 s 460640 6598 473160 19088 6 flash_io1
port 4 nsew signal tristate
rlabel metal5 s 515440 6598 527960 19088 6 gpio
port 5 nsew signal bidirectional
rlabel metal5 s 698512 101240 711002 113760 6 mprj_io[0]
port 6 nsew signal bidirectional
rlabel metal5 s 698512 684440 711002 696960 6 mprj_io[10]
port 7 nsew signal bidirectional
rlabel metal5 s 698512 729440 711002 741960 6 mprj_io[11]
port 8 nsew signal bidirectional
rlabel metal5 s 698512 774440 711002 786960 6 mprj_io[12]
port 9 nsew signal bidirectional
rlabel metal5 s 698512 863640 711002 876160 6 mprj_io[13]
port 10 nsew signal bidirectional
rlabel metal5 s 698512 952840 711002 965360 6 mprj_io[14]
port 11 nsew signal bidirectional
rlabel metal5 s 628240 1018512 640760 1031002 6 mprj_io[15]
port 12 nsew signal bidirectional
rlabel metal5 s 526440 1018512 538960 1031002 6 mprj_io[16]
port 13 nsew signal bidirectional
rlabel metal5 s 475040 1018512 487560 1031002 6 mprj_io[17]
port 14 nsew signal bidirectional
rlabel metal5 s 386040 1018512 398560 1031002 6 mprj_io[18]
port 15 nsew signal bidirectional
rlabel metal5 s 284240 1018512 296760 1031002 6 mprj_io[19]
port 16 nsew signal bidirectional
rlabel metal5 s 698512 146440 711002 158960 6 mprj_io[1]
port 17 nsew signal bidirectional
rlabel metal5 s 232640 1018512 245160 1031002 6 mprj_io[20]
port 18 nsew signal bidirectional
rlabel metal5 s 181240 1018512 193760 1031002 6 mprj_io[21]
port 19 nsew signal bidirectional
rlabel metal5 s 129840 1018512 142360 1031002 6 mprj_io[22]
port 20 nsew signal bidirectional
rlabel metal5 s 78440 1018512 90960 1031002 6 mprj_io[23]
port 21 nsew signal bidirectional
rlabel metal5 s 6598 956440 19088 968960 6 mprj_io[24]
port 22 nsew signal bidirectional
rlabel metal5 s 6598 786640 19088 799160 6 mprj_io[25]
port 23 nsew signal bidirectional
rlabel metal5 s 6598 743440 19088 755960 6 mprj_io[26]
port 24 nsew signal bidirectional
rlabel metal5 s 6598 700240 19088 712760 6 mprj_io[27]
port 25 nsew signal bidirectional
rlabel metal5 s 6598 657040 19088 669560 6 mprj_io[28]
port 26 nsew signal bidirectional
rlabel metal5 s 6598 613840 19088 626360 6 mprj_io[29]
port 27 nsew signal bidirectional
rlabel metal5 s 698512 191440 711002 203960 6 mprj_io[2]
port 28 nsew signal bidirectional
rlabel metal5 s 6598 570640 19088 583160 6 mprj_io[30]
port 29 nsew signal bidirectional
rlabel metal5 s 6598 527440 19088 539960 6 mprj_io[31]
port 30 nsew signal bidirectional
rlabel metal5 s 6598 399840 19088 412360 6 mprj_io[32]
port 31 nsew signal bidirectional
rlabel metal5 s 6598 356640 19088 369160 6 mprj_io[33]
port 32 nsew signal bidirectional
rlabel metal5 s 6598 313440 19088 325960 6 mprj_io[34]
port 33 nsew signal bidirectional
rlabel metal5 s 6598 270240 19088 282760 6 mprj_io[35]
port 34 nsew signal bidirectional
rlabel metal5 s 6598 227040 19088 239560 6 mprj_io[36]
port 35 nsew signal bidirectional
rlabel metal5 s 6598 183840 19088 196360 6 mprj_io[37]
port 36 nsew signal bidirectional
rlabel metal5 s 698512 236640 711002 249160 6 mprj_io[3]
port 37 nsew signal bidirectional
rlabel metal5 s 698512 281640 711002 294160 6 mprj_io[4]
port 38 nsew signal bidirectional
rlabel metal5 s 698512 326640 711002 339160 6 mprj_io[5]
port 39 nsew signal bidirectional
rlabel metal5 s 698512 371840 711002 384360 6 mprj_io[6]
port 40 nsew signal bidirectional
rlabel metal5 s 698512 549040 711002 561560 6 mprj_io[7]
port 41 nsew signal bidirectional
rlabel metal5 s 698512 594240 711002 606760 6 mprj_io[8]
port 42 nsew signal bidirectional
rlabel metal5 s 698512 639240 711002 651760 6 mprj_io[9]
port 43 nsew signal bidirectional
rlabel metal5 s 136713 7143 144150 18309 6 resetb
port 44 nsew signal input
rlabel metal5 s 6167 70054 19620 80934 6 vccd
port 45 nsew signal bidirectional
rlabel metal5 s 697980 909666 711433 920546 6 vccd1
port 46 nsew signal bidirectional
rlabel metal5 s 6167 914054 19620 924934 6 vccd2
port 47 nsew signal bidirectional
rlabel metal5 s 624222 6811 636390 18976 6 vdda
port 48 nsew signal bidirectional
rlabel metal5 s 698624 819822 710789 831990 6 vdda1
port 49 nsew signal bidirectional
rlabel metal5 s 698624 505222 710789 517390 6 vdda1_2
port 50 nsew signal bidirectional
rlabel metal5 s 6811 484410 18976 496578 6 vdda2
port 51 nsew signal bidirectional
rlabel metal5 s 6811 111610 18976 123778 6 vddio
port 52 nsew signal bidirectional
rlabel metal5 s 6811 871210 18976 883378 6 vddio_2
port 53 nsew signal bidirectional
rlabel metal5 s 80222 6811 92390 18976 6 vssa
port 54 nsew signal bidirectional
rlabel metal5 s 577010 1018624 589178 1030789 6 vssa1
port 55 nsew signal bidirectional
rlabel metal5 s 698624 417022 710789 429190 6 vssa1_2
port 56 nsew signal bidirectional
rlabel metal5 s 6811 829010 18976 841178 6 vssa2
port 57 nsew signal bidirectional
rlabel metal5 s 243266 6167 254146 19620 6 vssd
port 58 nsew signal bidirectional
rlabel metal5 s 697980 461866 711433 472746 6 vssd1
port 59 nsew signal bidirectional
rlabel metal5 s 6167 442854 19620 453734 6 vssd2
port 60 nsew signal bidirectional
rlabel metal5 s 570422 6811 582590 18976 6 vssio
port 61 nsew signal bidirectional
rlabel metal5 s 334810 1018624 346978 1030789 6 vssio_2
port 62 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
