VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO housekeeping
  CLASS BLOCK ;
  FOREIGN housekeeping ;
  ORIGIN 0.000 0.000 ;
  SIZE 370.230 BY 550.950 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 538.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 103.080 364.560 104.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 256.260 364.560 257.860 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 409.440 364.560 411.040 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 538.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.490 364.560 28.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.670 364.560 181.270 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 332.850 364.560 334.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 486.030 364.560 487.630 ;
    END
  END VPWR
  PIN debug_in
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END debug_in
  PIN debug_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END debug_mode
  PIN debug_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END debug_oeb
  PIN debug_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END debug_out
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END irq[2]
  PIN mask_rev_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END mask_rev_in[0]
  PIN mask_rev_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END mask_rev_in[10]
  PIN mask_rev_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 0.000 266.250 4.000 ;
    END
  END mask_rev_in[11]
  PIN mask_rev_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END mask_rev_in[12]
  PIN mask_rev_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END mask_rev_in[13]
  PIN mask_rev_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END mask_rev_in[14]
  PIN mask_rev_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END mask_rev_in[15]
  PIN mask_rev_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END mask_rev_in[16]
  PIN mask_rev_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END mask_rev_in[17]
  PIN mask_rev_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END mask_rev_in[18]
  PIN mask_rev_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END mask_rev_in[19]
  PIN mask_rev_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 0.000 229.450 4.000 ;
    END
  END mask_rev_in[1]
  PIN mask_rev_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 0.000 299.370 4.000 ;
    END
  END mask_rev_in[20]
  PIN mask_rev_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END mask_rev_in[21]
  PIN mask_rev_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 4.000 ;
    END
  END mask_rev_in[22]
  PIN mask_rev_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 0.000 310.410 4.000 ;
    END
  END mask_rev_in[23]
  PIN mask_rev_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END mask_rev_in[24]
  PIN mask_rev_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END mask_rev_in[25]
  PIN mask_rev_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 0.000 321.450 4.000 ;
    END
  END mask_rev_in[26]
  PIN mask_rev_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END mask_rev_in[27]
  PIN mask_rev_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END mask_rev_in[28]
  PIN mask_rev_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END mask_rev_in[29]
  PIN mask_rev_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 0.000 233.130 4.000 ;
    END
  END mask_rev_in[2]
  PIN mask_rev_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END mask_rev_in[30]
  PIN mask_rev_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 4.000 ;
    END
  END mask_rev_in[31]
  PIN mask_rev_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END mask_rev_in[3]
  PIN mask_rev_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END mask_rev_in[4]
  PIN mask_rev_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 4.000 ;
    END
  END mask_rev_in[5]
  PIN mask_rev_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 4.000 ;
    END
  END mask_rev_in[6]
  PIN mask_rev_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END mask_rev_in[7]
  PIN mask_rev_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END mask_rev_in[8]
  PIN mask_rev_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END mask_rev_in[9]
  PIN mgmt_gpio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 54.440 370.230 55.040 ;
    END
  END mgmt_gpio_in[0]
  PIN mgmt_gpio_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 299.240 370.230 299.840 ;
    END
  END mgmt_gpio_in[10]
  PIN mgmt_gpio_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 323.720 370.230 324.320 ;
    END
  END mgmt_gpio_in[11]
  PIN mgmt_gpio_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 348.200 370.230 348.800 ;
    END
  END mgmt_gpio_in[12]
  PIN mgmt_gpio_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 372.680 370.230 373.280 ;
    END
  END mgmt_gpio_in[13]
  PIN mgmt_gpio_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 397.160 370.230 397.760 ;
    END
  END mgmt_gpio_in[14]
  PIN mgmt_gpio_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 421.640 370.230 422.240 ;
    END
  END mgmt_gpio_in[15]
  PIN mgmt_gpio_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 446.120 370.230 446.720 ;
    END
  END mgmt_gpio_in[16]
  PIN mgmt_gpio_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 470.600 370.230 471.200 ;
    END
  END mgmt_gpio_in[17]
  PIN mgmt_gpio_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 495.080 370.230 495.680 ;
    END
  END mgmt_gpio_in[18]
  PIN mgmt_gpio_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 519.560 370.230 520.160 ;
    END
  END mgmt_gpio_in[19]
  PIN mgmt_gpio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 78.920 370.230 79.520 ;
    END
  END mgmt_gpio_in[1]
  PIN mgmt_gpio_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 546.950 214.270 550.950 ;
    END
  END mgmt_gpio_in[20]
  PIN mgmt_gpio_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 546.950 222.550 550.950 ;
    END
  END mgmt_gpio_in[21]
  PIN mgmt_gpio_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 546.950 230.830 550.950 ;
    END
  END mgmt_gpio_in[22]
  PIN mgmt_gpio_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 546.950 239.110 550.950 ;
    END
  END mgmt_gpio_in[23]
  PIN mgmt_gpio_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 546.950 247.390 550.950 ;
    END
  END mgmt_gpio_in[24]
  PIN mgmt_gpio_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 546.950 255.670 550.950 ;
    END
  END mgmt_gpio_in[25]
  PIN mgmt_gpio_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 546.950 263.950 550.950 ;
    END
  END mgmt_gpio_in[26]
  PIN mgmt_gpio_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 546.950 272.230 550.950 ;
    END
  END mgmt_gpio_in[27]
  PIN mgmt_gpio_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 546.950 280.510 550.950 ;
    END
  END mgmt_gpio_in[28]
  PIN mgmt_gpio_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 546.950 288.790 550.950 ;
    END
  END mgmt_gpio_in[29]
  PIN mgmt_gpio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 103.400 370.230 104.000 ;
    END
  END mgmt_gpio_in[2]
  PIN mgmt_gpio_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 546.950 297.070 550.950 ;
    END
  END mgmt_gpio_in[30]
  PIN mgmt_gpio_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 546.950 305.350 550.950 ;
    END
  END mgmt_gpio_in[31]
  PIN mgmt_gpio_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 546.950 313.630 550.950 ;
    END
  END mgmt_gpio_in[32]
  PIN mgmt_gpio_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 546.950 321.910 550.950 ;
    END
  END mgmt_gpio_in[33]
  PIN mgmt_gpio_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 546.950 330.190 550.950 ;
    END
  END mgmt_gpio_in[34]
  PIN mgmt_gpio_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 546.950 338.470 550.950 ;
    END
  END mgmt_gpio_in[35]
  PIN mgmt_gpio_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 546.950 346.750 550.950 ;
    END
  END mgmt_gpio_in[36]
  PIN mgmt_gpio_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 546.950 355.030 550.950 ;
    END
  END mgmt_gpio_in[37]
  PIN mgmt_gpio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 127.880 370.230 128.480 ;
    END
  END mgmt_gpio_in[3]
  PIN mgmt_gpio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 152.360 370.230 152.960 ;
    END
  END mgmt_gpio_in[4]
  PIN mgmt_gpio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 176.840 370.230 177.440 ;
    END
  END mgmt_gpio_in[5]
  PIN mgmt_gpio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 201.320 370.230 201.920 ;
    END
  END mgmt_gpio_in[6]
  PIN mgmt_gpio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 225.800 370.230 226.400 ;
    END
  END mgmt_gpio_in[7]
  PIN mgmt_gpio_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 250.280 370.230 250.880 ;
    END
  END mgmt_gpio_in[8]
  PIN mgmt_gpio_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 274.760 370.230 275.360 ;
    END
  END mgmt_gpio_in[9]
  PIN mgmt_gpio_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 62.600 370.230 63.200 ;
    END
  END mgmt_gpio_oeb[0]
  PIN mgmt_gpio_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 307.400 370.230 308.000 ;
    END
  END mgmt_gpio_oeb[10]
  PIN mgmt_gpio_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 331.880 370.230 332.480 ;
    END
  END mgmt_gpio_oeb[11]
  PIN mgmt_gpio_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 356.360 370.230 356.960 ;
    END
  END mgmt_gpio_oeb[12]
  PIN mgmt_gpio_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 380.840 370.230 381.440 ;
    END
  END mgmt_gpio_oeb[13]
  PIN mgmt_gpio_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 405.320 370.230 405.920 ;
    END
  END mgmt_gpio_oeb[14]
  PIN mgmt_gpio_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 429.800 370.230 430.400 ;
    END
  END mgmt_gpio_oeb[15]
  PIN mgmt_gpio_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 454.280 370.230 454.880 ;
    END
  END mgmt_gpio_oeb[16]
  PIN mgmt_gpio_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 478.760 370.230 479.360 ;
    END
  END mgmt_gpio_oeb[17]
  PIN mgmt_gpio_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 503.240 370.230 503.840 ;
    END
  END mgmt_gpio_oeb[18]
  PIN mgmt_gpio_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 527.720 370.230 528.320 ;
    END
  END mgmt_gpio_oeb[19]
  PIN mgmt_gpio_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 87.080 370.230 87.680 ;
    END
  END mgmt_gpio_oeb[1]
  PIN mgmt_gpio_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 546.950 217.030 550.950 ;
    END
  END mgmt_gpio_oeb[20]
  PIN mgmt_gpio_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 546.950 225.310 550.950 ;
    END
  END mgmt_gpio_oeb[21]
  PIN mgmt_gpio_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 546.950 233.590 550.950 ;
    END
  END mgmt_gpio_oeb[22]
  PIN mgmt_gpio_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 546.950 241.870 550.950 ;
    END
  END mgmt_gpio_oeb[23]
  PIN mgmt_gpio_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 546.950 250.150 550.950 ;
    END
  END mgmt_gpio_oeb[24]
  PIN mgmt_gpio_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 546.950 258.430 550.950 ;
    END
  END mgmt_gpio_oeb[25]
  PIN mgmt_gpio_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 546.950 266.710 550.950 ;
    END
  END mgmt_gpio_oeb[26]
  PIN mgmt_gpio_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 546.950 274.990 550.950 ;
    END
  END mgmt_gpio_oeb[27]
  PIN mgmt_gpio_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 546.950 283.270 550.950 ;
    END
  END mgmt_gpio_oeb[28]
  PIN mgmt_gpio_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 546.950 291.550 550.950 ;
    END
  END mgmt_gpio_oeb[29]
  PIN mgmt_gpio_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 111.560 370.230 112.160 ;
    END
  END mgmt_gpio_oeb[2]
  PIN mgmt_gpio_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 546.950 299.830 550.950 ;
    END
  END mgmt_gpio_oeb[30]
  PIN mgmt_gpio_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 546.950 308.110 550.950 ;
    END
  END mgmt_gpio_oeb[31]
  PIN mgmt_gpio_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 546.950 316.390 550.950 ;
    END
  END mgmt_gpio_oeb[32]
  PIN mgmt_gpio_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 546.950 324.670 550.950 ;
    END
  END mgmt_gpio_oeb[33]
  PIN mgmt_gpio_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 546.950 332.950 550.950 ;
    END
  END mgmt_gpio_oeb[34]
  PIN mgmt_gpio_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 546.950 341.230 550.950 ;
    END
  END mgmt_gpio_oeb[35]
  PIN mgmt_gpio_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 546.950 349.510 550.950 ;
    END
  END mgmt_gpio_oeb[36]
  PIN mgmt_gpio_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 546.950 357.790 550.950 ;
    END
  END mgmt_gpio_oeb[37]
  PIN mgmt_gpio_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 136.040 370.230 136.640 ;
    END
  END mgmt_gpio_oeb[3]
  PIN mgmt_gpio_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 160.520 370.230 161.120 ;
    END
  END mgmt_gpio_oeb[4]
  PIN mgmt_gpio_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 185.000 370.230 185.600 ;
    END
  END mgmt_gpio_oeb[5]
  PIN mgmt_gpio_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 209.480 370.230 210.080 ;
    END
  END mgmt_gpio_oeb[6]
  PIN mgmt_gpio_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 233.960 370.230 234.560 ;
    END
  END mgmt_gpio_oeb[7]
  PIN mgmt_gpio_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 258.440 370.230 259.040 ;
    END
  END mgmt_gpio_oeb[8]
  PIN mgmt_gpio_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 282.920 370.230 283.520 ;
    END
  END mgmt_gpio_oeb[9]
  PIN mgmt_gpio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 70.760 370.230 71.360 ;
    END
  END mgmt_gpio_out[0]
  PIN mgmt_gpio_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 315.560 370.230 316.160 ;
    END
  END mgmt_gpio_out[10]
  PIN mgmt_gpio_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 340.040 370.230 340.640 ;
    END
  END mgmt_gpio_out[11]
  PIN mgmt_gpio_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 364.520 370.230 365.120 ;
    END
  END mgmt_gpio_out[12]
  PIN mgmt_gpio_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 389.000 370.230 389.600 ;
    END
  END mgmt_gpio_out[13]
  PIN mgmt_gpio_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 413.480 370.230 414.080 ;
    END
  END mgmt_gpio_out[14]
  PIN mgmt_gpio_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 437.960 370.230 438.560 ;
    END
  END mgmt_gpio_out[15]
  PIN mgmt_gpio_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 462.440 370.230 463.040 ;
    END
  END mgmt_gpio_out[16]
  PIN mgmt_gpio_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 486.920 370.230 487.520 ;
    END
  END mgmt_gpio_out[17]
  PIN mgmt_gpio_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 511.400 370.230 512.000 ;
    END
  END mgmt_gpio_out[18]
  PIN mgmt_gpio_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 535.880 370.230 536.480 ;
    END
  END mgmt_gpio_out[19]
  PIN mgmt_gpio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 95.240 370.230 95.840 ;
    END
  END mgmt_gpio_out[1]
  PIN mgmt_gpio_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 546.950 219.790 550.950 ;
    END
  END mgmt_gpio_out[20]
  PIN mgmt_gpio_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 546.950 228.070 550.950 ;
    END
  END mgmt_gpio_out[21]
  PIN mgmt_gpio_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 546.950 236.350 550.950 ;
    END
  END mgmt_gpio_out[22]
  PIN mgmt_gpio_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 546.950 244.630 550.950 ;
    END
  END mgmt_gpio_out[23]
  PIN mgmt_gpio_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 546.950 252.910 550.950 ;
    END
  END mgmt_gpio_out[24]
  PIN mgmt_gpio_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 546.950 261.190 550.950 ;
    END
  END mgmt_gpio_out[25]
  PIN mgmt_gpio_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 546.950 269.470 550.950 ;
    END
  END mgmt_gpio_out[26]
  PIN mgmt_gpio_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 546.950 277.750 550.950 ;
    END
  END mgmt_gpio_out[27]
  PIN mgmt_gpio_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 546.950 286.030 550.950 ;
    END
  END mgmt_gpio_out[28]
  PIN mgmt_gpio_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 546.950 294.310 550.950 ;
    END
  END mgmt_gpio_out[29]
  PIN mgmt_gpio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 119.720 370.230 120.320 ;
    END
  END mgmt_gpio_out[2]
  PIN mgmt_gpio_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 546.950 302.590 550.950 ;
    END
  END mgmt_gpio_out[30]
  PIN mgmt_gpio_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 546.950 310.870 550.950 ;
    END
  END mgmt_gpio_out[31]
  PIN mgmt_gpio_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 546.950 319.150 550.950 ;
    END
  END mgmt_gpio_out[32]
  PIN mgmt_gpio_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 546.950 327.430 550.950 ;
    END
  END mgmt_gpio_out[33]
  PIN mgmt_gpio_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 546.950 335.710 550.950 ;
    END
  END mgmt_gpio_out[34]
  PIN mgmt_gpio_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 546.950 343.990 550.950 ;
    END
  END mgmt_gpio_out[35]
  PIN mgmt_gpio_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 546.950 352.270 550.950 ;
    END
  END mgmt_gpio_out[36]
  PIN mgmt_gpio_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 546.950 360.550 550.950 ;
    END
  END mgmt_gpio_out[37]
  PIN mgmt_gpio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 144.200 370.230 144.800 ;
    END
  END mgmt_gpio_out[3]
  PIN mgmt_gpio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 168.680 370.230 169.280 ;
    END
  END mgmt_gpio_out[4]
  PIN mgmt_gpio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 193.160 370.230 193.760 ;
    END
  END mgmt_gpio_out[5]
  PIN mgmt_gpio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 217.640 370.230 218.240 ;
    END
  END mgmt_gpio_out[6]
  PIN mgmt_gpio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 242.120 370.230 242.720 ;
    END
  END mgmt_gpio_out[7]
  PIN mgmt_gpio_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 266.600 370.230 267.200 ;
    END
  END mgmt_gpio_out[8]
  PIN mgmt_gpio_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 291.080 370.230 291.680 ;
    END
  END mgmt_gpio_out[9]
  PIN pad_flash_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END pad_flash_clk
  PIN pad_flash_clk_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END pad_flash_clk_oeb
  PIN pad_flash_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END pad_flash_csb
  PIN pad_flash_csb_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END pad_flash_csb_oeb
  PIN pad_flash_io0_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END pad_flash_io0_di
  PIN pad_flash_io0_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END pad_flash_io0_do
  PIN pad_flash_io0_ieb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END pad_flash_io0_ieb
  PIN pad_flash_io0_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END pad_flash_io0_oeb
  PIN pad_flash_io1_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END pad_flash_io1_di
  PIN pad_flash_io1_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END pad_flash_io1_do
  PIN pad_flash_io1_ieb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END pad_flash_io1_ieb
  PIN pad_flash_io1_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END pad_flash_io1_oeb
  PIN pll90_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 4.000 ;
    END
  END pll90_sel[0]
  PIN pll90_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END pll90_sel[1]
  PIN pll90_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END pll90_sel[2]
  PIN pll_bypass
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END pll_bypass
  PIN pll_dco_ena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END pll_dco_ena
  PIN pll_div[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END pll_div[0]
  PIN pll_div[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END pll_div[1]
  PIN pll_div[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END pll_div[2]
  PIN pll_div[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END pll_div[3]
  PIN pll_div[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END pll_div[4]
  PIN pll_ena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END pll_ena
  PIN pll_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END pll_sel[0]
  PIN pll_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END pll_sel[1]
  PIN pll_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END pll_sel[2]
  PIN pll_trim[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END pll_trim[0]
  PIN pll_trim[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END pll_trim[10]
  PIN pll_trim[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END pll_trim[11]
  PIN pll_trim[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END pll_trim[12]
  PIN pll_trim[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END pll_trim[13]
  PIN pll_trim[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END pll_trim[14]
  PIN pll_trim[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END pll_trim[15]
  PIN pll_trim[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END pll_trim[16]
  PIN pll_trim[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END pll_trim[17]
  PIN pll_trim[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END pll_trim[18]
  PIN pll_trim[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 4.000 ;
    END
  END pll_trim[19]
  PIN pll_trim[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END pll_trim[1]
  PIN pll_trim[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END pll_trim[20]
  PIN pll_trim[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 0.000 196.330 4.000 ;
    END
  END pll_trim[21]
  PIN pll_trim[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END pll_trim[22]
  PIN pll_trim[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END pll_trim[23]
  PIN pll_trim[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END pll_trim[24]
  PIN pll_trim[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 0.000 211.050 4.000 ;
    END
  END pll_trim[25]
  PIN pll_trim[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END pll_trim[2]
  PIN pll_trim[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END pll_trim[3]
  PIN pll_trim[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END pll_trim[4]
  PIN pll_trim[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END pll_trim[5]
  PIN pll_trim[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END pll_trim[6]
  PIN pll_trim[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END pll_trim[7]
  PIN pll_trim[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END pll_trim[8]
  PIN pll_trim[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END pll_trim[9]
  PIN porb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END porb
  PIN pwr_ctrl_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 4.000 ;
    END
  END pwr_ctrl_out[0]
  PIN pwr_ctrl_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.930 0.000 347.210 4.000 ;
    END
  END pwr_ctrl_out[1]
  PIN pwr_ctrl_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END pwr_ctrl_out[2]
  PIN pwr_ctrl_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END pwr_ctrl_out[3]
  PIN qspi_enabled
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END qspi_enabled
  PIN reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END reset
  PIN ser_rx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END ser_rx
  PIN ser_tx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END ser_tx
  PIN serial_clock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 13.640 370.230 14.240 ;
    END
  END serial_clock
  PIN serial_data_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 38.120 370.230 38.720 ;
    END
  END serial_data_1
  PIN serial_data_2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 46.280 370.230 46.880 ;
    END
  END serial_data_2
  PIN serial_load
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 29.960 370.230 30.560 ;
    END
  END serial_load
  PIN serial_resetn
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.230 21.800 370.230 22.400 ;
    END
  END serial_resetn
  PIN spi_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END spi_csb
  PIN spi_enabled
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END spi_enabled
  PIN spi_sck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END spi_sck
  PIN spi_sdi
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END spi_sdi
  PIN spi_sdo
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END spi_sdo
  PIN spi_sdoenb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END spi_sdoenb
  PIN spimemio_flash_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 4.000 434.480 ;
    END
  END spimemio_flash_clk
  PIN spimemio_flash_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END spimemio_flash_csb
  PIN spimemio_flash_io0_di
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.200 4.000 450.800 ;
    END
  END spimemio_flash_io0_di
  PIN spimemio_flash_io0_do
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 4.000 458.960 ;
    END
  END spimemio_flash_io0_do
  PIN spimemio_flash_io0_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 4.000 467.120 ;
    END
  END spimemio_flash_io0_oeb
  PIN spimemio_flash_io1_di
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.680 4.000 475.280 ;
    END
  END spimemio_flash_io1_di
  PIN spimemio_flash_io1_do
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END spimemio_flash_io1_do
  PIN spimemio_flash_io1_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END spimemio_flash_io1_oeb
  PIN spimemio_flash_io2_di
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END spimemio_flash_io2_di
  PIN spimemio_flash_io2_do
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END spimemio_flash_io2_do
  PIN spimemio_flash_io2_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END spimemio_flash_io2_oeb
  PIN spimemio_flash_io3_di
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END spimemio_flash_io3_di
  PIN spimemio_flash_io3_do
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END spimemio_flash_io3_do
  PIN spimemio_flash_io3_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.960 4.000 540.560 ;
    END
  END spimemio_flash_io3_oeb
  PIN trap
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END trap
  PIN uart_enabled
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END uart_enabled
  PIN user_clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END user_clock
  PIN usr1_vcc_pwrgood
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 546.950 203.230 550.950 ;
    END
  END usr1_vcc_pwrgood
  PIN usr1_vdd_pwrgood
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 546.950 208.750 550.950 ;
    END
  END usr1_vdd_pwrgood
  PIN usr2_vcc_pwrgood
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 546.950 205.990 550.950 ;
    END
  END usr2_vcc_pwrgood
  PIN usr2_vdd_pwrgood
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 546.950 211.510 550.950 ;
    END
  END usr2_vdd_pwrgood
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 546.950 10.030 550.950 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 546.950 37.630 550.950 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 546.950 40.390 550.950 ;
    END
  END wb_adr_i[11]
  PIN wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 546.950 43.150 550.950 ;
    END
  END wb_adr_i[12]
  PIN wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 546.950 45.910 550.950 ;
    END
  END wb_adr_i[13]
  PIN wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 546.950 48.670 550.950 ;
    END
  END wb_adr_i[14]
  PIN wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 546.950 51.430 550.950 ;
    END
  END wb_adr_i[15]
  PIN wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 546.950 54.190 550.950 ;
    END
  END wb_adr_i[16]
  PIN wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 546.950 56.950 550.950 ;
    END
  END wb_adr_i[17]
  PIN wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 546.950 59.710 550.950 ;
    END
  END wb_adr_i[18]
  PIN wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 546.950 62.470 550.950 ;
    END
  END wb_adr_i[19]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 546.950 12.790 550.950 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 546.950 65.230 550.950 ;
    END
  END wb_adr_i[20]
  PIN wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 546.950 67.990 550.950 ;
    END
  END wb_adr_i[21]
  PIN wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 546.950 70.750 550.950 ;
    END
  END wb_adr_i[22]
  PIN wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 546.950 73.510 550.950 ;
    END
  END wb_adr_i[23]
  PIN wb_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 546.950 76.270 550.950 ;
    END
  END wb_adr_i[24]
  PIN wb_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 546.950 79.030 550.950 ;
    END
  END wb_adr_i[25]
  PIN wb_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 546.950 81.790 550.950 ;
    END
  END wb_adr_i[26]
  PIN wb_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 546.950 84.550 550.950 ;
    END
  END wb_adr_i[27]
  PIN wb_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 546.950 87.310 550.950 ;
    END
  END wb_adr_i[28]
  PIN wb_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 546.950 90.070 550.950 ;
    END
  END wb_adr_i[29]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 546.950 15.550 550.950 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 546.950 92.830 550.950 ;
    END
  END wb_adr_i[30]
  PIN wb_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 546.950 95.590 550.950 ;
    END
  END wb_adr_i[31]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 546.950 18.310 550.950 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 546.950 21.070 550.950 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 546.950 23.830 550.950 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 546.950 26.590 550.950 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 546.950 29.350 550.950 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 546.950 32.110 550.950 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 546.950 34.870 550.950 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 546.950 200.470 550.950 ;
    END
  END wb_cyc_i
  PIN wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 546.950 98.350 550.950 ;
    END
  END wb_dat_i[0]
  PIN wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 546.950 125.950 550.950 ;
    END
  END wb_dat_i[10]
  PIN wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 546.950 128.710 550.950 ;
    END
  END wb_dat_i[11]
  PIN wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 546.950 131.470 550.950 ;
    END
  END wb_dat_i[12]
  PIN wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 546.950 134.230 550.950 ;
    END
  END wb_dat_i[13]
  PIN wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 546.950 136.990 550.950 ;
    END
  END wb_dat_i[14]
  PIN wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 546.950 139.750 550.950 ;
    END
  END wb_dat_i[15]
  PIN wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 546.950 142.510 550.950 ;
    END
  END wb_dat_i[16]
  PIN wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 546.950 145.270 550.950 ;
    END
  END wb_dat_i[17]
  PIN wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 546.950 148.030 550.950 ;
    END
  END wb_dat_i[18]
  PIN wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 546.950 150.790 550.950 ;
    END
  END wb_dat_i[19]
  PIN wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 546.950 101.110 550.950 ;
    END
  END wb_dat_i[1]
  PIN wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 546.950 153.550 550.950 ;
    END
  END wb_dat_i[20]
  PIN wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 546.950 156.310 550.950 ;
    END
  END wb_dat_i[21]
  PIN wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 546.950 159.070 550.950 ;
    END
  END wb_dat_i[22]
  PIN wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 546.950 161.830 550.950 ;
    END
  END wb_dat_i[23]
  PIN wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 546.950 164.590 550.950 ;
    END
  END wb_dat_i[24]
  PIN wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 546.950 167.350 550.950 ;
    END
  END wb_dat_i[25]
  PIN wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 546.950 170.110 550.950 ;
    END
  END wb_dat_i[26]
  PIN wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 546.950 172.870 550.950 ;
    END
  END wb_dat_i[27]
  PIN wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 546.950 175.630 550.950 ;
    END
  END wb_dat_i[28]
  PIN wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 546.950 178.390 550.950 ;
    END
  END wb_dat_i[29]
  PIN wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 546.950 103.870 550.950 ;
    END
  END wb_dat_i[2]
  PIN wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 546.950 181.150 550.950 ;
    END
  END wb_dat_i[30]
  PIN wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 546.950 183.910 550.950 ;
    END
  END wb_dat_i[31]
  PIN wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 546.950 106.630 550.950 ;
    END
  END wb_dat_i[3]
  PIN wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 546.950 109.390 550.950 ;
    END
  END wb_dat_i[4]
  PIN wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 546.950 112.150 550.950 ;
    END
  END wb_dat_i[5]
  PIN wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 546.950 114.910 550.950 ;
    END
  END wb_dat_i[6]
  PIN wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 546.950 117.670 550.950 ;
    END
  END wb_dat_i[7]
  PIN wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 546.950 120.430 550.950 ;
    END
  END wb_dat_i[8]
  PIN wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 546.950 123.190 550.950 ;
    END
  END wb_dat_i[9]
  PIN wb_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END wb_dat_o[0]
  PIN wb_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END wb_dat_o[10]
  PIN wb_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END wb_dat_o[11]
  PIN wb_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END wb_dat_o[12]
  PIN wb_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END wb_dat_o[13]
  PIN wb_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END wb_dat_o[14]
  PIN wb_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END wb_dat_o[15]
  PIN wb_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END wb_dat_o[16]
  PIN wb_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END wb_dat_o[17]
  PIN wb_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END wb_dat_o[18]
  PIN wb_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END wb_dat_o[19]
  PIN wb_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END wb_dat_o[1]
  PIN wb_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END wb_dat_o[20]
  PIN wb_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END wb_dat_o[21]
  PIN wb_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END wb_dat_o[22]
  PIN wb_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END wb_dat_o[23]
  PIN wb_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END wb_dat_o[24]
  PIN wb_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END wb_dat_o[25]
  PIN wb_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END wb_dat_o[26]
  PIN wb_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END wb_dat_o[27]
  PIN wb_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END wb_dat_o[28]
  PIN wb_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 4.000 410.000 ;
    END
  END wb_dat_o[29]
  PIN wb_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END wb_dat_o[2]
  PIN wb_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END wb_dat_o[30]
  PIN wb_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END wb_dat_o[31]
  PIN wb_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END wb_dat_o[3]
  PIN wb_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END wb_dat_o[4]
  PIN wb_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END wb_dat_o[5]
  PIN wb_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END wb_dat_o[6]
  PIN wb_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END wb_dat_o[7]
  PIN wb_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END wb_dat_o[8]
  PIN wb_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END wb_dat_o[9]
  PIN wb_rstn_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END wb_rstn_i
  PIN wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 546.950 186.670 550.950 ;
    END
  END wb_sel_i[0]
  PIN wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 546.950 189.430 550.950 ;
    END
  END wb_sel_i[1]
  PIN wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 546.950 192.190 550.950 ;
    END
  END wb_sel_i[2]
  PIN wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 546.950 194.950 550.950 ;
    END
  END wb_sel_i[3]
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 546.950 197.710 550.950 ;
    END
  END wb_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 364.320 538.645 ;
      LAYER met1 ;
        RECT 5.130 6.160 367.930 542.260 ;
      LAYER met2 ;
        RECT 5.160 546.670 9.470 547.130 ;
        RECT 10.310 546.670 12.230 547.130 ;
        RECT 13.070 546.670 14.990 547.130 ;
        RECT 15.830 546.670 17.750 547.130 ;
        RECT 18.590 546.670 20.510 547.130 ;
        RECT 21.350 546.670 23.270 547.130 ;
        RECT 24.110 546.670 26.030 547.130 ;
        RECT 26.870 546.670 28.790 547.130 ;
        RECT 29.630 546.670 31.550 547.130 ;
        RECT 32.390 546.670 34.310 547.130 ;
        RECT 35.150 546.670 37.070 547.130 ;
        RECT 37.910 546.670 39.830 547.130 ;
        RECT 40.670 546.670 42.590 547.130 ;
        RECT 43.430 546.670 45.350 547.130 ;
        RECT 46.190 546.670 48.110 547.130 ;
        RECT 48.950 546.670 50.870 547.130 ;
        RECT 51.710 546.670 53.630 547.130 ;
        RECT 54.470 546.670 56.390 547.130 ;
        RECT 57.230 546.670 59.150 547.130 ;
        RECT 59.990 546.670 61.910 547.130 ;
        RECT 62.750 546.670 64.670 547.130 ;
        RECT 65.510 546.670 67.430 547.130 ;
        RECT 68.270 546.670 70.190 547.130 ;
        RECT 71.030 546.670 72.950 547.130 ;
        RECT 73.790 546.670 75.710 547.130 ;
        RECT 76.550 546.670 78.470 547.130 ;
        RECT 79.310 546.670 81.230 547.130 ;
        RECT 82.070 546.670 83.990 547.130 ;
        RECT 84.830 546.670 86.750 547.130 ;
        RECT 87.590 546.670 89.510 547.130 ;
        RECT 90.350 546.670 92.270 547.130 ;
        RECT 93.110 546.670 95.030 547.130 ;
        RECT 95.870 546.670 97.790 547.130 ;
        RECT 98.630 546.670 100.550 547.130 ;
        RECT 101.390 546.670 103.310 547.130 ;
        RECT 104.150 546.670 106.070 547.130 ;
        RECT 106.910 546.670 108.830 547.130 ;
        RECT 109.670 546.670 111.590 547.130 ;
        RECT 112.430 546.670 114.350 547.130 ;
        RECT 115.190 546.670 117.110 547.130 ;
        RECT 117.950 546.670 119.870 547.130 ;
        RECT 120.710 546.670 122.630 547.130 ;
        RECT 123.470 546.670 125.390 547.130 ;
        RECT 126.230 546.670 128.150 547.130 ;
        RECT 128.990 546.670 130.910 547.130 ;
        RECT 131.750 546.670 133.670 547.130 ;
        RECT 134.510 546.670 136.430 547.130 ;
        RECT 137.270 546.670 139.190 547.130 ;
        RECT 140.030 546.670 141.950 547.130 ;
        RECT 142.790 546.670 144.710 547.130 ;
        RECT 145.550 546.670 147.470 547.130 ;
        RECT 148.310 546.670 150.230 547.130 ;
        RECT 151.070 546.670 152.990 547.130 ;
        RECT 153.830 546.670 155.750 547.130 ;
        RECT 156.590 546.670 158.510 547.130 ;
        RECT 159.350 546.670 161.270 547.130 ;
        RECT 162.110 546.670 164.030 547.130 ;
        RECT 164.870 546.670 166.790 547.130 ;
        RECT 167.630 546.670 169.550 547.130 ;
        RECT 170.390 546.670 172.310 547.130 ;
        RECT 173.150 546.670 175.070 547.130 ;
        RECT 175.910 546.670 177.830 547.130 ;
        RECT 178.670 546.670 180.590 547.130 ;
        RECT 181.430 546.670 183.350 547.130 ;
        RECT 184.190 546.670 186.110 547.130 ;
        RECT 186.950 546.670 188.870 547.130 ;
        RECT 189.710 546.670 191.630 547.130 ;
        RECT 192.470 546.670 194.390 547.130 ;
        RECT 195.230 546.670 197.150 547.130 ;
        RECT 197.990 546.670 199.910 547.130 ;
        RECT 200.750 546.670 202.670 547.130 ;
        RECT 203.510 546.670 205.430 547.130 ;
        RECT 206.270 546.670 208.190 547.130 ;
        RECT 209.030 546.670 210.950 547.130 ;
        RECT 211.790 546.670 213.710 547.130 ;
        RECT 214.550 546.670 216.470 547.130 ;
        RECT 217.310 546.670 219.230 547.130 ;
        RECT 220.070 546.670 221.990 547.130 ;
        RECT 222.830 546.670 224.750 547.130 ;
        RECT 225.590 546.670 227.510 547.130 ;
        RECT 228.350 546.670 230.270 547.130 ;
        RECT 231.110 546.670 233.030 547.130 ;
        RECT 233.870 546.670 235.790 547.130 ;
        RECT 236.630 546.670 238.550 547.130 ;
        RECT 239.390 546.670 241.310 547.130 ;
        RECT 242.150 546.670 244.070 547.130 ;
        RECT 244.910 546.670 246.830 547.130 ;
        RECT 247.670 546.670 249.590 547.130 ;
        RECT 250.430 546.670 252.350 547.130 ;
        RECT 253.190 546.670 255.110 547.130 ;
        RECT 255.950 546.670 257.870 547.130 ;
        RECT 258.710 546.670 260.630 547.130 ;
        RECT 261.470 546.670 263.390 547.130 ;
        RECT 264.230 546.670 266.150 547.130 ;
        RECT 266.990 546.670 268.910 547.130 ;
        RECT 269.750 546.670 271.670 547.130 ;
        RECT 272.510 546.670 274.430 547.130 ;
        RECT 275.270 546.670 277.190 547.130 ;
        RECT 278.030 546.670 279.950 547.130 ;
        RECT 280.790 546.670 282.710 547.130 ;
        RECT 283.550 546.670 285.470 547.130 ;
        RECT 286.310 546.670 288.230 547.130 ;
        RECT 289.070 546.670 290.990 547.130 ;
        RECT 291.830 546.670 293.750 547.130 ;
        RECT 294.590 546.670 296.510 547.130 ;
        RECT 297.350 546.670 299.270 547.130 ;
        RECT 300.110 546.670 302.030 547.130 ;
        RECT 302.870 546.670 304.790 547.130 ;
        RECT 305.630 546.670 307.550 547.130 ;
        RECT 308.390 546.670 310.310 547.130 ;
        RECT 311.150 546.670 313.070 547.130 ;
        RECT 313.910 546.670 315.830 547.130 ;
        RECT 316.670 546.670 318.590 547.130 ;
        RECT 319.430 546.670 321.350 547.130 ;
        RECT 322.190 546.670 324.110 547.130 ;
        RECT 324.950 546.670 326.870 547.130 ;
        RECT 327.710 546.670 329.630 547.130 ;
        RECT 330.470 546.670 332.390 547.130 ;
        RECT 333.230 546.670 335.150 547.130 ;
        RECT 335.990 546.670 337.910 547.130 ;
        RECT 338.750 546.670 340.670 547.130 ;
        RECT 341.510 546.670 343.430 547.130 ;
        RECT 344.270 546.670 346.190 547.130 ;
        RECT 347.030 546.670 348.950 547.130 ;
        RECT 349.790 546.670 351.710 547.130 ;
        RECT 352.550 546.670 354.470 547.130 ;
        RECT 355.310 546.670 357.230 547.130 ;
        RECT 358.070 546.670 359.990 547.130 ;
        RECT 360.830 546.670 367.900 547.130 ;
        RECT 5.160 4.280 367.900 546.670 ;
        RECT 5.160 3.670 15.450 4.280 ;
        RECT 16.290 3.670 19.130 4.280 ;
        RECT 19.970 3.670 22.810 4.280 ;
        RECT 23.650 3.670 26.490 4.280 ;
        RECT 27.330 3.670 30.170 4.280 ;
        RECT 31.010 3.670 33.850 4.280 ;
        RECT 34.690 3.670 37.530 4.280 ;
        RECT 38.370 3.670 41.210 4.280 ;
        RECT 42.050 3.670 44.890 4.280 ;
        RECT 45.730 3.670 48.570 4.280 ;
        RECT 49.410 3.670 52.250 4.280 ;
        RECT 53.090 3.670 55.930 4.280 ;
        RECT 56.770 3.670 59.610 4.280 ;
        RECT 60.450 3.670 63.290 4.280 ;
        RECT 64.130 3.670 66.970 4.280 ;
        RECT 67.810 3.670 70.650 4.280 ;
        RECT 71.490 3.670 74.330 4.280 ;
        RECT 75.170 3.670 78.010 4.280 ;
        RECT 78.850 3.670 81.690 4.280 ;
        RECT 82.530 3.670 85.370 4.280 ;
        RECT 86.210 3.670 89.050 4.280 ;
        RECT 89.890 3.670 92.730 4.280 ;
        RECT 93.570 3.670 96.410 4.280 ;
        RECT 97.250 3.670 100.090 4.280 ;
        RECT 100.930 3.670 103.770 4.280 ;
        RECT 104.610 3.670 107.450 4.280 ;
        RECT 108.290 3.670 111.130 4.280 ;
        RECT 111.970 3.670 114.810 4.280 ;
        RECT 115.650 3.670 118.490 4.280 ;
        RECT 119.330 3.670 122.170 4.280 ;
        RECT 123.010 3.670 125.850 4.280 ;
        RECT 126.690 3.670 129.530 4.280 ;
        RECT 130.370 3.670 133.210 4.280 ;
        RECT 134.050 3.670 136.890 4.280 ;
        RECT 137.730 3.670 140.570 4.280 ;
        RECT 141.410 3.670 144.250 4.280 ;
        RECT 145.090 3.670 147.930 4.280 ;
        RECT 148.770 3.670 151.610 4.280 ;
        RECT 152.450 3.670 155.290 4.280 ;
        RECT 156.130 3.670 158.970 4.280 ;
        RECT 159.810 3.670 162.650 4.280 ;
        RECT 163.490 3.670 166.330 4.280 ;
        RECT 167.170 3.670 170.010 4.280 ;
        RECT 170.850 3.670 173.690 4.280 ;
        RECT 174.530 3.670 177.370 4.280 ;
        RECT 178.210 3.670 181.050 4.280 ;
        RECT 181.890 3.670 184.730 4.280 ;
        RECT 185.570 3.670 188.410 4.280 ;
        RECT 189.250 3.670 192.090 4.280 ;
        RECT 192.930 3.670 195.770 4.280 ;
        RECT 196.610 3.670 199.450 4.280 ;
        RECT 200.290 3.670 203.130 4.280 ;
        RECT 203.970 3.670 206.810 4.280 ;
        RECT 207.650 3.670 210.490 4.280 ;
        RECT 211.330 3.670 214.170 4.280 ;
        RECT 215.010 3.670 217.850 4.280 ;
        RECT 218.690 3.670 221.530 4.280 ;
        RECT 222.370 3.670 225.210 4.280 ;
        RECT 226.050 3.670 228.890 4.280 ;
        RECT 229.730 3.670 232.570 4.280 ;
        RECT 233.410 3.670 236.250 4.280 ;
        RECT 237.090 3.670 239.930 4.280 ;
        RECT 240.770 3.670 243.610 4.280 ;
        RECT 244.450 3.670 247.290 4.280 ;
        RECT 248.130 3.670 250.970 4.280 ;
        RECT 251.810 3.670 254.650 4.280 ;
        RECT 255.490 3.670 258.330 4.280 ;
        RECT 259.170 3.670 262.010 4.280 ;
        RECT 262.850 3.670 265.690 4.280 ;
        RECT 266.530 3.670 269.370 4.280 ;
        RECT 270.210 3.670 273.050 4.280 ;
        RECT 273.890 3.670 276.730 4.280 ;
        RECT 277.570 3.670 280.410 4.280 ;
        RECT 281.250 3.670 284.090 4.280 ;
        RECT 284.930 3.670 287.770 4.280 ;
        RECT 288.610 3.670 291.450 4.280 ;
        RECT 292.290 3.670 295.130 4.280 ;
        RECT 295.970 3.670 298.810 4.280 ;
        RECT 299.650 3.670 302.490 4.280 ;
        RECT 303.330 3.670 306.170 4.280 ;
        RECT 307.010 3.670 309.850 4.280 ;
        RECT 310.690 3.670 313.530 4.280 ;
        RECT 314.370 3.670 317.210 4.280 ;
        RECT 318.050 3.670 320.890 4.280 ;
        RECT 321.730 3.670 324.570 4.280 ;
        RECT 325.410 3.670 328.250 4.280 ;
        RECT 329.090 3.670 331.930 4.280 ;
        RECT 332.770 3.670 335.610 4.280 ;
        RECT 336.450 3.670 339.290 4.280 ;
        RECT 340.130 3.670 342.970 4.280 ;
        RECT 343.810 3.670 346.650 4.280 ;
        RECT 347.490 3.670 350.330 4.280 ;
        RECT 351.170 3.670 354.010 4.280 ;
        RECT 354.850 3.670 367.900 4.280 ;
      LAYER met3 ;
        RECT 4.400 539.560 367.015 540.425 ;
        RECT 4.000 536.880 367.015 539.560 ;
        RECT 4.000 535.480 365.830 536.880 ;
        RECT 4.000 532.800 367.015 535.480 ;
        RECT 4.400 531.400 367.015 532.800 ;
        RECT 4.000 528.720 367.015 531.400 ;
        RECT 4.000 527.320 365.830 528.720 ;
        RECT 4.000 524.640 367.015 527.320 ;
        RECT 4.400 523.240 367.015 524.640 ;
        RECT 4.000 520.560 367.015 523.240 ;
        RECT 4.000 519.160 365.830 520.560 ;
        RECT 4.000 516.480 367.015 519.160 ;
        RECT 4.400 515.080 367.015 516.480 ;
        RECT 4.000 512.400 367.015 515.080 ;
        RECT 4.000 511.000 365.830 512.400 ;
        RECT 4.000 508.320 367.015 511.000 ;
        RECT 4.400 506.920 367.015 508.320 ;
        RECT 4.000 504.240 367.015 506.920 ;
        RECT 4.000 502.840 365.830 504.240 ;
        RECT 4.000 500.160 367.015 502.840 ;
        RECT 4.400 498.760 367.015 500.160 ;
        RECT 4.000 496.080 367.015 498.760 ;
        RECT 4.000 494.680 365.830 496.080 ;
        RECT 4.000 492.000 367.015 494.680 ;
        RECT 4.400 490.600 367.015 492.000 ;
        RECT 4.000 487.920 367.015 490.600 ;
        RECT 4.000 486.520 365.830 487.920 ;
        RECT 4.000 483.840 367.015 486.520 ;
        RECT 4.400 482.440 367.015 483.840 ;
        RECT 4.000 479.760 367.015 482.440 ;
        RECT 4.000 478.360 365.830 479.760 ;
        RECT 4.000 475.680 367.015 478.360 ;
        RECT 4.400 474.280 367.015 475.680 ;
        RECT 4.000 471.600 367.015 474.280 ;
        RECT 4.000 470.200 365.830 471.600 ;
        RECT 4.000 467.520 367.015 470.200 ;
        RECT 4.400 466.120 367.015 467.520 ;
        RECT 4.000 463.440 367.015 466.120 ;
        RECT 4.000 462.040 365.830 463.440 ;
        RECT 4.000 459.360 367.015 462.040 ;
        RECT 4.400 457.960 367.015 459.360 ;
        RECT 4.000 455.280 367.015 457.960 ;
        RECT 4.000 453.880 365.830 455.280 ;
        RECT 4.000 451.200 367.015 453.880 ;
        RECT 4.400 449.800 367.015 451.200 ;
        RECT 4.000 447.120 367.015 449.800 ;
        RECT 4.000 445.720 365.830 447.120 ;
        RECT 4.000 443.040 367.015 445.720 ;
        RECT 4.400 441.640 367.015 443.040 ;
        RECT 4.000 438.960 367.015 441.640 ;
        RECT 4.000 437.560 365.830 438.960 ;
        RECT 4.000 434.880 367.015 437.560 ;
        RECT 4.400 433.480 367.015 434.880 ;
        RECT 4.000 430.800 367.015 433.480 ;
        RECT 4.000 429.400 365.830 430.800 ;
        RECT 4.000 426.720 367.015 429.400 ;
        RECT 4.400 425.320 367.015 426.720 ;
        RECT 4.000 422.640 367.015 425.320 ;
        RECT 4.000 421.240 365.830 422.640 ;
        RECT 4.000 418.560 367.015 421.240 ;
        RECT 4.400 417.160 367.015 418.560 ;
        RECT 4.000 414.480 367.015 417.160 ;
        RECT 4.000 413.080 365.830 414.480 ;
        RECT 4.000 410.400 367.015 413.080 ;
        RECT 4.400 409.000 367.015 410.400 ;
        RECT 4.000 406.320 367.015 409.000 ;
        RECT 4.000 404.920 365.830 406.320 ;
        RECT 4.000 402.240 367.015 404.920 ;
        RECT 4.400 400.840 367.015 402.240 ;
        RECT 4.000 398.160 367.015 400.840 ;
        RECT 4.000 396.760 365.830 398.160 ;
        RECT 4.000 394.080 367.015 396.760 ;
        RECT 4.400 392.680 367.015 394.080 ;
        RECT 4.000 390.000 367.015 392.680 ;
        RECT 4.000 388.600 365.830 390.000 ;
        RECT 4.000 385.920 367.015 388.600 ;
        RECT 4.400 384.520 367.015 385.920 ;
        RECT 4.000 381.840 367.015 384.520 ;
        RECT 4.000 380.440 365.830 381.840 ;
        RECT 4.000 377.760 367.015 380.440 ;
        RECT 4.400 376.360 367.015 377.760 ;
        RECT 4.000 373.680 367.015 376.360 ;
        RECT 4.000 372.280 365.830 373.680 ;
        RECT 4.000 369.600 367.015 372.280 ;
        RECT 4.400 368.200 367.015 369.600 ;
        RECT 4.000 365.520 367.015 368.200 ;
        RECT 4.000 364.120 365.830 365.520 ;
        RECT 4.000 361.440 367.015 364.120 ;
        RECT 4.400 360.040 367.015 361.440 ;
        RECT 4.000 357.360 367.015 360.040 ;
        RECT 4.000 355.960 365.830 357.360 ;
        RECT 4.000 353.280 367.015 355.960 ;
        RECT 4.400 351.880 367.015 353.280 ;
        RECT 4.000 349.200 367.015 351.880 ;
        RECT 4.000 347.800 365.830 349.200 ;
        RECT 4.000 345.120 367.015 347.800 ;
        RECT 4.400 343.720 367.015 345.120 ;
        RECT 4.000 341.040 367.015 343.720 ;
        RECT 4.000 339.640 365.830 341.040 ;
        RECT 4.000 336.960 367.015 339.640 ;
        RECT 4.400 335.560 367.015 336.960 ;
        RECT 4.000 332.880 367.015 335.560 ;
        RECT 4.000 331.480 365.830 332.880 ;
        RECT 4.000 328.800 367.015 331.480 ;
        RECT 4.400 327.400 367.015 328.800 ;
        RECT 4.000 324.720 367.015 327.400 ;
        RECT 4.000 323.320 365.830 324.720 ;
        RECT 4.000 320.640 367.015 323.320 ;
        RECT 4.400 319.240 367.015 320.640 ;
        RECT 4.000 316.560 367.015 319.240 ;
        RECT 4.000 315.160 365.830 316.560 ;
        RECT 4.000 312.480 367.015 315.160 ;
        RECT 4.400 311.080 367.015 312.480 ;
        RECT 4.000 308.400 367.015 311.080 ;
        RECT 4.000 307.000 365.830 308.400 ;
        RECT 4.000 304.320 367.015 307.000 ;
        RECT 4.400 302.920 367.015 304.320 ;
        RECT 4.000 300.240 367.015 302.920 ;
        RECT 4.000 298.840 365.830 300.240 ;
        RECT 4.000 296.160 367.015 298.840 ;
        RECT 4.400 294.760 367.015 296.160 ;
        RECT 4.000 292.080 367.015 294.760 ;
        RECT 4.000 290.680 365.830 292.080 ;
        RECT 4.000 288.000 367.015 290.680 ;
        RECT 4.400 286.600 367.015 288.000 ;
        RECT 4.000 283.920 367.015 286.600 ;
        RECT 4.000 282.520 365.830 283.920 ;
        RECT 4.000 279.840 367.015 282.520 ;
        RECT 4.400 278.440 367.015 279.840 ;
        RECT 4.000 275.760 367.015 278.440 ;
        RECT 4.000 274.360 365.830 275.760 ;
        RECT 4.000 271.680 367.015 274.360 ;
        RECT 4.400 270.280 367.015 271.680 ;
        RECT 4.000 267.600 367.015 270.280 ;
        RECT 4.000 266.200 365.830 267.600 ;
        RECT 4.000 263.520 367.015 266.200 ;
        RECT 4.400 262.120 367.015 263.520 ;
        RECT 4.000 259.440 367.015 262.120 ;
        RECT 4.000 258.040 365.830 259.440 ;
        RECT 4.000 255.360 367.015 258.040 ;
        RECT 4.400 253.960 367.015 255.360 ;
        RECT 4.000 251.280 367.015 253.960 ;
        RECT 4.000 249.880 365.830 251.280 ;
        RECT 4.000 247.200 367.015 249.880 ;
        RECT 4.400 245.800 367.015 247.200 ;
        RECT 4.000 243.120 367.015 245.800 ;
        RECT 4.000 241.720 365.830 243.120 ;
        RECT 4.000 239.040 367.015 241.720 ;
        RECT 4.400 237.640 367.015 239.040 ;
        RECT 4.000 234.960 367.015 237.640 ;
        RECT 4.000 233.560 365.830 234.960 ;
        RECT 4.000 230.880 367.015 233.560 ;
        RECT 4.400 229.480 367.015 230.880 ;
        RECT 4.000 226.800 367.015 229.480 ;
        RECT 4.000 225.400 365.830 226.800 ;
        RECT 4.000 222.720 367.015 225.400 ;
        RECT 4.400 221.320 367.015 222.720 ;
        RECT 4.000 218.640 367.015 221.320 ;
        RECT 4.000 217.240 365.830 218.640 ;
        RECT 4.000 214.560 367.015 217.240 ;
        RECT 4.400 213.160 367.015 214.560 ;
        RECT 4.000 210.480 367.015 213.160 ;
        RECT 4.000 209.080 365.830 210.480 ;
        RECT 4.000 206.400 367.015 209.080 ;
        RECT 4.400 205.000 367.015 206.400 ;
        RECT 4.000 202.320 367.015 205.000 ;
        RECT 4.000 200.920 365.830 202.320 ;
        RECT 4.000 198.240 367.015 200.920 ;
        RECT 4.400 196.840 367.015 198.240 ;
        RECT 4.000 194.160 367.015 196.840 ;
        RECT 4.000 192.760 365.830 194.160 ;
        RECT 4.000 190.080 367.015 192.760 ;
        RECT 4.400 188.680 367.015 190.080 ;
        RECT 4.000 186.000 367.015 188.680 ;
        RECT 4.000 184.600 365.830 186.000 ;
        RECT 4.000 181.920 367.015 184.600 ;
        RECT 4.400 180.520 367.015 181.920 ;
        RECT 4.000 177.840 367.015 180.520 ;
        RECT 4.000 176.440 365.830 177.840 ;
        RECT 4.000 173.760 367.015 176.440 ;
        RECT 4.400 172.360 367.015 173.760 ;
        RECT 4.000 169.680 367.015 172.360 ;
        RECT 4.000 168.280 365.830 169.680 ;
        RECT 4.000 165.600 367.015 168.280 ;
        RECT 4.400 164.200 367.015 165.600 ;
        RECT 4.000 161.520 367.015 164.200 ;
        RECT 4.000 160.120 365.830 161.520 ;
        RECT 4.000 157.440 367.015 160.120 ;
        RECT 4.400 156.040 367.015 157.440 ;
        RECT 4.000 153.360 367.015 156.040 ;
        RECT 4.000 151.960 365.830 153.360 ;
        RECT 4.000 149.280 367.015 151.960 ;
        RECT 4.400 147.880 367.015 149.280 ;
        RECT 4.000 145.200 367.015 147.880 ;
        RECT 4.000 143.800 365.830 145.200 ;
        RECT 4.000 141.120 367.015 143.800 ;
        RECT 4.400 139.720 367.015 141.120 ;
        RECT 4.000 137.040 367.015 139.720 ;
        RECT 4.000 135.640 365.830 137.040 ;
        RECT 4.000 132.960 367.015 135.640 ;
        RECT 4.400 131.560 367.015 132.960 ;
        RECT 4.000 128.880 367.015 131.560 ;
        RECT 4.000 127.480 365.830 128.880 ;
        RECT 4.000 124.800 367.015 127.480 ;
        RECT 4.400 123.400 367.015 124.800 ;
        RECT 4.000 120.720 367.015 123.400 ;
        RECT 4.000 119.320 365.830 120.720 ;
        RECT 4.000 116.640 367.015 119.320 ;
        RECT 4.400 115.240 367.015 116.640 ;
        RECT 4.000 112.560 367.015 115.240 ;
        RECT 4.000 111.160 365.830 112.560 ;
        RECT 4.000 108.480 367.015 111.160 ;
        RECT 4.400 107.080 367.015 108.480 ;
        RECT 4.000 104.400 367.015 107.080 ;
        RECT 4.000 103.000 365.830 104.400 ;
        RECT 4.000 100.320 367.015 103.000 ;
        RECT 4.400 98.920 367.015 100.320 ;
        RECT 4.000 96.240 367.015 98.920 ;
        RECT 4.000 94.840 365.830 96.240 ;
        RECT 4.000 92.160 367.015 94.840 ;
        RECT 4.400 90.760 367.015 92.160 ;
        RECT 4.000 88.080 367.015 90.760 ;
        RECT 4.000 86.680 365.830 88.080 ;
        RECT 4.000 84.000 367.015 86.680 ;
        RECT 4.400 82.600 367.015 84.000 ;
        RECT 4.000 79.920 367.015 82.600 ;
        RECT 4.000 78.520 365.830 79.920 ;
        RECT 4.000 75.840 367.015 78.520 ;
        RECT 4.400 74.440 367.015 75.840 ;
        RECT 4.000 71.760 367.015 74.440 ;
        RECT 4.000 70.360 365.830 71.760 ;
        RECT 4.000 67.680 367.015 70.360 ;
        RECT 4.400 66.280 367.015 67.680 ;
        RECT 4.000 63.600 367.015 66.280 ;
        RECT 4.000 62.200 365.830 63.600 ;
        RECT 4.000 59.520 367.015 62.200 ;
        RECT 4.400 58.120 367.015 59.520 ;
        RECT 4.000 55.440 367.015 58.120 ;
        RECT 4.000 54.040 365.830 55.440 ;
        RECT 4.000 51.360 367.015 54.040 ;
        RECT 4.400 49.960 367.015 51.360 ;
        RECT 4.000 47.280 367.015 49.960 ;
        RECT 4.000 45.880 365.830 47.280 ;
        RECT 4.000 43.200 367.015 45.880 ;
        RECT 4.400 41.800 367.015 43.200 ;
        RECT 4.000 39.120 367.015 41.800 ;
        RECT 4.000 37.720 365.830 39.120 ;
        RECT 4.000 35.040 367.015 37.720 ;
        RECT 4.400 33.640 367.015 35.040 ;
        RECT 4.000 30.960 367.015 33.640 ;
        RECT 4.000 29.560 365.830 30.960 ;
        RECT 4.000 26.880 367.015 29.560 ;
        RECT 4.400 25.480 367.015 26.880 ;
        RECT 4.000 22.800 367.015 25.480 ;
        RECT 4.000 21.400 365.830 22.800 ;
        RECT 4.000 18.720 367.015 21.400 ;
        RECT 4.400 17.320 367.015 18.720 ;
        RECT 4.000 14.640 367.015 17.320 ;
        RECT 4.000 13.240 365.830 14.640 ;
        RECT 4.000 10.560 367.015 13.240 ;
        RECT 4.400 9.695 367.015 10.560 ;
      LAYER met4 ;
        RECT 13.175 34.855 20.640 531.585 ;
        RECT 23.040 34.855 23.940 531.585 ;
        RECT 26.340 34.855 174.240 531.585 ;
        RECT 176.640 34.855 177.540 531.585 ;
        RECT 179.940 34.855 327.840 531.585 ;
        RECT 330.240 34.855 331.140 531.585 ;
        RECT 333.540 34.855 359.425 531.585 ;
      LAYER met5 ;
        RECT 130.300 272.900 346.260 288.100 ;
  END
END housekeeping
END LIBRARY

