magic
tech sky130A
magscale 1 2
timestamp 1686190293
<< checkpaint >>
rect 40504 1532674 43088 1535246
rect 40504 1443474 43088 1446046
rect 40504 1354274 43088 1356846
rect 40504 1309274 43088 1311846
rect 40504 1264274 43088 1266846
rect 40504 1219074 43088 1221646
rect 40504 1174074 43088 1176646
rect 40504 1128874 43088 1131446
rect -1260 -1260 718860 1038860
rect 674512 -42446 677096 -39874
rect 674512 -170046 677096 -167474
rect 674512 -213246 677096 -210674
rect 674512 -256446 677096 -253874
rect 674512 -299646 677096 -297074
rect 674512 -342846 677096 -340274
rect 674512 -386046 677096 -383474
<< error_p >>
rect 149223 18082 150855 18116
<< metal5 >>
rect 78440 1018512 90960 1031002
rect 129840 1018512 142360 1031002
rect 181240 1018512 193760 1031002
rect 232640 1018512 245160 1031002
rect 284240 1018512 296760 1031002
rect 334810 1018624 346978 1030788
rect 386040 1018512 398560 1031002
rect 475040 1018512 487560 1031002
rect 526440 1018512 538960 1031002
rect 577010 1018624 589178 1030788
rect 628240 1018512 640760 1031002
rect 6598 956440 19088 968960
rect 698512 952840 711002 965360
rect 6167 914054 19619 924934
rect 697980 909666 711432 920546
rect 6811 871210 18975 883378
rect 698512 863640 711002 876160
rect 6811 829010 18975 841178
rect 698624 819822 710788 831990
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 698624 505222 710788 517390
rect 6811 484410 18975 496578
rect 697980 461866 711432 472746
rect 6167 442854 19619 453734
rect 698624 417022 710788 429190
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6811 111610 18975 123778
rect 698512 101240 711002 113760
rect 6167 70054 19619 80934
rect 80222 6811 92390 18975
rect 136713 7143 144149 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19619
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18975
rect 624222 6811 636390 18975
use chip_io_openframe  chip_io_openframe_0
timestamp 1686190293
transform 1 0 0 0 1 0
box 0 0 717600 1037600
use openframe_project_wrapper  openframe_project_wrapper_0
timestamp 1686190293
transform 1 0 42137 0 1 42137
box -444 -444 633770 953770
<< labels >>
flabel metal5 s 187640 6598 200160 19088 0 FreeSans 16000 0 0 0 gpio[38]
port 57 nsew
flabel metal5 s 296240 6598 308760 19088 0 FreeSans 16000 0 0 0 gpio[39]
port 58 nsew
flabel metal5 s 351040 6598 363560 19088 0 FreeSans 16000 0 0 0 gpio[40]
port 59 nsew
flabel metal5 s 405840 6598 418360 19088 0 FreeSans 16000 0 0 0 gpio[41]
port 60 nsew
flabel metal5 s 460640 6598 473160 19088 0 FreeSans 16000 0 0 0 gpio[42]
port 61 nsew
flabel metal5 s 515440 6598 527960 19088 0 FreeSans 16000 0 0 0 gpio[43]
port 62 nsew
flabel metal5 s 624222 6811 636390 18975 0 FreeSans 16000 0 0 0 vdda
port 5 nsew
flabel metal5 s 80222 6811 92390 18975 0 FreeSans 16000 0 0 0 vssa
port 6 nsew
flabel metal5 s 243266 6167 254146 19619 0 FreeSans 16000 0 0 0 vssd
port 8 nsew
flabel metal5 s 570422 6811 582590 18975 0 FreeSans 16000 0 0 0 vssio
port 3 nsew
flabel metal5 s 136713 7143 144149 18309 0 FreeSans 16000 0 0 0 resetb
port 63 nsew
flabel metal5 s 334810 1018624 346978 1030788 0 FreeSans 16000 0 0 0 vssio_2
port 4 nsew
flabel metal5 s 628240 1018512 640760 1031002 0 FreeSans 16000 0 0 0 gpio[15]
port 34 nsew
flabel metal5 s 526440 1018512 538960 1031002 0 FreeSans 16000 0 0 0 gpio[16]
port 35 nsew
flabel metal5 s 475040 1018512 487560 1031002 0 FreeSans 16000 0 0 0 gpio[17]
port 36 nsew
flabel metal5 s 386040 1018512 398560 1031002 0 FreeSans 16000 0 0 0 gpio[18]
port 37 nsew
flabel metal5 s 284240 1018512 296760 1031002 0 FreeSans 16000 0 0 0 gpio[19]
port 38 nsew
flabel metal5 s 232640 1018512 245160 1031002 0 FreeSans 16000 0 0 0 gpio[20]
port 39 nsew
flabel metal5 s 181240 1018512 193760 1031002 0 FreeSans 16000 0 0 0 gpio[21]
port 40 nsew
flabel metal5 s 129840 1018512 142360 1031002 0 FreeSans 16000 0 0 0 gpio[22]
port 41 nsew
flabel metal5 s 78440 1018512 90960 1031002 0 FreeSans 16000 0 0 0 gpio[23]
port 42 nsew
flabel metal5 s 577010 1018624 589178 1030788 0 FreeSans 16000 0 0 0 vssa1
port 11 nsew
flabel metal5 s 698512 684440 711002 696960 0 FreeSans 16000 0 0 0 gpio[10]
port 29 nsew
flabel metal5 s 698512 729440 711002 741960 0 FreeSans 16000 0 0 0 gpio[11]
port 30 nsew
flabel metal5 s 698512 774440 711002 786960 0 FreeSans 16000 0 0 0 gpio[12]
port 31 nsew
flabel metal5 s 698512 863640 711002 876160 0 FreeSans 16000 0 0 0 gpio[13]
port 32 nsew
flabel metal5 s 698512 146440 711002 158960 0 FreeSans 16000 0 0 0 gpio[1]
port 20 nsew
flabel metal5 s 698512 191440 711002 203960 0 FreeSans 16000 0 0 0 gpio[2]
port 21 nsew
flabel metal5 s 698512 236640 711002 249160 0 FreeSans 16000 0 0 0 gpio[3]
port 22 nsew
flabel metal5 s 698512 281640 711002 294160 0 FreeSans 16000 0 0 0 gpio[4]
port 23 nsew
flabel metal5 s 698512 326640 711002 339160 0 FreeSans 16000 0 0 0 gpio[5]
port 24 nsew
flabel metal5 s 698512 371840 711002 384360 0 FreeSans 16000 0 0 0 gpio[6]
port 25 nsew
flabel metal5 s 698512 549040 711002 561560 0 FreeSans 16000 0 0 0 gpio[7]
port 26 nsew
flabel metal5 s 698512 594240 711002 606760 0 FreeSans 16000 0 0 0 gpio[8]
port 27 nsew
flabel metal5 s 698512 639240 711002 651760 0 FreeSans 16000 0 0 0 gpio[9]
port 28 nsew
flabel metal5 s 697980 909666 711432 920546 0 FreeSans 16000 0 0 0 vccd1
port 14 nsew
flabel metal5 s 698624 819822 710788 831990 0 FreeSans 16000 0 0 0 vdda1
port 9 nsew
flabel metal5 s 698624 505222 710788 517390 0 FreeSans 16000 0 0 0 vdda1_2
port 10 nsew
flabel metal5 s 698624 417022 710788 429190 0 FreeSans 16000 0 0 0 vssa1_2
port 12 nsew
flabel metal5 s 697980 461866 711432 472746 0 FreeSans 16000 0 0 0 vssd1
port 16 nsew
flabel metal5 s 698512 101240 711002 113760 0 FreeSans 16000 0 0 0 gpio[0]
port 19 nsew
flabel metal5 s 698512 952840 711002 965360 0 FreeSans 16000 0 0 0 gpio[14]
port 33 nsew
flabel metal5 s 6167 70054 19619 80934 0 FreeSans 16000 0 0 0 vccd
port 7 nsew
flabel metal5 s 6811 111610 18975 123778 0 FreeSans 16000 0 0 0 vddio
port 1 nsew
flabel metal5 s 6811 871210 18975 883378 0 FreeSans 16000 0 0 0 vddio_2
port 2 nsew
flabel metal5 s 6598 613840 19088 626360 0 FreeSans 16000 0 0 0 gpio[29]
port 48 nsew
flabel metal5 s 6598 570640 19088 583160 0 FreeSans 16000 0 0 0 gpio[30]
port 49 nsew
flabel metal5 s 6598 527440 19088 539960 0 FreeSans 16000 0 0 0 gpio[31]
port 50 nsew
flabel metal5 s 6598 399840 19088 412360 0 FreeSans 16000 0 0 0 gpio[32]
port 51 nsew
flabel metal5 s 6598 356640 19088 369160 0 FreeSans 16000 0 0 0 gpio[33]
port 52 nsew
flabel metal5 s 6598 313440 19088 325960 0 FreeSans 16000 0 0 0 gpio[34]
port 53 nsew
flabel metal5 s 6598 270240 19088 282760 0 FreeSans 16000 0 0 0 gpio[35]
port 54 nsew
flabel metal5 s 6598 227040 19088 239560 0 FreeSans 16000 0 0 0 gpio[36]
port 55 nsew
flabel metal5 s 6598 956440 19088 968960 0 FreeSans 16000 0 0 0 gpio[24]
port 43 nsew
flabel metal5 s 6598 786640 19088 799160 0 FreeSans 16000 0 0 0 gpio[25]
port 44 nsew
flabel metal5 s 6598 743440 19088 755960 0 FreeSans 16000 0 0 0 gpio[26]
port 45 nsew
flabel metal5 s 6598 700240 19088 712760 0 FreeSans 16000 0 0 0 gpio[27]
port 46 nsew
flabel metal5 s 6598 657040 19088 669560 0 FreeSans 16000 0 0 0 gpio[28]
port 47 nsew
flabel metal5 s 6167 914054 19619 924934 0 FreeSans 16000 0 0 0 vccd2
port 15 nsew
flabel metal5 s 6811 484410 18975 496578 0 FreeSans 16000 0 0 0 vdda2
port 2569 nsew
flabel metal5 s 6811 829010 18975 841178 0 FreeSans 16000 0 0 0 vssa2
port 13 nsew
flabel metal5 s 6167 442854 19619 453734 0 FreeSans 16000 0 0 0 vssd2
port 17 nsew
flabel metal5 s 6598 183840 19088 196360 0 FreeSans 16000 0 0 0 gpio[37]
port 56 nsew
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
