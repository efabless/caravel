VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravel_power_routing
  CLASS BLOCK ;
  FOREIGN caravel_power_routing ;
  ORIGIN 0.000 0.000 ;
  SIZE 3528.960 BY 4988.980 ;
  PIN vccd_core
    PORT
      LAYER met3 ;
        RECT 167.170 221.255 199.110 244.220 ;
        RECT 167.170 171.780 199.110 195.000 ;
      LAYER via3 ;
        RECT 179.775 221.710 198.095 244.030 ;
        RECT 179.655 172.190 197.975 194.510 ;
      LAYER met4 ;
        RECT 190.820 982.830 285.690 997.830 ;
        RECT 635.190 982.830 637.470 997.820 ;
        RECT 710.440 982.830 712.720 997.820 ;
        RECT 785.690 982.830 787.970 997.820 ;
        RECT 860.940 982.830 863.220 997.820 ;
        RECT 936.190 982.830 938.470 997.820 ;
        RECT 1011.440 982.830 1013.720 997.820 ;
        RECT 1086.690 982.830 1088.970 997.820 ;
        RECT 1161.940 982.830 1164.220 997.820 ;
        RECT 1237.190 982.830 1239.470 997.820 ;
        RECT 1312.440 982.830 1314.720 997.820 ;
        RECT 1387.690 982.830 1389.970 997.820 ;
        RECT 1462.940 982.830 1465.220 997.820 ;
        RECT 1538.190 982.830 1540.470 997.820 ;
        RECT 1613.440 982.830 1615.720 997.820 ;
        RECT 1688.690 982.830 1690.970 997.820 ;
        RECT 1763.940 982.830 1766.220 997.820 ;
        RECT 1839.190 982.830 1841.470 997.820 ;
        RECT 1914.440 982.830 1916.720 997.820 ;
        RECT 1989.690 982.830 1991.970 997.820 ;
        RECT 2064.940 982.830 2067.220 997.820 ;
        RECT 2140.190 982.830 2142.470 997.820 ;
        RECT 2215.440 982.830 2217.720 997.820 ;
        RECT 2290.690 982.830 2292.970 997.820 ;
        RECT 2365.940 982.830 2368.220 997.820 ;
        RECT 2441.190 982.830 2443.470 997.820 ;
        RECT 190.880 817.990 203.880 982.830 ;
        RECT 2891.730 878.020 2954.700 893.020 ;
        RECT 3105.110 878.140 3110.430 892.800 ;
        RECT 2953.100 868.960 2954.700 878.020 ;
        RECT 3106.700 868.920 3108.300 878.140 ;
        RECT 2892.370 818.140 2905.760 819.880 ;
        RECT 190.880 814.790 231.610 817.990 ;
        RECT 2892.370 816.540 2934.770 818.140 ;
        RECT 2892.370 815.460 2905.760 816.540 ;
        RECT 190.880 714.210 203.880 814.790 ;
        RECT 179.210 696.130 203.880 714.210 ;
        RECT 183.120 684.790 231.120 687.990 ;
        RECT 2892.370 664.960 2905.760 666.680 ;
        RECT 2892.370 663.360 2934.770 664.960 ;
        RECT 2892.370 662.260 2905.760 663.360 ;
        RECT 182.780 554.790 230.780 557.990 ;
        RECT 2892.370 511.780 2905.760 513.480 ;
        RECT 2892.370 510.180 2934.770 511.780 ;
        RECT 2892.370 509.060 2905.760 510.180 ;
        RECT 182.780 424.790 230.780 427.990 ;
        RECT 2892.370 358.600 2905.760 358.880 ;
        RECT 2892.370 357.000 2934.770 358.600 ;
        RECT 2892.370 354.460 2905.760 357.000 ;
        RECT 182.780 294.790 230.780 297.990 ;
        RECT 179.210 221.270 198.780 244.470 ;
        RECT 3131.660 235.120 3133.260 240.810 ;
        RECT 3171.660 235.580 3173.260 240.500 ;
        RECT 3130.250 221.490 3134.940 235.120 ;
        RECT 3170.380 221.170 3174.500 235.580 ;
        RECT 3119.330 201.020 3120.930 217.370 ;
        RECT 3134.830 201.020 3136.430 217.370 ;
        RECT 3150.330 201.020 3151.930 217.370 ;
        RECT 3165.830 201.020 3167.430 217.370 ;
        RECT 3181.330 201.020 3182.930 217.370 ;
        RECT 179.180 171.750 198.750 194.950 ;
        RECT 179.200 164.790 231.700 167.990 ;
        RECT 179.260 71.610 262.570 91.110 ;
        RECT 686.510 80.180 693.580 83.940 ;
        RECT 689.190 78.690 690.090 80.180 ;
        RECT 3276.240 65.455 3317.020 67.100 ;
      LAYER via4 ;
        RECT 252.660 984.175 284.240 996.555 ;
        RECT 635.590 996.130 636.770 997.310 ;
        RECT 635.590 994.530 636.770 995.710 ;
        RECT 635.590 992.930 636.770 994.110 ;
        RECT 635.590 991.330 636.770 992.510 ;
        RECT 635.590 989.730 636.770 990.910 ;
        RECT 635.590 988.130 636.770 989.310 ;
        RECT 635.590 986.530 636.770 987.710 ;
        RECT 635.590 984.930 636.770 986.110 ;
        RECT 635.590 983.330 636.770 984.510 ;
        RECT 710.840 996.130 712.020 997.310 ;
        RECT 710.840 994.530 712.020 995.710 ;
        RECT 710.840 992.930 712.020 994.110 ;
        RECT 710.840 991.330 712.020 992.510 ;
        RECT 710.840 989.730 712.020 990.910 ;
        RECT 710.840 988.130 712.020 989.310 ;
        RECT 710.840 986.530 712.020 987.710 ;
        RECT 710.840 984.930 712.020 986.110 ;
        RECT 710.840 983.330 712.020 984.510 ;
        RECT 786.090 996.130 787.270 997.310 ;
        RECT 786.090 994.530 787.270 995.710 ;
        RECT 786.090 992.930 787.270 994.110 ;
        RECT 786.090 991.330 787.270 992.510 ;
        RECT 786.090 989.730 787.270 990.910 ;
        RECT 786.090 988.130 787.270 989.310 ;
        RECT 786.090 986.530 787.270 987.710 ;
        RECT 786.090 984.930 787.270 986.110 ;
        RECT 786.090 983.330 787.270 984.510 ;
        RECT 861.340 996.130 862.520 997.310 ;
        RECT 861.340 994.530 862.520 995.710 ;
        RECT 861.340 992.930 862.520 994.110 ;
        RECT 861.340 991.330 862.520 992.510 ;
        RECT 861.340 989.730 862.520 990.910 ;
        RECT 861.340 988.130 862.520 989.310 ;
        RECT 861.340 986.530 862.520 987.710 ;
        RECT 861.340 984.930 862.520 986.110 ;
        RECT 861.340 983.330 862.520 984.510 ;
        RECT 936.590 996.130 937.770 997.310 ;
        RECT 936.590 994.530 937.770 995.710 ;
        RECT 936.590 992.930 937.770 994.110 ;
        RECT 936.590 991.330 937.770 992.510 ;
        RECT 936.590 989.730 937.770 990.910 ;
        RECT 936.590 988.130 937.770 989.310 ;
        RECT 936.590 986.530 937.770 987.710 ;
        RECT 936.590 984.930 937.770 986.110 ;
        RECT 936.590 983.330 937.770 984.510 ;
        RECT 1011.840 996.130 1013.020 997.310 ;
        RECT 1011.840 994.530 1013.020 995.710 ;
        RECT 1011.840 992.930 1013.020 994.110 ;
        RECT 1011.840 991.330 1013.020 992.510 ;
        RECT 1011.840 989.730 1013.020 990.910 ;
        RECT 1011.840 988.130 1013.020 989.310 ;
        RECT 1011.840 986.530 1013.020 987.710 ;
        RECT 1011.840 984.930 1013.020 986.110 ;
        RECT 1011.840 983.330 1013.020 984.510 ;
        RECT 1087.090 996.130 1088.270 997.310 ;
        RECT 1087.090 994.530 1088.270 995.710 ;
        RECT 1087.090 992.930 1088.270 994.110 ;
        RECT 1087.090 991.330 1088.270 992.510 ;
        RECT 1087.090 989.730 1088.270 990.910 ;
        RECT 1087.090 988.130 1088.270 989.310 ;
        RECT 1087.090 986.530 1088.270 987.710 ;
        RECT 1087.090 984.930 1088.270 986.110 ;
        RECT 1087.090 983.330 1088.270 984.510 ;
        RECT 1162.340 996.130 1163.520 997.310 ;
        RECT 1162.340 994.530 1163.520 995.710 ;
        RECT 1162.340 992.930 1163.520 994.110 ;
        RECT 1162.340 991.330 1163.520 992.510 ;
        RECT 1162.340 989.730 1163.520 990.910 ;
        RECT 1162.340 988.130 1163.520 989.310 ;
        RECT 1162.340 986.530 1163.520 987.710 ;
        RECT 1162.340 984.930 1163.520 986.110 ;
        RECT 1162.340 983.330 1163.520 984.510 ;
        RECT 1237.590 996.130 1238.770 997.310 ;
        RECT 1237.590 994.530 1238.770 995.710 ;
        RECT 1237.590 992.930 1238.770 994.110 ;
        RECT 1237.590 991.330 1238.770 992.510 ;
        RECT 1237.590 989.730 1238.770 990.910 ;
        RECT 1237.590 988.130 1238.770 989.310 ;
        RECT 1237.590 986.530 1238.770 987.710 ;
        RECT 1237.590 984.930 1238.770 986.110 ;
        RECT 1237.590 983.330 1238.770 984.510 ;
        RECT 1312.840 996.130 1314.020 997.310 ;
        RECT 1312.840 994.530 1314.020 995.710 ;
        RECT 1312.840 992.930 1314.020 994.110 ;
        RECT 1312.840 991.330 1314.020 992.510 ;
        RECT 1312.840 989.730 1314.020 990.910 ;
        RECT 1312.840 988.130 1314.020 989.310 ;
        RECT 1312.840 986.530 1314.020 987.710 ;
        RECT 1312.840 984.930 1314.020 986.110 ;
        RECT 1312.840 983.330 1314.020 984.510 ;
        RECT 1388.090 996.130 1389.270 997.310 ;
        RECT 1388.090 994.530 1389.270 995.710 ;
        RECT 1388.090 992.930 1389.270 994.110 ;
        RECT 1388.090 991.330 1389.270 992.510 ;
        RECT 1388.090 989.730 1389.270 990.910 ;
        RECT 1388.090 988.130 1389.270 989.310 ;
        RECT 1388.090 986.530 1389.270 987.710 ;
        RECT 1388.090 984.930 1389.270 986.110 ;
        RECT 1388.090 983.330 1389.270 984.510 ;
        RECT 1463.340 996.130 1464.520 997.310 ;
        RECT 1463.340 994.530 1464.520 995.710 ;
        RECT 1463.340 992.930 1464.520 994.110 ;
        RECT 1463.340 991.330 1464.520 992.510 ;
        RECT 1463.340 989.730 1464.520 990.910 ;
        RECT 1463.340 988.130 1464.520 989.310 ;
        RECT 1463.340 986.530 1464.520 987.710 ;
        RECT 1463.340 984.930 1464.520 986.110 ;
        RECT 1463.340 983.330 1464.520 984.510 ;
        RECT 1538.590 996.130 1539.770 997.310 ;
        RECT 1538.590 994.530 1539.770 995.710 ;
        RECT 1538.590 992.930 1539.770 994.110 ;
        RECT 1538.590 991.330 1539.770 992.510 ;
        RECT 1538.590 989.730 1539.770 990.910 ;
        RECT 1538.590 988.130 1539.770 989.310 ;
        RECT 1538.590 986.530 1539.770 987.710 ;
        RECT 1538.590 984.930 1539.770 986.110 ;
        RECT 1538.590 983.330 1539.770 984.510 ;
        RECT 1613.840 996.130 1615.020 997.310 ;
        RECT 1613.840 994.530 1615.020 995.710 ;
        RECT 1613.840 992.930 1615.020 994.110 ;
        RECT 1613.840 991.330 1615.020 992.510 ;
        RECT 1613.840 989.730 1615.020 990.910 ;
        RECT 1613.840 988.130 1615.020 989.310 ;
        RECT 1613.840 986.530 1615.020 987.710 ;
        RECT 1613.840 984.930 1615.020 986.110 ;
        RECT 1613.840 983.330 1615.020 984.510 ;
        RECT 1689.090 996.130 1690.270 997.310 ;
        RECT 1689.090 994.530 1690.270 995.710 ;
        RECT 1689.090 992.930 1690.270 994.110 ;
        RECT 1689.090 991.330 1690.270 992.510 ;
        RECT 1689.090 989.730 1690.270 990.910 ;
        RECT 1689.090 988.130 1690.270 989.310 ;
        RECT 1689.090 986.530 1690.270 987.710 ;
        RECT 1689.090 984.930 1690.270 986.110 ;
        RECT 1689.090 983.330 1690.270 984.510 ;
        RECT 1764.340 996.130 1765.520 997.310 ;
        RECT 1764.340 994.530 1765.520 995.710 ;
        RECT 1764.340 992.930 1765.520 994.110 ;
        RECT 1764.340 991.330 1765.520 992.510 ;
        RECT 1764.340 989.730 1765.520 990.910 ;
        RECT 1764.340 988.130 1765.520 989.310 ;
        RECT 1764.340 986.530 1765.520 987.710 ;
        RECT 1764.340 984.930 1765.520 986.110 ;
        RECT 1764.340 983.330 1765.520 984.510 ;
        RECT 1839.590 996.130 1840.770 997.310 ;
        RECT 1839.590 994.530 1840.770 995.710 ;
        RECT 1839.590 992.930 1840.770 994.110 ;
        RECT 1839.590 991.330 1840.770 992.510 ;
        RECT 1839.590 989.730 1840.770 990.910 ;
        RECT 1839.590 988.130 1840.770 989.310 ;
        RECT 1839.590 986.530 1840.770 987.710 ;
        RECT 1839.590 984.930 1840.770 986.110 ;
        RECT 1839.590 983.330 1840.770 984.510 ;
        RECT 1914.840 996.130 1916.020 997.310 ;
        RECT 1914.840 994.530 1916.020 995.710 ;
        RECT 1914.840 992.930 1916.020 994.110 ;
        RECT 1914.840 991.330 1916.020 992.510 ;
        RECT 1914.840 989.730 1916.020 990.910 ;
        RECT 1914.840 988.130 1916.020 989.310 ;
        RECT 1914.840 986.530 1916.020 987.710 ;
        RECT 1914.840 984.930 1916.020 986.110 ;
        RECT 1914.840 983.330 1916.020 984.510 ;
        RECT 1990.090 996.130 1991.270 997.310 ;
        RECT 1990.090 994.530 1991.270 995.710 ;
        RECT 1990.090 992.930 1991.270 994.110 ;
        RECT 1990.090 991.330 1991.270 992.510 ;
        RECT 1990.090 989.730 1991.270 990.910 ;
        RECT 1990.090 988.130 1991.270 989.310 ;
        RECT 1990.090 986.530 1991.270 987.710 ;
        RECT 1990.090 984.930 1991.270 986.110 ;
        RECT 1990.090 983.330 1991.270 984.510 ;
        RECT 2065.340 996.130 2066.520 997.310 ;
        RECT 2065.340 994.530 2066.520 995.710 ;
        RECT 2065.340 992.930 2066.520 994.110 ;
        RECT 2065.340 991.330 2066.520 992.510 ;
        RECT 2065.340 989.730 2066.520 990.910 ;
        RECT 2065.340 988.130 2066.520 989.310 ;
        RECT 2065.340 986.530 2066.520 987.710 ;
        RECT 2065.340 984.930 2066.520 986.110 ;
        RECT 2065.340 983.330 2066.520 984.510 ;
        RECT 2140.590 996.130 2141.770 997.310 ;
        RECT 2140.590 994.530 2141.770 995.710 ;
        RECT 2140.590 992.930 2141.770 994.110 ;
        RECT 2140.590 991.330 2141.770 992.510 ;
        RECT 2140.590 989.730 2141.770 990.910 ;
        RECT 2140.590 988.130 2141.770 989.310 ;
        RECT 2140.590 986.530 2141.770 987.710 ;
        RECT 2140.590 984.930 2141.770 986.110 ;
        RECT 2140.590 983.330 2141.770 984.510 ;
        RECT 2215.840 996.130 2217.020 997.310 ;
        RECT 2215.840 994.530 2217.020 995.710 ;
        RECT 2215.840 992.930 2217.020 994.110 ;
        RECT 2215.840 991.330 2217.020 992.510 ;
        RECT 2215.840 989.730 2217.020 990.910 ;
        RECT 2215.840 988.130 2217.020 989.310 ;
        RECT 2215.840 986.530 2217.020 987.710 ;
        RECT 2215.840 984.930 2217.020 986.110 ;
        RECT 2215.840 983.330 2217.020 984.510 ;
        RECT 2291.090 996.130 2292.270 997.310 ;
        RECT 2291.090 994.530 2292.270 995.710 ;
        RECT 2291.090 992.930 2292.270 994.110 ;
        RECT 2291.090 991.330 2292.270 992.510 ;
        RECT 2291.090 989.730 2292.270 990.910 ;
        RECT 2291.090 988.130 2292.270 989.310 ;
        RECT 2291.090 986.530 2292.270 987.710 ;
        RECT 2291.090 984.930 2292.270 986.110 ;
        RECT 2291.090 983.330 2292.270 984.510 ;
        RECT 2366.340 996.130 2367.520 997.310 ;
        RECT 2366.340 994.530 2367.520 995.710 ;
        RECT 2366.340 992.930 2367.520 994.110 ;
        RECT 2366.340 991.330 2367.520 992.510 ;
        RECT 2366.340 989.730 2367.520 990.910 ;
        RECT 2366.340 988.130 2367.520 989.310 ;
        RECT 2366.340 986.530 2367.520 987.710 ;
        RECT 2366.340 984.930 2367.520 986.110 ;
        RECT 2366.340 983.330 2367.520 984.510 ;
        RECT 2441.590 996.130 2442.770 997.310 ;
        RECT 2441.590 994.530 2442.770 995.710 ;
        RECT 2441.590 992.930 2442.770 994.110 ;
        RECT 2441.590 991.330 2442.770 992.510 ;
        RECT 2441.590 989.730 2442.770 990.910 ;
        RECT 2441.590 988.130 2442.770 989.310 ;
        RECT 2441.590 986.530 2442.770 987.710 ;
        RECT 2441.590 984.930 2442.770 986.110 ;
        RECT 2441.590 983.330 2442.770 984.510 ;
        RECT 2892.940 879.475 2905.320 891.855 ;
        RECT 2937.210 879.475 2949.590 891.855 ;
        RECT 3106.405 879.290 3109.185 891.670 ;
        RECT 227.755 815.880 228.935 817.060 ;
        RECT 229.355 815.880 230.535 817.060 ;
        RECT 2893.805 816.325 2904.585 819.105 ;
        RECT 2930.080 816.735 2931.260 817.915 ;
        RECT 2931.680 816.735 2932.860 817.915 ;
        RECT 2933.280 816.735 2934.460 817.915 ;
        RECT 180.325 697.445 197.505 713.025 ;
        RECT 184.175 685.790 185.355 686.970 ;
        RECT 185.775 685.790 186.955 686.970 ;
        RECT 187.375 685.790 188.555 686.970 ;
        RECT 188.975 685.790 190.155 686.970 ;
        RECT 190.575 685.790 191.755 686.970 ;
        RECT 192.175 685.790 193.355 686.970 ;
        RECT 193.775 685.790 194.955 686.970 ;
        RECT 195.375 685.790 196.555 686.970 ;
        RECT 196.975 685.790 198.155 686.970 ;
        RECT 227.215 685.810 228.395 686.990 ;
        RECT 228.815 685.810 229.995 686.990 ;
        RECT 2893.805 663.125 2904.585 665.905 ;
        RECT 2929.995 663.595 2931.175 664.775 ;
        RECT 2931.595 663.595 2932.775 664.775 ;
        RECT 2933.195 663.595 2934.375 664.775 ;
        RECT 184.245 555.820 185.425 557.000 ;
        RECT 185.845 555.820 187.025 557.000 ;
        RECT 187.445 555.820 188.625 557.000 ;
        RECT 189.045 555.820 190.225 557.000 ;
        RECT 190.645 555.820 191.825 557.000 ;
        RECT 192.245 555.820 193.425 557.000 ;
        RECT 193.845 555.820 195.025 557.000 ;
        RECT 195.445 555.820 196.625 557.000 ;
        RECT 197.045 555.820 198.225 557.000 ;
        RECT 226.885 555.770 228.065 556.950 ;
        RECT 228.485 555.770 229.665 556.950 ;
        RECT 2893.805 509.925 2904.585 512.705 ;
        RECT 2929.945 510.395 2931.125 511.575 ;
        RECT 2931.545 510.395 2932.725 511.575 ;
        RECT 2933.145 510.395 2934.325 511.575 ;
        RECT 184.195 425.800 185.375 426.980 ;
        RECT 185.795 425.800 186.975 426.980 ;
        RECT 187.395 425.800 188.575 426.980 ;
        RECT 188.995 425.800 190.175 426.980 ;
        RECT 190.595 425.800 191.775 426.980 ;
        RECT 192.195 425.800 193.375 426.980 ;
        RECT 193.795 425.800 194.975 426.980 ;
        RECT 195.395 425.800 196.575 426.980 ;
        RECT 196.995 425.800 198.175 426.980 ;
        RECT 226.865 425.800 228.045 426.980 ;
        RECT 228.465 425.800 229.645 426.980 ;
        RECT 2893.805 355.325 2904.585 358.105 ;
        RECT 2930.005 357.210 2931.185 358.390 ;
        RECT 2931.605 357.210 2932.785 358.390 ;
        RECT 2933.205 357.210 2934.385 358.390 ;
        RECT 184.175 295.790 185.355 296.970 ;
        RECT 185.775 295.790 186.955 296.970 ;
        RECT 187.375 295.790 188.555 296.970 ;
        RECT 188.975 295.790 190.155 296.970 ;
        RECT 190.575 295.790 191.755 296.970 ;
        RECT 192.175 295.790 193.355 296.970 ;
        RECT 193.775 295.790 194.955 296.970 ;
        RECT 195.375 295.790 196.555 296.970 ;
        RECT 196.975 295.790 198.155 296.970 ;
        RECT 226.885 295.780 228.065 296.960 ;
        RECT 228.485 295.780 229.665 296.960 ;
        RECT 180.345 221.880 197.525 243.860 ;
        RECT 3131.160 222.865 3133.940 233.645 ;
        RECT 3171.050 222.200 3173.830 234.580 ;
        RECT 3119.485 215.285 3120.665 216.465 ;
        RECT 3119.485 213.685 3120.665 214.865 ;
        RECT 3119.485 212.085 3120.665 213.265 ;
        RECT 3135.045 215.355 3136.225 216.535 ;
        RECT 3135.045 213.755 3136.225 214.935 ;
        RECT 3135.045 212.155 3136.225 213.335 ;
        RECT 3150.495 215.335 3151.675 216.515 ;
        RECT 3150.495 213.735 3151.675 214.915 ;
        RECT 3150.495 212.135 3151.675 213.315 ;
        RECT 3165.965 215.335 3167.145 216.515 ;
        RECT 3165.965 213.735 3167.145 214.915 ;
        RECT 3165.965 212.135 3167.145 213.315 ;
        RECT 3181.505 215.395 3182.685 216.575 ;
        RECT 3181.505 213.795 3182.685 214.975 ;
        RECT 3181.505 212.195 3182.685 213.375 ;
        RECT 180.225 172.360 197.405 194.340 ;
        RECT 180.365 165.760 181.545 166.940 ;
        RECT 181.965 165.760 183.145 166.940 ;
        RECT 183.565 165.760 184.745 166.940 ;
        RECT 185.165 165.760 186.345 166.940 ;
        RECT 186.765 165.760 187.945 166.940 ;
        RECT 188.365 165.760 189.545 166.940 ;
        RECT 189.965 165.760 191.145 166.940 ;
        RECT 191.565 165.760 192.745 166.940 ;
        RECT 193.165 165.760 194.345 166.940 ;
        RECT 194.765 165.760 195.945 166.940 ;
        RECT 196.365 165.760 197.545 166.940 ;
        RECT 227.875 165.790 229.055 166.970 ;
        RECT 229.475 165.790 230.655 166.970 ;
        RECT 180.290 72.890 197.470 90.070 ;
        RECT 243.140 72.720 260.320 89.900 ;
        RECT 687.005 80.680 692.985 83.460 ;
        RECT 3302.500 65.690 3303.680 66.870 ;
        RECT 3304.100 65.690 3305.280 66.870 ;
        RECT 3305.700 65.690 3306.880 66.870 ;
        RECT 3307.300 65.690 3308.480 66.870 ;
        RECT 3308.900 65.690 3310.080 66.870 ;
        RECT 3310.500 65.690 3311.680 66.870 ;
        RECT 3312.100 65.690 3313.280 66.870 ;
        RECT 3313.700 65.690 3314.880 66.870 ;
        RECT 3315.300 65.690 3316.480 66.870 ;
      LAYER met5 ;
        RECT 251.370 982.830 2906.760 997.830 ;
        RECT 2891.760 817.990 2906.760 982.830 ;
        RECT 3212.930 959.860 3226.680 961.460 ;
        RECT 3221.010 941.460 3226.680 959.860 ;
        RECT 3213.090 939.860 3226.680 941.460 ;
        RECT 3221.010 893.020 3226.680 939.860 ;
        RECT 2936.150 878.020 3317.020 893.020 ;
        RECT 3302.020 818.140 3317.020 878.020 ;
        RECT 226.610 814.790 235.970 817.990 ;
        RECT 2843.120 814.790 2906.760 817.990 ;
        RECT 2929.770 816.540 2937.860 818.140 ;
        RECT 3296.080 816.540 3317.020 818.140 ;
        RECT 178.730 70.870 198.730 714.870 ;
        RECT 2891.760 687.990 2906.760 814.790 ;
        RECT 226.120 684.790 236.090 687.990 ;
        RECT 2843.120 684.790 2906.760 687.990 ;
        RECT 2891.760 557.990 2906.760 684.790 ;
        RECT 3302.020 664.960 3317.020 816.540 ;
        RECT 2929.650 663.360 2937.860 664.960 ;
        RECT 3295.920 663.360 3317.020 664.960 ;
        RECT 225.780 554.790 236.220 557.990 ;
        RECT 2843.120 554.790 2906.760 557.990 ;
        RECT 2891.760 427.990 2906.760 554.790 ;
        RECT 3302.020 511.780 3317.020 663.360 ;
        RECT 2929.590 510.180 2937.860 511.780 ;
        RECT 3295.710 510.180 3317.020 511.780 ;
        RECT 225.780 424.790 236.220 427.990 ;
        RECT 2843.120 424.790 2906.760 427.990 ;
        RECT 2891.760 297.990 2906.760 424.790 ;
        RECT 3302.020 358.600 3317.020 510.180 ;
        RECT 2929.590 357.000 2937.860 358.600 ;
        RECT 3295.770 357.000 3317.020 358.600 ;
        RECT 225.780 294.790 236.220 297.990 ;
        RECT 2843.120 294.790 2906.760 297.990 ;
        RECT 3187.610 297.870 3202.610 298.440 ;
        RECT 3179.420 296.270 3202.610 297.870 ;
        RECT 3302.020 297.530 3317.020 357.000 ;
        RECT 2891.760 167.990 2906.760 294.790 ;
        RECT 3187.610 257.870 3202.610 296.270 ;
        RECT 3282.500 295.930 3317.020 297.530 ;
        RECT 3302.020 289.370 3317.020 295.930 ;
        RECT 3282.310 287.770 3317.020 289.370 ;
        RECT 3302.020 281.210 3317.020 287.770 ;
        RECT 3282.410 279.610 3317.020 281.210 ;
        RECT 3179.730 256.270 3202.610 257.870 ;
        RECT 3187.610 235.910 3202.610 256.270 ;
        RECT 3302.020 235.910 3317.020 279.610 ;
        RECT 3129.900 220.910 3317.020 235.910 ;
        RECT 3196.170 216.840 3205.310 220.910 ;
        RECT 3118.820 211.840 3205.310 216.840 ;
        RECT 3201.310 197.930 3205.310 211.840 ;
        RECT 3197.570 196.330 3205.310 197.930 ;
        RECT 3201.310 181.030 3205.310 196.330 ;
        RECT 3197.400 179.430 3205.310 181.030 ;
        RECT 226.700 164.790 235.750 167.990 ;
        RECT 2843.660 164.790 2906.760 167.990 ;
        RECT 2891.760 91.610 2906.760 164.790 ;
        RECT 3201.310 164.130 3205.310 179.430 ;
        RECT 3198.010 162.530 3205.310 164.130 ;
        RECT 241.760 71.610 2906.760 91.610 ;
        RECT 3302.020 65.390 3317.020 220.910 ;
    END
  END vccd_core
  PIN vssd_core
    PORT
      LAYER met1 ;
        RECT 3210.410 64.190 3218.240 66.440 ;
        RECT 3210.410 63.490 3220.690 64.190 ;
        RECT 3210.410 63.450 3218.240 63.490 ;
      LAYER via ;
        RECT 3210.835 63.870 3217.815 66.050 ;
      LAYER met2 ;
        RECT 3210.410 64.190 3218.240 66.440 ;
        RECT 3210.410 63.490 3220.690 64.190 ;
        RECT 3210.410 63.450 3218.240 63.490 ;
      LAYER via2 ;
        RECT 3210.785 63.820 3217.865 66.100 ;
      LAYER met3 ;
        RECT 3210.410 64.720 3218.240 66.440 ;
        RECT 1178.340 27.630 1200.135 63.930 ;
        RECT 1226.390 27.630 1248.400 63.930 ;
        RECT 3210.410 63.490 3220.680 64.720 ;
        RECT 3210.410 63.450 3218.240 63.490 ;
      LAYER via3 ;
        RECT 1178.645 44.785 1199.765 63.505 ;
        RECT 1226.905 44.855 1248.025 63.575 ;
        RECT 3210.765 63.800 3217.885 66.120 ;
      LAYER met4 ;
        RECT 208.820 1002.830 286.140 1017.830 ;
        RECT 672.110 1002.740 674.510 1017.870 ;
        RECT 747.510 1002.740 749.910 1017.870 ;
        RECT 822.760 1002.740 825.160 1017.870 ;
        RECT 897.810 1002.740 900.210 1017.870 ;
        RECT 1048.510 1002.740 1050.910 1017.870 ;
        RECT 1123.760 1002.740 1126.160 1017.870 ;
        RECT 1199.010 1002.740 1201.410 1017.870 ;
        RECT 1274.260 1002.740 1276.660 1017.870 ;
        RECT 1349.510 1002.740 1351.910 1017.870 ;
        RECT 1424.760 1002.740 1427.160 1017.870 ;
        RECT 1499.810 1002.740 1502.210 1017.870 ;
        RECT 1575.760 1002.740 1578.160 1017.870 ;
        RECT 1650.510 1002.740 1652.910 1017.870 ;
        RECT 1726.260 1002.740 1728.660 1017.870 ;
        RECT 1801.010 1002.740 1803.410 1017.870 ;
        RECT 1875.260 1002.740 1877.660 1017.870 ;
        RECT 1951.110 1002.740 1953.510 1017.870 ;
        RECT 2026.760 1002.740 2029.160 1017.870 ;
        RECT 2102.010 1002.740 2104.410 1017.870 ;
        RECT 2177.260 1002.740 2179.660 1017.870 ;
        RECT 2252.510 1002.740 2254.910 1017.870 ;
        RECT 2327.760 1002.740 2330.160 1017.870 ;
        RECT 2403.010 1002.740 2405.410 1017.870 ;
        RECT 2478.260 1002.740 2480.660 1017.870 ;
        RECT 2881.200 869.810 2926.830 873.010 ;
        RECT 2880.250 749.810 2926.830 753.010 ;
        RECT 2870.250 619.810 2926.830 623.010 ;
        RECT 2870.250 489.810 2926.830 493.010 ;
        RECT 2870.250 359.810 2926.830 363.010 ;
        RECT 2956.400 324.300 2958.000 342.080 ;
        RECT 3110.000 324.520 3111.600 341.690 ;
        RECT 2953.600 310.280 2960.650 324.300 ;
        RECT 3107.810 310.750 3114.400 324.520 ;
        RECT 3150.290 312.670 3154.860 324.290 ;
        RECT 3151.660 302.740 3153.260 312.670 ;
        RECT 2870.250 229.810 2926.830 233.010 ;
        RECT 3127.080 201.020 3128.680 217.370 ;
        RECT 3142.580 201.020 3144.180 217.370 ;
        RECT 3158.080 201.020 3159.680 217.370 ;
        RECT 3173.580 201.020 3175.180 217.370 ;
        RECT 3189.080 201.020 3190.680 217.370 ;
        RECT 682.690 57.480 683.590 66.780 ;
        RECT 678.770 57.470 684.220 57.480 ;
        RECT 676.770 51.150 684.220 57.470 ;
        RECT 1178.290 44.420 1200.170 63.960 ;
        RECT 1226.400 44.440 1248.390 63.920 ;
        RECT 3210.410 63.450 3218.240 66.440 ;
      LAYER via4 ;
        RECT 210.345 1004.195 222.725 1016.575 ;
        RECT 252.165 1004.225 285.345 1016.605 ;
        RECT 672.490 1016.125 673.670 1017.305 ;
        RECT 672.490 1014.525 673.670 1015.705 ;
        RECT 672.490 1012.925 673.670 1014.105 ;
        RECT 672.490 1011.325 673.670 1012.505 ;
        RECT 672.490 1009.725 673.670 1010.905 ;
        RECT 672.490 1008.125 673.670 1009.305 ;
        RECT 672.490 1006.525 673.670 1007.705 ;
        RECT 672.490 1004.925 673.670 1006.105 ;
        RECT 672.490 1003.325 673.670 1004.505 ;
        RECT 747.890 1016.125 749.070 1017.305 ;
        RECT 747.890 1014.525 749.070 1015.705 ;
        RECT 747.890 1012.925 749.070 1014.105 ;
        RECT 747.890 1011.325 749.070 1012.505 ;
        RECT 747.890 1009.725 749.070 1010.905 ;
        RECT 747.890 1008.125 749.070 1009.305 ;
        RECT 747.890 1006.525 749.070 1007.705 ;
        RECT 747.890 1004.925 749.070 1006.105 ;
        RECT 747.890 1003.325 749.070 1004.505 ;
        RECT 823.140 1016.125 824.320 1017.305 ;
        RECT 823.140 1014.525 824.320 1015.705 ;
        RECT 823.140 1012.925 824.320 1014.105 ;
        RECT 823.140 1011.325 824.320 1012.505 ;
        RECT 823.140 1009.725 824.320 1010.905 ;
        RECT 823.140 1008.125 824.320 1009.305 ;
        RECT 823.140 1006.525 824.320 1007.705 ;
        RECT 823.140 1004.925 824.320 1006.105 ;
        RECT 823.140 1003.325 824.320 1004.505 ;
        RECT 898.190 1016.125 899.370 1017.305 ;
        RECT 898.190 1014.525 899.370 1015.705 ;
        RECT 898.190 1012.925 899.370 1014.105 ;
        RECT 898.190 1011.325 899.370 1012.505 ;
        RECT 898.190 1009.725 899.370 1010.905 ;
        RECT 898.190 1008.125 899.370 1009.305 ;
        RECT 898.190 1006.525 899.370 1007.705 ;
        RECT 898.190 1004.925 899.370 1006.105 ;
        RECT 898.190 1003.325 899.370 1004.505 ;
        RECT 1048.890 1016.125 1050.070 1017.305 ;
        RECT 1048.890 1014.525 1050.070 1015.705 ;
        RECT 1048.890 1012.925 1050.070 1014.105 ;
        RECT 1048.890 1011.325 1050.070 1012.505 ;
        RECT 1048.890 1009.725 1050.070 1010.905 ;
        RECT 1048.890 1008.125 1050.070 1009.305 ;
        RECT 1048.890 1006.525 1050.070 1007.705 ;
        RECT 1048.890 1004.925 1050.070 1006.105 ;
        RECT 1048.890 1003.325 1050.070 1004.505 ;
        RECT 1124.140 1016.125 1125.320 1017.305 ;
        RECT 1124.140 1014.525 1125.320 1015.705 ;
        RECT 1124.140 1012.925 1125.320 1014.105 ;
        RECT 1124.140 1011.325 1125.320 1012.505 ;
        RECT 1124.140 1009.725 1125.320 1010.905 ;
        RECT 1124.140 1008.125 1125.320 1009.305 ;
        RECT 1124.140 1006.525 1125.320 1007.705 ;
        RECT 1124.140 1004.925 1125.320 1006.105 ;
        RECT 1124.140 1003.325 1125.320 1004.505 ;
        RECT 1199.390 1016.125 1200.570 1017.305 ;
        RECT 1199.390 1014.525 1200.570 1015.705 ;
        RECT 1199.390 1012.925 1200.570 1014.105 ;
        RECT 1199.390 1011.325 1200.570 1012.505 ;
        RECT 1199.390 1009.725 1200.570 1010.905 ;
        RECT 1199.390 1008.125 1200.570 1009.305 ;
        RECT 1199.390 1006.525 1200.570 1007.705 ;
        RECT 1199.390 1004.925 1200.570 1006.105 ;
        RECT 1199.390 1003.325 1200.570 1004.505 ;
        RECT 1274.640 1016.125 1275.820 1017.305 ;
        RECT 1274.640 1014.525 1275.820 1015.705 ;
        RECT 1274.640 1012.925 1275.820 1014.105 ;
        RECT 1274.640 1011.325 1275.820 1012.505 ;
        RECT 1274.640 1009.725 1275.820 1010.905 ;
        RECT 1274.640 1008.125 1275.820 1009.305 ;
        RECT 1274.640 1006.525 1275.820 1007.705 ;
        RECT 1274.640 1004.925 1275.820 1006.105 ;
        RECT 1274.640 1003.325 1275.820 1004.505 ;
        RECT 1349.890 1016.125 1351.070 1017.305 ;
        RECT 1349.890 1014.525 1351.070 1015.705 ;
        RECT 1349.890 1012.925 1351.070 1014.105 ;
        RECT 1349.890 1011.325 1351.070 1012.505 ;
        RECT 1349.890 1009.725 1351.070 1010.905 ;
        RECT 1349.890 1008.125 1351.070 1009.305 ;
        RECT 1349.890 1006.525 1351.070 1007.705 ;
        RECT 1349.890 1004.925 1351.070 1006.105 ;
        RECT 1349.890 1003.325 1351.070 1004.505 ;
        RECT 1425.140 1016.125 1426.320 1017.305 ;
        RECT 1425.140 1014.525 1426.320 1015.705 ;
        RECT 1425.140 1012.925 1426.320 1014.105 ;
        RECT 1425.140 1011.325 1426.320 1012.505 ;
        RECT 1425.140 1009.725 1426.320 1010.905 ;
        RECT 1425.140 1008.125 1426.320 1009.305 ;
        RECT 1425.140 1006.525 1426.320 1007.705 ;
        RECT 1425.140 1004.925 1426.320 1006.105 ;
        RECT 1425.140 1003.325 1426.320 1004.505 ;
        RECT 1500.190 1016.125 1501.370 1017.305 ;
        RECT 1500.190 1014.525 1501.370 1015.705 ;
        RECT 1500.190 1012.925 1501.370 1014.105 ;
        RECT 1500.190 1011.325 1501.370 1012.505 ;
        RECT 1500.190 1009.725 1501.370 1010.905 ;
        RECT 1500.190 1008.125 1501.370 1009.305 ;
        RECT 1500.190 1006.525 1501.370 1007.705 ;
        RECT 1500.190 1004.925 1501.370 1006.105 ;
        RECT 1500.190 1003.325 1501.370 1004.505 ;
        RECT 1576.140 1016.125 1577.320 1017.305 ;
        RECT 1576.140 1014.525 1577.320 1015.705 ;
        RECT 1576.140 1012.925 1577.320 1014.105 ;
        RECT 1576.140 1011.325 1577.320 1012.505 ;
        RECT 1576.140 1009.725 1577.320 1010.905 ;
        RECT 1576.140 1008.125 1577.320 1009.305 ;
        RECT 1576.140 1006.525 1577.320 1007.705 ;
        RECT 1576.140 1004.925 1577.320 1006.105 ;
        RECT 1576.140 1003.325 1577.320 1004.505 ;
        RECT 1650.890 1016.125 1652.070 1017.305 ;
        RECT 1650.890 1014.525 1652.070 1015.705 ;
        RECT 1650.890 1012.925 1652.070 1014.105 ;
        RECT 1650.890 1011.325 1652.070 1012.505 ;
        RECT 1650.890 1009.725 1652.070 1010.905 ;
        RECT 1650.890 1008.125 1652.070 1009.305 ;
        RECT 1650.890 1006.525 1652.070 1007.705 ;
        RECT 1650.890 1004.925 1652.070 1006.105 ;
        RECT 1650.890 1003.325 1652.070 1004.505 ;
        RECT 1726.640 1016.125 1727.820 1017.305 ;
        RECT 1726.640 1014.525 1727.820 1015.705 ;
        RECT 1726.640 1012.925 1727.820 1014.105 ;
        RECT 1726.640 1011.325 1727.820 1012.505 ;
        RECT 1726.640 1009.725 1727.820 1010.905 ;
        RECT 1726.640 1008.125 1727.820 1009.305 ;
        RECT 1726.640 1006.525 1727.820 1007.705 ;
        RECT 1726.640 1004.925 1727.820 1006.105 ;
        RECT 1726.640 1003.325 1727.820 1004.505 ;
        RECT 1801.390 1016.125 1802.570 1017.305 ;
        RECT 1801.390 1014.525 1802.570 1015.705 ;
        RECT 1801.390 1012.925 1802.570 1014.105 ;
        RECT 1801.390 1011.325 1802.570 1012.505 ;
        RECT 1801.390 1009.725 1802.570 1010.905 ;
        RECT 1801.390 1008.125 1802.570 1009.305 ;
        RECT 1801.390 1006.525 1802.570 1007.705 ;
        RECT 1801.390 1004.925 1802.570 1006.105 ;
        RECT 1801.390 1003.325 1802.570 1004.505 ;
        RECT 1875.640 1016.125 1876.820 1017.305 ;
        RECT 1875.640 1014.525 1876.820 1015.705 ;
        RECT 1875.640 1012.925 1876.820 1014.105 ;
        RECT 1875.640 1011.325 1876.820 1012.505 ;
        RECT 1875.640 1009.725 1876.820 1010.905 ;
        RECT 1875.640 1008.125 1876.820 1009.305 ;
        RECT 1875.640 1006.525 1876.820 1007.705 ;
        RECT 1875.640 1004.925 1876.820 1006.105 ;
        RECT 1875.640 1003.325 1876.820 1004.505 ;
        RECT 1951.490 1016.125 1952.670 1017.305 ;
        RECT 1951.490 1014.525 1952.670 1015.705 ;
        RECT 1951.490 1012.925 1952.670 1014.105 ;
        RECT 1951.490 1011.325 1952.670 1012.505 ;
        RECT 1951.490 1009.725 1952.670 1010.905 ;
        RECT 1951.490 1008.125 1952.670 1009.305 ;
        RECT 1951.490 1006.525 1952.670 1007.705 ;
        RECT 1951.490 1004.925 1952.670 1006.105 ;
        RECT 1951.490 1003.325 1952.670 1004.505 ;
        RECT 2027.140 1016.125 2028.320 1017.305 ;
        RECT 2027.140 1014.525 2028.320 1015.705 ;
        RECT 2027.140 1012.925 2028.320 1014.105 ;
        RECT 2027.140 1011.325 2028.320 1012.505 ;
        RECT 2027.140 1009.725 2028.320 1010.905 ;
        RECT 2027.140 1008.125 2028.320 1009.305 ;
        RECT 2027.140 1006.525 2028.320 1007.705 ;
        RECT 2027.140 1004.925 2028.320 1006.105 ;
        RECT 2027.140 1003.325 2028.320 1004.505 ;
        RECT 2102.390 1016.125 2103.570 1017.305 ;
        RECT 2102.390 1014.525 2103.570 1015.705 ;
        RECT 2102.390 1012.925 2103.570 1014.105 ;
        RECT 2102.390 1011.325 2103.570 1012.505 ;
        RECT 2102.390 1009.725 2103.570 1010.905 ;
        RECT 2102.390 1008.125 2103.570 1009.305 ;
        RECT 2102.390 1006.525 2103.570 1007.705 ;
        RECT 2102.390 1004.925 2103.570 1006.105 ;
        RECT 2102.390 1003.325 2103.570 1004.505 ;
        RECT 2177.640 1016.125 2178.820 1017.305 ;
        RECT 2177.640 1014.525 2178.820 1015.705 ;
        RECT 2177.640 1012.925 2178.820 1014.105 ;
        RECT 2177.640 1011.325 2178.820 1012.505 ;
        RECT 2177.640 1009.725 2178.820 1010.905 ;
        RECT 2177.640 1008.125 2178.820 1009.305 ;
        RECT 2177.640 1006.525 2178.820 1007.705 ;
        RECT 2177.640 1004.925 2178.820 1006.105 ;
        RECT 2177.640 1003.325 2178.820 1004.505 ;
        RECT 2252.890 1016.125 2254.070 1017.305 ;
        RECT 2252.890 1014.525 2254.070 1015.705 ;
        RECT 2252.890 1012.925 2254.070 1014.105 ;
        RECT 2252.890 1011.325 2254.070 1012.505 ;
        RECT 2252.890 1009.725 2254.070 1010.905 ;
        RECT 2252.890 1008.125 2254.070 1009.305 ;
        RECT 2252.890 1006.525 2254.070 1007.705 ;
        RECT 2252.890 1004.925 2254.070 1006.105 ;
        RECT 2252.890 1003.325 2254.070 1004.505 ;
        RECT 2328.140 1016.125 2329.320 1017.305 ;
        RECT 2328.140 1014.525 2329.320 1015.705 ;
        RECT 2328.140 1012.925 2329.320 1014.105 ;
        RECT 2328.140 1011.325 2329.320 1012.505 ;
        RECT 2328.140 1009.725 2329.320 1010.905 ;
        RECT 2328.140 1008.125 2329.320 1009.305 ;
        RECT 2328.140 1006.525 2329.320 1007.705 ;
        RECT 2328.140 1004.925 2329.320 1006.105 ;
        RECT 2328.140 1003.325 2329.320 1004.505 ;
        RECT 2403.390 1016.125 2404.570 1017.305 ;
        RECT 2403.390 1014.525 2404.570 1015.705 ;
        RECT 2403.390 1012.925 2404.570 1014.105 ;
        RECT 2403.390 1011.325 2404.570 1012.505 ;
        RECT 2403.390 1009.725 2404.570 1010.905 ;
        RECT 2403.390 1008.125 2404.570 1009.305 ;
        RECT 2403.390 1006.525 2404.570 1007.705 ;
        RECT 2403.390 1004.925 2404.570 1006.105 ;
        RECT 2403.390 1003.325 2404.570 1004.505 ;
        RECT 2478.640 1016.125 2479.820 1017.305 ;
        RECT 2478.640 1014.525 2479.820 1015.705 ;
        RECT 2478.640 1012.925 2479.820 1014.105 ;
        RECT 2478.640 1011.325 2479.820 1012.505 ;
        RECT 2478.640 1009.725 2479.820 1010.905 ;
        RECT 2478.640 1008.125 2479.820 1009.305 ;
        RECT 2478.640 1006.525 2479.820 1007.705 ;
        RECT 2478.640 1004.925 2479.820 1006.105 ;
        RECT 2478.640 1003.325 2479.820 1004.505 ;
        RECT 2881.890 870.830 2883.070 872.010 ;
        RECT 2883.490 870.830 2884.670 872.010 ;
        RECT 2885.090 870.830 2886.270 872.010 ;
        RECT 2886.690 870.830 2887.870 872.010 ;
        RECT 2912.355 870.830 2913.535 872.010 ;
        RECT 2913.955 870.830 2915.135 872.010 ;
        RECT 2915.555 870.830 2916.735 872.010 ;
        RECT 2917.155 870.830 2918.335 872.010 ;
        RECT 2918.755 870.830 2919.935 872.010 ;
        RECT 2920.355 870.830 2921.535 872.010 ;
        RECT 2921.955 870.830 2923.135 872.010 ;
        RECT 2923.555 870.830 2924.735 872.010 ;
        RECT 2925.155 870.830 2926.335 872.010 ;
        RECT 2880.910 750.770 2882.090 751.950 ;
        RECT 2882.510 750.770 2883.690 751.950 ;
        RECT 2912.355 750.750 2913.535 751.930 ;
        RECT 2913.955 750.750 2915.135 751.930 ;
        RECT 2915.555 750.750 2916.735 751.930 ;
        RECT 2917.155 750.750 2918.335 751.930 ;
        RECT 2918.755 750.750 2919.935 751.930 ;
        RECT 2920.355 750.750 2921.535 751.930 ;
        RECT 2921.955 750.750 2923.135 751.930 ;
        RECT 2923.555 750.750 2924.735 751.930 ;
        RECT 2925.155 750.750 2926.335 751.930 ;
        RECT 2871.100 620.790 2872.280 621.970 ;
        RECT 2872.700 620.790 2873.880 621.970 ;
        RECT 2874.300 620.790 2875.480 621.970 ;
        RECT 2875.900 620.790 2877.080 621.970 ;
        RECT 2877.500 620.790 2878.680 621.970 ;
        RECT 2879.100 620.790 2880.280 621.970 ;
        RECT 2880.700 620.790 2881.880 621.970 ;
        RECT 2882.300 620.790 2883.480 621.970 ;
        RECT 2912.225 620.810 2913.405 621.990 ;
        RECT 2913.825 620.810 2915.005 621.990 ;
        RECT 2915.425 620.810 2916.605 621.990 ;
        RECT 2917.025 620.810 2918.205 621.990 ;
        RECT 2918.625 620.810 2919.805 621.990 ;
        RECT 2920.225 620.810 2921.405 621.990 ;
        RECT 2921.825 620.810 2923.005 621.990 ;
        RECT 2923.425 620.810 2924.605 621.990 ;
        RECT 2925.025 620.810 2926.205 621.990 ;
        RECT 2871.150 490.760 2872.330 491.940 ;
        RECT 2872.750 490.760 2873.930 491.940 ;
        RECT 2874.350 490.760 2875.530 491.940 ;
        RECT 2875.950 490.760 2877.130 491.940 ;
        RECT 2877.550 490.760 2878.730 491.940 ;
        RECT 2879.150 490.760 2880.330 491.940 ;
        RECT 2880.750 490.760 2881.930 491.940 ;
        RECT 2882.350 490.760 2883.530 491.940 ;
        RECT 2912.355 490.730 2913.535 491.910 ;
        RECT 2913.955 490.730 2915.135 491.910 ;
        RECT 2915.555 490.730 2916.735 491.910 ;
        RECT 2917.155 490.730 2918.335 491.910 ;
        RECT 2918.755 490.730 2919.935 491.910 ;
        RECT 2920.355 490.730 2921.535 491.910 ;
        RECT 2921.955 490.730 2923.135 491.910 ;
        RECT 2923.555 490.730 2924.735 491.910 ;
        RECT 2925.155 490.730 2926.335 491.910 ;
        RECT 2871.160 360.790 2872.340 361.970 ;
        RECT 2872.760 360.790 2873.940 361.970 ;
        RECT 2874.360 360.790 2875.540 361.970 ;
        RECT 2875.960 360.790 2877.140 361.970 ;
        RECT 2877.560 360.790 2878.740 361.970 ;
        RECT 2879.160 360.790 2880.340 361.970 ;
        RECT 2880.760 360.790 2881.940 361.970 ;
        RECT 2882.360 360.790 2883.540 361.970 ;
        RECT 2912.375 360.790 2913.555 361.970 ;
        RECT 2913.975 360.790 2915.155 361.970 ;
        RECT 2915.575 360.790 2916.755 361.970 ;
        RECT 2917.175 360.790 2918.355 361.970 ;
        RECT 2918.775 360.790 2919.955 361.970 ;
        RECT 2920.375 360.790 2921.555 361.970 ;
        RECT 2921.975 360.790 2923.155 361.970 ;
        RECT 2923.575 360.790 2924.755 361.970 ;
        RECT 2925.175 360.790 2926.355 361.970 ;
        RECT 2954.950 311.135 2959.330 323.515 ;
        RECT 3109.005 311.445 3113.385 323.825 ;
        RECT 3151.185 313.925 3153.965 323.105 ;
        RECT 2871.130 230.840 2872.310 232.020 ;
        RECT 2872.730 230.840 2873.910 232.020 ;
        RECT 2874.330 230.840 2875.510 232.020 ;
        RECT 2875.930 230.840 2877.110 232.020 ;
        RECT 2877.530 230.840 2878.710 232.020 ;
        RECT 2879.130 230.840 2880.310 232.020 ;
        RECT 2880.730 230.840 2881.910 232.020 ;
        RECT 2882.330 230.840 2883.510 232.020 ;
        RECT 2912.345 230.850 2913.525 232.030 ;
        RECT 2913.945 230.850 2915.125 232.030 ;
        RECT 2915.545 230.850 2916.725 232.030 ;
        RECT 2917.145 230.850 2918.325 232.030 ;
        RECT 2918.745 230.850 2919.925 232.030 ;
        RECT 2920.345 230.850 2921.525 232.030 ;
        RECT 2921.945 230.850 2923.125 232.030 ;
        RECT 2923.545 230.850 2924.725 232.030 ;
        RECT 2925.145 230.850 2926.325 232.030 ;
        RECT 3127.245 208.275 3128.425 209.455 ;
        RECT 3127.245 206.675 3128.425 207.855 ;
        RECT 3127.245 205.075 3128.425 206.255 ;
        RECT 3142.715 208.295 3143.895 209.475 ;
        RECT 3142.715 206.695 3143.895 207.875 ;
        RECT 3142.715 205.095 3143.895 206.275 ;
        RECT 3158.255 208.315 3159.435 209.495 ;
        RECT 3158.255 206.715 3159.435 207.895 ;
        RECT 3158.255 205.115 3159.435 206.295 ;
        RECT 3173.775 208.275 3174.955 209.455 ;
        RECT 3173.775 206.675 3174.955 207.855 ;
        RECT 3173.775 205.075 3174.955 206.255 ;
        RECT 3189.285 208.405 3190.465 209.585 ;
        RECT 3189.285 206.805 3190.465 207.985 ;
        RECT 3189.285 205.205 3190.465 206.385 ;
        RECT 3211.335 64.370 3212.515 65.550 ;
        RECT 3212.935 64.370 3214.115 65.550 ;
        RECT 3214.535 64.370 3215.715 65.550 ;
        RECT 3216.135 64.370 3217.315 65.550 ;
        RECT 677.530 52.090 683.510 56.470 ;
        RECT 1179.015 44.755 1199.395 63.535 ;
        RECT 1227.275 44.825 1247.655 63.605 ;
      LAYER met5 ;
        RECT 209.070 882.990 224.070 1018.560 ;
        RECT 251.330 1002.830 2926.840 1017.830 ;
        RECT 2911.840 960.920 2926.840 1002.830 ;
        RECT 2911.840 951.460 3171.720 960.920 ;
        RECT 2911.840 950.910 3179.880 951.460 ;
        RECT 209.070 879.790 236.050 882.990 ;
        RECT 2843.120 879.790 2884.440 882.990 ;
        RECT 209.070 752.990 224.070 879.790 ;
        RECT 2881.240 873.010 2884.440 879.790 ;
        RECT 2881.240 869.810 2888.600 873.010 ;
        RECT 209.070 749.790 235.950 752.990 ;
        RECT 2843.120 749.790 2884.440 752.990 ;
        RECT 209.070 664.440 224.070 749.790 ;
        RECT 204.070 622.990 224.070 664.440 ;
        RECT 2911.840 741.550 2926.840 950.910 ;
        RECT 3167.220 949.860 3179.880 950.910 ;
        RECT 2911.840 739.950 2937.860 741.550 ;
        RECT 204.070 619.790 235.990 622.990 ;
        RECT 2843.120 619.790 2884.440 622.990 ;
        RECT 204.070 492.990 224.070 619.790 ;
        RECT 2911.840 588.370 2926.840 739.950 ;
        RECT 2911.840 586.770 2937.860 588.370 ;
        RECT 204.070 489.790 235.920 492.990 ;
        RECT 2843.120 489.790 2884.440 492.990 ;
        RECT 204.070 362.990 224.070 489.790 ;
        RECT 2911.840 435.190 2926.840 586.770 ;
        RECT 2911.840 433.590 2937.940 435.190 ;
        RECT 204.070 359.790 236.000 362.990 ;
        RECT 2843.120 359.790 2884.440 362.990 ;
        RECT 204.070 232.990 224.070 359.790 ;
        RECT 2911.840 325.280 2926.840 433.590 ;
        RECT 2911.840 310.280 3258.530 325.280 ;
        RECT 204.070 229.790 235.730 232.990 ;
        RECT 2843.120 229.790 2884.440 232.990 ;
        RECT 204.070 64.440 224.070 229.790 ;
        RECT 2911.840 66.440 2926.840 310.280 ;
        RECT 3094.010 277.870 3109.010 310.280 ;
        RECT 3224.860 293.450 3239.860 310.280 ;
        RECT 3224.860 291.850 3258.660 293.450 ;
        RECT 3224.860 285.290 3239.860 291.850 ;
        RECT 3224.860 283.690 3258.810 285.290 ;
        RECT 3224.860 283.110 3239.860 283.690 ;
        RECT 3094.010 276.270 3116.700 277.870 ;
        RECT 3094.010 275.560 3109.010 276.270 ;
        RECT 3097.980 209.840 3105.060 275.560 ;
        RECT 3097.980 204.840 3190.830 209.840 ;
        RECT 3097.980 189.480 3101.980 204.840 ;
        RECT 3097.980 187.880 3104.730 189.480 ;
        RECT 3097.980 172.580 3101.980 187.880 ;
        RECT 3097.980 170.980 3104.120 172.580 ;
        RECT 2911.840 64.440 3218.230 66.440 ;
        RECT 204.070 63.440 3218.230 64.440 ;
        RECT 204.070 44.440 2926.870 63.440 ;
    END
  END vssd_core
  PIN vccd2_core
    PORT
      LAYER met4 ;
        RECT 276.800 1173.190 279.900 1209.880 ;
        RECT 276.800 1170.090 296.150 1173.190 ;
        RECT 293.050 1037.830 296.150 1170.090 ;
        RECT 190.870 1022.830 296.150 1037.830 ;
        RECT 944.300 1022.830 945.960 1037.820 ;
        RECT 994.900 1022.830 996.560 1037.820 ;
        RECT 190.870 1002.830 203.900 1022.830 ;
        RECT 293.050 1022.500 296.150 1022.830 ;
        RECT 3232.580 1021.830 3235.680 1209.880 ;
      LAYER via4 ;
        RECT 191.930 1003.635 202.710 1036.815 ;
        RECT 252.720 1024.195 285.900 1036.575 ;
        RECT 293.955 1036.150 295.135 1037.330 ;
        RECT 293.955 1034.550 295.135 1035.730 ;
        RECT 293.955 1032.950 295.135 1034.130 ;
        RECT 293.955 1031.350 295.135 1032.530 ;
        RECT 293.955 1029.750 295.135 1030.930 ;
        RECT 293.955 1028.150 295.135 1029.330 ;
        RECT 293.955 1026.550 295.135 1027.730 ;
        RECT 293.955 1024.950 295.135 1026.130 ;
        RECT 293.955 1023.350 295.135 1024.530 ;
        RECT 944.540 1036.185 945.720 1037.365 ;
        RECT 944.540 1034.585 945.720 1035.765 ;
        RECT 944.540 1032.985 945.720 1034.165 ;
        RECT 944.540 1031.385 945.720 1032.565 ;
        RECT 944.540 1029.785 945.720 1030.965 ;
        RECT 944.540 1028.185 945.720 1029.365 ;
        RECT 944.540 1026.585 945.720 1027.765 ;
        RECT 944.540 1024.985 945.720 1026.165 ;
        RECT 944.540 1023.385 945.720 1024.565 ;
        RECT 995.140 1036.185 996.320 1037.365 ;
        RECT 995.140 1034.585 996.320 1035.765 ;
        RECT 995.140 1032.985 996.320 1034.165 ;
        RECT 995.140 1031.385 996.320 1032.565 ;
        RECT 995.140 1029.785 996.320 1030.965 ;
        RECT 995.140 1028.185 996.320 1029.365 ;
        RECT 995.140 1026.585 996.320 1027.765 ;
        RECT 995.140 1024.985 996.320 1026.165 ;
        RECT 995.140 1023.385 996.320 1024.565 ;
        RECT 3233.495 1036.175 3234.675 1037.355 ;
        RECT 3233.495 1034.575 3234.675 1035.755 ;
        RECT 3233.495 1032.975 3234.675 1034.155 ;
        RECT 3233.495 1031.375 3234.675 1032.555 ;
        RECT 3233.495 1029.775 3234.675 1030.955 ;
        RECT 3233.495 1028.175 3234.675 1029.355 ;
        RECT 3233.495 1026.575 3234.675 1027.755 ;
        RECT 3233.495 1024.975 3234.675 1026.155 ;
        RECT 3233.495 1023.375 3234.675 1024.555 ;
      LAYER met5 ;
        RECT 191.160 1003.160 203.480 1037.290 ;
        RECT 251.280 1022.830 3236.420 1037.830 ;
    END
  END vccd2_core
  PIN vssd2_core
    PORT
      LAYER met4 ;
        RECT 272.000 1168.390 275.100 1205.110 ;
        RECT 272.000 1165.290 291.350 1168.390 ;
        RECT 288.250 1057.830 291.350 1165.290 ;
        RECT 174.810 1042.830 291.350 1057.830 ;
        RECT 965.200 1042.830 966.860 1057.820 ;
        RECT 1015.500 1042.840 1017.160 1057.830 ;
        RECT 174.810 1021.830 187.950 1042.830 ;
        RECT 288.250 1042.290 291.350 1042.830 ;
        RECT 3237.380 1042.310 3240.480 1205.080 ;
      LAYER via4 ;
        RECT 175.990 1022.485 186.770 1057.265 ;
        RECT 252.645 1044.025 285.825 1056.405 ;
        RECT 289.205 1056.170 290.385 1057.350 ;
        RECT 289.205 1054.570 290.385 1055.750 ;
        RECT 289.205 1052.970 290.385 1054.150 ;
        RECT 289.205 1051.370 290.385 1052.550 ;
        RECT 289.205 1049.770 290.385 1050.950 ;
        RECT 289.205 1048.170 290.385 1049.350 ;
        RECT 289.205 1046.570 290.385 1047.750 ;
        RECT 289.205 1044.970 290.385 1046.150 ;
        RECT 289.205 1043.370 290.385 1044.550 ;
        RECT 965.440 1056.185 966.620 1057.365 ;
        RECT 965.440 1054.585 966.620 1055.765 ;
        RECT 965.440 1052.985 966.620 1054.165 ;
        RECT 965.440 1051.385 966.620 1052.565 ;
        RECT 965.440 1049.785 966.620 1050.965 ;
        RECT 965.440 1048.185 966.620 1049.365 ;
        RECT 965.440 1046.585 966.620 1047.765 ;
        RECT 965.440 1044.985 966.620 1046.165 ;
        RECT 965.440 1043.385 966.620 1044.565 ;
        RECT 1015.740 1056.195 1016.920 1057.375 ;
        RECT 1015.740 1054.595 1016.920 1055.775 ;
        RECT 1015.740 1052.995 1016.920 1054.175 ;
        RECT 1015.740 1051.395 1016.920 1052.575 ;
        RECT 1015.740 1049.795 1016.920 1050.975 ;
        RECT 1015.740 1048.195 1016.920 1049.375 ;
        RECT 1015.740 1046.595 1016.920 1047.775 ;
        RECT 1015.740 1044.995 1016.920 1046.175 ;
        RECT 1015.740 1043.395 1016.920 1044.575 ;
        RECT 3238.285 1056.185 3239.465 1057.365 ;
        RECT 3238.285 1054.585 3239.465 1055.765 ;
        RECT 3238.285 1052.985 3239.465 1054.165 ;
        RECT 3238.285 1051.385 3239.465 1052.565 ;
        RECT 3238.285 1049.785 3239.465 1050.965 ;
        RECT 3238.285 1048.185 3239.465 1049.365 ;
        RECT 3238.285 1046.585 3239.465 1047.765 ;
        RECT 3238.285 1044.985 3239.465 1046.165 ;
        RECT 3238.285 1043.385 3239.465 1044.565 ;
      LAYER met5 ;
        RECT 175.220 1022.310 187.540 1057.440 ;
        RECT 251.280 1042.830 3241.000 1057.830 ;
    END
  END vssd2_core
  PIN vdda2_core
    PORT
      LAYER met3 ;
        RECT 169.510 2295.890 231.350 2319.790 ;
        RECT 169.510 2245.995 231.350 2269.895 ;
      LAYER via3 ;
        RECT 221.870 2296.795 230.190 2319.115 ;
        RECT 221.810 2246.845 230.130 2269.165 ;
      LAYER met4 ;
        RECT 220.860 4774.180 252.060 4777.240 ;
        RECT 220.750 2295.920 230.870 2319.870 ;
        RECT 220.880 2245.970 231.000 2269.920 ;
        RECT 220.820 1193.690 230.880 1197.690 ;
        RECT 220.820 1190.630 251.920 1193.690 ;
        RECT 257.600 1153.990 260.700 1190.710 ;
        RECT 257.600 1150.890 276.950 1153.990 ;
        RECT 273.850 1117.830 276.950 1150.890 ;
        RECT 220.740 1102.830 276.950 1117.830 ;
        RECT 273.850 1102.610 276.950 1102.830 ;
        RECT 1892.820 1102.760 1898.430 1117.850 ;
        RECT 1968.320 1102.760 1973.930 1117.850 ;
        RECT 3251.780 1102.430 3254.880 1190.680 ;
      LAYER via4 ;
        RECT 221.290 4775.125 222.470 4776.305 ;
        RECT 222.890 4775.125 224.070 4776.305 ;
        RECT 224.490 4775.125 225.670 4776.305 ;
        RECT 226.090 4775.125 227.270 4776.305 ;
        RECT 227.690 4775.125 228.870 4776.305 ;
        RECT 229.290 4775.125 230.470 4776.305 ;
        RECT 249.055 4775.150 250.235 4776.330 ;
        RECT 250.655 4775.150 251.835 4776.330 ;
        RECT 222.240 2296.965 229.820 2318.945 ;
        RECT 222.180 2247.015 229.760 2268.995 ;
        RECT 221.255 1191.180 230.435 1197.160 ;
        RECT 248.900 1190.785 251.680 1193.565 ;
        RECT 222.245 1104.345 229.825 1116.725 ;
        RECT 252.710 1104.040 271.490 1116.420 ;
        RECT 274.790 1116.130 275.970 1117.310 ;
        RECT 274.790 1114.530 275.970 1115.710 ;
        RECT 274.790 1112.930 275.970 1114.110 ;
        RECT 274.790 1111.330 275.970 1112.510 ;
        RECT 274.790 1109.730 275.970 1110.910 ;
        RECT 274.790 1108.130 275.970 1109.310 ;
        RECT 274.790 1106.530 275.970 1107.710 ;
        RECT 274.790 1104.930 275.970 1106.110 ;
        RECT 274.790 1103.330 275.970 1104.510 ;
        RECT 1893.465 1103.350 1897.845 1117.330 ;
        RECT 1968.965 1103.350 1973.345 1117.330 ;
        RECT 3252.695 1116.095 3253.875 1117.275 ;
        RECT 3252.695 1114.495 3253.875 1115.675 ;
        RECT 3252.695 1112.895 3253.875 1114.075 ;
        RECT 3252.695 1111.295 3253.875 1112.475 ;
        RECT 3252.695 1109.695 3253.875 1110.875 ;
        RECT 3252.695 1108.095 3253.875 1109.275 ;
        RECT 3252.695 1106.495 3253.875 1107.675 ;
        RECT 3252.695 1104.895 3253.875 1106.075 ;
        RECT 3252.695 1103.295 3253.875 1104.475 ;
      LAYER met5 ;
        RECT 220.880 1102.990 230.880 4782.830 ;
        RECT 248.770 4774.140 257.650 4777.240 ;
        RECT 248.660 1190.620 257.620 1193.720 ;
        RECT 251.740 1102.830 3255.270 1117.830 ;
    END
  END vdda2_core
  PIN vssa2_core
    PORT
      LAYER met3 ;
        RECT 169.150 4018.890 219.900 4042.790 ;
        RECT 169.150 3968.995 219.900 3992.895 ;
      LAYER via3 ;
        RECT 209.535 4019.650 218.255 4041.970 ;
        RECT 209.535 3969.990 218.255 3992.310 ;
      LAYER met4 ;
        RECT 208.870 4778.960 252.800 4782.050 ;
        RECT 208.850 4018.790 219.000 4042.810 ;
        RECT 208.850 3969.010 219.000 3993.030 ;
        RECT 208.850 1185.910 252.970 1188.940 ;
        RECT 208.850 1185.790 255.900 1185.910 ;
        RECT 208.850 1181.790 218.900 1185.790 ;
        RECT 252.750 1137.830 255.900 1185.790 ;
        RECT 208.740 1122.830 267.240 1137.830 ;
        RECT 1929.610 1122.840 1934.120 1137.750 ;
        RECT 2005.210 1122.840 2009.720 1137.750 ;
        RECT 3256.580 1122.450 3259.680 1185.910 ;
      LAYER via4 ;
        RECT 209.260 4779.945 210.440 4781.125 ;
        RECT 210.860 4779.945 212.040 4781.125 ;
        RECT 212.460 4779.945 213.640 4781.125 ;
        RECT 214.060 4779.945 215.240 4781.125 ;
        RECT 215.660 4779.945 216.840 4781.125 ;
        RECT 217.260 4779.945 218.440 4781.125 ;
        RECT 249.035 4779.950 250.215 4781.130 ;
        RECT 250.635 4779.950 251.815 4781.130 ;
        RECT 210.105 4019.820 217.685 4041.800 ;
        RECT 210.105 3970.160 217.685 3992.140 ;
        RECT 209.285 1182.415 218.465 1188.395 ;
        RECT 249.170 1185.970 251.950 1188.750 ;
        RECT 210.245 1124.345 217.825 1136.725 ;
        RECT 252.665 1124.040 266.645 1136.420 ;
        RECT 1930.475 1124.065 1933.255 1136.445 ;
        RECT 2006.075 1124.065 2008.855 1136.445 ;
        RECT 3257.505 1136.185 3258.685 1137.365 ;
        RECT 3257.505 1134.585 3258.685 1135.765 ;
        RECT 3257.505 1132.985 3258.685 1134.165 ;
        RECT 3257.505 1131.385 3258.685 1132.565 ;
        RECT 3257.505 1129.785 3258.685 1130.965 ;
        RECT 3257.505 1128.185 3258.685 1129.365 ;
        RECT 3257.505 1126.585 3258.685 1127.765 ;
        RECT 3257.505 1124.985 3258.685 1126.165 ;
        RECT 3257.505 1123.385 3258.685 1124.565 ;
      LAYER met5 ;
        RECT 208.880 1122.920 218.880 4782.830 ;
        RECT 248.770 4778.940 252.870 4782.040 ;
        RECT 248.660 1185.820 252.840 1188.920 ;
        RECT 251.740 1122.830 3260.340 1137.830 ;
    END
  END vssa2_core
  PIN vssd1_core
    PORT
      LAYER met3 ;
        RECT 535.800 4808.010 541.800 4982.910 ;
        RECT 792.800 4808.010 798.800 4982.910 ;
        RECT 1049.800 4808.010 1055.800 4982.910 ;
        RECT 1306.800 4808.010 1312.800 4982.910 ;
        RECT 1564.800 4808.010 1570.800 4982.910 ;
        RECT 1816.800 4808.010 1822.800 4982.910 ;
        RECT 2153.800 4808.010 2159.800 4982.910 ;
        RECT 2538.800 4808.010 2544.800 4982.910 ;
        RECT 2795.800 4808.010 2801.800 4982.910 ;
        RECT 6.070 4571.410 252.940 4572.410 ;
        RECT 6.070 4566.410 284.610 4571.410 ;
        RECT 247.050 4565.410 284.610 4566.410 ;
        RECT 6.070 3937.410 284.610 3943.410 ;
        RECT 6.070 3721.410 284.610 3727.410 ;
        RECT 6.070 3505.410 284.610 3511.410 ;
        RECT 6.070 3289.410 284.610 3295.410 ;
        RECT 6.070 3073.410 284.610 3079.410 ;
        RECT 6.070 2857.410 284.610 2863.410 ;
        RECT 6.070 2641.410 284.610 2647.410 ;
        RECT 6.070 2003.410 284.610 2009.410 ;
        RECT 6.070 1787.410 284.610 1793.410 ;
        RECT 6.070 1571.410 284.610 1577.410 ;
        RECT 6.070 1355.410 284.610 1361.410 ;
        RECT 6.070 1139.410 238.970 1145.410 ;
        RECT 6.070 923.410 238.970 929.410 ;
      LAYER via3 ;
        RECT 536.055 4979.030 541.575 4982.150 ;
        RECT 536.225 4808.565 541.345 4813.685 ;
        RECT 793.055 4979.030 798.575 4982.150 ;
        RECT 793.225 4808.565 798.345 4813.685 ;
        RECT 1050.055 4979.030 1055.575 4982.150 ;
        RECT 1050.225 4808.565 1055.345 4813.685 ;
        RECT 1307.055 4979.030 1312.575 4982.150 ;
        RECT 1307.225 4808.565 1312.345 4813.685 ;
        RECT 1565.055 4979.030 1570.575 4982.150 ;
        RECT 1565.225 4808.565 1570.345 4813.685 ;
        RECT 1817.055 4979.030 1822.575 4982.150 ;
        RECT 1817.225 4808.565 1822.345 4813.685 ;
        RECT 2154.055 4979.030 2159.575 4982.150 ;
        RECT 2154.225 4808.565 2159.345 4813.685 ;
        RECT 2539.055 4979.030 2544.575 4982.150 ;
        RECT 2539.225 4808.565 2544.345 4813.685 ;
        RECT 2796.055 4979.030 2801.575 4982.150 ;
        RECT 2796.225 4808.565 2801.345 4813.685 ;
        RECT 6.830 4566.665 9.950 4572.185 ;
        RECT 233.295 4566.835 238.415 4571.955 ;
        RECT 281.945 4565.585 284.265 4571.105 ;
        RECT 6.830 3937.665 9.950 3943.185 ;
        RECT 233.295 3937.835 238.415 3942.955 ;
        RECT 281.945 3937.585 284.265 3943.105 ;
        RECT 6.830 3721.665 9.950 3727.185 ;
        RECT 233.295 3721.835 238.415 3726.955 ;
        RECT 281.945 3721.585 284.265 3727.105 ;
        RECT 6.830 3505.665 9.950 3511.185 ;
        RECT 233.295 3505.835 238.415 3510.955 ;
        RECT 281.945 3505.585 284.265 3511.105 ;
        RECT 6.830 3289.665 9.950 3295.185 ;
        RECT 233.295 3289.835 238.415 3294.955 ;
        RECT 281.945 3289.585 284.265 3295.105 ;
        RECT 6.830 3073.665 9.950 3079.185 ;
        RECT 233.295 3073.835 238.415 3078.955 ;
        RECT 281.945 3073.585 284.265 3079.105 ;
        RECT 6.830 2857.665 9.950 2863.185 ;
        RECT 233.295 2857.835 238.415 2862.955 ;
        RECT 281.945 2857.585 284.265 2863.105 ;
        RECT 6.830 2641.665 9.950 2647.185 ;
        RECT 233.295 2641.835 238.415 2646.955 ;
        RECT 281.945 2641.585 284.265 2647.105 ;
        RECT 6.830 2003.665 9.950 2009.185 ;
        RECT 233.295 2003.835 238.415 2008.955 ;
        RECT 281.945 2003.585 284.265 2009.105 ;
        RECT 6.830 1787.665 9.950 1793.185 ;
        RECT 233.295 1787.835 238.415 1792.955 ;
        RECT 281.945 1787.585 284.265 1793.105 ;
        RECT 6.830 1571.665 9.950 1577.185 ;
        RECT 233.295 1571.835 238.415 1576.955 ;
        RECT 281.945 1571.585 284.265 1577.105 ;
        RECT 6.830 1355.665 9.950 1361.185 ;
        RECT 233.295 1355.835 238.415 1360.955 ;
        RECT 281.945 1355.585 284.265 1361.105 ;
        RECT 6.830 1139.665 9.950 1145.185 ;
        RECT 233.295 1139.835 238.415 1144.955 ;
        RECT 6.830 923.665 9.950 929.185 ;
        RECT 233.295 923.835 238.415 928.955 ;
      LAYER met4 ;
        RECT 475.270 4978.560 542.100 4982.560 ;
        RECT 732.270 4978.560 799.100 4982.560 ;
        RECT 989.270 4978.560 1056.100 4982.560 ;
        RECT 1246.270 4978.560 1313.100 4982.560 ;
        RECT 1504.270 4978.560 1571.100 4982.560 ;
        RECT 1756.270 4978.560 1823.100 4982.560 ;
        RECT 2093.270 4978.560 2160.100 4982.560 ;
        RECT 2478.270 4978.560 2545.100 4982.560 ;
        RECT 2735.270 4978.560 2802.100 4982.560 ;
        RECT 535.760 4808.160 541.830 4814.190 ;
        RECT 792.760 4808.160 798.830 4814.190 ;
        RECT 1049.760 4808.160 1055.830 4814.190 ;
        RECT 1306.760 4808.160 1312.830 4814.190 ;
        RECT 1564.760 4808.160 1570.830 4814.190 ;
        RECT 1816.760 4808.160 1822.830 4814.190 ;
        RECT 2153.760 4808.160 2159.830 4814.190 ;
        RECT 2538.760 4808.160 2544.830 4814.190 ;
        RECT 2795.760 4808.160 2801.830 4814.190 ;
        RECT 3323.970 4813.960 3337.020 4813.980 ;
        RECT 3323.930 4807.960 3353.160 4813.960 ;
        RECT 3323.970 4781.500 3337.020 4807.960 ;
        RECT 232.870 4750.140 251.910 4753.240 ;
        RECT 6.420 4505.880 10.420 4572.710 ;
        RECT 232.790 4566.370 238.820 4572.440 ;
        RECT 281.800 4565.570 284.410 4571.120 ;
        RECT 6.420 3876.880 10.420 3943.710 ;
        RECT 232.790 3937.370 238.820 3943.440 ;
        RECT 281.800 3937.570 284.410 3943.120 ;
        RECT 6.420 3660.880 10.420 3727.710 ;
        RECT 232.790 3721.370 238.820 3727.440 ;
        RECT 281.800 3721.570 284.410 3727.120 ;
        RECT 6.420 3444.880 10.420 3511.710 ;
        RECT 232.790 3505.370 238.820 3511.440 ;
        RECT 281.800 3505.570 284.410 3511.120 ;
        RECT 6.420 3228.880 10.420 3295.710 ;
        RECT 232.790 3289.370 238.820 3295.440 ;
        RECT 281.800 3289.570 284.410 3295.120 ;
        RECT 6.420 3012.880 10.420 3079.710 ;
        RECT 232.790 3073.370 238.820 3079.440 ;
        RECT 281.800 3073.570 284.410 3079.120 ;
        RECT 6.420 2796.880 10.420 2863.710 ;
        RECT 232.790 2857.370 238.820 2863.440 ;
        RECT 281.800 2857.570 284.410 2863.120 ;
        RECT 6.420 2580.880 10.420 2647.710 ;
        RECT 232.790 2641.370 238.820 2647.440 ;
        RECT 281.800 2641.570 284.410 2647.120 ;
        RECT 6.420 1942.880 10.420 2009.710 ;
        RECT 232.790 2003.370 238.820 2009.440 ;
        RECT 281.800 2003.570 284.410 2009.120 ;
        RECT 6.420 1726.880 10.420 1793.710 ;
        RECT 232.790 1787.370 238.820 1793.440 ;
        RECT 281.800 1787.570 284.410 1793.120 ;
        RECT 6.420 1510.880 10.420 1577.710 ;
        RECT 232.790 1571.370 238.820 1577.440 ;
        RECT 281.800 1571.570 284.410 1577.120 ;
        RECT 6.420 1294.880 10.420 1361.710 ;
        RECT 232.790 1355.370 238.820 1361.440 ;
        RECT 281.800 1355.570 284.410 1361.120 ;
        RECT 232.800 1217.730 238.890 1220.730 ;
        RECT 232.800 1214.610 251.970 1217.730 ;
        RECT 281.600 1177.990 284.700 1214.670 ;
        RECT 281.600 1174.890 300.950 1177.990 ;
        RECT 6.420 1078.880 10.420 1145.710 ;
        RECT 232.790 1139.370 238.820 1145.440 ;
        RECT 232.780 1082.830 286.350 1097.830 ;
        RECT 297.850 1082.430 300.950 1174.890 ;
        RECT 1353.500 1082.850 1356.190 1097.860 ;
        RECT 1428.500 1082.850 1431.190 1097.860 ;
        RECT 1503.700 1082.850 1506.390 1097.860 ;
        RECT 1579.300 1082.850 1581.990 1097.860 ;
        RECT 3227.780 1082.460 3230.880 1214.720 ;
        RECT 6.420 862.880 10.420 929.710 ;
        RECT 232.790 923.370 238.820 929.440 ;
      LAYER via4 ;
        RECT 475.685 4980.785 476.865 4981.965 ;
        RECT 492.600 4980.785 493.780 4981.965 ;
        RECT 509.480 4980.775 510.660 4981.955 ;
        RECT 475.685 4979.185 476.865 4980.365 ;
        RECT 492.600 4979.185 493.780 4980.365 ;
        RECT 509.480 4979.175 510.660 4980.355 ;
        RECT 732.685 4980.785 733.865 4981.965 ;
        RECT 749.600 4980.785 750.780 4981.965 ;
        RECT 766.480 4980.775 767.660 4981.955 ;
        RECT 732.685 4979.185 733.865 4980.365 ;
        RECT 749.600 4979.185 750.780 4980.365 ;
        RECT 766.480 4979.175 767.660 4980.355 ;
        RECT 989.685 4980.785 990.865 4981.965 ;
        RECT 1006.600 4980.785 1007.780 4981.965 ;
        RECT 1023.480 4980.775 1024.660 4981.955 ;
        RECT 989.685 4979.185 990.865 4980.365 ;
        RECT 1006.600 4979.185 1007.780 4980.365 ;
        RECT 1023.480 4979.175 1024.660 4980.355 ;
        RECT 1246.685 4980.785 1247.865 4981.965 ;
        RECT 1263.600 4980.785 1264.780 4981.965 ;
        RECT 1280.480 4980.775 1281.660 4981.955 ;
        RECT 1246.685 4979.185 1247.865 4980.365 ;
        RECT 1263.600 4979.185 1264.780 4980.365 ;
        RECT 1280.480 4979.175 1281.660 4980.355 ;
        RECT 1504.685 4980.785 1505.865 4981.965 ;
        RECT 1521.600 4980.785 1522.780 4981.965 ;
        RECT 1538.480 4980.775 1539.660 4981.955 ;
        RECT 1504.685 4979.185 1505.865 4980.365 ;
        RECT 1521.600 4979.185 1522.780 4980.365 ;
        RECT 1538.480 4979.175 1539.660 4980.355 ;
        RECT 1756.685 4980.785 1757.865 4981.965 ;
        RECT 1773.600 4980.785 1774.780 4981.965 ;
        RECT 1790.480 4980.775 1791.660 4981.955 ;
        RECT 1756.685 4979.185 1757.865 4980.365 ;
        RECT 1773.600 4979.185 1774.780 4980.365 ;
        RECT 1790.480 4979.175 1791.660 4980.355 ;
        RECT 2093.685 4980.785 2094.865 4981.965 ;
        RECT 2110.600 4980.785 2111.780 4981.965 ;
        RECT 2127.480 4980.775 2128.660 4981.955 ;
        RECT 2093.685 4979.185 2094.865 4980.365 ;
        RECT 2110.600 4979.185 2111.780 4980.365 ;
        RECT 2127.480 4979.175 2128.660 4980.355 ;
        RECT 2478.685 4980.785 2479.865 4981.965 ;
        RECT 2495.600 4980.785 2496.780 4981.965 ;
        RECT 2512.480 4980.775 2513.660 4981.955 ;
        RECT 2478.685 4979.185 2479.865 4980.365 ;
        RECT 2495.600 4979.185 2496.780 4980.365 ;
        RECT 2512.480 4979.175 2513.660 4980.355 ;
        RECT 2735.685 4980.785 2736.865 4981.965 ;
        RECT 2752.600 4980.785 2753.780 4981.965 ;
        RECT 2769.480 4980.775 2770.660 4981.955 ;
        RECT 2735.685 4979.185 2736.865 4980.365 ;
        RECT 2752.600 4979.185 2753.780 4980.365 ;
        RECT 2769.480 4979.175 2770.660 4980.355 ;
        RECT 536.595 4808.935 540.975 4813.315 ;
        RECT 793.595 4808.935 797.975 4813.315 ;
        RECT 1050.595 4808.935 1054.975 4813.315 ;
        RECT 1307.595 4808.935 1311.975 4813.315 ;
        RECT 1565.595 4808.935 1569.975 4813.315 ;
        RECT 1817.595 4808.935 1821.975 4813.315 ;
        RECT 2154.595 4808.935 2158.975 4813.315 ;
        RECT 2539.595 4808.935 2543.975 4813.315 ;
        RECT 2796.595 4808.935 2800.975 4813.315 ;
        RECT 3325.070 4808.840 3351.850 4813.220 ;
        RECT 3325.100 4782.320 3335.880 4793.100 ;
        RECT 233.685 4751.105 234.865 4752.285 ;
        RECT 235.285 4751.105 236.465 4752.285 ;
        RECT 236.885 4751.105 238.065 4752.285 ;
        RECT 248.945 4750.305 251.725 4753.085 ;
        RECT 233.665 4567.205 238.045 4571.585 ;
        RECT 7.025 4540.095 8.205 4541.275 ;
        RECT 8.625 4540.095 9.805 4541.275 ;
        RECT 7.030 4523.195 8.210 4524.375 ;
        RECT 8.630 4523.195 9.810 4524.375 ;
        RECT 7.015 4506.295 8.195 4507.475 ;
        RECT 8.615 4506.295 9.795 4507.475 ;
        RECT 233.665 3938.205 238.045 3942.585 ;
        RECT 7.025 3911.095 8.205 3912.275 ;
        RECT 8.625 3911.095 9.805 3912.275 ;
        RECT 7.030 3894.195 8.210 3895.375 ;
        RECT 8.630 3894.195 9.810 3895.375 ;
        RECT 7.015 3877.295 8.195 3878.475 ;
        RECT 8.615 3877.295 9.795 3878.475 ;
        RECT 233.665 3722.205 238.045 3726.585 ;
        RECT 7.025 3695.095 8.205 3696.275 ;
        RECT 8.625 3695.095 9.805 3696.275 ;
        RECT 7.030 3678.195 8.210 3679.375 ;
        RECT 8.630 3678.195 9.810 3679.375 ;
        RECT 7.015 3661.295 8.195 3662.475 ;
        RECT 8.615 3661.295 9.795 3662.475 ;
        RECT 233.665 3506.205 238.045 3510.585 ;
        RECT 7.025 3479.095 8.205 3480.275 ;
        RECT 8.625 3479.095 9.805 3480.275 ;
        RECT 7.030 3462.195 8.210 3463.375 ;
        RECT 8.630 3462.195 9.810 3463.375 ;
        RECT 7.015 3445.295 8.195 3446.475 ;
        RECT 8.615 3445.295 9.795 3446.475 ;
        RECT 233.665 3290.205 238.045 3294.585 ;
        RECT 7.025 3263.095 8.205 3264.275 ;
        RECT 8.625 3263.095 9.805 3264.275 ;
        RECT 7.030 3246.195 8.210 3247.375 ;
        RECT 8.630 3246.195 9.810 3247.375 ;
        RECT 7.015 3229.295 8.195 3230.475 ;
        RECT 8.615 3229.295 9.795 3230.475 ;
        RECT 233.665 3074.205 238.045 3078.585 ;
        RECT 7.025 3047.095 8.205 3048.275 ;
        RECT 8.625 3047.095 9.805 3048.275 ;
        RECT 7.030 3030.195 8.210 3031.375 ;
        RECT 8.630 3030.195 9.810 3031.375 ;
        RECT 7.015 3013.295 8.195 3014.475 ;
        RECT 8.615 3013.295 9.795 3014.475 ;
        RECT 233.665 2858.205 238.045 2862.585 ;
        RECT 7.025 2831.095 8.205 2832.275 ;
        RECT 8.625 2831.095 9.805 2832.275 ;
        RECT 7.030 2814.195 8.210 2815.375 ;
        RECT 8.630 2814.195 9.810 2815.375 ;
        RECT 7.015 2797.295 8.195 2798.475 ;
        RECT 8.615 2797.295 9.795 2798.475 ;
        RECT 233.665 2642.205 238.045 2646.585 ;
        RECT 7.025 2615.095 8.205 2616.275 ;
        RECT 8.625 2615.095 9.805 2616.275 ;
        RECT 7.030 2598.195 8.210 2599.375 ;
        RECT 8.630 2598.195 9.810 2599.375 ;
        RECT 7.015 2581.295 8.195 2582.475 ;
        RECT 8.615 2581.295 9.795 2582.475 ;
        RECT 233.665 2004.205 238.045 2008.585 ;
        RECT 7.025 1977.095 8.205 1978.275 ;
        RECT 8.625 1977.095 9.805 1978.275 ;
        RECT 7.030 1960.195 8.210 1961.375 ;
        RECT 8.630 1960.195 9.810 1961.375 ;
        RECT 7.015 1943.295 8.195 1944.475 ;
        RECT 8.615 1943.295 9.795 1944.475 ;
        RECT 233.665 1788.205 238.045 1792.585 ;
        RECT 7.025 1761.095 8.205 1762.275 ;
        RECT 8.625 1761.095 9.805 1762.275 ;
        RECT 7.030 1744.195 8.210 1745.375 ;
        RECT 8.630 1744.195 9.810 1745.375 ;
        RECT 7.015 1727.295 8.195 1728.475 ;
        RECT 8.615 1727.295 9.795 1728.475 ;
        RECT 233.665 1572.205 238.045 1576.585 ;
        RECT 7.025 1545.095 8.205 1546.275 ;
        RECT 8.625 1545.095 9.805 1546.275 ;
        RECT 7.030 1528.195 8.210 1529.375 ;
        RECT 8.630 1528.195 9.810 1529.375 ;
        RECT 7.015 1511.295 8.195 1512.475 ;
        RECT 8.615 1511.295 9.795 1512.475 ;
        RECT 233.665 1356.205 238.045 1360.585 ;
        RECT 7.025 1329.095 8.205 1330.275 ;
        RECT 8.625 1329.095 9.805 1330.275 ;
        RECT 7.030 1312.195 8.210 1313.375 ;
        RECT 8.630 1312.195 9.810 1313.375 ;
        RECT 7.015 1295.295 8.195 1296.475 ;
        RECT 8.615 1295.295 9.795 1296.475 ;
        RECT 233.655 1215.550 238.035 1219.930 ;
        RECT 248.920 1214.795 251.700 1217.575 ;
        RECT 233.665 1140.205 238.045 1144.585 ;
        RECT 7.025 1113.095 8.205 1114.275 ;
        RECT 8.625 1113.095 9.805 1114.275 ;
        RECT 7.030 1096.195 8.210 1097.375 ;
        RECT 8.630 1096.195 9.810 1097.375 ;
        RECT 233.700 1083.360 238.080 1097.340 ;
        RECT 251.050 1083.370 285.830 1097.350 ;
        RECT 298.765 1096.110 299.945 1097.290 ;
        RECT 298.765 1094.510 299.945 1095.690 ;
        RECT 298.765 1092.910 299.945 1094.090 ;
        RECT 298.765 1091.310 299.945 1092.490 ;
        RECT 298.765 1089.710 299.945 1090.890 ;
        RECT 298.765 1088.110 299.945 1089.290 ;
        RECT 298.765 1086.510 299.945 1087.690 ;
        RECT 298.765 1084.910 299.945 1086.090 ;
        RECT 298.765 1083.310 299.945 1084.490 ;
        RECT 1354.025 1096.200 1355.205 1097.380 ;
        RECT 1354.025 1094.600 1355.205 1095.780 ;
        RECT 1354.025 1093.000 1355.205 1094.180 ;
        RECT 1354.025 1091.400 1355.205 1092.580 ;
        RECT 1354.025 1089.800 1355.205 1090.980 ;
        RECT 1354.025 1088.200 1355.205 1089.380 ;
        RECT 1354.025 1086.600 1355.205 1087.780 ;
        RECT 1354.025 1085.000 1355.205 1086.180 ;
        RECT 1354.025 1083.400 1355.205 1084.580 ;
        RECT 1429.025 1096.200 1430.205 1097.380 ;
        RECT 1429.025 1094.600 1430.205 1095.780 ;
        RECT 1429.025 1093.000 1430.205 1094.180 ;
        RECT 1429.025 1091.400 1430.205 1092.580 ;
        RECT 1429.025 1089.800 1430.205 1090.980 ;
        RECT 1429.025 1088.200 1430.205 1089.380 ;
        RECT 1429.025 1086.600 1430.205 1087.780 ;
        RECT 1429.025 1085.000 1430.205 1086.180 ;
        RECT 1429.025 1083.400 1430.205 1084.580 ;
        RECT 1504.225 1096.200 1505.405 1097.380 ;
        RECT 1504.225 1094.600 1505.405 1095.780 ;
        RECT 1504.225 1093.000 1505.405 1094.180 ;
        RECT 1504.225 1091.400 1505.405 1092.580 ;
        RECT 1504.225 1089.800 1505.405 1090.980 ;
        RECT 1504.225 1088.200 1505.405 1089.380 ;
        RECT 1504.225 1086.600 1505.405 1087.780 ;
        RECT 1504.225 1085.000 1505.405 1086.180 ;
        RECT 1504.225 1083.400 1505.405 1084.580 ;
        RECT 1579.825 1096.200 1581.005 1097.380 ;
        RECT 1579.825 1094.600 1581.005 1095.780 ;
        RECT 1579.825 1093.000 1581.005 1094.180 ;
        RECT 1579.825 1091.400 1581.005 1092.580 ;
        RECT 1579.825 1089.800 1581.005 1090.980 ;
        RECT 1579.825 1088.200 1581.005 1089.380 ;
        RECT 1579.825 1086.600 1581.005 1087.780 ;
        RECT 1579.825 1085.000 1581.005 1086.180 ;
        RECT 1579.825 1083.400 1581.005 1084.580 ;
        RECT 3227.960 1083.305 3230.740 1097.285 ;
        RECT 7.015 1079.295 8.195 1080.475 ;
        RECT 8.615 1079.295 9.795 1080.475 ;
        RECT 233.665 924.205 238.045 928.585 ;
        RECT 7.025 897.095 8.205 898.275 ;
        RECT 8.625 897.095 9.805 898.275 ;
        RECT 7.030 880.195 8.210 881.375 ;
        RECT 8.630 880.195 9.810 881.375 ;
        RECT 7.015 863.295 8.195 864.475 ;
        RECT 8.615 863.295 9.795 864.475 ;
      LAYER met5 ;
        RECT 475.400 4978.480 477.150 4982.640 ;
        RECT 475.480 4976.020 477.080 4978.480 ;
        RECT 492.290 4978.440 494.020 4982.820 ;
        RECT 509.230 4978.470 510.960 4982.850 ;
        RECT 732.400 4978.480 734.150 4982.640 ;
        RECT 492.380 4976.180 493.980 4978.440 ;
        RECT 509.280 4976.180 510.880 4978.470 ;
        RECT 732.480 4976.020 734.080 4978.480 ;
        RECT 749.290 4978.440 751.020 4982.820 ;
        RECT 766.230 4978.470 767.960 4982.850 ;
        RECT 989.400 4978.480 991.150 4982.640 ;
        RECT 749.380 4976.180 750.980 4978.440 ;
        RECT 766.280 4976.180 767.880 4978.470 ;
        RECT 989.480 4976.020 991.080 4978.480 ;
        RECT 1006.290 4978.440 1008.020 4982.820 ;
        RECT 1023.230 4978.470 1024.960 4982.850 ;
        RECT 1246.400 4978.480 1248.150 4982.640 ;
        RECT 1006.380 4976.180 1007.980 4978.440 ;
        RECT 1023.280 4976.180 1024.880 4978.470 ;
        RECT 1246.480 4976.020 1248.080 4978.480 ;
        RECT 1263.290 4978.440 1265.020 4982.820 ;
        RECT 1280.230 4978.470 1281.960 4982.850 ;
        RECT 1504.400 4978.480 1506.150 4982.640 ;
        RECT 1263.380 4976.180 1264.980 4978.440 ;
        RECT 1280.280 4976.180 1281.880 4978.470 ;
        RECT 1504.480 4976.020 1506.080 4978.480 ;
        RECT 1521.290 4978.440 1523.020 4982.820 ;
        RECT 1538.230 4978.470 1539.960 4982.850 ;
        RECT 1756.400 4978.480 1758.150 4982.640 ;
        RECT 1521.380 4976.180 1522.980 4978.440 ;
        RECT 1538.280 4976.180 1539.880 4978.470 ;
        RECT 1756.480 4976.020 1758.080 4978.480 ;
        RECT 1773.290 4978.440 1775.020 4982.820 ;
        RECT 1790.230 4978.470 1791.960 4982.850 ;
        RECT 2093.400 4978.480 2095.150 4982.640 ;
        RECT 1773.380 4976.180 1774.980 4978.440 ;
        RECT 1790.280 4976.180 1791.880 4978.470 ;
        RECT 2093.480 4976.020 2095.080 4978.480 ;
        RECT 2110.290 4978.440 2112.020 4982.820 ;
        RECT 2127.230 4978.470 2128.960 4982.850 ;
        RECT 2478.400 4978.480 2480.150 4982.640 ;
        RECT 2110.380 4976.180 2111.980 4978.440 ;
        RECT 2127.280 4976.180 2128.880 4978.470 ;
        RECT 2478.480 4976.020 2480.080 4978.480 ;
        RECT 2495.290 4978.440 2497.020 4982.820 ;
        RECT 2512.230 4978.470 2513.960 4982.850 ;
        RECT 2735.400 4978.480 2737.150 4982.640 ;
        RECT 2495.380 4976.180 2496.980 4978.440 ;
        RECT 2512.280 4976.180 2513.880 4978.470 ;
        RECT 2735.480 4976.020 2737.080 4978.480 ;
        RECT 2752.290 4978.440 2754.020 4982.820 ;
        RECT 2769.230 4978.470 2770.960 4982.850 ;
        RECT 2752.380 4976.180 2753.980 4978.440 ;
        RECT 2769.280 4976.180 2770.880 4978.470 ;
        RECT 232.880 4808.010 3353.190 4814.010 ;
        RECT 6.285 4541.490 10.480 4541.595 ;
        RECT 6.190 4539.890 12.800 4541.490 ;
        RECT 6.285 4539.790 10.480 4539.890 ;
        RECT 6.375 4524.590 10.570 4524.705 ;
        RECT 6.220 4522.990 12.800 4524.590 ;
        RECT 6.375 4522.900 10.570 4522.990 ;
        RECT 6.275 4507.690 10.750 4507.765 ;
        RECT 6.275 4506.090 12.960 4507.690 ;
        RECT 6.275 4506.010 10.750 4506.090 ;
        RECT 6.285 3912.490 10.480 3912.595 ;
        RECT 6.190 3910.890 12.800 3912.490 ;
        RECT 6.285 3910.790 10.480 3910.890 ;
        RECT 6.375 3895.590 10.570 3895.705 ;
        RECT 6.220 3893.990 12.800 3895.590 ;
        RECT 6.375 3893.900 10.570 3893.990 ;
        RECT 6.275 3878.690 10.750 3878.765 ;
        RECT 6.275 3877.090 12.960 3878.690 ;
        RECT 6.275 3877.010 10.750 3877.090 ;
        RECT 6.285 3696.490 10.480 3696.595 ;
        RECT 6.190 3694.890 12.800 3696.490 ;
        RECT 6.285 3694.790 10.480 3694.890 ;
        RECT 6.375 3679.590 10.570 3679.705 ;
        RECT 6.220 3677.990 12.800 3679.590 ;
        RECT 6.375 3677.900 10.570 3677.990 ;
        RECT 6.275 3662.690 10.750 3662.765 ;
        RECT 6.275 3661.090 12.960 3662.690 ;
        RECT 6.275 3661.010 10.750 3661.090 ;
        RECT 6.285 3480.490 10.480 3480.595 ;
        RECT 6.190 3478.890 12.800 3480.490 ;
        RECT 6.285 3478.790 10.480 3478.890 ;
        RECT 6.375 3463.590 10.570 3463.705 ;
        RECT 6.220 3461.990 12.800 3463.590 ;
        RECT 6.375 3461.900 10.570 3461.990 ;
        RECT 6.275 3446.690 10.750 3446.765 ;
        RECT 6.275 3445.090 12.960 3446.690 ;
        RECT 6.275 3445.010 10.750 3445.090 ;
        RECT 6.285 3264.490 10.480 3264.595 ;
        RECT 6.190 3262.890 12.800 3264.490 ;
        RECT 6.285 3262.790 10.480 3262.890 ;
        RECT 6.375 3247.590 10.570 3247.705 ;
        RECT 6.220 3245.990 12.800 3247.590 ;
        RECT 6.375 3245.900 10.570 3245.990 ;
        RECT 6.275 3230.690 10.750 3230.765 ;
        RECT 6.275 3229.090 12.960 3230.690 ;
        RECT 6.275 3229.010 10.750 3229.090 ;
        RECT 6.285 3048.490 10.480 3048.595 ;
        RECT 6.190 3046.890 12.800 3048.490 ;
        RECT 6.285 3046.790 10.480 3046.890 ;
        RECT 6.375 3031.590 10.570 3031.705 ;
        RECT 6.220 3029.990 12.800 3031.590 ;
        RECT 6.375 3029.900 10.570 3029.990 ;
        RECT 6.275 3014.690 10.750 3014.765 ;
        RECT 6.275 3013.090 12.960 3014.690 ;
        RECT 6.275 3013.010 10.750 3013.090 ;
        RECT 6.285 2832.490 10.480 2832.595 ;
        RECT 6.190 2830.890 12.800 2832.490 ;
        RECT 6.285 2830.790 10.480 2830.890 ;
        RECT 6.375 2815.590 10.570 2815.705 ;
        RECT 6.220 2813.990 12.800 2815.590 ;
        RECT 6.375 2813.900 10.570 2813.990 ;
        RECT 6.275 2798.690 10.750 2798.765 ;
        RECT 6.275 2797.090 12.960 2798.690 ;
        RECT 6.275 2797.010 10.750 2797.090 ;
        RECT 6.285 2616.490 10.480 2616.595 ;
        RECT 6.190 2614.890 12.800 2616.490 ;
        RECT 6.285 2614.790 10.480 2614.890 ;
        RECT 6.375 2599.590 10.570 2599.705 ;
        RECT 6.220 2597.990 12.800 2599.590 ;
        RECT 6.375 2597.900 10.570 2597.990 ;
        RECT 6.275 2582.690 10.750 2582.765 ;
        RECT 6.275 2581.090 12.960 2582.690 ;
        RECT 6.275 2581.010 10.750 2581.090 ;
        RECT 6.285 1978.490 10.480 1978.595 ;
        RECT 6.190 1976.890 12.800 1978.490 ;
        RECT 6.285 1976.790 10.480 1976.890 ;
        RECT 6.375 1961.590 10.570 1961.705 ;
        RECT 6.220 1959.990 12.800 1961.590 ;
        RECT 6.375 1959.900 10.570 1959.990 ;
        RECT 6.275 1944.690 10.750 1944.765 ;
        RECT 6.275 1943.090 12.960 1944.690 ;
        RECT 6.275 1943.010 10.750 1943.090 ;
        RECT 6.285 1762.490 10.480 1762.595 ;
        RECT 6.190 1760.890 12.800 1762.490 ;
        RECT 6.285 1760.790 10.480 1760.890 ;
        RECT 6.375 1745.590 10.570 1745.705 ;
        RECT 6.220 1743.990 12.800 1745.590 ;
        RECT 6.375 1743.900 10.570 1743.990 ;
        RECT 6.275 1728.690 10.750 1728.765 ;
        RECT 6.275 1727.090 12.960 1728.690 ;
        RECT 6.275 1727.010 10.750 1727.090 ;
        RECT 6.285 1546.490 10.480 1546.595 ;
        RECT 6.190 1544.890 12.800 1546.490 ;
        RECT 6.285 1544.790 10.480 1544.890 ;
        RECT 6.375 1529.590 10.570 1529.705 ;
        RECT 6.220 1527.990 12.800 1529.590 ;
        RECT 6.375 1527.900 10.570 1527.990 ;
        RECT 6.275 1512.690 10.750 1512.765 ;
        RECT 6.275 1511.090 12.960 1512.690 ;
        RECT 6.275 1511.010 10.750 1511.090 ;
        RECT 6.285 1330.490 10.480 1330.595 ;
        RECT 6.190 1328.890 12.800 1330.490 ;
        RECT 6.285 1328.790 10.480 1328.890 ;
        RECT 6.375 1313.590 10.570 1313.705 ;
        RECT 6.220 1311.990 12.800 1313.590 ;
        RECT 6.375 1311.900 10.570 1311.990 ;
        RECT 6.275 1296.690 10.750 1296.765 ;
        RECT 6.275 1295.090 12.960 1296.690 ;
        RECT 6.275 1295.010 10.750 1295.090 ;
        RECT 6.285 1114.490 10.480 1114.595 ;
        RECT 6.190 1112.890 12.800 1114.490 ;
        RECT 6.285 1112.790 10.480 1112.890 ;
        RECT 6.375 1097.590 10.570 1097.705 ;
        RECT 6.220 1095.990 12.800 1097.590 ;
        RECT 6.375 1095.900 10.570 1095.990 ;
        RECT 6.275 1080.690 10.750 1080.765 ;
        RECT 6.275 1079.090 12.960 1080.690 ;
        RECT 6.275 1079.010 10.750 1079.090 ;
        RECT 232.880 919.210 238.880 4808.010 ;
        RECT 3324.770 4782.270 3336.210 4793.150 ;
        RECT 248.770 4750.140 281.680 4753.240 ;
        RECT 248.660 1214.620 281.650 1217.720 ;
        RECT 250.520 1082.830 3324.820 1097.830 ;
        RECT 6.285 898.490 10.480 898.595 ;
        RECT 6.190 896.890 12.800 898.490 ;
        RECT 6.285 896.790 10.480 896.890 ;
        RECT 6.375 881.590 10.570 881.705 ;
        RECT 6.220 879.990 12.800 881.590 ;
        RECT 6.375 879.900 10.570 879.990 ;
        RECT 6.275 864.690 10.750 864.765 ;
        RECT 6.275 863.090 12.960 864.690 ;
        RECT 6.275 863.010 10.750 863.090 ;
    END
  END vssd1_core
  PIN vccd1_core
    PORT
      LAYER met3 ;
        RECT 543.800 4799.790 549.800 4988.980 ;
        RECT 800.800 4799.790 806.800 4988.980 ;
        RECT 1057.800 4799.790 1063.800 4988.980 ;
        RECT 1314.800 4799.790 1320.800 4988.980 ;
        RECT 1572.800 4799.790 1578.800 4988.980 ;
        RECT 1824.800 4799.790 1830.800 4988.980 ;
        RECT 2161.800 4799.790 2167.800 4988.980 ;
        RECT 2546.800 4799.790 2552.800 4988.980 ;
        RECT 2803.800 4799.790 2809.800 4988.980 ;
        RECT 0.000 4578.910 260.980 4580.410 ;
        RECT 0.000 4574.410 289.500 4578.910 ;
        RECT 255.080 4572.910 289.500 4574.410 ;
        RECT 0.000 3945.410 289.500 3951.410 ;
        RECT 250.280 3735.410 289.500 3741.410 ;
        RECT 0.000 3729.410 256.740 3735.410 ;
        RECT 0.000 3513.410 289.500 3519.410 ;
        RECT 0.000 3297.410 289.500 3303.410 ;
        RECT 0.000 3081.410 289.500 3087.410 ;
        RECT 0.000 2865.410 289.500 2871.410 ;
        RECT 0.000 2649.410 289.500 2655.410 ;
        RECT 0.000 2011.410 289.500 2017.410 ;
        RECT 0.000 1795.410 289.500 1801.410 ;
        RECT 249.730 1585.410 289.500 1589.410 ;
        RECT 0.000 1583.410 289.500 1585.410 ;
        RECT 0.000 1579.410 256.210 1583.410 ;
        RECT 0.000 1363.410 289.500 1369.410 ;
        RECT 0.000 1147.410 247.190 1153.410 ;
        RECT 0.000 931.410 247.190 937.410 ;
      LAYER via3 ;
        RECT 544.035 4985.020 549.555 4988.140 ;
        RECT 544.315 4800.595 549.435 4805.715 ;
        RECT 801.035 4985.020 806.555 4988.140 ;
        RECT 801.315 4800.595 806.435 4805.715 ;
        RECT 1058.035 4985.020 1063.555 4988.140 ;
        RECT 1058.315 4800.595 1063.435 4805.715 ;
        RECT 1315.035 4985.020 1320.555 4988.140 ;
        RECT 1315.315 4800.595 1320.435 4805.715 ;
        RECT 1573.035 4985.020 1578.555 4988.140 ;
        RECT 1573.315 4800.595 1578.435 4805.715 ;
        RECT 1825.035 4985.020 1830.555 4988.140 ;
        RECT 1825.315 4800.595 1830.435 4805.715 ;
        RECT 2162.035 4985.020 2167.555 4988.140 ;
        RECT 2162.315 4800.595 2167.435 4805.715 ;
        RECT 2547.035 4985.020 2552.555 4988.140 ;
        RECT 2547.315 4800.595 2552.435 4805.715 ;
        RECT 2804.035 4985.020 2809.555 4988.140 ;
        RECT 2804.315 4800.595 2809.435 4805.715 ;
        RECT 0.840 4574.645 3.960 4580.165 ;
        RECT 241.265 4574.925 246.385 4580.045 ;
        RECT 286.785 4573.125 289.105 4578.645 ;
        RECT 0.840 3945.645 3.960 3951.165 ;
        RECT 241.265 3945.925 246.385 3951.045 ;
        RECT 286.785 3945.625 289.105 3951.145 ;
        RECT 286.785 3735.625 289.105 3741.145 ;
        RECT 0.840 3729.645 3.960 3735.165 ;
        RECT 241.265 3729.925 246.385 3735.045 ;
        RECT 0.840 3513.645 3.960 3519.165 ;
        RECT 241.265 3513.925 246.385 3519.045 ;
        RECT 286.785 3513.625 289.105 3519.145 ;
        RECT 0.840 3297.645 3.960 3303.165 ;
        RECT 241.265 3297.925 246.385 3303.045 ;
        RECT 286.785 3297.625 289.105 3303.145 ;
        RECT 0.840 3081.645 3.960 3087.165 ;
        RECT 241.265 3081.925 246.385 3087.045 ;
        RECT 286.785 3081.625 289.105 3087.145 ;
        RECT 0.840 2865.645 3.960 2871.165 ;
        RECT 241.265 2865.925 246.385 2871.045 ;
        RECT 286.785 2865.625 289.105 2871.145 ;
        RECT 0.840 2649.645 3.960 2655.165 ;
        RECT 241.265 2649.925 246.385 2655.045 ;
        RECT 286.785 2649.625 289.105 2655.145 ;
        RECT 0.840 2011.645 3.960 2017.165 ;
        RECT 241.265 2011.925 246.385 2017.045 ;
        RECT 286.785 2011.625 289.105 2017.145 ;
        RECT 0.840 1795.645 3.960 1801.165 ;
        RECT 241.265 1795.925 246.385 1801.045 ;
        RECT 286.785 1795.625 289.105 1801.145 ;
        RECT 0.840 1579.645 3.960 1585.165 ;
        RECT 241.265 1579.925 246.385 1585.045 ;
        RECT 286.785 1583.625 289.105 1589.145 ;
        RECT 0.840 1363.645 3.960 1369.165 ;
        RECT 241.265 1363.925 246.385 1369.045 ;
        RECT 286.785 1363.625 289.105 1369.145 ;
        RECT 0.840 1147.645 3.960 1153.165 ;
        RECT 241.265 1147.925 246.385 1153.045 ;
        RECT 0.840 931.645 3.960 937.165 ;
        RECT 241.265 931.925 246.385 937.045 ;
      LAYER met4 ;
        RECT 466.620 4984.560 550.240 4988.560 ;
        RECT 723.620 4984.560 807.240 4988.560 ;
        RECT 980.620 4984.560 1064.240 4988.560 ;
        RECT 1237.620 4984.560 1321.240 4988.560 ;
        RECT 1495.620 4984.560 1579.240 4988.560 ;
        RECT 1747.620 4984.560 1831.240 4988.560 ;
        RECT 2084.620 4984.560 2168.240 4988.560 ;
        RECT 2469.620 4984.560 2553.240 4988.560 ;
        RECT 2726.620 4984.560 2810.240 4988.560 ;
        RECT 543.760 4800.140 549.830 4806.170 ;
        RECT 800.760 4800.140 806.830 4806.170 ;
        RECT 1057.760 4800.140 1063.830 4806.170 ;
        RECT 1314.760 4800.140 1320.830 4806.170 ;
        RECT 1572.760 4800.140 1578.830 4806.170 ;
        RECT 1824.760 4800.140 1830.830 4806.170 ;
        RECT 2161.760 4800.140 2167.830 4806.170 ;
        RECT 2546.760 4800.140 2552.830 4806.170 ;
        RECT 2803.760 4800.140 2809.830 4806.170 ;
        RECT 0.420 4497.230 4.420 4580.850 ;
        RECT 240.810 4574.370 246.840 4580.440 ;
        RECT 286.640 4573.110 289.250 4578.660 ;
        RECT 0.420 3868.230 4.420 3951.850 ;
        RECT 240.810 3945.370 246.840 3951.440 ;
        RECT 286.640 3945.610 289.250 3951.160 ;
        RECT 0.420 3652.230 4.420 3735.850 ;
        RECT 286.640 3735.610 289.250 3741.160 ;
        RECT 240.810 3729.370 246.840 3735.440 ;
        RECT 0.420 3436.230 4.420 3519.850 ;
        RECT 240.810 3513.370 246.840 3519.440 ;
        RECT 286.640 3513.610 289.250 3519.160 ;
        RECT 0.420 3220.230 4.420 3303.850 ;
        RECT 240.810 3297.370 246.840 3303.440 ;
        RECT 286.640 3297.610 289.250 3303.160 ;
        RECT 0.420 3004.230 4.420 3087.850 ;
        RECT 240.810 3081.370 246.840 3087.440 ;
        RECT 286.640 3081.610 289.250 3087.160 ;
        RECT 0.420 2788.230 4.420 2871.850 ;
        RECT 240.810 2865.370 246.840 2871.440 ;
        RECT 286.640 2865.610 289.250 2871.160 ;
        RECT 0.420 2572.230 4.420 2655.850 ;
        RECT 240.810 2649.370 246.840 2655.440 ;
        RECT 286.640 2649.610 289.250 2655.160 ;
        RECT 0.420 1934.230 4.420 2017.850 ;
        RECT 240.810 2011.370 246.840 2017.440 ;
        RECT 286.640 2011.610 289.250 2017.160 ;
        RECT 0.420 1718.230 4.420 1801.850 ;
        RECT 240.810 1795.370 246.840 1801.440 ;
        RECT 286.640 1795.610 289.250 1801.160 ;
        RECT 0.420 1502.230 4.420 1585.850 ;
        RECT 240.810 1579.370 246.840 1585.440 ;
        RECT 286.640 1583.610 289.250 1589.160 ;
        RECT 0.420 1286.230 4.420 1369.850 ;
        RECT 240.810 1363.370 246.840 1369.440 ;
        RECT 286.640 1363.610 289.250 1369.160 ;
        RECT 286.400 1182.790 289.500 1219.460 ;
        RECT 286.400 1179.690 305.750 1182.790 ;
        RECT 0.420 1070.230 4.420 1153.850 ;
        RECT 240.810 1147.370 246.840 1153.440 ;
        RECT 302.650 1062.240 305.750 1179.690 ;
        RECT 1316.710 1062.840 1318.950 1077.120 ;
        RECT 1391.660 1062.840 1393.900 1077.120 ;
        RECT 1466.660 1062.840 1468.900 1077.120 ;
        RECT 1542.960 1062.840 1545.200 1077.120 ;
        RECT 3222.980 1061.980 3226.080 1219.490 ;
        RECT 3304.340 1062.830 3353.240 1077.880 ;
        RECT 0.420 854.230 4.420 937.850 ;
        RECT 240.810 931.370 246.840 937.440 ;
      LAYER via4 ;
        RECT 467.245 4986.755 468.425 4987.935 ;
        RECT 484.180 4986.775 485.360 4987.955 ;
        RECT 501.030 4986.765 502.210 4987.945 ;
        RECT 467.245 4985.155 468.425 4986.335 ;
        RECT 484.180 4985.175 485.360 4986.355 ;
        RECT 501.030 4985.165 502.210 4986.345 ;
        RECT 724.245 4986.755 725.425 4987.935 ;
        RECT 741.180 4986.775 742.360 4987.955 ;
        RECT 758.030 4986.765 759.210 4987.945 ;
        RECT 724.245 4985.155 725.425 4986.335 ;
        RECT 741.180 4985.175 742.360 4986.355 ;
        RECT 758.030 4985.165 759.210 4986.345 ;
        RECT 981.245 4986.755 982.425 4987.935 ;
        RECT 998.180 4986.775 999.360 4987.955 ;
        RECT 1015.030 4986.765 1016.210 4987.945 ;
        RECT 981.245 4985.155 982.425 4986.335 ;
        RECT 998.180 4985.175 999.360 4986.355 ;
        RECT 1015.030 4985.165 1016.210 4986.345 ;
        RECT 1238.245 4986.755 1239.425 4987.935 ;
        RECT 1255.180 4986.775 1256.360 4987.955 ;
        RECT 1272.030 4986.765 1273.210 4987.945 ;
        RECT 1238.245 4985.155 1239.425 4986.335 ;
        RECT 1255.180 4985.175 1256.360 4986.355 ;
        RECT 1272.030 4985.165 1273.210 4986.345 ;
        RECT 1496.245 4986.755 1497.425 4987.935 ;
        RECT 1513.180 4986.775 1514.360 4987.955 ;
        RECT 1530.030 4986.765 1531.210 4987.945 ;
        RECT 1496.245 4985.155 1497.425 4986.335 ;
        RECT 1513.180 4985.175 1514.360 4986.355 ;
        RECT 1530.030 4985.165 1531.210 4986.345 ;
        RECT 1748.245 4986.755 1749.425 4987.935 ;
        RECT 1765.180 4986.775 1766.360 4987.955 ;
        RECT 1782.030 4986.765 1783.210 4987.945 ;
        RECT 1748.245 4985.155 1749.425 4986.335 ;
        RECT 1765.180 4985.175 1766.360 4986.355 ;
        RECT 1782.030 4985.165 1783.210 4986.345 ;
        RECT 2085.245 4986.755 2086.425 4987.935 ;
        RECT 2102.180 4986.775 2103.360 4987.955 ;
        RECT 2119.030 4986.765 2120.210 4987.945 ;
        RECT 2085.245 4985.155 2086.425 4986.335 ;
        RECT 2102.180 4985.175 2103.360 4986.355 ;
        RECT 2119.030 4985.165 2120.210 4986.345 ;
        RECT 2470.245 4986.755 2471.425 4987.935 ;
        RECT 2487.180 4986.775 2488.360 4987.955 ;
        RECT 2504.030 4986.765 2505.210 4987.945 ;
        RECT 2470.245 4985.155 2471.425 4986.335 ;
        RECT 2487.180 4985.175 2488.360 4986.355 ;
        RECT 2504.030 4985.165 2505.210 4986.345 ;
        RECT 2727.245 4986.755 2728.425 4987.935 ;
        RECT 2744.180 4986.775 2745.360 4987.955 ;
        RECT 2761.030 4986.765 2762.210 4987.945 ;
        RECT 2727.245 4985.155 2728.425 4986.335 ;
        RECT 2744.180 4985.175 2745.360 4986.355 ;
        RECT 2761.030 4985.165 2762.210 4986.345 ;
        RECT 544.685 4800.965 549.065 4805.345 ;
        RECT 801.685 4800.965 806.065 4805.345 ;
        RECT 1058.685 4800.965 1063.065 4805.345 ;
        RECT 1315.685 4800.965 1320.065 4805.345 ;
        RECT 1573.685 4800.965 1578.065 4805.345 ;
        RECT 1825.685 4800.965 1830.065 4805.345 ;
        RECT 2162.685 4800.965 2167.065 4805.345 ;
        RECT 2547.685 4800.965 2552.065 4805.345 ;
        RECT 2804.685 4800.965 2809.065 4805.345 ;
        RECT 241.635 4575.295 246.015 4579.675 ;
        RECT 1.010 4531.635 2.190 4532.815 ;
        RECT 2.610 4531.635 3.790 4532.815 ;
        RECT 1.040 4514.805 2.220 4515.985 ;
        RECT 2.640 4514.805 3.820 4515.985 ;
        RECT 1.045 4497.855 2.225 4499.035 ;
        RECT 2.645 4497.855 3.825 4499.035 ;
        RECT 241.635 3946.295 246.015 3950.675 ;
        RECT 1.010 3902.635 2.190 3903.815 ;
        RECT 2.610 3902.635 3.790 3903.815 ;
        RECT 1.040 3885.805 2.220 3886.985 ;
        RECT 2.640 3885.805 3.820 3886.985 ;
        RECT 1.045 3868.855 2.225 3870.035 ;
        RECT 2.645 3868.855 3.825 3870.035 ;
        RECT 241.635 3730.295 246.015 3734.675 ;
        RECT 1.010 3686.635 2.190 3687.815 ;
        RECT 2.610 3686.635 3.790 3687.815 ;
        RECT 1.040 3669.805 2.220 3670.985 ;
        RECT 2.640 3669.805 3.820 3670.985 ;
        RECT 1.045 3652.855 2.225 3654.035 ;
        RECT 2.645 3652.855 3.825 3654.035 ;
        RECT 241.635 3514.295 246.015 3518.675 ;
        RECT 1.010 3470.635 2.190 3471.815 ;
        RECT 2.610 3470.635 3.790 3471.815 ;
        RECT 1.040 3453.805 2.220 3454.985 ;
        RECT 2.640 3453.805 3.820 3454.985 ;
        RECT 1.045 3436.855 2.225 3438.035 ;
        RECT 2.645 3436.855 3.825 3438.035 ;
        RECT 241.635 3298.295 246.015 3302.675 ;
        RECT 1.010 3254.635 2.190 3255.815 ;
        RECT 2.610 3254.635 3.790 3255.815 ;
        RECT 1.040 3237.805 2.220 3238.985 ;
        RECT 2.640 3237.805 3.820 3238.985 ;
        RECT 1.045 3220.855 2.225 3222.035 ;
        RECT 2.645 3220.855 3.825 3222.035 ;
        RECT 241.635 3082.295 246.015 3086.675 ;
        RECT 1.010 3038.635 2.190 3039.815 ;
        RECT 2.610 3038.635 3.790 3039.815 ;
        RECT 1.040 3021.805 2.220 3022.985 ;
        RECT 2.640 3021.805 3.820 3022.985 ;
        RECT 1.045 3004.855 2.225 3006.035 ;
        RECT 2.645 3004.855 3.825 3006.035 ;
        RECT 241.635 2866.295 246.015 2870.675 ;
        RECT 1.010 2822.635 2.190 2823.815 ;
        RECT 2.610 2822.635 3.790 2823.815 ;
        RECT 1.040 2805.805 2.220 2806.985 ;
        RECT 2.640 2805.805 3.820 2806.985 ;
        RECT 1.045 2788.855 2.225 2790.035 ;
        RECT 2.645 2788.855 3.825 2790.035 ;
        RECT 241.635 2650.295 246.015 2654.675 ;
        RECT 1.010 2606.635 2.190 2607.815 ;
        RECT 2.610 2606.635 3.790 2607.815 ;
        RECT 1.040 2589.805 2.220 2590.985 ;
        RECT 2.640 2589.805 3.820 2590.985 ;
        RECT 1.045 2572.855 2.225 2574.035 ;
        RECT 2.645 2572.855 3.825 2574.035 ;
        RECT 241.635 2012.295 246.015 2016.675 ;
        RECT 1.010 1968.635 2.190 1969.815 ;
        RECT 2.610 1968.635 3.790 1969.815 ;
        RECT 1.040 1951.805 2.220 1952.985 ;
        RECT 2.640 1951.805 3.820 1952.985 ;
        RECT 1.045 1934.855 2.225 1936.035 ;
        RECT 2.645 1934.855 3.825 1936.035 ;
        RECT 241.635 1796.295 246.015 1800.675 ;
        RECT 1.010 1752.635 2.190 1753.815 ;
        RECT 2.610 1752.635 3.790 1753.815 ;
        RECT 1.040 1735.805 2.220 1736.985 ;
        RECT 2.640 1735.805 3.820 1736.985 ;
        RECT 1.045 1718.855 2.225 1720.035 ;
        RECT 2.645 1718.855 3.825 1720.035 ;
        RECT 241.635 1580.295 246.015 1584.675 ;
        RECT 1.010 1536.635 2.190 1537.815 ;
        RECT 2.610 1536.635 3.790 1537.815 ;
        RECT 1.040 1519.805 2.220 1520.985 ;
        RECT 2.640 1519.805 3.820 1520.985 ;
        RECT 1.045 1502.855 2.225 1504.035 ;
        RECT 2.645 1502.855 3.825 1504.035 ;
        RECT 241.635 1364.295 246.015 1368.675 ;
        RECT 1.010 1320.635 2.190 1321.815 ;
        RECT 2.610 1320.635 3.790 1321.815 ;
        RECT 1.040 1303.805 2.220 1304.985 ;
        RECT 2.640 1303.805 3.820 1304.985 ;
        RECT 1.045 1286.855 2.225 1288.035 ;
        RECT 2.645 1286.855 3.825 1288.035 ;
        RECT 241.635 1148.295 246.015 1152.675 ;
        RECT 1.010 1104.635 2.190 1105.815 ;
        RECT 2.610 1104.635 3.790 1105.815 ;
        RECT 1.040 1087.805 2.220 1088.985 ;
        RECT 2.640 1087.805 3.820 1088.985 ;
        RECT 1.045 1070.855 2.225 1072.035 ;
        RECT 2.645 1070.855 3.825 1072.035 ;
        RECT 303.585 1076.170 304.765 1077.350 ;
        RECT 303.585 1074.570 304.765 1075.750 ;
        RECT 303.585 1072.970 304.765 1074.150 ;
        RECT 303.585 1071.370 304.765 1072.550 ;
        RECT 303.585 1069.770 304.765 1070.950 ;
        RECT 303.585 1068.170 304.765 1069.350 ;
        RECT 303.585 1066.570 304.765 1067.750 ;
        RECT 303.585 1064.970 304.765 1066.150 ;
        RECT 303.585 1063.370 304.765 1064.550 ;
        RECT 1317.240 1075.205 1318.420 1076.385 ;
        RECT 1317.240 1073.605 1318.420 1074.785 ;
        RECT 1317.240 1072.005 1318.420 1073.185 ;
        RECT 1317.240 1070.405 1318.420 1071.585 ;
        RECT 1317.240 1068.805 1318.420 1069.985 ;
        RECT 1317.240 1067.205 1318.420 1068.385 ;
        RECT 1317.240 1065.605 1318.420 1066.785 ;
        RECT 1317.240 1064.005 1318.420 1065.185 ;
        RECT 1392.190 1075.205 1393.370 1076.385 ;
        RECT 1392.190 1073.605 1393.370 1074.785 ;
        RECT 1392.190 1072.005 1393.370 1073.185 ;
        RECT 1392.190 1070.405 1393.370 1071.585 ;
        RECT 1392.190 1068.805 1393.370 1069.985 ;
        RECT 1392.190 1067.205 1393.370 1068.385 ;
        RECT 1392.190 1065.605 1393.370 1066.785 ;
        RECT 1392.190 1064.005 1393.370 1065.185 ;
        RECT 1467.190 1075.205 1468.370 1076.385 ;
        RECT 1467.190 1073.605 1468.370 1074.785 ;
        RECT 1467.190 1072.005 1468.370 1073.185 ;
        RECT 1467.190 1070.405 1468.370 1071.585 ;
        RECT 1467.190 1068.805 1468.370 1069.985 ;
        RECT 1467.190 1067.205 1468.370 1068.385 ;
        RECT 1467.190 1065.605 1468.370 1066.785 ;
        RECT 1467.190 1064.005 1468.370 1065.185 ;
        RECT 1543.490 1075.205 1544.670 1076.385 ;
        RECT 1543.490 1073.605 1544.670 1074.785 ;
        RECT 1543.490 1072.005 1544.670 1073.185 ;
        RECT 1543.490 1070.405 1544.670 1071.585 ;
        RECT 1543.490 1068.805 1544.670 1069.985 ;
        RECT 1543.490 1067.205 1544.670 1068.385 ;
        RECT 1543.490 1065.605 1544.670 1066.785 ;
        RECT 1543.490 1064.005 1544.670 1065.185 ;
        RECT 3223.130 1063.395 3225.910 1077.375 ;
        RECT 3305.450 1064.185 3317.830 1076.565 ;
        RECT 3341.020 1064.090 3351.800 1076.470 ;
        RECT 241.635 932.295 246.015 936.675 ;
        RECT 1.010 888.635 2.190 889.815 ;
        RECT 2.610 888.635 3.790 889.815 ;
        RECT 1.040 871.805 2.220 872.985 ;
        RECT 2.640 871.805 3.820 872.985 ;
        RECT 1.045 854.855 2.225 856.035 ;
        RECT 2.645 854.855 3.825 856.035 ;
      LAYER met5 ;
        RECT 466.950 4984.470 468.700 4988.630 ;
        RECT 483.900 4984.510 485.630 4988.890 ;
        RECT 467.030 4976.020 468.630 4984.470 ;
        RECT 483.930 4976.180 485.530 4984.510 ;
        RECT 500.720 4984.490 502.450 4988.870 ;
        RECT 500.830 4976.180 502.430 4984.490 ;
        RECT 723.950 4984.470 725.700 4988.630 ;
        RECT 740.900 4984.510 742.630 4988.890 ;
        RECT 724.030 4976.020 725.630 4984.470 ;
        RECT 740.930 4976.180 742.530 4984.510 ;
        RECT 757.720 4984.490 759.450 4988.870 ;
        RECT 757.830 4976.180 759.430 4984.490 ;
        RECT 980.950 4984.470 982.700 4988.630 ;
        RECT 997.900 4984.510 999.630 4988.890 ;
        RECT 981.030 4976.020 982.630 4984.470 ;
        RECT 997.930 4976.180 999.530 4984.510 ;
        RECT 1014.720 4984.490 1016.450 4988.870 ;
        RECT 1014.830 4976.180 1016.430 4984.490 ;
        RECT 1237.950 4984.470 1239.700 4988.630 ;
        RECT 1254.900 4984.510 1256.630 4988.890 ;
        RECT 1238.030 4976.020 1239.630 4984.470 ;
        RECT 1254.930 4976.180 1256.530 4984.510 ;
        RECT 1271.720 4984.490 1273.450 4988.870 ;
        RECT 1271.830 4976.180 1273.430 4984.490 ;
        RECT 1495.950 4984.470 1497.700 4988.630 ;
        RECT 1512.900 4984.510 1514.630 4988.890 ;
        RECT 1496.030 4976.020 1497.630 4984.470 ;
        RECT 1512.930 4976.180 1514.530 4984.510 ;
        RECT 1529.720 4984.490 1531.450 4988.870 ;
        RECT 1529.830 4976.180 1531.430 4984.490 ;
        RECT 1747.950 4984.470 1749.700 4988.630 ;
        RECT 1764.900 4984.510 1766.630 4988.890 ;
        RECT 1748.030 4976.020 1749.630 4984.470 ;
        RECT 1764.930 4976.180 1766.530 4984.510 ;
        RECT 1781.720 4984.490 1783.450 4988.870 ;
        RECT 1781.830 4976.180 1783.430 4984.490 ;
        RECT 2084.950 4984.470 2086.700 4988.630 ;
        RECT 2101.900 4984.510 2103.630 4988.890 ;
        RECT 2085.030 4976.020 2086.630 4984.470 ;
        RECT 2101.930 4976.180 2103.530 4984.510 ;
        RECT 2118.720 4984.490 2120.450 4988.870 ;
        RECT 2118.830 4976.180 2120.430 4984.490 ;
        RECT 2469.950 4984.470 2471.700 4988.630 ;
        RECT 2486.900 4984.510 2488.630 4988.890 ;
        RECT 2470.030 4976.020 2471.630 4984.470 ;
        RECT 2486.930 4976.180 2488.530 4984.510 ;
        RECT 2503.720 4984.490 2505.450 4988.870 ;
        RECT 2503.830 4976.180 2505.430 4984.490 ;
        RECT 2726.950 4984.470 2728.700 4988.630 ;
        RECT 2743.900 4984.510 2745.630 4988.890 ;
        RECT 2727.030 4976.020 2728.630 4984.470 ;
        RECT 2743.930 4976.180 2745.530 4984.510 ;
        RECT 2760.720 4984.490 2762.450 4988.870 ;
        RECT 2760.830 4976.180 2762.430 4984.490 ;
        RECT 240.880 4800.010 3352.990 4806.010 ;
        RECT 240.880 4748.440 246.880 4800.010 ;
        RECT 3339.990 4793.980 3352.990 4800.010 ;
        RECT 240.880 4745.340 286.470 4748.440 ;
        RECT 0.330 4533.040 4.525 4533.200 ;
        RECT 0.130 4531.440 12.800 4533.040 ;
        RECT 0.330 4531.395 4.525 4531.440 ;
        RECT 0.060 4516.140 4.535 4516.270 ;
        RECT 0.060 4514.540 12.800 4516.140 ;
        RECT 0.060 4514.530 4.535 4514.540 ;
        RECT 0.315 4499.240 4.790 4499.350 ;
        RECT 0.315 4497.640 12.960 4499.240 ;
        RECT 0.315 4497.540 4.790 4497.640 ;
        RECT 0.330 3904.040 4.525 3904.200 ;
        RECT 0.130 3902.440 12.800 3904.040 ;
        RECT 0.330 3902.395 4.525 3902.440 ;
        RECT 0.060 3887.140 4.535 3887.270 ;
        RECT 0.060 3885.540 12.800 3887.140 ;
        RECT 0.060 3885.530 4.535 3885.540 ;
        RECT 0.315 3870.240 4.790 3870.350 ;
        RECT 0.315 3868.640 12.960 3870.240 ;
        RECT 0.315 3868.540 4.790 3868.640 ;
        RECT 0.330 3688.040 4.525 3688.200 ;
        RECT 0.130 3686.440 12.800 3688.040 ;
        RECT 0.330 3686.395 4.525 3686.440 ;
        RECT 0.060 3671.140 4.535 3671.270 ;
        RECT 0.060 3669.540 12.800 3671.140 ;
        RECT 0.060 3669.530 4.535 3669.540 ;
        RECT 0.315 3654.240 4.790 3654.350 ;
        RECT 0.315 3652.640 12.960 3654.240 ;
        RECT 0.315 3652.540 4.790 3652.640 ;
        RECT 0.330 3472.040 4.525 3472.200 ;
        RECT 0.130 3470.440 12.800 3472.040 ;
        RECT 0.330 3470.395 4.525 3470.440 ;
        RECT 0.060 3455.140 4.535 3455.270 ;
        RECT 0.060 3453.540 12.800 3455.140 ;
        RECT 0.060 3453.530 4.535 3453.540 ;
        RECT 0.315 3438.240 4.790 3438.350 ;
        RECT 0.315 3436.640 12.960 3438.240 ;
        RECT 0.315 3436.540 4.790 3436.640 ;
        RECT 0.330 3256.040 4.525 3256.200 ;
        RECT 0.130 3254.440 12.800 3256.040 ;
        RECT 0.330 3254.395 4.525 3254.440 ;
        RECT 0.060 3239.140 4.535 3239.270 ;
        RECT 0.060 3237.540 12.800 3239.140 ;
        RECT 0.060 3237.530 4.535 3237.540 ;
        RECT 0.315 3222.240 4.790 3222.350 ;
        RECT 0.315 3220.640 12.960 3222.240 ;
        RECT 0.315 3220.540 4.790 3220.640 ;
        RECT 0.330 3040.040 4.525 3040.200 ;
        RECT 0.130 3038.440 12.800 3040.040 ;
        RECT 0.330 3038.395 4.525 3038.440 ;
        RECT 0.060 3023.140 4.535 3023.270 ;
        RECT 0.060 3021.540 12.800 3023.140 ;
        RECT 0.060 3021.530 4.535 3021.540 ;
        RECT 0.315 3006.240 4.790 3006.350 ;
        RECT 0.315 3004.640 12.960 3006.240 ;
        RECT 0.315 3004.540 4.790 3004.640 ;
        RECT 0.330 2824.040 4.525 2824.200 ;
        RECT 0.130 2822.440 12.800 2824.040 ;
        RECT 0.330 2822.395 4.525 2822.440 ;
        RECT 0.060 2807.140 4.535 2807.270 ;
        RECT 0.060 2805.540 12.800 2807.140 ;
        RECT 0.060 2805.530 4.535 2805.540 ;
        RECT 0.315 2790.240 4.790 2790.350 ;
        RECT 0.315 2788.640 12.960 2790.240 ;
        RECT 0.315 2788.540 4.790 2788.640 ;
        RECT 0.330 2608.040 4.525 2608.200 ;
        RECT 0.130 2606.440 12.800 2608.040 ;
        RECT 0.330 2606.395 4.525 2606.440 ;
        RECT 0.060 2591.140 4.535 2591.270 ;
        RECT 0.060 2589.540 12.800 2591.140 ;
        RECT 0.060 2589.530 4.535 2589.540 ;
        RECT 0.315 2574.240 4.790 2574.350 ;
        RECT 0.315 2572.640 12.960 2574.240 ;
        RECT 0.315 2572.540 4.790 2572.640 ;
        RECT 0.330 1970.040 4.525 1970.200 ;
        RECT 0.130 1968.440 12.800 1970.040 ;
        RECT 0.330 1968.395 4.525 1968.440 ;
        RECT 0.060 1953.140 4.535 1953.270 ;
        RECT 0.060 1951.540 12.800 1953.140 ;
        RECT 0.060 1951.530 4.535 1951.540 ;
        RECT 0.315 1936.240 4.790 1936.350 ;
        RECT 0.315 1934.640 12.960 1936.240 ;
        RECT 0.315 1934.540 4.790 1934.640 ;
        RECT 0.330 1754.040 4.525 1754.200 ;
        RECT 0.130 1752.440 12.800 1754.040 ;
        RECT 0.330 1752.395 4.525 1752.440 ;
        RECT 0.060 1737.140 4.535 1737.270 ;
        RECT 0.060 1735.540 12.800 1737.140 ;
        RECT 0.060 1735.530 4.535 1735.540 ;
        RECT 0.315 1720.240 4.790 1720.350 ;
        RECT 0.315 1718.640 12.960 1720.240 ;
        RECT 0.315 1718.540 4.790 1718.640 ;
        RECT 0.330 1538.040 4.525 1538.200 ;
        RECT 0.130 1536.440 12.800 1538.040 ;
        RECT 0.330 1536.395 4.525 1536.440 ;
        RECT 0.060 1521.140 4.535 1521.270 ;
        RECT 0.060 1519.540 12.800 1521.140 ;
        RECT 0.060 1519.530 4.535 1519.540 ;
        RECT 0.315 1504.240 4.790 1504.350 ;
        RECT 0.315 1502.640 12.960 1504.240 ;
        RECT 0.315 1502.540 4.790 1502.640 ;
        RECT 0.330 1322.040 4.525 1322.200 ;
        RECT 0.130 1320.440 12.800 1322.040 ;
        RECT 0.330 1320.395 4.525 1320.440 ;
        RECT 0.060 1305.140 4.535 1305.270 ;
        RECT 0.060 1303.540 12.800 1305.140 ;
        RECT 0.060 1303.530 4.535 1303.540 ;
        RECT 0.315 1288.240 4.790 1288.350 ;
        RECT 0.315 1286.640 12.960 1288.240 ;
        RECT 0.315 1286.540 4.790 1286.640 ;
        RECT 240.880 1222.520 246.880 4745.340 ;
        RECT 240.880 1219.420 286.450 1222.520 ;
        RECT 0.330 1106.040 4.525 1106.200 ;
        RECT 0.130 1104.440 12.800 1106.040 ;
        RECT 0.330 1104.395 4.525 1104.440 ;
        RECT 0.060 1089.140 4.535 1089.270 ;
        RECT 0.060 1087.540 12.800 1089.140 ;
        RECT 0.060 1087.530 4.535 1087.540 ;
        RECT 240.880 1077.830 246.880 1219.420 ;
        RECT 0.315 1072.240 4.790 1072.350 ;
        RECT 0.315 1070.640 12.960 1072.240 ;
        RECT 0.315 1070.540 4.790 1070.640 ;
        RECT 240.880 1062.830 3319.340 1077.830 ;
        RECT 3340.670 1063.580 3352.150 1076.980 ;
        RECT 240.880 927.210 246.880 1062.830 ;
        RECT 0.330 890.040 4.525 890.200 ;
        RECT 0.130 888.440 12.800 890.040 ;
        RECT 0.330 888.395 4.525 888.440 ;
        RECT 0.060 873.140 4.535 873.270 ;
        RECT 0.060 871.540 12.800 873.140 ;
        RECT 0.060 871.530 4.535 871.540 ;
        RECT 0.315 856.240 4.790 856.350 ;
        RECT 0.315 854.640 12.960 856.240 ;
        RECT 0.315 854.540 4.790 854.640 ;
    END
  END vccd1_core
  PIN vssa1_core
    PORT
      LAYER met3 ;
        RECT 2848.390 4805.660 2872.285 4818.890 ;
        RECT 2898.280 4805.660 2922.180 4818.890 ;
        RECT 3289.460 1959.240 3358.450 1983.005 ;
        RECT 3289.460 1958.310 3305.440 1959.240 ;
        RECT 3289.460 1909.210 3358.450 1933.110 ;
      LAYER via3 ;
        RECT 2848.960 4806.215 2871.680 4815.735 ;
        RECT 2898.810 4806.245 2921.530 4815.765 ;
        RECT 3290.615 1958.925 3302.535 1982.445 ;
        RECT 3290.530 1909.935 3302.450 1932.655 ;
      LAYER met4 ;
        RECT 2848.290 4784.440 2872.280 4816.150 ;
        RECT 2898.240 4784.510 2922.230 4816.220 ;
        RECT 3289.930 1958.360 3302.950 1982.950 ;
        RECT 3289.980 1909.300 3303.060 1933.120 ;
        RECT 262.400 1162.540 265.500 1195.460 ;
        RECT 1923.750 1162.870 1927.680 1177.850 ;
        RECT 1999.000 1162.870 2002.930 1177.850 ;
        RECT 1926.760 1141.540 1927.660 1162.870 ;
        RECT 2002.010 1141.540 2002.910 1162.870 ;
        RECT 3246.980 1162.430 3250.080 1195.520 ;
      LAYER via4 ;
        RECT 2849.265 4785.605 2871.245 4796.385 ;
        RECT 2899.245 4785.675 2921.225 4796.455 ;
        RECT 3291.185 1959.695 3301.965 1981.675 ;
        RECT 3291.100 1910.305 3301.880 1932.285 ;
        RECT 263.335 1176.140 264.515 1177.320 ;
        RECT 263.335 1174.540 264.515 1175.720 ;
        RECT 263.335 1172.940 264.515 1174.120 ;
        RECT 263.335 1171.340 264.515 1172.520 ;
        RECT 263.335 1169.740 264.515 1170.920 ;
        RECT 263.335 1168.140 264.515 1169.320 ;
        RECT 263.335 1166.540 264.515 1167.720 ;
        RECT 263.335 1164.940 264.515 1166.120 ;
        RECT 263.335 1163.340 264.515 1164.520 ;
        RECT 1924.345 1163.325 1927.125 1177.305 ;
        RECT 1999.595 1163.325 2002.375 1177.305 ;
        RECT 3247.925 1176.125 3249.105 1177.305 ;
        RECT 3247.925 1174.525 3249.105 1175.705 ;
        RECT 3247.925 1172.925 3249.105 1174.105 ;
        RECT 3247.925 1171.325 3249.105 1172.505 ;
        RECT 3247.925 1169.725 3249.105 1170.905 ;
        RECT 3247.925 1168.125 3249.105 1169.305 ;
        RECT 3247.925 1166.525 3249.105 1167.705 ;
        RECT 3247.925 1164.925 3249.105 1166.105 ;
        RECT 3247.925 1163.325 3249.105 1164.505 ;
      LAYER met5 ;
        RECT 2848.090 4784.480 3302.990 4797.480 ;
        RECT 3289.990 4772.440 3302.990 4784.480 ;
        RECT 3250.080 4769.340 3302.990 4772.440 ;
        RECT 3289.990 1198.520 3302.990 4769.340 ;
        RECT 3250.020 1195.420 3302.990 1198.520 ;
        RECT 3289.990 1177.830 3302.990 1195.420 ;
        RECT 261.830 1162.830 3302.990 1177.830 ;
    END
  END vssa1_core
  PIN vdda1_core
    PORT
      LAYER met3 ;
        RECT 3305.750 3973.105 3358.980 3997.005 ;
        RECT 3305.750 3923.210 3358.980 3947.110 ;
        RECT 3305.200 2400.105 3358.390 2424.005 ;
        RECT 3305.200 2350.210 3358.390 2374.110 ;
      LAYER via3 ;
        RECT 3306.470 3973.730 3318.390 3996.450 ;
        RECT 3306.400 3923.760 3318.320 3946.480 ;
        RECT 3306.735 2400.935 3318.255 2423.255 ;
        RECT 3306.805 2350.985 3318.325 2373.305 ;
      LAYER met4 ;
        RECT 3261.790 4764.560 3319.020 4767.680 ;
        RECT 3305.900 3973.100 3318.900 3997.050 ;
        RECT 3305.960 3923.230 3318.960 3947.180 ;
        RECT 3305.920 2400.100 3318.960 2423.980 ;
        RECT 3305.980 2350.250 3319.020 2374.130 ;
        RECT 267.200 1163.590 270.300 1200.260 ;
        RECT 267.200 1160.490 286.550 1163.590 ;
        RECT 283.450 1142.510 286.550 1160.490 ;
        RECT 1889.860 1157.810 1890.760 1157.880 ;
        RECT 1965.110 1157.810 1966.010 1157.880 ;
        RECT 1886.720 1144.770 1890.760 1157.810 ;
        RECT 1961.970 1144.770 1966.010 1157.810 ;
        RECT 1889.860 1141.720 1890.760 1144.770 ;
        RECT 1965.110 1141.720 1966.010 1144.770 ;
        RECT 3242.180 1142.310 3245.280 1200.280 ;
        RECT 3264.640 1200.190 3318.950 1203.370 ;
        RECT 3305.970 1196.190 3318.950 1200.190 ;
      LAYER via4 ;
        RECT 3262.775 4765.530 3263.955 4766.710 ;
        RECT 3264.375 4765.530 3265.555 4766.710 ;
        RECT 3265.975 4765.530 3267.155 4766.710 ;
        RECT 3267.575 4765.530 3268.755 4766.710 ;
        RECT 3269.175 4765.530 3270.355 4766.710 ;
        RECT 3270.775 4765.530 3271.955 4766.710 ;
        RECT 3272.375 4765.530 3273.555 4766.710 ;
        RECT 3273.975 4765.530 3275.155 4766.710 ;
        RECT 3275.575 4765.530 3276.755 4766.710 ;
        RECT 3277.175 4765.530 3278.355 4766.710 ;
        RECT 3278.775 4765.530 3279.955 4766.710 ;
        RECT 3280.375 4765.530 3281.555 4766.710 ;
        RECT 3281.975 4765.530 3283.155 4766.710 ;
        RECT 3283.575 4765.530 3284.755 4766.710 ;
        RECT 3306.295 4765.555 3307.475 4766.735 ;
        RECT 3307.895 4765.555 3309.075 4766.735 ;
        RECT 3309.495 4765.555 3310.675 4766.735 ;
        RECT 3311.095 4765.555 3312.275 4766.735 ;
        RECT 3312.695 4765.555 3313.875 4766.735 ;
        RECT 3314.295 4765.555 3315.475 4766.735 ;
        RECT 3315.895 4765.555 3317.075 4766.735 ;
        RECT 3317.495 4765.555 3318.675 4766.735 ;
        RECT 3307.040 3974.100 3317.820 3996.080 ;
        RECT 3306.970 3924.130 3317.750 3946.110 ;
        RECT 3307.105 2401.105 3317.885 2423.085 ;
        RECT 3307.175 2351.155 3317.955 2373.135 ;
        RECT 3265.815 1201.145 3266.995 1202.325 ;
        RECT 3267.415 1201.145 3268.595 1202.325 ;
        RECT 3269.015 1201.145 3270.195 1202.325 ;
        RECT 3270.615 1201.145 3271.795 1202.325 ;
        RECT 3272.215 1201.145 3273.395 1202.325 ;
        RECT 3273.815 1201.145 3274.995 1202.325 ;
        RECT 3275.415 1201.145 3276.595 1202.325 ;
        RECT 3277.015 1201.145 3278.195 1202.325 ;
        RECT 3278.615 1201.145 3279.795 1202.325 ;
        RECT 3280.215 1201.145 3281.395 1202.325 ;
        RECT 3281.815 1201.145 3282.995 1202.325 ;
        RECT 3283.415 1201.145 3284.595 1202.325 ;
        RECT 284.375 1156.120 285.555 1157.300 ;
        RECT 284.375 1154.520 285.555 1155.700 ;
        RECT 284.375 1152.920 285.555 1154.100 ;
        RECT 284.375 1151.320 285.555 1152.500 ;
        RECT 284.375 1149.720 285.555 1150.900 ;
        RECT 284.375 1148.120 285.555 1149.300 ;
        RECT 284.375 1146.520 285.555 1147.700 ;
        RECT 284.375 1144.920 285.555 1146.100 ;
        RECT 1887.325 1145.760 1890.105 1156.540 ;
        RECT 1962.575 1145.760 1965.355 1156.540 ;
        RECT 284.375 1143.320 285.555 1144.500 ;
        RECT 3307.130 1196.780 3317.910 1202.760 ;
        RECT 3243.135 1156.115 3244.315 1157.295 ;
        RECT 3243.135 1154.515 3244.315 1155.695 ;
        RECT 3243.135 1152.915 3244.315 1154.095 ;
        RECT 3243.135 1151.315 3244.315 1152.495 ;
        RECT 3243.135 1149.715 3244.315 1150.895 ;
        RECT 3243.135 1148.115 3244.315 1149.295 ;
        RECT 3243.135 1146.515 3244.315 1147.695 ;
        RECT 3243.135 1144.915 3244.315 1146.095 ;
        RECT 3243.135 1143.315 3244.315 1144.495 ;
      LAYER met5 ;
        RECT 3245.280 4764.540 3285.780 4767.640 ;
        RECT 3245.190 1200.220 3285.680 1203.320 ;
        RECT 3305.990 1157.830 3318.990 4768.330 ;
        RECT 282.560 1142.830 3318.990 1157.830 ;
    END
  END vdda1_core
  OBS
      LAYER met3 ;
        RECT 519.390 4827.130 525.390 4923.980 ;
        RECT 527.390 4860.080 533.390 4929.950 ;
        RECT 776.390 4827.130 782.390 4923.980 ;
        RECT 784.390 4860.080 790.390 4929.950 ;
        RECT 1033.390 4827.130 1039.390 4923.980 ;
        RECT 1041.390 4860.080 1047.390 4929.950 ;
        RECT 1290.390 4827.130 1296.390 4923.980 ;
        RECT 1298.390 4860.080 1304.390 4929.950 ;
        RECT 1548.390 4827.130 1554.390 4923.980 ;
        RECT 1556.390 4860.080 1562.390 4929.950 ;
        RECT 1800.390 4827.130 1806.390 4923.980 ;
        RECT 1808.390 4860.080 1814.390 4929.950 ;
        RECT 2137.390 4827.130 2143.390 4923.980 ;
        RECT 2145.390 4860.080 2151.390 4929.950 ;
        RECT 2522.390 4827.130 2528.390 4923.980 ;
        RECT 2530.390 4860.080 2536.390 4929.950 ;
        RECT 2779.390 4827.130 2785.390 4923.980 ;
        RECT 2787.390 4860.080 2793.390 4929.950 ;
        RECT 190.880 4590.120 279.870 4596.120 ;
        RECT 174.810 4582.120 275.050 4588.120 ;
        RECT 59.030 4558.000 128.200 4564.000 ;
        RECT 3222.970 4556.410 3528.910 4562.410 ;
        RECT 65.000 4550.000 161.150 4556.000 ;
        RECT 3227.790 4548.410 3522.840 4554.410 ;
        RECT 3399.460 4540.000 3469.880 4546.000 ;
        RECT 3366.510 4532.000 3463.910 4538.000 ;
        RECT 3222.970 4330.410 3349.040 4336.410 ;
        RECT 3227.790 4322.410 3333.270 4328.410 ;
        RECT 3222.970 4105.410 3346.210 4111.410 ;
        RECT 3227.790 4097.410 3333.430 4103.410 ;
        RECT 190.880 3961.120 279.870 3967.120 ;
        RECT 174.810 3953.120 275.050 3959.120 ;
        RECT 59.030 3929.000 128.200 3935.000 ;
        RECT 65.000 3921.000 161.150 3927.000 ;
        RECT 190.880 3753.120 279.870 3759.120 ;
        RECT 174.810 3745.120 275.050 3751.120 ;
        RECT 59.030 3713.000 128.200 3719.000 ;
        RECT 65.000 3705.000 161.150 3711.000 ;
        RECT 3222.970 3664.410 3528.960 3670.410 ;
        RECT 3227.790 3656.410 3522.890 3662.410 ;
        RECT 3399.510 3648.000 3469.930 3654.000 ;
        RECT 3366.560 3640.000 3463.960 3646.000 ;
        RECT 190.880 3529.120 279.870 3535.120 ;
        RECT 174.810 3521.120 275.050 3527.120 ;
        RECT 59.030 3497.000 128.200 3503.000 ;
        RECT 65.000 3489.000 161.150 3495.000 ;
        RECT 3222.970 3439.410 3528.960 3445.410 ;
        RECT 3227.790 3431.410 3522.890 3437.410 ;
        RECT 3399.510 3423.000 3469.930 3429.000 ;
        RECT 3366.560 3415.000 3463.960 3421.000 ;
        RECT 190.880 3313.120 279.870 3319.120 ;
        RECT 174.810 3305.120 275.050 3311.120 ;
        RECT 59.030 3281.000 128.200 3287.000 ;
        RECT 65.000 3273.000 161.150 3279.000 ;
        RECT 3222.970 3213.410 3528.960 3219.410 ;
        RECT 3227.790 3205.410 3522.890 3211.410 ;
        RECT 3399.510 3197.000 3469.930 3203.000 ;
        RECT 3366.560 3189.000 3463.960 3195.000 ;
        RECT 190.880 3097.120 279.870 3103.120 ;
        RECT 174.810 3089.120 275.050 3095.120 ;
        RECT 59.030 3065.000 128.200 3071.000 ;
        RECT 65.000 3057.000 161.150 3063.000 ;
        RECT 3222.970 2988.410 3528.960 2994.410 ;
        RECT 3266.440 2980.410 3522.890 2986.410 ;
        RECT 3227.790 2974.410 3272.890 2980.410 ;
        RECT 3399.510 2972.000 3469.930 2978.000 ;
        RECT 3366.560 2964.000 3463.960 2970.000 ;
        RECT 190.880 2886.420 279.870 2892.420 ;
        RECT 174.810 2878.420 275.050 2884.420 ;
        RECT 59.030 2849.000 128.200 2855.000 ;
        RECT 65.000 2841.000 161.150 2847.000 ;
        RECT 3222.970 2762.410 3528.960 2768.410 ;
        RECT 3227.790 2754.410 3522.890 2760.410 ;
        RECT 3399.510 2746.000 3469.930 2752.000 ;
        RECT 3366.560 2738.000 3463.960 2744.000 ;
        RECT 190.880 2665.120 279.870 2671.120 ;
        RECT 174.810 2657.120 275.050 2663.120 ;
        RECT 59.030 2633.000 128.200 2639.000 ;
        RECT 65.000 2625.000 161.150 2631.000 ;
        RECT 3222.970 2537.410 3528.960 2543.410 ;
        RECT 3227.790 2529.410 3522.890 2535.410 ;
        RECT 3399.510 2521.000 3469.930 2527.000 ;
        RECT 3366.560 2513.000 3463.960 2519.000 ;
        RECT 3222.970 2323.410 3268.680 2326.410 ;
        RECT 3222.970 2320.410 3528.960 2323.410 ;
        RECT 3262.730 2317.410 3528.960 2320.410 ;
        RECT 3227.790 2309.410 3522.890 2315.410 ;
        RECT 3399.510 2301.000 3469.930 2307.000 ;
        RECT 3366.560 2293.000 3463.960 2299.000 ;
        RECT 190.880 2027.120 279.870 2033.120 ;
        RECT 174.810 2019.120 275.050 2025.120 ;
        RECT 59.030 1995.000 128.200 2001.000 ;
        RECT 65.000 1987.000 161.150 1993.000 ;
        RECT 3222.970 1876.410 3528.960 1882.410 ;
        RECT 3227.790 1868.410 3522.890 1874.410 ;
        RECT 3399.510 1860.000 3469.930 1866.000 ;
        RECT 3366.560 1852.000 3463.960 1858.000 ;
        RECT 190.880 1811.120 279.870 1817.120 ;
        RECT 174.810 1803.120 275.050 1809.120 ;
        RECT 59.030 1779.000 128.200 1785.000 ;
        RECT 65.000 1771.000 161.150 1777.000 ;
        RECT 3222.970 1657.410 3298.210 1663.410 ;
        RECT 3292.210 1656.410 3298.210 1657.410 ;
        RECT 3292.210 1650.410 3528.960 1656.410 ;
        RECT 3227.790 1642.410 3522.890 1648.410 ;
        RECT 3399.510 1634.000 3469.930 1640.000 ;
        RECT 3366.560 1626.000 3463.960 1632.000 ;
        RECT 190.880 1600.120 279.870 1606.120 ;
        RECT 174.810 1592.120 275.050 1598.120 ;
        RECT 59.030 1563.000 128.200 1569.000 ;
        RECT 65.000 1555.000 161.150 1561.000 ;
        RECT 3222.970 1425.410 3528.960 1431.410 ;
        RECT 3227.790 1417.410 3522.890 1423.410 ;
        RECT 3399.510 1409.000 3469.930 1415.000 ;
        RECT 3366.560 1401.000 3463.960 1407.000 ;
        RECT 190.880 1379.120 279.870 1385.120 ;
        RECT 174.810 1371.120 275.050 1377.120 ;
        RECT 59.030 1347.000 128.200 1353.000 ;
        RECT 65.000 1339.000 161.150 1345.000 ;
        RECT 3346.270 1200.410 3528.960 1206.410 ;
        RECT 3327.990 1192.410 3522.890 1198.410 ;
        RECT 3399.510 1184.000 3469.930 1190.000 ;
        RECT 3366.560 1176.000 3463.960 1182.000 ;
        RECT 59.030 1131.000 128.200 1137.000 ;
        RECT 65.000 1123.000 161.150 1129.000 ;
        RECT 3346.270 974.410 3528.960 980.410 ;
        RECT 3327.990 966.410 3522.890 972.410 ;
        RECT 3399.510 958.000 3469.930 964.000 ;
        RECT 3366.560 950.000 3463.960 956.000 ;
        RECT 59.030 915.000 128.200 921.000 ;
        RECT 65.000 907.000 161.150 913.000 ;
        RECT 3346.270 749.410 3528.960 755.410 ;
        RECT 3327.990 741.410 3522.890 747.410 ;
        RECT 3399.510 733.000 3469.930 739.000 ;
        RECT 3366.560 725.000 3463.960 731.000 ;
        RECT 3346.270 523.410 3528.960 529.410 ;
        RECT 3327.990 515.410 3522.890 521.410 ;
        RECT 3399.510 507.000 3469.930 513.000 ;
        RECT 3366.560 499.000 3463.960 505.000 ;
        RECT 710.230 0.000 714.520 34.410 ;
        RECT 717.890 6.070 722.180 36.535 ;
        RECT 3179.660 0.100 3188.360 50.630 ;
        RECT 3237.200 9.540 3254.440 56.280 ;
      LAYER via3 ;
        RECT 527.640 4926.025 533.160 4929.545 ;
        RECT 519.650 4920.005 525.170 4923.525 ;
        RECT 784.640 4926.025 790.160 4929.545 ;
        RECT 527.795 4860.645 532.915 4864.165 ;
        RECT 776.650 4920.005 782.170 4923.525 ;
        RECT 519.940 4827.935 525.060 4831.455 ;
        RECT 1041.640 4926.025 1047.160 4929.545 ;
        RECT 784.795 4860.645 789.915 4864.165 ;
        RECT 1033.650 4920.005 1039.170 4923.525 ;
        RECT 776.940 4827.935 782.060 4831.455 ;
        RECT 1298.640 4926.025 1304.160 4929.545 ;
        RECT 1041.795 4860.645 1046.915 4864.165 ;
        RECT 1290.650 4920.005 1296.170 4923.525 ;
        RECT 1033.940 4827.935 1039.060 4831.455 ;
        RECT 1556.640 4926.025 1562.160 4929.545 ;
        RECT 1298.795 4860.645 1303.915 4864.165 ;
        RECT 1548.650 4920.005 1554.170 4923.525 ;
        RECT 1290.940 4827.935 1296.060 4831.455 ;
        RECT 1808.640 4926.025 1814.160 4929.545 ;
        RECT 1556.795 4860.645 1561.915 4864.165 ;
        RECT 1800.650 4920.005 1806.170 4923.525 ;
        RECT 1548.940 4827.935 1554.060 4831.455 ;
        RECT 2145.640 4926.025 2151.160 4929.545 ;
        RECT 1808.795 4860.645 1813.915 4864.165 ;
        RECT 2137.650 4920.005 2143.170 4923.525 ;
        RECT 1800.940 4827.935 1806.060 4831.455 ;
        RECT 2530.640 4926.025 2536.160 4929.545 ;
        RECT 2145.795 4860.645 2150.915 4864.165 ;
        RECT 2522.650 4920.005 2528.170 4923.525 ;
        RECT 2137.940 4827.935 2143.060 4831.455 ;
        RECT 2787.640 4926.025 2793.160 4929.545 ;
        RECT 2530.795 4860.645 2535.915 4864.165 ;
        RECT 2779.650 4920.005 2785.170 4923.525 ;
        RECT 2522.940 4827.935 2528.060 4831.455 ;
        RECT 2787.795 4860.645 2792.915 4864.165 ;
        RECT 2779.940 4827.935 2785.060 4831.455 ;
        RECT 191.460 4590.455 203.380 4595.575 ;
        RECT 277.195 4590.340 279.515 4595.860 ;
        RECT 175.410 4582.545 187.330 4587.665 ;
        RECT 272.375 4582.380 274.695 4587.900 ;
        RECT 59.435 4558.250 62.955 4563.770 ;
        RECT 124.115 4558.405 127.635 4563.525 ;
        RECT 3223.170 4556.665 3225.890 4562.185 ;
        RECT 3347.025 4556.925 3352.145 4562.045 ;
        RECT 3524.950 4556.645 3528.070 4562.165 ;
        RECT 65.455 4550.260 68.975 4555.780 ;
        RECT 156.825 4550.550 160.345 4555.670 ;
        RECT 3227.960 4548.645 3230.680 4554.165 ;
        RECT 3328.495 4548.835 3333.615 4553.955 ;
        RECT 3518.960 4548.665 3522.080 4554.185 ;
        RECT 3400.025 4540.405 3403.545 4545.525 ;
        RECT 3465.955 4540.250 3469.475 4545.770 ;
        RECT 3367.315 4532.550 3370.835 4537.670 ;
        RECT 3459.935 4532.260 3463.455 4537.780 ;
        RECT 3223.170 4330.665 3225.890 4336.185 ;
        RECT 3343.715 4330.905 3348.435 4336.025 ;
        RECT 3227.960 4322.645 3230.680 4328.165 ;
        RECT 3327.735 4322.865 3332.855 4327.985 ;
        RECT 3223.170 4105.665 3225.890 4111.185 ;
        RECT 3340.570 4105.860 3345.690 4110.980 ;
        RECT 3227.960 4097.645 3230.680 4103.165 ;
        RECT 3327.850 4097.850 3332.970 4102.970 ;
        RECT 191.460 3961.455 203.380 3966.575 ;
        RECT 277.195 3961.340 279.515 3966.860 ;
        RECT 175.410 3953.545 187.330 3958.665 ;
        RECT 272.375 3953.380 274.695 3958.900 ;
        RECT 59.435 3929.250 62.955 3934.770 ;
        RECT 124.115 3929.405 127.635 3934.525 ;
        RECT 65.455 3921.260 68.975 3926.780 ;
        RECT 156.825 3921.550 160.345 3926.670 ;
        RECT 191.460 3753.455 203.380 3758.575 ;
        RECT 277.195 3753.340 279.515 3758.860 ;
        RECT 175.410 3745.545 187.330 3750.665 ;
        RECT 272.375 3745.380 274.695 3750.900 ;
        RECT 59.435 3713.250 62.955 3718.770 ;
        RECT 124.115 3713.405 127.635 3718.525 ;
        RECT 65.455 3705.260 68.975 3710.780 ;
        RECT 156.825 3705.550 160.345 3710.670 ;
        RECT 3223.170 3664.665 3225.890 3670.185 ;
        RECT 3347.075 3664.925 3352.195 3670.045 ;
        RECT 3525.000 3664.645 3528.120 3670.165 ;
        RECT 3227.960 3656.645 3230.680 3662.165 ;
        RECT 3328.545 3656.835 3333.665 3661.955 ;
        RECT 3519.010 3656.665 3522.130 3662.185 ;
        RECT 3400.075 3648.405 3403.595 3653.525 ;
        RECT 3466.005 3648.250 3469.525 3653.770 ;
        RECT 3367.365 3640.550 3370.885 3645.670 ;
        RECT 3459.985 3640.260 3463.505 3645.780 ;
        RECT 191.460 3529.455 203.380 3534.575 ;
        RECT 277.195 3529.340 279.515 3534.860 ;
        RECT 175.410 3521.545 187.330 3526.665 ;
        RECT 272.375 3521.380 274.695 3526.900 ;
        RECT 59.435 3497.250 62.955 3502.770 ;
        RECT 124.115 3497.405 127.635 3502.525 ;
        RECT 65.455 3489.260 68.975 3494.780 ;
        RECT 156.825 3489.550 160.345 3494.670 ;
        RECT 3223.170 3439.665 3225.890 3445.185 ;
        RECT 3347.075 3439.925 3352.195 3445.045 ;
        RECT 3525.000 3439.645 3528.120 3445.165 ;
        RECT 3227.960 3431.645 3230.680 3437.165 ;
        RECT 3328.545 3431.835 3333.665 3436.955 ;
        RECT 3519.010 3431.665 3522.130 3437.185 ;
        RECT 3400.075 3423.405 3403.595 3428.525 ;
        RECT 3466.005 3423.250 3469.525 3428.770 ;
        RECT 3367.365 3415.550 3370.885 3420.670 ;
        RECT 3459.985 3415.260 3463.505 3420.780 ;
        RECT 191.460 3313.455 203.380 3318.575 ;
        RECT 277.195 3313.340 279.515 3318.860 ;
        RECT 175.410 3305.545 187.330 3310.665 ;
        RECT 272.375 3305.380 274.695 3310.900 ;
        RECT 59.435 3281.250 62.955 3286.770 ;
        RECT 124.115 3281.405 127.635 3286.525 ;
        RECT 65.455 3273.260 68.975 3278.780 ;
        RECT 156.825 3273.550 160.345 3278.670 ;
        RECT 3223.170 3213.665 3225.890 3219.185 ;
        RECT 3347.075 3213.925 3352.195 3219.045 ;
        RECT 3525.000 3213.645 3528.120 3219.165 ;
        RECT 3227.960 3205.645 3230.680 3211.165 ;
        RECT 3328.545 3205.835 3333.665 3210.955 ;
        RECT 3519.010 3205.665 3522.130 3211.185 ;
        RECT 3400.075 3197.405 3403.595 3202.525 ;
        RECT 3466.005 3197.250 3469.525 3202.770 ;
        RECT 3367.365 3189.550 3370.885 3194.670 ;
        RECT 3459.985 3189.260 3463.505 3194.780 ;
        RECT 191.460 3097.455 203.380 3102.575 ;
        RECT 277.195 3097.340 279.515 3102.860 ;
        RECT 175.410 3089.545 187.330 3094.665 ;
        RECT 272.375 3089.380 274.695 3094.900 ;
        RECT 59.435 3065.250 62.955 3070.770 ;
        RECT 124.115 3065.405 127.635 3070.525 ;
        RECT 65.455 3057.260 68.975 3062.780 ;
        RECT 156.825 3057.550 160.345 3062.670 ;
        RECT 3223.170 2988.665 3225.890 2994.185 ;
        RECT 3347.075 2988.925 3352.195 2994.045 ;
        RECT 3525.000 2988.645 3528.120 2994.165 ;
        RECT 3328.545 2980.835 3333.665 2985.955 ;
        RECT 3519.010 2980.665 3522.130 2986.185 ;
        RECT 3227.960 2974.645 3230.680 2980.165 ;
        RECT 3400.075 2972.405 3403.595 2977.525 ;
        RECT 3466.005 2972.250 3469.525 2977.770 ;
        RECT 3367.365 2964.550 3370.885 2969.670 ;
        RECT 3459.985 2964.260 3463.505 2969.780 ;
        RECT 191.460 2886.755 203.380 2891.875 ;
        RECT 277.195 2886.640 279.515 2892.160 ;
        RECT 175.410 2878.845 187.330 2883.965 ;
        RECT 272.375 2878.680 274.695 2884.200 ;
        RECT 59.435 2849.250 62.955 2854.770 ;
        RECT 124.115 2849.405 127.635 2854.525 ;
        RECT 65.455 2841.260 68.975 2846.780 ;
        RECT 156.825 2841.550 160.345 2846.670 ;
        RECT 3223.170 2762.665 3225.890 2768.185 ;
        RECT 3347.075 2762.925 3352.195 2768.045 ;
        RECT 3525.000 2762.645 3528.120 2768.165 ;
        RECT 3227.960 2754.645 3230.680 2760.165 ;
        RECT 3328.545 2754.835 3333.665 2759.955 ;
        RECT 3519.010 2754.665 3522.130 2760.185 ;
        RECT 3400.075 2746.405 3403.595 2751.525 ;
        RECT 3466.005 2746.250 3469.525 2751.770 ;
        RECT 3367.365 2738.550 3370.885 2743.670 ;
        RECT 3459.985 2738.260 3463.505 2743.780 ;
        RECT 191.460 2665.455 203.380 2670.575 ;
        RECT 277.195 2665.340 279.515 2670.860 ;
        RECT 175.410 2657.545 187.330 2662.665 ;
        RECT 272.375 2657.380 274.695 2662.900 ;
        RECT 59.435 2633.250 62.955 2638.770 ;
        RECT 124.115 2633.405 127.635 2638.525 ;
        RECT 65.455 2625.260 68.975 2630.780 ;
        RECT 156.825 2625.550 160.345 2630.670 ;
        RECT 3223.170 2537.665 3225.890 2543.185 ;
        RECT 3347.075 2537.925 3352.195 2543.045 ;
        RECT 3525.000 2537.645 3528.120 2543.165 ;
        RECT 3227.960 2529.645 3230.680 2535.165 ;
        RECT 3328.545 2529.835 3333.665 2534.955 ;
        RECT 3519.010 2529.665 3522.130 2535.185 ;
        RECT 3400.075 2521.405 3403.595 2526.525 ;
        RECT 3466.005 2521.250 3469.525 2526.770 ;
        RECT 3367.365 2513.550 3370.885 2518.670 ;
        RECT 3459.985 2513.260 3463.505 2518.780 ;
        RECT 3223.170 2320.665 3225.890 2326.185 ;
        RECT 3347.075 2317.925 3352.195 2323.045 ;
        RECT 3525.000 2317.645 3528.120 2323.165 ;
        RECT 3227.960 2309.645 3230.680 2315.165 ;
        RECT 3328.545 2309.835 3333.665 2314.955 ;
        RECT 3519.010 2309.665 3522.130 2315.185 ;
        RECT 3400.075 2301.405 3403.595 2306.525 ;
        RECT 3466.005 2301.250 3469.525 2306.770 ;
        RECT 3367.365 2293.550 3370.885 2298.670 ;
        RECT 3459.985 2293.260 3463.505 2298.780 ;
        RECT 191.460 2027.455 203.380 2032.575 ;
        RECT 277.195 2027.340 279.515 2032.860 ;
        RECT 175.410 2019.545 187.330 2024.665 ;
        RECT 272.375 2019.380 274.695 2024.900 ;
        RECT 59.435 1995.250 62.955 2000.770 ;
        RECT 124.115 1995.405 127.635 2000.525 ;
        RECT 65.455 1987.260 68.975 1992.780 ;
        RECT 156.825 1987.550 160.345 1992.670 ;
        RECT 3223.170 1876.665 3225.890 1882.185 ;
        RECT 3347.075 1876.925 3352.195 1882.045 ;
        RECT 3525.000 1876.645 3528.120 1882.165 ;
        RECT 3227.960 1868.645 3230.680 1874.165 ;
        RECT 3328.545 1868.835 3333.665 1873.955 ;
        RECT 3519.010 1868.665 3522.130 1874.185 ;
        RECT 3400.075 1860.405 3403.595 1865.525 ;
        RECT 3466.005 1860.250 3469.525 1865.770 ;
        RECT 3367.365 1852.550 3370.885 1857.670 ;
        RECT 3459.985 1852.260 3463.505 1857.780 ;
        RECT 191.460 1811.455 203.380 1816.575 ;
        RECT 277.195 1811.340 279.515 1816.860 ;
        RECT 175.410 1803.545 187.330 1808.665 ;
        RECT 272.375 1803.380 274.695 1808.900 ;
        RECT 59.435 1779.250 62.955 1784.770 ;
        RECT 124.115 1779.405 127.635 1784.525 ;
        RECT 65.455 1771.260 68.975 1776.780 ;
        RECT 156.825 1771.550 160.345 1776.670 ;
        RECT 3223.170 1657.665 3225.890 1663.185 ;
        RECT 3347.075 1650.925 3352.195 1656.045 ;
        RECT 3525.000 1650.645 3528.120 1656.165 ;
        RECT 3227.960 1642.645 3230.680 1648.165 ;
        RECT 3328.545 1642.835 3333.665 1647.955 ;
        RECT 3519.010 1642.665 3522.130 1648.185 ;
        RECT 3400.075 1634.405 3403.595 1639.525 ;
        RECT 3466.005 1634.250 3469.525 1639.770 ;
        RECT 3367.365 1626.550 3370.885 1631.670 ;
        RECT 3459.985 1626.260 3463.505 1631.780 ;
        RECT 191.460 1600.455 203.380 1605.575 ;
        RECT 277.195 1600.340 279.515 1605.860 ;
        RECT 175.410 1592.545 187.330 1597.665 ;
        RECT 272.375 1592.380 274.695 1597.900 ;
        RECT 59.435 1563.250 62.955 1568.770 ;
        RECT 124.115 1563.405 127.635 1568.525 ;
        RECT 65.455 1555.260 68.975 1560.780 ;
        RECT 156.825 1555.550 160.345 1560.670 ;
        RECT 3223.170 1425.665 3225.890 1431.185 ;
        RECT 3347.075 1425.925 3352.195 1431.045 ;
        RECT 3525.000 1425.645 3528.120 1431.165 ;
        RECT 3227.960 1417.645 3230.680 1423.165 ;
        RECT 3328.545 1417.835 3333.665 1422.955 ;
        RECT 3519.010 1417.665 3522.130 1423.185 ;
        RECT 3400.075 1409.405 3403.595 1414.525 ;
        RECT 3466.005 1409.250 3469.525 1414.770 ;
        RECT 3367.365 1401.550 3370.885 1406.670 ;
        RECT 3459.985 1401.260 3463.505 1406.780 ;
        RECT 191.460 1379.455 203.380 1384.575 ;
        RECT 277.195 1379.340 279.515 1384.860 ;
        RECT 175.410 1371.545 187.330 1376.665 ;
        RECT 272.375 1371.380 274.695 1376.900 ;
        RECT 59.435 1347.250 62.955 1352.770 ;
        RECT 124.115 1347.405 127.635 1352.525 ;
        RECT 65.455 1339.260 68.975 1344.780 ;
        RECT 156.825 1339.550 160.345 1344.670 ;
        RECT 3347.075 1200.925 3352.195 1206.045 ;
        RECT 3525.000 1200.645 3528.120 1206.165 ;
        RECT 3328.545 1192.835 3333.665 1197.955 ;
        RECT 3519.010 1192.665 3522.130 1198.185 ;
        RECT 3400.075 1184.405 3403.595 1189.525 ;
        RECT 3466.005 1184.250 3469.525 1189.770 ;
        RECT 3367.365 1176.550 3370.885 1181.670 ;
        RECT 3459.985 1176.260 3463.505 1181.780 ;
        RECT 59.435 1131.250 62.955 1136.770 ;
        RECT 124.115 1131.405 127.635 1136.525 ;
        RECT 65.455 1123.260 68.975 1128.780 ;
        RECT 156.825 1123.550 160.345 1128.670 ;
        RECT 3347.075 974.925 3352.195 980.045 ;
        RECT 3525.000 974.645 3528.120 980.165 ;
        RECT 3328.545 966.835 3333.665 971.955 ;
        RECT 3519.010 966.665 3522.130 972.185 ;
        RECT 3400.075 958.405 3403.595 963.525 ;
        RECT 3466.005 958.250 3469.525 963.770 ;
        RECT 3367.365 950.550 3370.885 955.670 ;
        RECT 3459.985 950.260 3463.505 955.780 ;
        RECT 59.435 915.250 62.955 920.770 ;
        RECT 124.115 915.405 127.635 920.525 ;
        RECT 65.455 907.260 68.975 912.780 ;
        RECT 156.825 907.550 160.345 912.670 ;
        RECT 3347.075 749.925 3352.195 755.045 ;
        RECT 3525.000 749.645 3528.120 755.165 ;
        RECT 3328.545 741.835 3333.665 746.955 ;
        RECT 3519.010 741.665 3522.130 747.185 ;
        RECT 3400.075 733.405 3403.595 738.525 ;
        RECT 3466.005 733.250 3469.525 738.770 ;
        RECT 3367.365 725.550 3370.885 730.670 ;
        RECT 3459.985 725.260 3463.505 730.780 ;
        RECT 3347.075 523.925 3352.195 529.045 ;
        RECT 3525.000 523.645 3528.120 529.165 ;
        RECT 3328.545 515.835 3333.665 520.955 ;
        RECT 3519.010 515.665 3522.130 521.185 ;
        RECT 3400.075 507.405 3403.595 512.525 ;
        RECT 3466.005 507.250 3469.525 512.770 ;
        RECT 3367.365 499.550 3370.885 504.670 ;
        RECT 3459.985 499.260 3463.505 504.780 ;
        RECT 3179.865 41.605 3188.185 50.325 ;
        RECT 718.075 35.480 721.995 36.200 ;
        RECT 710.415 33.500 714.335 34.220 ;
        RECT 718.100 6.445 722.020 10.365 ;
        RECT 710.430 0.405 714.350 4.325 ;
        RECT 3237.805 43.690 3253.725 55.610 ;
        RECT 3180.080 0.610 3188.000 4.130 ;
      LAYER met4 ;
        RECT 470.000 4925.740 533.440 4929.740 ;
        RECT 727.000 4925.740 790.440 4929.740 ;
        RECT 984.000 4925.740 1047.440 4929.740 ;
        RECT 1241.000 4925.740 1304.440 4929.740 ;
        RECT 1499.000 4925.740 1562.440 4929.740 ;
        RECT 1751.000 4925.740 1814.440 4929.740 ;
        RECT 2088.000 4925.740 2151.440 4929.740 ;
        RECT 2473.000 4925.740 2536.440 4929.740 ;
        RECT 2730.000 4925.740 2793.440 4929.740 ;
        RECT 461.630 4919.740 526.550 4923.740 ;
        RECT 718.630 4919.740 783.550 4923.740 ;
        RECT 975.630 4919.740 1040.550 4923.740 ;
        RECT 1232.630 4919.740 1297.550 4923.740 ;
        RECT 1490.630 4919.740 1555.550 4923.740 ;
        RECT 1742.630 4919.740 1807.550 4923.740 ;
        RECT 2079.630 4919.740 2144.550 4923.740 ;
        RECT 2464.630 4919.740 2529.550 4923.740 ;
        RECT 2721.630 4919.740 2786.550 4923.740 ;
        RECT 527.660 4860.520 533.050 4864.290 ;
        RECT 784.660 4860.520 790.050 4864.290 ;
        RECT 1041.660 4860.520 1047.050 4864.290 ;
        RECT 1298.660 4860.520 1304.050 4864.290 ;
        RECT 1556.660 4860.520 1562.050 4864.290 ;
        RECT 1808.660 4860.520 1814.050 4864.290 ;
        RECT 2145.660 4860.520 2151.050 4864.290 ;
        RECT 2530.660 4860.520 2536.050 4864.290 ;
        RECT 2787.660 4860.520 2793.050 4864.290 ;
        RECT 519.790 4827.790 525.210 4831.600 ;
        RECT 776.790 4827.790 782.210 4831.600 ;
        RECT 1033.790 4827.790 1039.210 4831.600 ;
        RECT 1290.790 4827.790 1296.210 4831.600 ;
        RECT 1548.790 4827.790 1554.210 4831.600 ;
        RECT 1800.790 4827.790 1806.210 4831.600 ;
        RECT 2137.790 4827.790 2143.210 4831.600 ;
        RECT 2522.790 4827.790 2528.210 4831.600 ;
        RECT 2779.790 4827.790 2785.210 4831.600 ;
        RECT 174.855 4759.770 251.960 4762.840 ;
        RECT 190.890 4754.870 252.090 4758.130 ;
        RECT 3261.470 4750.140 3337.040 4753.350 ;
        RECT 3261.330 4745.300 3353.010 4748.510 ;
        RECT 190.890 4590.110 203.850 4596.130 ;
        RECT 277.010 4590.300 279.700 4595.900 ;
        RECT 174.860 4582.130 187.830 4588.110 ;
        RECT 272.190 4582.340 274.880 4587.940 ;
        RECT 59.240 4500.610 63.240 4564.050 ;
        RECT 123.990 4558.270 127.760 4563.660 ;
        RECT 65.240 4492.240 69.240 4557.160 ;
        RECT 3223.160 4556.620 3225.900 4562.230 ;
        RECT 3346.570 4556.370 3352.600 4562.440 ;
        RECT 156.680 4550.400 160.490 4555.820 ;
        RECT 3227.900 4548.560 3230.740 4554.250 ;
        RECT 3328.090 4548.370 3334.120 4554.440 ;
        RECT 3399.900 4540.270 3403.670 4545.660 ;
        RECT 3367.170 4532.400 3370.980 4537.820 ;
        RECT 3459.670 4474.240 3463.670 4539.160 ;
        RECT 3465.670 4482.610 3469.670 4546.050 ;
        RECT 3518.490 4487.880 3522.490 4554.710 ;
        RECT 3524.490 4479.230 3528.490 4562.850 ;
        RECT 3223.160 4330.620 3225.900 4336.230 ;
        RECT 3343.040 4330.410 3349.040 4336.410 ;
        RECT 3227.900 4322.560 3230.740 4328.250 ;
        RECT 3327.270 4322.410 3333.270 4328.410 ;
        RECT 3223.160 4105.620 3225.900 4111.230 ;
        RECT 3340.160 4105.410 3346.160 4111.410 ;
        RECT 3227.900 4097.560 3230.740 4103.250 ;
        RECT 3327.430 4097.410 3333.430 4103.410 ;
        RECT 190.890 3961.110 203.850 3967.130 ;
        RECT 277.010 3961.300 279.700 3966.900 ;
        RECT 174.860 3953.130 187.830 3959.110 ;
        RECT 272.190 3953.340 274.880 3958.940 ;
        RECT 59.240 3871.610 63.240 3935.050 ;
        RECT 123.990 3929.270 127.760 3934.660 ;
        RECT 65.240 3863.240 69.240 3928.160 ;
        RECT 156.680 3921.400 160.490 3926.820 ;
        RECT 190.890 3753.110 203.850 3759.130 ;
        RECT 277.010 3753.300 279.700 3758.900 ;
        RECT 174.860 3745.130 187.830 3751.110 ;
        RECT 272.190 3745.340 274.880 3750.940 ;
        RECT 59.240 3655.610 63.240 3719.050 ;
        RECT 123.990 3713.270 127.760 3718.660 ;
        RECT 65.240 3647.240 69.240 3712.160 ;
        RECT 156.680 3705.400 160.490 3710.820 ;
        RECT 3223.160 3664.620 3225.900 3670.230 ;
        RECT 3346.620 3664.370 3352.650 3670.440 ;
        RECT 3227.900 3656.560 3230.740 3662.250 ;
        RECT 3328.140 3656.370 3334.170 3662.440 ;
        RECT 3399.950 3648.270 3403.720 3653.660 ;
        RECT 3367.220 3640.400 3371.030 3645.820 ;
        RECT 3459.720 3582.240 3463.720 3647.160 ;
        RECT 3465.720 3590.610 3469.720 3654.050 ;
        RECT 3518.540 3595.880 3522.540 3662.710 ;
        RECT 3524.540 3587.230 3528.540 3670.850 ;
        RECT 190.890 3529.110 203.850 3535.130 ;
        RECT 277.010 3529.300 279.700 3534.900 ;
        RECT 174.860 3521.130 187.830 3527.110 ;
        RECT 272.190 3521.340 274.880 3526.940 ;
        RECT 59.240 3439.610 63.240 3503.050 ;
        RECT 123.990 3497.270 127.760 3502.660 ;
        RECT 65.240 3431.240 69.240 3496.160 ;
        RECT 156.680 3489.400 160.490 3494.820 ;
        RECT 3223.160 3439.620 3225.900 3445.230 ;
        RECT 3346.620 3439.370 3352.650 3445.440 ;
        RECT 3227.900 3431.560 3230.740 3437.250 ;
        RECT 3328.140 3431.370 3334.170 3437.440 ;
        RECT 3399.950 3423.270 3403.720 3428.660 ;
        RECT 3367.220 3415.400 3371.030 3420.820 ;
        RECT 3459.720 3357.240 3463.720 3422.160 ;
        RECT 3465.720 3365.610 3469.720 3429.050 ;
        RECT 3518.540 3370.880 3522.540 3437.710 ;
        RECT 3524.540 3362.230 3528.540 3445.850 ;
        RECT 190.890 3313.110 203.850 3319.130 ;
        RECT 277.010 3313.300 279.700 3318.900 ;
        RECT 174.860 3305.130 187.830 3311.110 ;
        RECT 272.190 3305.340 274.880 3310.940 ;
        RECT 59.240 3223.610 63.240 3287.050 ;
        RECT 123.990 3281.270 127.760 3286.660 ;
        RECT 65.240 3215.240 69.240 3280.160 ;
        RECT 156.680 3273.400 160.490 3278.820 ;
        RECT 3223.160 3213.620 3225.900 3219.230 ;
        RECT 3346.620 3213.370 3352.650 3219.440 ;
        RECT 3227.900 3205.560 3230.740 3211.250 ;
        RECT 3328.140 3205.370 3334.170 3211.440 ;
        RECT 3399.950 3197.270 3403.720 3202.660 ;
        RECT 3367.220 3189.400 3371.030 3194.820 ;
        RECT 3459.720 3131.240 3463.720 3196.160 ;
        RECT 3465.720 3139.610 3469.720 3203.050 ;
        RECT 3518.540 3144.880 3522.540 3211.710 ;
        RECT 3524.540 3136.230 3528.540 3219.850 ;
        RECT 190.890 3097.110 203.850 3103.130 ;
        RECT 277.010 3097.300 279.700 3102.900 ;
        RECT 174.860 3089.130 187.830 3095.110 ;
        RECT 272.190 3089.340 274.880 3094.940 ;
        RECT 59.240 3007.610 63.240 3071.050 ;
        RECT 123.990 3065.270 127.760 3070.660 ;
        RECT 65.240 2999.240 69.240 3064.160 ;
        RECT 156.680 3057.400 160.490 3062.820 ;
        RECT 3223.160 2988.620 3225.900 2994.230 ;
        RECT 3346.620 2988.370 3352.650 2994.440 ;
        RECT 3328.140 2980.370 3334.170 2986.440 ;
        RECT 3227.900 2974.560 3230.740 2980.250 ;
        RECT 3399.950 2972.270 3403.720 2977.660 ;
        RECT 3367.220 2964.400 3371.030 2969.820 ;
        RECT 3459.720 2906.240 3463.720 2971.160 ;
        RECT 3465.720 2914.610 3469.720 2978.050 ;
        RECT 3518.540 2919.880 3522.540 2986.710 ;
        RECT 3524.540 2911.230 3528.540 2994.850 ;
        RECT 190.890 2886.410 203.850 2892.430 ;
        RECT 277.010 2886.600 279.700 2892.200 ;
        RECT 174.860 2878.430 187.830 2884.410 ;
        RECT 272.190 2878.640 274.880 2884.240 ;
        RECT 59.240 2791.610 63.240 2855.050 ;
        RECT 123.990 2849.270 127.760 2854.660 ;
        RECT 65.240 2783.240 69.240 2848.160 ;
        RECT 156.680 2841.400 160.490 2846.820 ;
        RECT 3223.160 2762.620 3225.900 2768.230 ;
        RECT 3346.620 2762.370 3352.650 2768.440 ;
        RECT 3227.900 2754.560 3230.740 2760.250 ;
        RECT 3328.140 2754.370 3334.170 2760.440 ;
        RECT 3399.950 2746.270 3403.720 2751.660 ;
        RECT 3367.220 2738.400 3371.030 2743.820 ;
        RECT 3459.720 2680.240 3463.720 2745.160 ;
        RECT 3465.720 2688.610 3469.720 2752.050 ;
        RECT 3518.540 2693.880 3522.540 2760.710 ;
        RECT 3524.540 2685.230 3528.540 2768.850 ;
        RECT 190.890 2665.110 203.850 2671.130 ;
        RECT 277.010 2665.300 279.700 2670.900 ;
        RECT 174.860 2657.130 187.830 2663.110 ;
        RECT 272.190 2657.340 274.880 2662.940 ;
        RECT 59.240 2575.610 63.240 2639.050 ;
        RECT 123.990 2633.270 127.760 2638.660 ;
        RECT 65.240 2567.240 69.240 2632.160 ;
        RECT 156.680 2625.400 160.490 2630.820 ;
        RECT 3223.160 2537.620 3225.900 2543.230 ;
        RECT 3346.620 2537.370 3352.650 2543.440 ;
        RECT 3227.900 2529.560 3230.740 2535.250 ;
        RECT 3328.140 2529.370 3334.170 2535.440 ;
        RECT 3399.950 2521.270 3403.720 2526.660 ;
        RECT 3367.220 2513.400 3371.030 2518.820 ;
        RECT 3459.720 2455.240 3463.720 2520.160 ;
        RECT 3465.720 2463.610 3469.720 2527.050 ;
        RECT 3518.540 2468.880 3522.540 2535.710 ;
        RECT 3524.540 2460.230 3528.540 2543.850 ;
        RECT 3223.160 2320.620 3225.900 2326.230 ;
        RECT 3346.620 2317.370 3352.650 2323.440 ;
        RECT 3227.900 2309.560 3230.740 2315.250 ;
        RECT 3328.140 2309.370 3334.170 2315.440 ;
        RECT 3399.950 2301.270 3403.720 2306.660 ;
        RECT 3367.220 2293.400 3371.030 2298.820 ;
        RECT 3459.720 2235.240 3463.720 2300.160 ;
        RECT 3465.720 2243.610 3469.720 2307.050 ;
        RECT 3518.540 2248.880 3522.540 2315.710 ;
        RECT 3524.540 2240.230 3528.540 2323.850 ;
        RECT 190.890 2027.110 203.850 2033.130 ;
        RECT 277.010 2027.300 279.700 2032.900 ;
        RECT 174.860 2019.130 187.830 2025.110 ;
        RECT 272.190 2019.340 274.880 2024.940 ;
        RECT 59.240 1937.610 63.240 2001.050 ;
        RECT 123.990 1995.270 127.760 2000.660 ;
        RECT 65.240 1929.240 69.240 1994.160 ;
        RECT 156.680 1987.400 160.490 1992.820 ;
        RECT 3223.160 1876.620 3225.900 1882.230 ;
        RECT 3346.620 1876.370 3352.650 1882.440 ;
        RECT 3227.900 1868.560 3230.740 1874.250 ;
        RECT 3328.140 1868.370 3334.170 1874.440 ;
        RECT 3399.950 1860.270 3403.720 1865.660 ;
        RECT 3367.220 1852.400 3371.030 1857.820 ;
        RECT 190.890 1811.110 203.850 1817.130 ;
        RECT 277.010 1811.300 279.700 1816.900 ;
        RECT 174.860 1803.130 187.830 1809.110 ;
        RECT 272.190 1803.340 274.880 1808.940 ;
        RECT 3459.720 1794.240 3463.720 1859.160 ;
        RECT 3465.720 1802.610 3469.720 1866.050 ;
        RECT 3518.540 1807.880 3522.540 1874.710 ;
        RECT 3524.540 1799.230 3528.540 1882.850 ;
        RECT 59.240 1721.610 63.240 1785.050 ;
        RECT 123.990 1779.270 127.760 1784.660 ;
        RECT 65.240 1713.240 69.240 1778.160 ;
        RECT 156.680 1771.400 160.490 1776.820 ;
        RECT 3223.160 1657.620 3225.900 1663.230 ;
        RECT 3346.620 1650.370 3352.650 1656.440 ;
        RECT 3227.900 1642.560 3230.740 1648.250 ;
        RECT 3328.140 1642.370 3334.170 1648.440 ;
        RECT 3399.950 1634.270 3403.720 1639.660 ;
        RECT 3367.220 1626.400 3371.030 1631.820 ;
        RECT 190.890 1600.110 203.850 1606.130 ;
        RECT 277.010 1600.300 279.700 1605.900 ;
        RECT 174.860 1592.130 187.830 1598.110 ;
        RECT 272.190 1592.340 274.880 1597.940 ;
        RECT 59.240 1505.610 63.240 1569.050 ;
        RECT 123.990 1563.270 127.760 1568.660 ;
        RECT 3459.720 1568.240 3463.720 1633.160 ;
        RECT 3465.720 1576.610 3469.720 1640.050 ;
        RECT 3518.540 1581.880 3522.540 1648.710 ;
        RECT 3524.540 1573.230 3528.540 1656.850 ;
        RECT 65.240 1497.240 69.240 1562.160 ;
        RECT 156.680 1555.400 160.490 1560.820 ;
        RECT 3223.160 1425.620 3225.900 1431.230 ;
        RECT 3346.620 1425.370 3352.650 1431.440 ;
        RECT 3227.900 1417.560 3230.740 1423.250 ;
        RECT 3328.140 1417.370 3334.170 1423.440 ;
        RECT 3399.950 1409.270 3403.720 1414.660 ;
        RECT 3367.220 1401.400 3371.030 1406.820 ;
        RECT 190.890 1379.110 203.850 1385.130 ;
        RECT 277.010 1379.300 279.700 1384.900 ;
        RECT 174.860 1371.130 187.830 1377.110 ;
        RECT 272.190 1371.340 274.880 1376.940 ;
        RECT 59.240 1289.610 63.240 1353.050 ;
        RECT 123.990 1347.270 127.760 1352.660 ;
        RECT 65.240 1281.240 69.240 1346.160 ;
        RECT 156.680 1339.400 160.490 1344.820 ;
        RECT 3459.720 1343.240 3463.720 1408.160 ;
        RECT 3465.720 1351.610 3469.720 1415.050 ;
        RECT 3518.540 1356.880 3522.540 1423.710 ;
        RECT 3524.540 1348.230 3528.540 1431.850 ;
        RECT 3264.300 1219.370 3353.030 1222.530 ;
        RECT 190.865 1212.920 203.900 1216.920 ;
        RECT 3264.170 1214.580 3337.140 1217.780 ;
        RECT 190.865 1209.790 252.050 1212.920 ;
        RECT 3323.980 1210.580 3337.140 1214.580 ;
        RECT 3339.970 1214.370 3353.030 1219.370 ;
        RECT 183.620 1205.030 252.130 1208.160 ;
        RECT 183.620 1176.890 187.940 1205.030 ;
        RECT 3346.620 1200.370 3352.650 1206.440 ;
        RECT 3328.140 1192.370 3334.170 1198.440 ;
        RECT 3399.950 1184.270 3403.720 1189.660 ;
        RECT 3367.220 1176.400 3371.030 1181.820 ;
        RECT 59.240 1073.610 63.240 1137.050 ;
        RECT 123.990 1131.270 127.760 1136.660 ;
        RECT 65.240 1065.240 69.240 1130.160 ;
        RECT 156.680 1123.400 160.490 1128.820 ;
        RECT 3459.720 1118.240 3463.720 1183.160 ;
        RECT 3465.720 1126.610 3469.720 1190.050 ;
        RECT 3518.540 1131.880 3522.540 1198.710 ;
        RECT 3524.540 1123.230 3528.540 1206.850 ;
        RECT 3346.620 974.370 3352.650 980.440 ;
        RECT 3328.140 966.370 3334.170 972.440 ;
        RECT 3399.950 958.270 3403.720 963.660 ;
        RECT 3367.220 950.400 3371.030 955.820 ;
        RECT 59.240 857.610 63.240 921.050 ;
        RECT 123.990 915.270 127.760 920.660 ;
        RECT 65.240 849.240 69.240 914.160 ;
        RECT 156.680 907.400 160.490 912.820 ;
        RECT 3459.720 892.240 3463.720 957.160 ;
        RECT 3465.720 900.610 3469.720 964.050 ;
        RECT 3518.540 905.880 3522.540 972.710 ;
        RECT 3524.540 897.230 3528.540 980.850 ;
        RECT 3346.620 749.370 3352.650 755.440 ;
        RECT 3328.140 741.370 3334.170 747.440 ;
        RECT 3399.950 733.270 3403.720 738.660 ;
        RECT 3367.220 725.400 3371.030 730.820 ;
        RECT 3459.720 667.240 3463.720 732.160 ;
        RECT 3465.720 675.610 3469.720 739.050 ;
        RECT 3518.540 680.880 3522.540 747.710 ;
        RECT 3524.540 672.230 3528.540 755.850 ;
        RECT 3346.620 523.370 3352.650 529.440 ;
        RECT 3328.140 515.370 3334.170 521.440 ;
        RECT 3399.950 507.270 3403.720 512.660 ;
        RECT 3367.220 499.400 3371.030 504.820 ;
        RECT 3459.720 441.240 3463.720 506.160 ;
        RECT 3465.720 449.610 3469.720 513.050 ;
        RECT 3518.540 454.880 3522.540 521.710 ;
        RECT 3524.540 446.230 3528.540 529.850 ;
        RECT 3179.570 68.635 3220.900 70.635 ;
        RECT 687.090 34.310 687.990 66.980 ;
        RECT 693.590 36.290 694.490 67.200 ;
        RECT 3179.570 41.320 3188.480 68.635 ;
        RECT 3237.050 42.940 3254.450 65.770 ;
        RECT 693.590 35.390 722.470 36.290 ;
        RECT 687.090 33.410 714.590 34.310 ;
        RECT 718.050 6.330 722.070 10.480 ;
        RECT 710.380 0.290 714.400 4.440 ;
        RECT 3180.020 0.440 3188.060 4.300 ;
      LAYER via4 ;
        RECT 470.430 4927.960 471.610 4929.140 ;
        RECT 487.340 4927.970 488.520 4929.150 ;
        RECT 504.250 4927.940 505.430 4929.120 ;
        RECT 528.285 4927.960 529.465 4929.140 ;
        RECT 470.430 4926.360 471.610 4927.540 ;
        RECT 487.340 4926.370 488.520 4927.550 ;
        RECT 504.250 4926.340 505.430 4927.520 ;
        RECT 528.285 4926.360 529.465 4927.540 ;
        RECT 727.430 4927.960 728.610 4929.140 ;
        RECT 744.340 4927.970 745.520 4929.150 ;
        RECT 761.250 4927.940 762.430 4929.120 ;
        RECT 785.285 4927.960 786.465 4929.140 ;
        RECT 727.430 4926.360 728.610 4927.540 ;
        RECT 744.340 4926.370 745.520 4927.550 ;
        RECT 761.250 4926.340 762.430 4927.520 ;
        RECT 785.285 4926.360 786.465 4927.540 ;
        RECT 984.430 4927.960 985.610 4929.140 ;
        RECT 1001.340 4927.970 1002.520 4929.150 ;
        RECT 1018.250 4927.940 1019.430 4929.120 ;
        RECT 1042.285 4927.960 1043.465 4929.140 ;
        RECT 984.430 4926.360 985.610 4927.540 ;
        RECT 1001.340 4926.370 1002.520 4927.550 ;
        RECT 1018.250 4926.340 1019.430 4927.520 ;
        RECT 1042.285 4926.360 1043.465 4927.540 ;
        RECT 1241.430 4927.960 1242.610 4929.140 ;
        RECT 1258.340 4927.970 1259.520 4929.150 ;
        RECT 1275.250 4927.940 1276.430 4929.120 ;
        RECT 1299.285 4927.960 1300.465 4929.140 ;
        RECT 1241.430 4926.360 1242.610 4927.540 ;
        RECT 1258.340 4926.370 1259.520 4927.550 ;
        RECT 1275.250 4926.340 1276.430 4927.520 ;
        RECT 1299.285 4926.360 1300.465 4927.540 ;
        RECT 1499.430 4927.960 1500.610 4929.140 ;
        RECT 1516.340 4927.970 1517.520 4929.150 ;
        RECT 1533.250 4927.940 1534.430 4929.120 ;
        RECT 1557.285 4927.960 1558.465 4929.140 ;
        RECT 1499.430 4926.360 1500.610 4927.540 ;
        RECT 1516.340 4926.370 1517.520 4927.550 ;
        RECT 1533.250 4926.340 1534.430 4927.520 ;
        RECT 1557.285 4926.360 1558.465 4927.540 ;
        RECT 1751.430 4927.960 1752.610 4929.140 ;
        RECT 1768.340 4927.970 1769.520 4929.150 ;
        RECT 1785.250 4927.940 1786.430 4929.120 ;
        RECT 1809.285 4927.960 1810.465 4929.140 ;
        RECT 1751.430 4926.360 1752.610 4927.540 ;
        RECT 1768.340 4926.370 1769.520 4927.550 ;
        RECT 1785.250 4926.340 1786.430 4927.520 ;
        RECT 1809.285 4926.360 1810.465 4927.540 ;
        RECT 2088.430 4927.960 2089.610 4929.140 ;
        RECT 2105.340 4927.970 2106.520 4929.150 ;
        RECT 2122.250 4927.940 2123.430 4929.120 ;
        RECT 2146.285 4927.960 2147.465 4929.140 ;
        RECT 2088.430 4926.360 2089.610 4927.540 ;
        RECT 2105.340 4926.370 2106.520 4927.550 ;
        RECT 2122.250 4926.340 2123.430 4927.520 ;
        RECT 2146.285 4926.360 2147.465 4927.540 ;
        RECT 2473.430 4927.960 2474.610 4929.140 ;
        RECT 2490.340 4927.970 2491.520 4929.150 ;
        RECT 2507.250 4927.940 2508.430 4929.120 ;
        RECT 2531.285 4927.960 2532.465 4929.140 ;
        RECT 2473.430 4926.360 2474.610 4927.540 ;
        RECT 2490.340 4926.370 2491.520 4927.550 ;
        RECT 2507.250 4926.340 2508.430 4927.520 ;
        RECT 2531.285 4926.360 2532.465 4927.540 ;
        RECT 2730.430 4927.960 2731.610 4929.140 ;
        RECT 2747.340 4927.970 2748.520 4929.150 ;
        RECT 2764.250 4927.940 2765.430 4929.120 ;
        RECT 2788.285 4927.960 2789.465 4929.140 ;
        RECT 2730.430 4926.360 2731.610 4927.540 ;
        RECT 2747.340 4926.370 2748.520 4927.550 ;
        RECT 2764.250 4926.340 2765.430 4927.520 ;
        RECT 2788.285 4926.360 2789.465 4927.540 ;
        RECT 462.000 4921.940 463.180 4923.120 ;
        RECT 478.900 4921.940 480.080 4923.120 ;
        RECT 495.800 4921.960 496.980 4923.140 ;
        RECT 524.765 4921.960 525.945 4923.140 ;
        RECT 462.000 4920.340 463.180 4921.520 ;
        RECT 478.900 4920.340 480.080 4921.520 ;
        RECT 495.800 4920.360 496.980 4921.540 ;
        RECT 524.765 4920.360 525.945 4921.540 ;
        RECT 719.000 4921.940 720.180 4923.120 ;
        RECT 735.900 4921.940 737.080 4923.120 ;
        RECT 752.800 4921.960 753.980 4923.140 ;
        RECT 781.765 4921.960 782.945 4923.140 ;
        RECT 719.000 4920.340 720.180 4921.520 ;
        RECT 735.900 4920.340 737.080 4921.520 ;
        RECT 752.800 4920.360 753.980 4921.540 ;
        RECT 781.765 4920.360 782.945 4921.540 ;
        RECT 976.000 4921.940 977.180 4923.120 ;
        RECT 992.900 4921.940 994.080 4923.120 ;
        RECT 1009.800 4921.960 1010.980 4923.140 ;
        RECT 1038.765 4921.960 1039.945 4923.140 ;
        RECT 976.000 4920.340 977.180 4921.520 ;
        RECT 992.900 4920.340 994.080 4921.520 ;
        RECT 1009.800 4920.360 1010.980 4921.540 ;
        RECT 1038.765 4920.360 1039.945 4921.540 ;
        RECT 1233.000 4921.940 1234.180 4923.120 ;
        RECT 1249.900 4921.940 1251.080 4923.120 ;
        RECT 1266.800 4921.960 1267.980 4923.140 ;
        RECT 1295.765 4921.960 1296.945 4923.140 ;
        RECT 1233.000 4920.340 1234.180 4921.520 ;
        RECT 1249.900 4920.340 1251.080 4921.520 ;
        RECT 1266.800 4920.360 1267.980 4921.540 ;
        RECT 1295.765 4920.360 1296.945 4921.540 ;
        RECT 1491.000 4921.940 1492.180 4923.120 ;
        RECT 1507.900 4921.940 1509.080 4923.120 ;
        RECT 1524.800 4921.960 1525.980 4923.140 ;
        RECT 1553.765 4921.960 1554.945 4923.140 ;
        RECT 1491.000 4920.340 1492.180 4921.520 ;
        RECT 1507.900 4920.340 1509.080 4921.520 ;
        RECT 1524.800 4920.360 1525.980 4921.540 ;
        RECT 1553.765 4920.360 1554.945 4921.540 ;
        RECT 1743.000 4921.940 1744.180 4923.120 ;
        RECT 1759.900 4921.940 1761.080 4923.120 ;
        RECT 1776.800 4921.960 1777.980 4923.140 ;
        RECT 1805.765 4921.960 1806.945 4923.140 ;
        RECT 1743.000 4920.340 1744.180 4921.520 ;
        RECT 1759.900 4920.340 1761.080 4921.520 ;
        RECT 1776.800 4920.360 1777.980 4921.540 ;
        RECT 1805.765 4920.360 1806.945 4921.540 ;
        RECT 2080.000 4921.940 2081.180 4923.120 ;
        RECT 2096.900 4921.940 2098.080 4923.120 ;
        RECT 2113.800 4921.960 2114.980 4923.140 ;
        RECT 2142.765 4921.960 2143.945 4923.140 ;
        RECT 2080.000 4920.340 2081.180 4921.520 ;
        RECT 2096.900 4920.340 2098.080 4921.520 ;
        RECT 2113.800 4920.360 2114.980 4921.540 ;
        RECT 2142.765 4920.360 2143.945 4921.540 ;
        RECT 2465.000 4921.940 2466.180 4923.120 ;
        RECT 2481.900 4921.940 2483.080 4923.120 ;
        RECT 2498.800 4921.960 2499.980 4923.140 ;
        RECT 2527.765 4921.960 2528.945 4923.140 ;
        RECT 2465.000 4920.340 2466.180 4921.520 ;
        RECT 2481.900 4920.340 2483.080 4921.520 ;
        RECT 2498.800 4920.360 2499.980 4921.540 ;
        RECT 2527.765 4920.360 2528.945 4921.540 ;
        RECT 2722.000 4921.940 2723.180 4923.120 ;
        RECT 2738.900 4921.940 2740.080 4923.120 ;
        RECT 2755.800 4921.960 2756.980 4923.140 ;
        RECT 2784.765 4921.960 2785.945 4923.140 ;
        RECT 2722.000 4920.340 2723.180 4921.520 ;
        RECT 2738.900 4920.340 2740.080 4921.520 ;
        RECT 2755.800 4920.360 2756.980 4921.540 ;
        RECT 2784.765 4920.360 2785.945 4921.540 ;
        RECT 175.220 4759.925 187.600 4762.705 ;
        RECT 248.955 4760.715 250.135 4761.895 ;
        RECT 250.555 4760.715 251.735 4761.895 ;
        RECT 191.235 4755.150 203.615 4757.930 ;
        RECT 249.030 4755.095 251.810 4757.875 ;
        RECT 3261.845 4751.100 3263.025 4752.280 ;
        RECT 3263.445 4751.100 3264.625 4752.280 ;
        RECT 3265.045 4751.100 3266.225 4752.280 ;
        RECT 3266.645 4751.100 3267.825 4752.280 ;
        RECT 3268.245 4751.100 3269.425 4752.280 ;
        RECT 3269.845 4751.100 3271.025 4752.280 ;
        RECT 3271.445 4751.100 3272.625 4752.280 ;
        RECT 3273.045 4751.100 3274.225 4752.280 ;
        RECT 3274.645 4751.100 3275.825 4752.280 ;
        RECT 3276.245 4751.100 3277.425 4752.280 ;
        RECT 3277.845 4751.100 3279.025 4752.280 ;
        RECT 3279.445 4751.100 3280.625 4752.280 ;
        RECT 3281.045 4751.100 3282.225 4752.280 ;
        RECT 3282.645 4751.100 3283.825 4752.280 ;
        RECT 3284.245 4751.100 3285.425 4752.280 ;
        RECT 3324.305 4750.325 3336.685 4753.105 ;
        RECT 3261.755 4746.320 3262.935 4747.500 ;
        RECT 3263.355 4746.320 3264.535 4747.500 ;
        RECT 3264.955 4746.320 3266.135 4747.500 ;
        RECT 3266.555 4746.320 3267.735 4747.500 ;
        RECT 3268.155 4746.320 3269.335 4747.500 ;
        RECT 3269.755 4746.320 3270.935 4747.500 ;
        RECT 3271.355 4746.320 3272.535 4747.500 ;
        RECT 3272.955 4746.320 3274.135 4747.500 ;
        RECT 3274.555 4746.320 3275.735 4747.500 ;
        RECT 3276.155 4746.320 3277.335 4747.500 ;
        RECT 3277.755 4746.320 3278.935 4747.500 ;
        RECT 3279.355 4746.320 3280.535 4747.500 ;
        RECT 3280.955 4746.320 3282.135 4747.500 ;
        RECT 3282.555 4746.320 3283.735 4747.500 ;
        RECT 3284.155 4746.320 3285.335 4747.500 ;
        RECT 3340.295 4745.515 3352.675 4748.295 ;
        RECT 192.030 4590.825 202.810 4595.205 ;
        RECT 175.980 4582.915 186.760 4587.295 ;
        RECT 59.840 4558.895 61.020 4560.075 ;
        RECT 61.440 4558.895 62.620 4560.075 ;
        RECT 59.860 4534.860 61.040 4536.040 ;
        RECT 61.460 4534.860 62.640 4536.040 ;
        RECT 59.830 4517.950 61.010 4519.130 ;
        RECT 61.430 4517.950 62.610 4519.130 ;
        RECT 59.840 4501.040 61.020 4502.220 ;
        RECT 61.440 4501.040 62.620 4502.220 ;
        RECT 3347.395 4557.295 3351.775 4561.675 ;
        RECT 65.840 4555.375 67.020 4556.555 ;
        RECT 67.440 4555.375 68.620 4556.555 ;
        RECT 3328.865 4549.205 3333.245 4553.585 ;
        RECT 3466.290 4540.895 3467.470 4542.075 ;
        RECT 3467.890 4540.895 3469.070 4542.075 ;
        RECT 3460.290 4537.375 3461.470 4538.555 ;
        RECT 3461.890 4537.375 3463.070 4538.555 ;
        RECT 65.840 4526.410 67.020 4527.590 ;
        RECT 67.440 4526.410 68.620 4527.590 ;
        RECT 65.860 4509.510 67.040 4510.690 ;
        RECT 67.460 4509.510 68.640 4510.690 ;
        RECT 65.860 4492.610 67.040 4493.790 ;
        RECT 67.460 4492.610 68.640 4493.790 ;
        RECT 3460.290 4508.410 3461.470 4509.590 ;
        RECT 3461.890 4508.410 3463.070 4509.590 ;
        RECT 3460.270 4491.510 3461.450 4492.690 ;
        RECT 3461.870 4491.510 3463.050 4492.690 ;
        RECT 3466.270 4516.860 3467.450 4518.040 ;
        RECT 3467.870 4516.860 3469.050 4518.040 ;
        RECT 3466.300 4499.950 3467.480 4501.130 ;
        RECT 3467.900 4499.950 3469.080 4501.130 ;
        RECT 3519.095 4522.085 3520.275 4523.265 ;
        RECT 3520.695 4522.085 3521.875 4523.265 ;
        RECT 3519.105 4505.165 3520.285 4506.345 ;
        RECT 3520.705 4505.165 3521.885 4506.345 ;
        RECT 3519.115 4488.295 3520.295 4489.475 ;
        RECT 3520.715 4488.295 3521.895 4489.475 ;
        RECT 3525.105 4513.605 3526.285 4514.785 ;
        RECT 3526.705 4513.605 3527.885 4514.785 ;
        RECT 3525.075 4496.805 3526.255 4497.985 ;
        RECT 3526.675 4496.805 3527.855 4497.985 ;
        RECT 3466.290 4483.040 3467.470 4484.220 ;
        RECT 3467.890 4483.040 3469.070 4484.220 ;
        RECT 3525.085 4479.855 3526.265 4481.035 ;
        RECT 3526.685 4479.855 3527.865 4481.035 ;
        RECT 3460.270 4474.610 3461.450 4475.790 ;
        RECT 3461.870 4474.610 3463.050 4475.790 ;
        RECT 3343.885 4331.275 3348.265 4335.655 ;
        RECT 3328.105 4323.235 3332.485 4327.615 ;
        RECT 3340.940 4106.230 3345.320 4110.610 ;
        RECT 3328.220 4098.220 3332.600 4102.600 ;
        RECT 192.030 3961.825 202.810 3966.205 ;
        RECT 175.980 3953.915 186.760 3958.295 ;
        RECT 59.840 3929.895 61.020 3931.075 ;
        RECT 61.440 3929.895 62.620 3931.075 ;
        RECT 59.860 3905.860 61.040 3907.040 ;
        RECT 61.460 3905.860 62.640 3907.040 ;
        RECT 59.830 3888.950 61.010 3890.130 ;
        RECT 61.430 3888.950 62.610 3890.130 ;
        RECT 59.840 3872.040 61.020 3873.220 ;
        RECT 61.440 3872.040 62.620 3873.220 ;
        RECT 65.840 3926.375 67.020 3927.555 ;
        RECT 67.440 3926.375 68.620 3927.555 ;
        RECT 65.840 3897.410 67.020 3898.590 ;
        RECT 67.440 3897.410 68.620 3898.590 ;
        RECT 65.860 3880.510 67.040 3881.690 ;
        RECT 67.460 3880.510 68.640 3881.690 ;
        RECT 65.860 3863.610 67.040 3864.790 ;
        RECT 67.460 3863.610 68.640 3864.790 ;
        RECT 192.030 3753.825 202.810 3758.205 ;
        RECT 175.980 3745.915 186.760 3750.295 ;
        RECT 59.840 3713.895 61.020 3715.075 ;
        RECT 61.440 3713.895 62.620 3715.075 ;
        RECT 59.860 3689.860 61.040 3691.040 ;
        RECT 61.460 3689.860 62.640 3691.040 ;
        RECT 59.830 3672.950 61.010 3674.130 ;
        RECT 61.430 3672.950 62.610 3674.130 ;
        RECT 59.840 3656.040 61.020 3657.220 ;
        RECT 61.440 3656.040 62.620 3657.220 ;
        RECT 65.840 3710.375 67.020 3711.555 ;
        RECT 67.440 3710.375 68.620 3711.555 ;
        RECT 65.840 3681.410 67.020 3682.590 ;
        RECT 67.440 3681.410 68.620 3682.590 ;
        RECT 65.860 3664.510 67.040 3665.690 ;
        RECT 67.460 3664.510 68.640 3665.690 ;
        RECT 3347.445 3665.295 3351.825 3669.675 ;
        RECT 3328.915 3657.205 3333.295 3661.585 ;
        RECT 65.860 3647.610 67.040 3648.790 ;
        RECT 67.460 3647.610 68.640 3648.790 ;
        RECT 3466.340 3648.895 3467.520 3650.075 ;
        RECT 3467.940 3648.895 3469.120 3650.075 ;
        RECT 3460.340 3645.375 3461.520 3646.555 ;
        RECT 3461.940 3645.375 3463.120 3646.555 ;
        RECT 3460.340 3616.410 3461.520 3617.590 ;
        RECT 3461.940 3616.410 3463.120 3617.590 ;
        RECT 3460.320 3599.510 3461.500 3600.690 ;
        RECT 3461.920 3599.510 3463.100 3600.690 ;
        RECT 3466.320 3624.860 3467.500 3626.040 ;
        RECT 3467.920 3624.860 3469.100 3626.040 ;
        RECT 3466.350 3607.950 3467.530 3609.130 ;
        RECT 3467.950 3607.950 3469.130 3609.130 ;
        RECT 3519.145 3630.085 3520.325 3631.265 ;
        RECT 3520.745 3630.085 3521.925 3631.265 ;
        RECT 3519.155 3613.165 3520.335 3614.345 ;
        RECT 3520.755 3613.165 3521.935 3614.345 ;
        RECT 3519.165 3596.295 3520.345 3597.475 ;
        RECT 3520.765 3596.295 3521.945 3597.475 ;
        RECT 3525.155 3621.605 3526.335 3622.785 ;
        RECT 3526.755 3621.605 3527.935 3622.785 ;
        RECT 3525.125 3604.805 3526.305 3605.985 ;
        RECT 3526.725 3604.805 3527.905 3605.985 ;
        RECT 3466.340 3591.040 3467.520 3592.220 ;
        RECT 3467.940 3591.040 3469.120 3592.220 ;
        RECT 3525.135 3587.855 3526.315 3589.035 ;
        RECT 3526.735 3587.855 3527.915 3589.035 ;
        RECT 3460.320 3582.610 3461.500 3583.790 ;
        RECT 3461.920 3582.610 3463.100 3583.790 ;
        RECT 192.030 3529.825 202.810 3534.205 ;
        RECT 175.980 3521.915 186.760 3526.295 ;
        RECT 59.840 3497.895 61.020 3499.075 ;
        RECT 61.440 3497.895 62.620 3499.075 ;
        RECT 59.860 3473.860 61.040 3475.040 ;
        RECT 61.460 3473.860 62.640 3475.040 ;
        RECT 59.830 3456.950 61.010 3458.130 ;
        RECT 61.430 3456.950 62.610 3458.130 ;
        RECT 59.840 3440.040 61.020 3441.220 ;
        RECT 61.440 3440.040 62.620 3441.220 ;
        RECT 65.840 3494.375 67.020 3495.555 ;
        RECT 67.440 3494.375 68.620 3495.555 ;
        RECT 65.840 3465.410 67.020 3466.590 ;
        RECT 67.440 3465.410 68.620 3466.590 ;
        RECT 65.860 3448.510 67.040 3449.690 ;
        RECT 67.460 3448.510 68.640 3449.690 ;
        RECT 3347.445 3440.295 3351.825 3444.675 ;
        RECT 65.860 3431.610 67.040 3432.790 ;
        RECT 67.460 3431.610 68.640 3432.790 ;
        RECT 3328.915 3432.205 3333.295 3436.585 ;
        RECT 3466.340 3423.895 3467.520 3425.075 ;
        RECT 3467.940 3423.895 3469.120 3425.075 ;
        RECT 3460.340 3420.375 3461.520 3421.555 ;
        RECT 3461.940 3420.375 3463.120 3421.555 ;
        RECT 3460.340 3391.410 3461.520 3392.590 ;
        RECT 3461.940 3391.410 3463.120 3392.590 ;
        RECT 3460.320 3374.510 3461.500 3375.690 ;
        RECT 3461.920 3374.510 3463.100 3375.690 ;
        RECT 3466.320 3399.860 3467.500 3401.040 ;
        RECT 3467.920 3399.860 3469.100 3401.040 ;
        RECT 3466.350 3382.950 3467.530 3384.130 ;
        RECT 3467.950 3382.950 3469.130 3384.130 ;
        RECT 3519.145 3405.085 3520.325 3406.265 ;
        RECT 3520.745 3405.085 3521.925 3406.265 ;
        RECT 3519.155 3388.165 3520.335 3389.345 ;
        RECT 3520.755 3388.165 3521.935 3389.345 ;
        RECT 3519.165 3371.295 3520.345 3372.475 ;
        RECT 3520.765 3371.295 3521.945 3372.475 ;
        RECT 3525.155 3396.605 3526.335 3397.785 ;
        RECT 3526.755 3396.605 3527.935 3397.785 ;
        RECT 3525.125 3379.805 3526.305 3380.985 ;
        RECT 3526.725 3379.805 3527.905 3380.985 ;
        RECT 3466.340 3366.040 3467.520 3367.220 ;
        RECT 3467.940 3366.040 3469.120 3367.220 ;
        RECT 3525.135 3362.855 3526.315 3364.035 ;
        RECT 3526.735 3362.855 3527.915 3364.035 ;
        RECT 3460.320 3357.610 3461.500 3358.790 ;
        RECT 3461.920 3357.610 3463.100 3358.790 ;
        RECT 192.030 3313.825 202.810 3318.205 ;
        RECT 175.980 3305.915 186.760 3310.295 ;
        RECT 59.840 3281.895 61.020 3283.075 ;
        RECT 61.440 3281.895 62.620 3283.075 ;
        RECT 59.860 3257.860 61.040 3259.040 ;
        RECT 61.460 3257.860 62.640 3259.040 ;
        RECT 59.830 3240.950 61.010 3242.130 ;
        RECT 61.430 3240.950 62.610 3242.130 ;
        RECT 59.840 3224.040 61.020 3225.220 ;
        RECT 61.440 3224.040 62.620 3225.220 ;
        RECT 65.840 3278.375 67.020 3279.555 ;
        RECT 67.440 3278.375 68.620 3279.555 ;
        RECT 65.840 3249.410 67.020 3250.590 ;
        RECT 67.440 3249.410 68.620 3250.590 ;
        RECT 65.860 3232.510 67.040 3233.690 ;
        RECT 67.460 3232.510 68.640 3233.690 ;
        RECT 65.860 3215.610 67.040 3216.790 ;
        RECT 67.460 3215.610 68.640 3216.790 ;
        RECT 3347.445 3214.295 3351.825 3218.675 ;
        RECT 3328.915 3206.205 3333.295 3210.585 ;
        RECT 3466.340 3197.895 3467.520 3199.075 ;
        RECT 3467.940 3197.895 3469.120 3199.075 ;
        RECT 3460.340 3194.375 3461.520 3195.555 ;
        RECT 3461.940 3194.375 3463.120 3195.555 ;
        RECT 3460.340 3165.410 3461.520 3166.590 ;
        RECT 3461.940 3165.410 3463.120 3166.590 ;
        RECT 3460.320 3148.510 3461.500 3149.690 ;
        RECT 3461.920 3148.510 3463.100 3149.690 ;
        RECT 3466.320 3173.860 3467.500 3175.040 ;
        RECT 3467.920 3173.860 3469.100 3175.040 ;
        RECT 3466.350 3156.950 3467.530 3158.130 ;
        RECT 3467.950 3156.950 3469.130 3158.130 ;
        RECT 3519.145 3179.085 3520.325 3180.265 ;
        RECT 3520.745 3179.085 3521.925 3180.265 ;
        RECT 3519.155 3162.165 3520.335 3163.345 ;
        RECT 3520.755 3162.165 3521.935 3163.345 ;
        RECT 3519.165 3145.295 3520.345 3146.475 ;
        RECT 3520.765 3145.295 3521.945 3146.475 ;
        RECT 3525.155 3170.605 3526.335 3171.785 ;
        RECT 3526.755 3170.605 3527.935 3171.785 ;
        RECT 3525.125 3153.805 3526.305 3154.985 ;
        RECT 3526.725 3153.805 3527.905 3154.985 ;
        RECT 3466.340 3140.040 3467.520 3141.220 ;
        RECT 3467.940 3140.040 3469.120 3141.220 ;
        RECT 3525.135 3136.855 3526.315 3138.035 ;
        RECT 3526.735 3136.855 3527.915 3138.035 ;
        RECT 3460.320 3131.610 3461.500 3132.790 ;
        RECT 3461.920 3131.610 3463.100 3132.790 ;
        RECT 192.030 3097.825 202.810 3102.205 ;
        RECT 175.980 3089.915 186.760 3094.295 ;
        RECT 59.840 3065.895 61.020 3067.075 ;
        RECT 61.440 3065.895 62.620 3067.075 ;
        RECT 59.860 3041.860 61.040 3043.040 ;
        RECT 61.460 3041.860 62.640 3043.040 ;
        RECT 59.830 3024.950 61.010 3026.130 ;
        RECT 61.430 3024.950 62.610 3026.130 ;
        RECT 59.840 3008.040 61.020 3009.220 ;
        RECT 61.440 3008.040 62.620 3009.220 ;
        RECT 65.840 3062.375 67.020 3063.555 ;
        RECT 67.440 3062.375 68.620 3063.555 ;
        RECT 65.840 3033.410 67.020 3034.590 ;
        RECT 67.440 3033.410 68.620 3034.590 ;
        RECT 65.860 3016.510 67.040 3017.690 ;
        RECT 67.460 3016.510 68.640 3017.690 ;
        RECT 65.860 2999.610 67.040 3000.790 ;
        RECT 67.460 2999.610 68.640 3000.790 ;
        RECT 3347.445 2989.295 3351.825 2993.675 ;
        RECT 3328.915 2981.205 3333.295 2985.585 ;
        RECT 3466.340 2972.895 3467.520 2974.075 ;
        RECT 3467.940 2972.895 3469.120 2974.075 ;
        RECT 3460.340 2969.375 3461.520 2970.555 ;
        RECT 3461.940 2969.375 3463.120 2970.555 ;
        RECT 3460.340 2940.410 3461.520 2941.590 ;
        RECT 3461.940 2940.410 3463.120 2941.590 ;
        RECT 3460.320 2923.510 3461.500 2924.690 ;
        RECT 3461.920 2923.510 3463.100 2924.690 ;
        RECT 3466.320 2948.860 3467.500 2950.040 ;
        RECT 3467.920 2948.860 3469.100 2950.040 ;
        RECT 3466.350 2931.950 3467.530 2933.130 ;
        RECT 3467.950 2931.950 3469.130 2933.130 ;
        RECT 3519.145 2954.085 3520.325 2955.265 ;
        RECT 3520.745 2954.085 3521.925 2955.265 ;
        RECT 3519.155 2937.165 3520.335 2938.345 ;
        RECT 3520.755 2937.165 3521.935 2938.345 ;
        RECT 3519.165 2920.295 3520.345 2921.475 ;
        RECT 3520.765 2920.295 3521.945 2921.475 ;
        RECT 3525.155 2945.605 3526.335 2946.785 ;
        RECT 3526.755 2945.605 3527.935 2946.785 ;
        RECT 3525.125 2928.805 3526.305 2929.985 ;
        RECT 3526.725 2928.805 3527.905 2929.985 ;
        RECT 3466.340 2915.040 3467.520 2916.220 ;
        RECT 3467.940 2915.040 3469.120 2916.220 ;
        RECT 3525.135 2911.855 3526.315 2913.035 ;
        RECT 3526.735 2911.855 3527.915 2913.035 ;
        RECT 3460.320 2906.610 3461.500 2907.790 ;
        RECT 3461.920 2906.610 3463.100 2907.790 ;
        RECT 192.030 2887.125 202.810 2891.505 ;
        RECT 175.980 2879.215 186.760 2883.595 ;
        RECT 59.840 2849.895 61.020 2851.075 ;
        RECT 61.440 2849.895 62.620 2851.075 ;
        RECT 59.860 2825.860 61.040 2827.040 ;
        RECT 61.460 2825.860 62.640 2827.040 ;
        RECT 59.830 2808.950 61.010 2810.130 ;
        RECT 61.430 2808.950 62.610 2810.130 ;
        RECT 59.840 2792.040 61.020 2793.220 ;
        RECT 61.440 2792.040 62.620 2793.220 ;
        RECT 65.840 2846.375 67.020 2847.555 ;
        RECT 67.440 2846.375 68.620 2847.555 ;
        RECT 65.840 2817.410 67.020 2818.590 ;
        RECT 67.440 2817.410 68.620 2818.590 ;
        RECT 65.860 2800.510 67.040 2801.690 ;
        RECT 67.460 2800.510 68.640 2801.690 ;
        RECT 65.860 2783.610 67.040 2784.790 ;
        RECT 67.460 2783.610 68.640 2784.790 ;
        RECT 3347.445 2763.295 3351.825 2767.675 ;
        RECT 3328.915 2755.205 3333.295 2759.585 ;
        RECT 3466.340 2746.895 3467.520 2748.075 ;
        RECT 3467.940 2746.895 3469.120 2748.075 ;
        RECT 3460.340 2743.375 3461.520 2744.555 ;
        RECT 3461.940 2743.375 3463.120 2744.555 ;
        RECT 3460.340 2714.410 3461.520 2715.590 ;
        RECT 3461.940 2714.410 3463.120 2715.590 ;
        RECT 3460.320 2697.510 3461.500 2698.690 ;
        RECT 3461.920 2697.510 3463.100 2698.690 ;
        RECT 3466.320 2722.860 3467.500 2724.040 ;
        RECT 3467.920 2722.860 3469.100 2724.040 ;
        RECT 3466.350 2705.950 3467.530 2707.130 ;
        RECT 3467.950 2705.950 3469.130 2707.130 ;
        RECT 3519.145 2728.085 3520.325 2729.265 ;
        RECT 3520.745 2728.085 3521.925 2729.265 ;
        RECT 3519.155 2711.165 3520.335 2712.345 ;
        RECT 3520.755 2711.165 3521.935 2712.345 ;
        RECT 3519.165 2694.295 3520.345 2695.475 ;
        RECT 3520.765 2694.295 3521.945 2695.475 ;
        RECT 3525.155 2719.605 3526.335 2720.785 ;
        RECT 3526.755 2719.605 3527.935 2720.785 ;
        RECT 3525.125 2702.805 3526.305 2703.985 ;
        RECT 3526.725 2702.805 3527.905 2703.985 ;
        RECT 3466.340 2689.040 3467.520 2690.220 ;
        RECT 3467.940 2689.040 3469.120 2690.220 ;
        RECT 3525.135 2685.855 3526.315 2687.035 ;
        RECT 3526.735 2685.855 3527.915 2687.035 ;
        RECT 3460.320 2680.610 3461.500 2681.790 ;
        RECT 3461.920 2680.610 3463.100 2681.790 ;
        RECT 192.030 2665.825 202.810 2670.205 ;
        RECT 175.980 2657.915 186.760 2662.295 ;
        RECT 59.840 2633.895 61.020 2635.075 ;
        RECT 61.440 2633.895 62.620 2635.075 ;
        RECT 59.860 2609.860 61.040 2611.040 ;
        RECT 61.460 2609.860 62.640 2611.040 ;
        RECT 59.830 2592.950 61.010 2594.130 ;
        RECT 61.430 2592.950 62.610 2594.130 ;
        RECT 59.840 2576.040 61.020 2577.220 ;
        RECT 61.440 2576.040 62.620 2577.220 ;
        RECT 65.840 2630.375 67.020 2631.555 ;
        RECT 67.440 2630.375 68.620 2631.555 ;
        RECT 65.840 2601.410 67.020 2602.590 ;
        RECT 67.440 2601.410 68.620 2602.590 ;
        RECT 65.860 2584.510 67.040 2585.690 ;
        RECT 67.460 2584.510 68.640 2585.690 ;
        RECT 65.860 2567.610 67.040 2568.790 ;
        RECT 67.460 2567.610 68.640 2568.790 ;
        RECT 3347.445 2538.295 3351.825 2542.675 ;
        RECT 3328.915 2530.205 3333.295 2534.585 ;
        RECT 3466.340 2521.895 3467.520 2523.075 ;
        RECT 3467.940 2521.895 3469.120 2523.075 ;
        RECT 3460.340 2518.375 3461.520 2519.555 ;
        RECT 3461.940 2518.375 3463.120 2519.555 ;
        RECT 3460.340 2489.410 3461.520 2490.590 ;
        RECT 3461.940 2489.410 3463.120 2490.590 ;
        RECT 3460.320 2472.510 3461.500 2473.690 ;
        RECT 3461.920 2472.510 3463.100 2473.690 ;
        RECT 3466.320 2497.860 3467.500 2499.040 ;
        RECT 3467.920 2497.860 3469.100 2499.040 ;
        RECT 3466.350 2480.950 3467.530 2482.130 ;
        RECT 3467.950 2480.950 3469.130 2482.130 ;
        RECT 3519.145 2503.085 3520.325 2504.265 ;
        RECT 3520.745 2503.085 3521.925 2504.265 ;
        RECT 3519.155 2486.165 3520.335 2487.345 ;
        RECT 3520.755 2486.165 3521.935 2487.345 ;
        RECT 3519.165 2469.295 3520.345 2470.475 ;
        RECT 3520.765 2469.295 3521.945 2470.475 ;
        RECT 3525.155 2494.605 3526.335 2495.785 ;
        RECT 3526.755 2494.605 3527.935 2495.785 ;
        RECT 3525.125 2477.805 3526.305 2478.985 ;
        RECT 3526.725 2477.805 3527.905 2478.985 ;
        RECT 3466.340 2464.040 3467.520 2465.220 ;
        RECT 3467.940 2464.040 3469.120 2465.220 ;
        RECT 3525.135 2460.855 3526.315 2462.035 ;
        RECT 3526.735 2460.855 3527.915 2462.035 ;
        RECT 3460.320 2455.610 3461.500 2456.790 ;
        RECT 3461.920 2455.610 3463.100 2456.790 ;
        RECT 3347.445 2318.295 3351.825 2322.675 ;
        RECT 3328.915 2310.205 3333.295 2314.585 ;
        RECT 3466.340 2301.895 3467.520 2303.075 ;
        RECT 3467.940 2301.895 3469.120 2303.075 ;
        RECT 3460.340 2298.375 3461.520 2299.555 ;
        RECT 3461.940 2298.375 3463.120 2299.555 ;
        RECT 3460.340 2269.410 3461.520 2270.590 ;
        RECT 3461.940 2269.410 3463.120 2270.590 ;
        RECT 3460.320 2252.510 3461.500 2253.690 ;
        RECT 3461.920 2252.510 3463.100 2253.690 ;
        RECT 3466.320 2277.860 3467.500 2279.040 ;
        RECT 3467.920 2277.860 3469.100 2279.040 ;
        RECT 3466.350 2260.950 3467.530 2262.130 ;
        RECT 3467.950 2260.950 3469.130 2262.130 ;
        RECT 3519.145 2283.085 3520.325 2284.265 ;
        RECT 3520.745 2283.085 3521.925 2284.265 ;
        RECT 3519.155 2266.165 3520.335 2267.345 ;
        RECT 3520.755 2266.165 3521.935 2267.345 ;
        RECT 3519.165 2249.295 3520.345 2250.475 ;
        RECT 3520.765 2249.295 3521.945 2250.475 ;
        RECT 3525.155 2274.605 3526.335 2275.785 ;
        RECT 3526.755 2274.605 3527.935 2275.785 ;
        RECT 3525.125 2257.805 3526.305 2258.985 ;
        RECT 3526.725 2257.805 3527.905 2258.985 ;
        RECT 3466.340 2244.040 3467.520 2245.220 ;
        RECT 3467.940 2244.040 3469.120 2245.220 ;
        RECT 3525.135 2240.855 3526.315 2242.035 ;
        RECT 3526.735 2240.855 3527.915 2242.035 ;
        RECT 3460.320 2235.610 3461.500 2236.790 ;
        RECT 3461.920 2235.610 3463.100 2236.790 ;
        RECT 192.030 2027.825 202.810 2032.205 ;
        RECT 175.980 2019.915 186.760 2024.295 ;
        RECT 59.840 1995.895 61.020 1997.075 ;
        RECT 61.440 1995.895 62.620 1997.075 ;
        RECT 59.860 1971.860 61.040 1973.040 ;
        RECT 61.460 1971.860 62.640 1973.040 ;
        RECT 59.830 1954.950 61.010 1956.130 ;
        RECT 61.430 1954.950 62.610 1956.130 ;
        RECT 59.840 1938.040 61.020 1939.220 ;
        RECT 61.440 1938.040 62.620 1939.220 ;
        RECT 65.840 1992.375 67.020 1993.555 ;
        RECT 67.440 1992.375 68.620 1993.555 ;
        RECT 65.840 1963.410 67.020 1964.590 ;
        RECT 67.440 1963.410 68.620 1964.590 ;
        RECT 65.860 1946.510 67.040 1947.690 ;
        RECT 67.460 1946.510 68.640 1947.690 ;
        RECT 65.860 1929.610 67.040 1930.790 ;
        RECT 67.460 1929.610 68.640 1930.790 ;
        RECT 3347.445 1877.295 3351.825 1881.675 ;
        RECT 3328.915 1869.205 3333.295 1873.585 ;
        RECT 3466.340 1860.895 3467.520 1862.075 ;
        RECT 3467.940 1860.895 3469.120 1862.075 ;
        RECT 3460.340 1857.375 3461.520 1858.555 ;
        RECT 3461.940 1857.375 3463.120 1858.555 ;
        RECT 3460.340 1828.410 3461.520 1829.590 ;
        RECT 3461.940 1828.410 3463.120 1829.590 ;
        RECT 192.030 1811.825 202.810 1816.205 ;
        RECT 3460.320 1811.510 3461.500 1812.690 ;
        RECT 3461.920 1811.510 3463.100 1812.690 ;
        RECT 175.980 1803.915 186.760 1808.295 ;
        RECT 3466.320 1836.860 3467.500 1838.040 ;
        RECT 3467.920 1836.860 3469.100 1838.040 ;
        RECT 3466.350 1819.950 3467.530 1821.130 ;
        RECT 3467.950 1819.950 3469.130 1821.130 ;
        RECT 3519.145 1842.085 3520.325 1843.265 ;
        RECT 3520.745 1842.085 3521.925 1843.265 ;
        RECT 3519.155 1825.165 3520.335 1826.345 ;
        RECT 3520.755 1825.165 3521.935 1826.345 ;
        RECT 3519.165 1808.295 3520.345 1809.475 ;
        RECT 3520.765 1808.295 3521.945 1809.475 ;
        RECT 3525.155 1833.605 3526.335 1834.785 ;
        RECT 3526.755 1833.605 3527.935 1834.785 ;
        RECT 3525.125 1816.805 3526.305 1817.985 ;
        RECT 3526.725 1816.805 3527.905 1817.985 ;
        RECT 3466.340 1803.040 3467.520 1804.220 ;
        RECT 3467.940 1803.040 3469.120 1804.220 ;
        RECT 3525.135 1799.855 3526.315 1801.035 ;
        RECT 3526.735 1799.855 3527.915 1801.035 ;
        RECT 3460.320 1794.610 3461.500 1795.790 ;
        RECT 3461.920 1794.610 3463.100 1795.790 ;
        RECT 59.840 1779.895 61.020 1781.075 ;
        RECT 61.440 1779.895 62.620 1781.075 ;
        RECT 59.860 1755.860 61.040 1757.040 ;
        RECT 61.460 1755.860 62.640 1757.040 ;
        RECT 59.830 1738.950 61.010 1740.130 ;
        RECT 61.430 1738.950 62.610 1740.130 ;
        RECT 59.840 1722.040 61.020 1723.220 ;
        RECT 61.440 1722.040 62.620 1723.220 ;
        RECT 65.840 1776.375 67.020 1777.555 ;
        RECT 67.440 1776.375 68.620 1777.555 ;
        RECT 65.840 1747.410 67.020 1748.590 ;
        RECT 67.440 1747.410 68.620 1748.590 ;
        RECT 65.860 1730.510 67.040 1731.690 ;
        RECT 67.460 1730.510 68.640 1731.690 ;
        RECT 65.860 1713.610 67.040 1714.790 ;
        RECT 67.460 1713.610 68.640 1714.790 ;
        RECT 3347.445 1651.295 3351.825 1655.675 ;
        RECT 3328.915 1643.205 3333.295 1647.585 ;
        RECT 3466.340 1634.895 3467.520 1636.075 ;
        RECT 3467.940 1634.895 3469.120 1636.075 ;
        RECT 3460.340 1631.375 3461.520 1632.555 ;
        RECT 3461.940 1631.375 3463.120 1632.555 ;
        RECT 192.030 1600.825 202.810 1605.205 ;
        RECT 3460.340 1602.410 3461.520 1603.590 ;
        RECT 3461.940 1602.410 3463.120 1603.590 ;
        RECT 175.980 1592.915 186.760 1597.295 ;
        RECT 3460.320 1585.510 3461.500 1586.690 ;
        RECT 3461.920 1585.510 3463.100 1586.690 ;
        RECT 3466.320 1610.860 3467.500 1612.040 ;
        RECT 3467.920 1610.860 3469.100 1612.040 ;
        RECT 3466.350 1593.950 3467.530 1595.130 ;
        RECT 3467.950 1593.950 3469.130 1595.130 ;
        RECT 3519.145 1616.085 3520.325 1617.265 ;
        RECT 3520.745 1616.085 3521.925 1617.265 ;
        RECT 3519.155 1599.165 3520.335 1600.345 ;
        RECT 3520.755 1599.165 3521.935 1600.345 ;
        RECT 3519.165 1582.295 3520.345 1583.475 ;
        RECT 3520.765 1582.295 3521.945 1583.475 ;
        RECT 3525.155 1607.605 3526.335 1608.785 ;
        RECT 3526.755 1607.605 3527.935 1608.785 ;
        RECT 3525.125 1590.805 3526.305 1591.985 ;
        RECT 3526.725 1590.805 3527.905 1591.985 ;
        RECT 3466.340 1577.040 3467.520 1578.220 ;
        RECT 3467.940 1577.040 3469.120 1578.220 ;
        RECT 3525.135 1573.855 3526.315 1575.035 ;
        RECT 3526.735 1573.855 3527.915 1575.035 ;
        RECT 59.840 1563.895 61.020 1565.075 ;
        RECT 61.440 1563.895 62.620 1565.075 ;
        RECT 3460.320 1568.610 3461.500 1569.790 ;
        RECT 3461.920 1568.610 3463.100 1569.790 ;
        RECT 59.860 1539.860 61.040 1541.040 ;
        RECT 61.460 1539.860 62.640 1541.040 ;
        RECT 59.830 1522.950 61.010 1524.130 ;
        RECT 61.430 1522.950 62.610 1524.130 ;
        RECT 59.840 1506.040 61.020 1507.220 ;
        RECT 61.440 1506.040 62.620 1507.220 ;
        RECT 65.840 1560.375 67.020 1561.555 ;
        RECT 67.440 1560.375 68.620 1561.555 ;
        RECT 65.840 1531.410 67.020 1532.590 ;
        RECT 67.440 1531.410 68.620 1532.590 ;
        RECT 65.860 1514.510 67.040 1515.690 ;
        RECT 67.460 1514.510 68.640 1515.690 ;
        RECT 65.860 1497.610 67.040 1498.790 ;
        RECT 67.460 1497.610 68.640 1498.790 ;
        RECT 3347.445 1426.295 3351.825 1430.675 ;
        RECT 3328.915 1418.205 3333.295 1422.585 ;
        RECT 3466.340 1409.895 3467.520 1411.075 ;
        RECT 3467.940 1409.895 3469.120 1411.075 ;
        RECT 3460.340 1406.375 3461.520 1407.555 ;
        RECT 3461.940 1406.375 3463.120 1407.555 ;
        RECT 192.030 1379.825 202.810 1384.205 ;
        RECT 3460.340 1377.410 3461.520 1378.590 ;
        RECT 3461.940 1377.410 3463.120 1378.590 ;
        RECT 175.980 1371.915 186.760 1376.295 ;
        RECT 3460.320 1360.510 3461.500 1361.690 ;
        RECT 3461.920 1360.510 3463.100 1361.690 ;
        RECT 59.840 1347.895 61.020 1349.075 ;
        RECT 61.440 1347.895 62.620 1349.075 ;
        RECT 59.860 1323.860 61.040 1325.040 ;
        RECT 61.460 1323.860 62.640 1325.040 ;
        RECT 59.830 1306.950 61.010 1308.130 ;
        RECT 61.430 1306.950 62.610 1308.130 ;
        RECT 59.840 1290.040 61.020 1291.220 ;
        RECT 61.440 1290.040 62.620 1291.220 ;
        RECT 65.840 1344.375 67.020 1345.555 ;
        RECT 67.440 1344.375 68.620 1345.555 ;
        RECT 3466.320 1385.860 3467.500 1387.040 ;
        RECT 3467.920 1385.860 3469.100 1387.040 ;
        RECT 3466.350 1368.950 3467.530 1370.130 ;
        RECT 3467.950 1368.950 3469.130 1370.130 ;
        RECT 3519.145 1391.085 3520.325 1392.265 ;
        RECT 3520.745 1391.085 3521.925 1392.265 ;
        RECT 3519.155 1374.165 3520.335 1375.345 ;
        RECT 3520.755 1374.165 3521.935 1375.345 ;
        RECT 3519.165 1357.295 3520.345 1358.475 ;
        RECT 3520.765 1357.295 3521.945 1358.475 ;
        RECT 3525.155 1382.605 3526.335 1383.785 ;
        RECT 3526.755 1382.605 3527.935 1383.785 ;
        RECT 3525.125 1365.805 3526.305 1366.985 ;
        RECT 3526.725 1365.805 3527.905 1366.985 ;
        RECT 3466.340 1352.040 3467.520 1353.220 ;
        RECT 3467.940 1352.040 3469.120 1353.220 ;
        RECT 3525.135 1348.855 3526.315 1350.035 ;
        RECT 3526.735 1348.855 3527.915 1350.035 ;
        RECT 3460.320 1343.610 3461.500 1344.790 ;
        RECT 3461.920 1343.610 3463.100 1344.790 ;
        RECT 65.840 1315.410 67.020 1316.590 ;
        RECT 67.440 1315.410 68.620 1316.590 ;
        RECT 65.860 1298.510 67.040 1299.690 ;
        RECT 67.460 1298.510 68.640 1299.690 ;
        RECT 65.860 1281.610 67.040 1282.790 ;
        RECT 67.460 1281.610 68.640 1282.790 ;
        RECT 3264.810 1220.375 3265.990 1221.555 ;
        RECT 3266.410 1220.375 3267.590 1221.555 ;
        RECT 3268.010 1220.375 3269.190 1221.555 ;
        RECT 3269.610 1220.375 3270.790 1221.555 ;
        RECT 3271.210 1220.375 3272.390 1221.555 ;
        RECT 3272.810 1220.375 3273.990 1221.555 ;
        RECT 3274.410 1220.375 3275.590 1221.555 ;
        RECT 3276.010 1220.375 3277.190 1221.555 ;
        RECT 3277.610 1220.375 3278.790 1221.555 ;
        RECT 3279.210 1220.375 3280.390 1221.555 ;
        RECT 3280.810 1220.375 3281.990 1221.555 ;
        RECT 3282.410 1220.375 3283.590 1221.555 ;
        RECT 3284.010 1220.375 3285.190 1221.555 ;
        RECT 191.175 1210.385 203.555 1216.365 ;
        RECT 3264.715 1215.650 3265.895 1216.830 ;
        RECT 3266.315 1215.650 3267.495 1216.830 ;
        RECT 3267.915 1215.650 3269.095 1216.830 ;
        RECT 3269.515 1215.650 3270.695 1216.830 ;
        RECT 3271.115 1215.650 3272.295 1216.830 ;
        RECT 3272.715 1215.650 3273.895 1216.830 ;
        RECT 3274.315 1215.650 3275.495 1216.830 ;
        RECT 3275.915 1215.650 3277.095 1216.830 ;
        RECT 3277.515 1215.650 3278.695 1216.830 ;
        RECT 3279.115 1215.650 3280.295 1216.830 ;
        RECT 3280.715 1215.650 3281.895 1216.830 ;
        RECT 3282.315 1215.650 3283.495 1216.830 ;
        RECT 3283.915 1215.650 3285.095 1216.830 ;
        RECT 248.970 1210.760 250.150 1211.940 ;
        RECT 250.570 1210.760 251.750 1211.940 ;
        RECT 3324.320 1211.220 3336.700 1217.200 ;
        RECT 3340.320 1214.650 3352.700 1222.230 ;
        RECT 184.395 1177.600 187.175 1207.580 ;
        RECT 249.010 1205.990 250.190 1207.170 ;
        RECT 250.610 1205.990 251.790 1207.170 ;
        RECT 3347.445 1201.295 3351.825 1205.675 ;
        RECT 3328.915 1193.205 3333.295 1197.585 ;
        RECT 3466.340 1184.895 3467.520 1186.075 ;
        RECT 3467.940 1184.895 3469.120 1186.075 ;
        RECT 3460.340 1181.375 3461.520 1182.555 ;
        RECT 3461.940 1181.375 3463.120 1182.555 ;
        RECT 3460.340 1152.410 3461.520 1153.590 ;
        RECT 3461.940 1152.410 3463.120 1153.590 ;
        RECT 59.840 1131.895 61.020 1133.075 ;
        RECT 61.440 1131.895 62.620 1133.075 ;
        RECT 3460.320 1135.510 3461.500 1136.690 ;
        RECT 3461.920 1135.510 3463.100 1136.690 ;
        RECT 59.860 1107.860 61.040 1109.040 ;
        RECT 61.460 1107.860 62.640 1109.040 ;
        RECT 59.830 1090.950 61.010 1092.130 ;
        RECT 61.430 1090.950 62.610 1092.130 ;
        RECT 59.840 1074.040 61.020 1075.220 ;
        RECT 61.440 1074.040 62.620 1075.220 ;
        RECT 65.840 1128.375 67.020 1129.555 ;
        RECT 67.440 1128.375 68.620 1129.555 ;
        RECT 3466.320 1160.860 3467.500 1162.040 ;
        RECT 3467.920 1160.860 3469.100 1162.040 ;
        RECT 3466.350 1143.950 3467.530 1145.130 ;
        RECT 3467.950 1143.950 3469.130 1145.130 ;
        RECT 3519.145 1166.085 3520.325 1167.265 ;
        RECT 3520.745 1166.085 3521.925 1167.265 ;
        RECT 3519.155 1149.165 3520.335 1150.345 ;
        RECT 3520.755 1149.165 3521.935 1150.345 ;
        RECT 3519.165 1132.295 3520.345 1133.475 ;
        RECT 3520.765 1132.295 3521.945 1133.475 ;
        RECT 3525.155 1157.605 3526.335 1158.785 ;
        RECT 3526.755 1157.605 3527.935 1158.785 ;
        RECT 3525.125 1140.805 3526.305 1141.985 ;
        RECT 3526.725 1140.805 3527.905 1141.985 ;
        RECT 3466.340 1127.040 3467.520 1128.220 ;
        RECT 3467.940 1127.040 3469.120 1128.220 ;
        RECT 3525.135 1123.855 3526.315 1125.035 ;
        RECT 3526.735 1123.855 3527.915 1125.035 ;
        RECT 3460.320 1118.610 3461.500 1119.790 ;
        RECT 3461.920 1118.610 3463.100 1119.790 ;
        RECT 65.840 1099.410 67.020 1100.590 ;
        RECT 67.440 1099.410 68.620 1100.590 ;
        RECT 65.860 1082.510 67.040 1083.690 ;
        RECT 67.460 1082.510 68.640 1083.690 ;
        RECT 65.860 1065.610 67.040 1066.790 ;
        RECT 67.460 1065.610 68.640 1066.790 ;
        RECT 3347.445 975.295 3351.825 979.675 ;
        RECT 3328.915 967.205 3333.295 971.585 ;
        RECT 3466.340 958.895 3467.520 960.075 ;
        RECT 3467.940 958.895 3469.120 960.075 ;
        RECT 3460.340 955.375 3461.520 956.555 ;
        RECT 3461.940 955.375 3463.120 956.555 ;
        RECT 3460.340 926.410 3461.520 927.590 ;
        RECT 3461.940 926.410 3463.120 927.590 ;
        RECT 59.840 915.895 61.020 917.075 ;
        RECT 61.440 915.895 62.620 917.075 ;
        RECT 59.860 891.860 61.040 893.040 ;
        RECT 61.460 891.860 62.640 893.040 ;
        RECT 59.830 874.950 61.010 876.130 ;
        RECT 61.430 874.950 62.610 876.130 ;
        RECT 59.840 858.040 61.020 859.220 ;
        RECT 61.440 858.040 62.620 859.220 ;
        RECT 65.840 912.375 67.020 913.555 ;
        RECT 67.440 912.375 68.620 913.555 ;
        RECT 3460.320 909.510 3461.500 910.690 ;
        RECT 3461.920 909.510 3463.100 910.690 ;
        RECT 3466.320 934.860 3467.500 936.040 ;
        RECT 3467.920 934.860 3469.100 936.040 ;
        RECT 3466.350 917.950 3467.530 919.130 ;
        RECT 3467.950 917.950 3469.130 919.130 ;
        RECT 3519.145 940.085 3520.325 941.265 ;
        RECT 3520.745 940.085 3521.925 941.265 ;
        RECT 3519.155 923.165 3520.335 924.345 ;
        RECT 3520.755 923.165 3521.935 924.345 ;
        RECT 3519.165 906.295 3520.345 907.475 ;
        RECT 3520.765 906.295 3521.945 907.475 ;
        RECT 3525.155 931.605 3526.335 932.785 ;
        RECT 3526.755 931.605 3527.935 932.785 ;
        RECT 3525.125 914.805 3526.305 915.985 ;
        RECT 3526.725 914.805 3527.905 915.985 ;
        RECT 3466.340 901.040 3467.520 902.220 ;
        RECT 3467.940 901.040 3469.120 902.220 ;
        RECT 3525.135 897.855 3526.315 899.035 ;
        RECT 3526.735 897.855 3527.915 899.035 ;
        RECT 3460.320 892.610 3461.500 893.790 ;
        RECT 3461.920 892.610 3463.100 893.790 ;
        RECT 65.840 883.410 67.020 884.590 ;
        RECT 67.440 883.410 68.620 884.590 ;
        RECT 65.860 866.510 67.040 867.690 ;
        RECT 67.460 866.510 68.640 867.690 ;
        RECT 65.860 849.610 67.040 850.790 ;
        RECT 67.460 849.610 68.640 850.790 ;
        RECT 3347.445 750.295 3351.825 754.675 ;
        RECT 3328.915 742.205 3333.295 746.585 ;
        RECT 3466.340 733.895 3467.520 735.075 ;
        RECT 3467.940 733.895 3469.120 735.075 ;
        RECT 3460.340 730.375 3461.520 731.555 ;
        RECT 3461.940 730.375 3463.120 731.555 ;
        RECT 3460.340 701.410 3461.520 702.590 ;
        RECT 3461.940 701.410 3463.120 702.590 ;
        RECT 3460.320 684.510 3461.500 685.690 ;
        RECT 3461.920 684.510 3463.100 685.690 ;
        RECT 3466.320 709.860 3467.500 711.040 ;
        RECT 3467.920 709.860 3469.100 711.040 ;
        RECT 3466.350 692.950 3467.530 694.130 ;
        RECT 3467.950 692.950 3469.130 694.130 ;
        RECT 3519.145 715.085 3520.325 716.265 ;
        RECT 3520.745 715.085 3521.925 716.265 ;
        RECT 3519.155 698.165 3520.335 699.345 ;
        RECT 3520.755 698.165 3521.935 699.345 ;
        RECT 3519.165 681.295 3520.345 682.475 ;
        RECT 3520.765 681.295 3521.945 682.475 ;
        RECT 3525.155 706.605 3526.335 707.785 ;
        RECT 3526.755 706.605 3527.935 707.785 ;
        RECT 3525.125 689.805 3526.305 690.985 ;
        RECT 3526.725 689.805 3527.905 690.985 ;
        RECT 3466.340 676.040 3467.520 677.220 ;
        RECT 3467.940 676.040 3469.120 677.220 ;
        RECT 3525.135 672.855 3526.315 674.035 ;
        RECT 3526.735 672.855 3527.915 674.035 ;
        RECT 3460.320 667.610 3461.500 668.790 ;
        RECT 3461.920 667.610 3463.100 668.790 ;
        RECT 3347.445 524.295 3351.825 528.675 ;
        RECT 3328.915 516.205 3333.295 520.585 ;
        RECT 3466.340 507.895 3467.520 509.075 ;
        RECT 3467.940 507.895 3469.120 509.075 ;
        RECT 3460.340 504.375 3461.520 505.555 ;
        RECT 3461.940 504.375 3463.120 505.555 ;
        RECT 3460.340 475.410 3461.520 476.590 ;
        RECT 3461.940 475.410 3463.120 476.590 ;
        RECT 3460.320 458.510 3461.500 459.690 ;
        RECT 3461.920 458.510 3463.100 459.690 ;
        RECT 3466.320 483.860 3467.500 485.040 ;
        RECT 3467.920 483.860 3469.100 485.040 ;
        RECT 3466.350 466.950 3467.530 468.130 ;
        RECT 3467.950 466.950 3469.130 468.130 ;
        RECT 3519.145 489.085 3520.325 490.265 ;
        RECT 3520.745 489.085 3521.925 490.265 ;
        RECT 3519.155 472.165 3520.335 473.345 ;
        RECT 3520.755 472.165 3521.935 473.345 ;
        RECT 3519.165 455.295 3520.345 456.475 ;
        RECT 3520.765 455.295 3521.945 456.475 ;
        RECT 3525.155 480.605 3526.335 481.785 ;
        RECT 3526.755 480.605 3527.935 481.785 ;
        RECT 3525.125 463.805 3526.305 464.985 ;
        RECT 3526.725 463.805 3527.905 464.985 ;
        RECT 3466.340 450.040 3467.520 451.220 ;
        RECT 3467.940 450.040 3469.120 451.220 ;
        RECT 3525.135 446.855 3526.315 448.035 ;
        RECT 3526.735 446.855 3527.915 448.035 ;
        RECT 3460.320 441.610 3461.500 442.790 ;
        RECT 3461.920 441.610 3463.100 442.790 ;
      LAYER met5 ;
        RECT 461.790 4923.960 463.390 4931.970 ;
        RECT 470.240 4929.950 471.840 4931.970 ;
        RECT 470.170 4925.570 471.900 4929.950 ;
        RECT 478.690 4923.970 480.290 4931.970 ;
        RECT 487.140 4930.030 488.740 4931.970 ;
        RECT 487.030 4925.650 488.790 4930.030 ;
        RECT 495.590 4923.980 497.190 4931.970 ;
        RECT 504.040 4929.890 505.640 4931.970 ;
        RECT 504.000 4925.510 505.730 4929.890 ;
        RECT 461.730 4919.580 463.460 4923.960 ;
        RECT 478.630 4919.590 480.360 4923.970 ;
        RECT 495.510 4919.600 497.240 4923.980 ;
        RECT 524.540 4923.850 526.140 4947.540 ;
        RECT 528.040 4930.110 529.640 4947.540 ;
        RECT 528.020 4925.730 529.750 4930.110 ;
        RECT 718.790 4923.960 720.390 4931.970 ;
        RECT 727.240 4929.950 728.840 4931.970 ;
        RECT 727.170 4925.570 728.900 4929.950 ;
        RECT 735.690 4923.970 737.290 4931.970 ;
        RECT 744.140 4930.030 745.740 4931.970 ;
        RECT 744.030 4925.650 745.790 4930.030 ;
        RECT 752.590 4923.980 754.190 4931.970 ;
        RECT 761.040 4929.890 762.640 4931.970 ;
        RECT 761.000 4925.510 762.730 4929.890 ;
        RECT 495.590 4919.590 497.190 4919.600 ;
        RECT 524.510 4919.470 526.240 4923.850 ;
        RECT 718.730 4919.580 720.460 4923.960 ;
        RECT 735.630 4919.590 737.360 4923.970 ;
        RECT 752.510 4919.600 754.240 4923.980 ;
        RECT 781.540 4923.850 783.140 4947.540 ;
        RECT 785.040 4930.110 786.640 4947.540 ;
        RECT 785.020 4925.730 786.750 4930.110 ;
        RECT 975.790 4923.960 977.390 4931.970 ;
        RECT 984.240 4929.950 985.840 4931.970 ;
        RECT 984.170 4925.570 985.900 4929.950 ;
        RECT 992.690 4923.970 994.290 4931.970 ;
        RECT 1001.140 4930.030 1002.740 4931.970 ;
        RECT 1001.030 4925.650 1002.790 4930.030 ;
        RECT 1009.590 4923.980 1011.190 4931.970 ;
        RECT 1018.040 4929.890 1019.640 4931.970 ;
        RECT 1018.000 4925.510 1019.730 4929.890 ;
        RECT 752.590 4919.590 754.190 4919.600 ;
        RECT 781.510 4919.470 783.240 4923.850 ;
        RECT 975.730 4919.580 977.460 4923.960 ;
        RECT 992.630 4919.590 994.360 4923.970 ;
        RECT 1009.510 4919.600 1011.240 4923.980 ;
        RECT 1038.540 4923.850 1040.140 4947.540 ;
        RECT 1042.040 4930.110 1043.640 4947.540 ;
        RECT 1042.020 4925.730 1043.750 4930.110 ;
        RECT 1232.790 4923.960 1234.390 4931.970 ;
        RECT 1241.240 4929.950 1242.840 4931.970 ;
        RECT 1241.170 4925.570 1242.900 4929.950 ;
        RECT 1249.690 4923.970 1251.290 4931.970 ;
        RECT 1258.140 4930.030 1259.740 4931.970 ;
        RECT 1258.030 4925.650 1259.790 4930.030 ;
        RECT 1266.590 4923.980 1268.190 4931.970 ;
        RECT 1275.040 4929.890 1276.640 4931.970 ;
        RECT 1275.000 4925.510 1276.730 4929.890 ;
        RECT 1009.590 4919.590 1011.190 4919.600 ;
        RECT 1038.510 4919.470 1040.240 4923.850 ;
        RECT 1232.730 4919.580 1234.460 4923.960 ;
        RECT 1249.630 4919.590 1251.360 4923.970 ;
        RECT 1266.510 4919.600 1268.240 4923.980 ;
        RECT 1295.540 4923.850 1297.140 4947.540 ;
        RECT 1299.040 4930.110 1300.640 4947.540 ;
        RECT 1299.020 4925.730 1300.750 4930.110 ;
        RECT 1490.790 4923.960 1492.390 4931.970 ;
        RECT 1499.240 4929.950 1500.840 4931.970 ;
        RECT 1499.170 4925.570 1500.900 4929.950 ;
        RECT 1507.690 4923.970 1509.290 4931.970 ;
        RECT 1516.140 4930.030 1517.740 4931.970 ;
        RECT 1516.030 4925.650 1517.790 4930.030 ;
        RECT 1524.590 4923.980 1526.190 4931.970 ;
        RECT 1533.040 4929.890 1534.640 4931.970 ;
        RECT 1533.000 4925.510 1534.730 4929.890 ;
        RECT 1266.590 4919.590 1268.190 4919.600 ;
        RECT 1295.510 4919.470 1297.240 4923.850 ;
        RECT 1490.730 4919.580 1492.460 4923.960 ;
        RECT 1507.630 4919.590 1509.360 4923.970 ;
        RECT 1524.510 4919.600 1526.240 4923.980 ;
        RECT 1553.540 4923.850 1555.140 4947.540 ;
        RECT 1557.040 4930.110 1558.640 4947.540 ;
        RECT 1557.020 4925.730 1558.750 4930.110 ;
        RECT 1742.790 4923.960 1744.390 4931.970 ;
        RECT 1751.240 4929.950 1752.840 4931.970 ;
        RECT 1751.170 4925.570 1752.900 4929.950 ;
        RECT 1759.690 4923.970 1761.290 4931.970 ;
        RECT 1768.140 4930.030 1769.740 4931.970 ;
        RECT 1768.030 4925.650 1769.790 4930.030 ;
        RECT 1776.590 4923.980 1778.190 4931.970 ;
        RECT 1785.040 4929.890 1786.640 4931.970 ;
        RECT 1785.000 4925.510 1786.730 4929.890 ;
        RECT 1524.590 4919.590 1526.190 4919.600 ;
        RECT 1553.510 4919.470 1555.240 4923.850 ;
        RECT 1742.730 4919.580 1744.460 4923.960 ;
        RECT 1759.630 4919.590 1761.360 4923.970 ;
        RECT 1776.510 4919.600 1778.240 4923.980 ;
        RECT 1805.540 4923.850 1807.140 4947.540 ;
        RECT 1809.040 4930.110 1810.640 4947.540 ;
        RECT 1809.020 4925.730 1810.750 4930.110 ;
        RECT 2079.790 4923.960 2081.390 4931.970 ;
        RECT 2088.240 4929.950 2089.840 4931.970 ;
        RECT 2088.170 4925.570 2089.900 4929.950 ;
        RECT 2096.690 4923.970 2098.290 4931.970 ;
        RECT 2105.140 4930.030 2106.740 4931.970 ;
        RECT 2105.030 4925.650 2106.790 4930.030 ;
        RECT 2113.590 4923.980 2115.190 4931.970 ;
        RECT 2122.040 4929.890 2123.640 4931.970 ;
        RECT 2122.000 4925.510 2123.730 4929.890 ;
        RECT 1776.590 4919.590 1778.190 4919.600 ;
        RECT 1805.510 4919.470 1807.240 4923.850 ;
        RECT 2079.730 4919.580 2081.460 4923.960 ;
        RECT 2096.630 4919.590 2098.360 4923.970 ;
        RECT 2113.510 4919.600 2115.240 4923.980 ;
        RECT 2142.540 4923.850 2144.140 4947.540 ;
        RECT 2146.040 4930.110 2147.640 4947.540 ;
        RECT 2146.020 4925.730 2147.750 4930.110 ;
        RECT 2464.790 4923.960 2466.390 4931.970 ;
        RECT 2473.240 4929.950 2474.840 4931.970 ;
        RECT 2473.170 4925.570 2474.900 4929.950 ;
        RECT 2481.690 4923.970 2483.290 4931.970 ;
        RECT 2490.140 4930.030 2491.740 4931.970 ;
        RECT 2490.030 4925.650 2491.790 4930.030 ;
        RECT 2498.590 4923.980 2500.190 4931.970 ;
        RECT 2507.040 4929.890 2508.640 4931.970 ;
        RECT 2507.000 4925.510 2508.730 4929.890 ;
        RECT 2113.590 4919.590 2115.190 4919.600 ;
        RECT 2142.510 4919.470 2144.240 4923.850 ;
        RECT 2464.730 4919.580 2466.460 4923.960 ;
        RECT 2481.630 4919.590 2483.360 4923.970 ;
        RECT 2498.510 4919.600 2500.240 4923.980 ;
        RECT 2527.540 4923.850 2529.140 4947.540 ;
        RECT 2531.040 4930.110 2532.640 4947.540 ;
        RECT 2531.020 4925.730 2532.750 4930.110 ;
        RECT 2721.790 4923.960 2723.390 4931.970 ;
        RECT 2730.240 4929.950 2731.840 4931.970 ;
        RECT 2730.170 4925.570 2731.900 4929.950 ;
        RECT 2738.690 4923.970 2740.290 4931.970 ;
        RECT 2747.140 4930.030 2748.740 4931.970 ;
        RECT 2747.030 4925.650 2748.790 4930.030 ;
        RECT 2755.590 4923.980 2757.190 4931.970 ;
        RECT 2764.040 4929.890 2765.640 4931.970 ;
        RECT 2764.000 4925.510 2765.730 4929.890 ;
        RECT 2498.590 4919.590 2500.190 4919.600 ;
        RECT 2527.510 4919.470 2529.240 4923.850 ;
        RECT 2721.730 4919.580 2723.460 4923.960 ;
        RECT 2738.630 4919.590 2740.360 4923.970 ;
        RECT 2755.510 4919.600 2757.240 4923.980 ;
        RECT 2784.540 4923.850 2786.140 4947.540 ;
        RECT 2788.040 4930.110 2789.640 4947.540 ;
        RECT 2788.020 4925.730 2789.750 4930.110 ;
        RECT 2755.590 4919.590 2757.190 4919.600 ;
        RECT 2784.510 4919.470 2786.240 4923.850 ;
        RECT 175.060 4759.890 187.760 4762.740 ;
        RECT 248.770 4759.740 272.070 4762.840 ;
        RECT 191.100 4755.090 203.750 4757.990 ;
        RECT 248.770 4754.940 276.880 4758.040 ;
        RECT 3230.790 4750.140 3285.780 4753.240 ;
        RECT 3324.180 4750.250 3336.810 4753.180 ;
        RECT 3226.030 4745.340 3285.780 4748.440 ;
        RECT 3340.170 4745.440 3352.800 4748.370 ;
        RECT 191.280 4590.380 203.560 4595.650 ;
        RECT 175.230 4582.470 187.510 4587.740 ;
        RECT 59.120 4560.280 63.315 4560.395 ;
        RECT 41.440 4558.680 63.315 4560.280 ;
        RECT 59.120 4558.590 63.315 4558.680 ;
        RECT 65.150 4556.780 69.345 4556.850 ;
        RECT 41.440 4555.180 69.500 4556.780 ;
        RECT 3346.880 4556.740 3352.290 4562.230 ;
        RECT 65.150 4555.045 69.345 4555.180 ;
        RECT 3328.350 4548.650 3333.760 4554.140 ;
        RECT 3465.630 4542.280 3469.760 4542.340 ;
        RECT 3465.630 4540.680 3487.470 4542.280 ;
        RECT 3465.630 4540.625 3469.760 4540.680 ;
        RECT 3459.575 4538.780 3463.705 4538.855 ;
        RECT 3459.410 4537.180 3487.470 4538.780 ;
        RECT 3459.575 4537.140 3463.705 4537.180 ;
        RECT 59.135 4536.250 63.345 4536.340 ;
        RECT 57.010 4534.650 63.430 4536.250 ;
        RECT 59.135 4534.540 63.345 4534.650 ;
        RECT 65.170 4527.800 69.380 4527.865 ;
        RECT 57.010 4526.200 69.390 4527.800 ;
        RECT 65.170 4526.120 69.380 4526.200 ;
        RECT 3518.420 4523.490 3522.605 4523.575 ;
        RECT 3516.110 4521.890 3522.720 4523.490 ;
        RECT 3518.420 4521.800 3522.605 4521.890 ;
        RECT 59.175 4519.350 63.385 4519.390 ;
        RECT 57.010 4517.750 63.385 4519.350 ;
        RECT 59.175 4517.645 63.385 4517.750 ;
        RECT 3465.470 4518.250 3469.795 4518.350 ;
        RECT 3465.470 4516.650 3471.900 4518.250 ;
        RECT 3465.470 4516.580 3469.795 4516.650 ;
        RECT 3524.425 4515.040 3528.610 4515.120 ;
        RECT 3516.110 4513.440 3528.780 4515.040 ;
        RECT 3524.425 4513.345 3528.610 4513.440 ;
        RECT 65.155 4510.900 69.365 4510.975 ;
        RECT 57.010 4509.300 69.390 4510.900 ;
        RECT 3459.485 4509.800 3463.810 4509.860 ;
        RECT 65.155 4509.230 69.365 4509.300 ;
        RECT 3459.485 4508.200 3471.900 4509.800 ;
        RECT 3459.485 4508.090 3463.810 4508.200 ;
        RECT 3518.395 4506.590 3522.580 4506.705 ;
        RECT 3516.110 4504.990 3522.690 4506.590 ;
        RECT 3518.395 4504.930 3522.580 4504.990 ;
        RECT 59.155 4502.450 63.365 4502.525 ;
        RECT 57.010 4500.850 63.400 4502.450 ;
        RECT 3465.585 4501.350 3469.910 4501.435 ;
        RECT 59.155 4500.780 63.365 4500.850 ;
        RECT 3465.585 4499.750 3471.900 4501.350 ;
        RECT 3465.585 4499.665 3469.910 4499.750 ;
        RECT 3524.370 4498.140 3528.780 4498.250 ;
        RECT 3516.110 4496.640 3528.780 4498.140 ;
        RECT 3516.110 4496.560 3528.775 4496.640 ;
        RECT 3516.110 4496.540 3528.770 4496.560 ;
        RECT 65.200 4494.000 69.410 4494.075 ;
        RECT 57.010 4492.400 69.410 4494.000 ;
        RECT 65.200 4492.330 69.410 4492.400 ;
        RECT 3459.490 4492.900 3463.815 4492.960 ;
        RECT 3459.490 4491.300 3471.900 4492.900 ;
        RECT 3459.490 4491.190 3463.815 4491.300 ;
        RECT 3518.400 4489.690 3522.580 4489.780 ;
        RECT 3515.950 4488.090 3522.580 4489.690 ;
        RECT 3518.400 4487.980 3522.580 4488.090 ;
        RECT 3465.490 4484.450 3469.815 4484.555 ;
        RECT 3465.490 4482.850 3471.900 4484.450 ;
        RECT 3465.490 4482.785 3469.815 4482.850 ;
        RECT 3524.365 4481.240 3528.550 4481.320 ;
        RECT 3515.950 4479.640 3528.550 4481.240 ;
        RECT 3524.365 4479.545 3528.550 4479.640 ;
        RECT 3459.520 4476.000 3463.845 4476.100 ;
        RECT 3459.520 4474.400 3471.900 4476.000 ;
        RECT 3459.520 4474.330 3463.845 4474.400 ;
        RECT 3343.560 4330.870 3348.590 4336.060 ;
        RECT 3327.720 4322.830 3332.870 4328.020 ;
        RECT 3340.470 4105.760 3345.790 4111.080 ;
        RECT 3327.740 4097.710 3333.080 4103.110 ;
        RECT 191.280 3961.380 203.560 3966.650 ;
        RECT 175.230 3953.470 187.510 3958.740 ;
        RECT 59.120 3931.280 63.315 3931.395 ;
        RECT 41.440 3929.680 63.315 3931.280 ;
        RECT 59.120 3929.590 63.315 3929.680 ;
        RECT 65.150 3927.780 69.345 3927.850 ;
        RECT 41.440 3926.180 69.500 3927.780 ;
        RECT 65.150 3926.045 69.345 3926.180 ;
        RECT 59.135 3907.250 63.345 3907.340 ;
        RECT 57.010 3905.650 63.430 3907.250 ;
        RECT 59.135 3905.540 63.345 3905.650 ;
        RECT 65.170 3898.800 69.380 3898.865 ;
        RECT 57.010 3897.200 69.390 3898.800 ;
        RECT 65.170 3897.120 69.380 3897.200 ;
        RECT 59.175 3890.350 63.385 3890.390 ;
        RECT 57.010 3888.750 63.385 3890.350 ;
        RECT 59.175 3888.645 63.385 3888.750 ;
        RECT 65.155 3881.900 69.365 3881.975 ;
        RECT 57.010 3880.300 69.390 3881.900 ;
        RECT 65.155 3880.230 69.365 3880.300 ;
        RECT 59.155 3873.450 63.365 3873.525 ;
        RECT 57.010 3871.850 63.400 3873.450 ;
        RECT 59.155 3871.780 63.365 3871.850 ;
        RECT 65.200 3865.000 69.410 3865.075 ;
        RECT 57.010 3863.400 69.410 3865.000 ;
        RECT 65.200 3863.330 69.410 3863.400 ;
        RECT 191.280 3753.380 203.560 3758.650 ;
        RECT 175.230 3745.470 187.510 3750.740 ;
        RECT 59.120 3715.280 63.315 3715.395 ;
        RECT 41.440 3713.680 63.315 3715.280 ;
        RECT 59.120 3713.590 63.315 3713.680 ;
        RECT 65.150 3711.780 69.345 3711.850 ;
        RECT 41.440 3710.180 69.500 3711.780 ;
        RECT 65.150 3710.045 69.345 3710.180 ;
        RECT 59.135 3691.250 63.345 3691.340 ;
        RECT 57.010 3689.650 63.430 3691.250 ;
        RECT 59.135 3689.540 63.345 3689.650 ;
        RECT 65.170 3682.800 69.380 3682.865 ;
        RECT 57.010 3681.200 69.390 3682.800 ;
        RECT 65.170 3681.120 69.380 3681.200 ;
        RECT 59.175 3674.350 63.385 3674.390 ;
        RECT 57.010 3672.750 63.385 3674.350 ;
        RECT 59.175 3672.645 63.385 3672.750 ;
        RECT 65.155 3665.900 69.365 3665.975 ;
        RECT 57.010 3664.300 69.390 3665.900 ;
        RECT 3346.930 3664.740 3352.340 3670.230 ;
        RECT 65.155 3664.230 69.365 3664.300 ;
        RECT 59.155 3657.450 63.365 3657.525 ;
        RECT 57.010 3655.850 63.400 3657.450 ;
        RECT 3328.400 3656.650 3333.810 3662.140 ;
        RECT 59.155 3655.780 63.365 3655.850 ;
        RECT 3465.680 3650.280 3469.810 3650.340 ;
        RECT 65.200 3649.000 69.410 3649.075 ;
        RECT 57.010 3647.400 69.410 3649.000 ;
        RECT 3465.680 3648.680 3487.520 3650.280 ;
        RECT 3465.680 3648.625 3469.810 3648.680 ;
        RECT 65.200 3647.330 69.410 3647.400 ;
        RECT 3459.625 3646.780 3463.755 3646.855 ;
        RECT 3459.460 3645.180 3487.520 3646.780 ;
        RECT 3459.625 3645.140 3463.755 3645.180 ;
        RECT 3518.470 3631.490 3522.655 3631.575 ;
        RECT 3516.160 3629.890 3522.770 3631.490 ;
        RECT 3518.470 3629.800 3522.655 3629.890 ;
        RECT 3465.520 3626.250 3469.845 3626.350 ;
        RECT 3465.520 3624.650 3471.950 3626.250 ;
        RECT 3465.520 3624.580 3469.845 3624.650 ;
        RECT 3524.475 3623.040 3528.660 3623.120 ;
        RECT 3516.160 3621.440 3528.830 3623.040 ;
        RECT 3524.475 3621.345 3528.660 3621.440 ;
        RECT 3459.535 3617.800 3463.860 3617.860 ;
        RECT 3459.535 3616.200 3471.950 3617.800 ;
        RECT 3459.535 3616.090 3463.860 3616.200 ;
        RECT 3518.445 3614.590 3522.630 3614.705 ;
        RECT 3516.160 3612.990 3522.740 3614.590 ;
        RECT 3518.445 3612.930 3522.630 3612.990 ;
        RECT 3465.635 3609.350 3469.960 3609.435 ;
        RECT 3465.635 3607.750 3471.950 3609.350 ;
        RECT 3465.635 3607.665 3469.960 3607.750 ;
        RECT 3524.420 3606.140 3528.830 3606.250 ;
        RECT 3516.160 3604.640 3528.830 3606.140 ;
        RECT 3516.160 3604.560 3528.825 3604.640 ;
        RECT 3516.160 3604.540 3528.820 3604.560 ;
        RECT 3459.540 3600.900 3463.865 3600.960 ;
        RECT 3459.540 3599.300 3471.950 3600.900 ;
        RECT 3459.540 3599.190 3463.865 3599.300 ;
        RECT 3518.450 3597.690 3522.630 3597.780 ;
        RECT 3516.000 3596.090 3522.630 3597.690 ;
        RECT 3518.450 3595.980 3522.630 3596.090 ;
        RECT 3465.540 3592.450 3469.865 3592.555 ;
        RECT 3465.540 3590.850 3471.950 3592.450 ;
        RECT 3465.540 3590.785 3469.865 3590.850 ;
        RECT 3524.415 3589.240 3528.600 3589.320 ;
        RECT 3516.000 3587.640 3528.600 3589.240 ;
        RECT 3524.415 3587.545 3528.600 3587.640 ;
        RECT 3459.570 3584.000 3463.895 3584.100 ;
        RECT 3459.570 3582.400 3471.950 3584.000 ;
        RECT 3459.570 3582.330 3463.895 3582.400 ;
        RECT 191.280 3529.380 203.560 3534.650 ;
        RECT 175.230 3521.470 187.510 3526.740 ;
        RECT 59.120 3499.280 63.315 3499.395 ;
        RECT 41.440 3497.680 63.315 3499.280 ;
        RECT 59.120 3497.590 63.315 3497.680 ;
        RECT 65.150 3495.780 69.345 3495.850 ;
        RECT 41.440 3494.180 69.500 3495.780 ;
        RECT 65.150 3494.045 69.345 3494.180 ;
        RECT 59.135 3475.250 63.345 3475.340 ;
        RECT 57.010 3473.650 63.430 3475.250 ;
        RECT 59.135 3473.540 63.345 3473.650 ;
        RECT 65.170 3466.800 69.380 3466.865 ;
        RECT 57.010 3465.200 69.390 3466.800 ;
        RECT 65.170 3465.120 69.380 3465.200 ;
        RECT 59.175 3458.350 63.385 3458.390 ;
        RECT 57.010 3456.750 63.385 3458.350 ;
        RECT 59.175 3456.645 63.385 3456.750 ;
        RECT 65.155 3449.900 69.365 3449.975 ;
        RECT 57.010 3448.300 69.390 3449.900 ;
        RECT 65.155 3448.230 69.365 3448.300 ;
        RECT 59.155 3441.450 63.365 3441.525 ;
        RECT 57.010 3439.850 63.400 3441.450 ;
        RECT 59.155 3439.780 63.365 3439.850 ;
        RECT 3346.930 3439.740 3352.340 3445.230 ;
        RECT 65.200 3433.000 69.410 3433.075 ;
        RECT 57.010 3431.400 69.410 3433.000 ;
        RECT 3328.400 3431.650 3333.810 3437.140 ;
        RECT 65.200 3431.330 69.410 3431.400 ;
        RECT 3465.680 3425.280 3469.810 3425.340 ;
        RECT 3465.680 3423.680 3487.520 3425.280 ;
        RECT 3465.680 3423.625 3469.810 3423.680 ;
        RECT 3459.625 3421.780 3463.755 3421.855 ;
        RECT 3459.460 3420.180 3487.520 3421.780 ;
        RECT 3459.625 3420.140 3463.755 3420.180 ;
        RECT 3518.470 3406.490 3522.655 3406.575 ;
        RECT 3516.160 3404.890 3522.770 3406.490 ;
        RECT 3518.470 3404.800 3522.655 3404.890 ;
        RECT 3465.520 3401.250 3469.845 3401.350 ;
        RECT 3465.520 3399.650 3471.950 3401.250 ;
        RECT 3465.520 3399.580 3469.845 3399.650 ;
        RECT 3524.475 3398.040 3528.660 3398.120 ;
        RECT 3516.160 3396.440 3528.830 3398.040 ;
        RECT 3524.475 3396.345 3528.660 3396.440 ;
        RECT 3459.535 3392.800 3463.860 3392.860 ;
        RECT 3459.535 3391.200 3471.950 3392.800 ;
        RECT 3459.535 3391.090 3463.860 3391.200 ;
        RECT 3518.445 3389.590 3522.630 3389.705 ;
        RECT 3516.160 3387.990 3522.740 3389.590 ;
        RECT 3518.445 3387.930 3522.630 3387.990 ;
        RECT 3465.635 3384.350 3469.960 3384.435 ;
        RECT 3465.635 3382.750 3471.950 3384.350 ;
        RECT 3465.635 3382.665 3469.960 3382.750 ;
        RECT 3524.420 3381.140 3528.830 3381.250 ;
        RECT 3516.160 3379.640 3528.830 3381.140 ;
        RECT 3516.160 3379.560 3528.825 3379.640 ;
        RECT 3516.160 3379.540 3528.820 3379.560 ;
        RECT 3459.540 3375.900 3463.865 3375.960 ;
        RECT 3459.540 3374.300 3471.950 3375.900 ;
        RECT 3459.540 3374.190 3463.865 3374.300 ;
        RECT 3518.450 3372.690 3522.630 3372.780 ;
        RECT 3516.000 3371.090 3522.630 3372.690 ;
        RECT 3518.450 3370.980 3522.630 3371.090 ;
        RECT 3465.540 3367.450 3469.865 3367.555 ;
        RECT 3465.540 3365.850 3471.950 3367.450 ;
        RECT 3465.540 3365.785 3469.865 3365.850 ;
        RECT 3524.415 3364.240 3528.600 3364.320 ;
        RECT 3516.000 3362.640 3528.600 3364.240 ;
        RECT 3524.415 3362.545 3528.600 3362.640 ;
        RECT 3459.570 3359.000 3463.895 3359.100 ;
        RECT 3459.570 3357.400 3471.950 3359.000 ;
        RECT 3459.570 3357.330 3463.895 3357.400 ;
        RECT 191.280 3313.380 203.560 3318.650 ;
        RECT 175.230 3305.470 187.510 3310.740 ;
        RECT 59.120 3283.280 63.315 3283.395 ;
        RECT 41.440 3281.680 63.315 3283.280 ;
        RECT 59.120 3281.590 63.315 3281.680 ;
        RECT 65.150 3279.780 69.345 3279.850 ;
        RECT 41.440 3278.180 69.500 3279.780 ;
        RECT 65.150 3278.045 69.345 3278.180 ;
        RECT 59.135 3259.250 63.345 3259.340 ;
        RECT 57.010 3257.650 63.430 3259.250 ;
        RECT 59.135 3257.540 63.345 3257.650 ;
        RECT 65.170 3250.800 69.380 3250.865 ;
        RECT 57.010 3249.200 69.390 3250.800 ;
        RECT 65.170 3249.120 69.380 3249.200 ;
        RECT 59.175 3242.350 63.385 3242.390 ;
        RECT 57.010 3240.750 63.385 3242.350 ;
        RECT 59.175 3240.645 63.385 3240.750 ;
        RECT 65.155 3233.900 69.365 3233.975 ;
        RECT 57.010 3232.300 69.390 3233.900 ;
        RECT 65.155 3232.230 69.365 3232.300 ;
        RECT 59.155 3225.450 63.365 3225.525 ;
        RECT 57.010 3223.850 63.400 3225.450 ;
        RECT 59.155 3223.780 63.365 3223.850 ;
        RECT 65.200 3217.000 69.410 3217.075 ;
        RECT 57.010 3215.400 69.410 3217.000 ;
        RECT 65.200 3215.330 69.410 3215.400 ;
        RECT 3346.930 3213.740 3352.340 3219.230 ;
        RECT 3328.400 3205.650 3333.810 3211.140 ;
        RECT 3465.680 3199.280 3469.810 3199.340 ;
        RECT 3465.680 3197.680 3487.520 3199.280 ;
        RECT 3465.680 3197.625 3469.810 3197.680 ;
        RECT 3459.625 3195.780 3463.755 3195.855 ;
        RECT 3459.460 3194.180 3487.520 3195.780 ;
        RECT 3459.625 3194.140 3463.755 3194.180 ;
        RECT 3518.470 3180.490 3522.655 3180.575 ;
        RECT 3516.160 3178.890 3522.770 3180.490 ;
        RECT 3518.470 3178.800 3522.655 3178.890 ;
        RECT 3465.520 3175.250 3469.845 3175.350 ;
        RECT 3465.520 3173.650 3471.950 3175.250 ;
        RECT 3465.520 3173.580 3469.845 3173.650 ;
        RECT 3524.475 3172.040 3528.660 3172.120 ;
        RECT 3516.160 3170.440 3528.830 3172.040 ;
        RECT 3524.475 3170.345 3528.660 3170.440 ;
        RECT 3459.535 3166.800 3463.860 3166.860 ;
        RECT 3459.535 3165.200 3471.950 3166.800 ;
        RECT 3459.535 3165.090 3463.860 3165.200 ;
        RECT 3518.445 3163.590 3522.630 3163.705 ;
        RECT 3516.160 3161.990 3522.740 3163.590 ;
        RECT 3518.445 3161.930 3522.630 3161.990 ;
        RECT 3465.635 3158.350 3469.960 3158.435 ;
        RECT 3465.635 3156.750 3471.950 3158.350 ;
        RECT 3465.635 3156.665 3469.960 3156.750 ;
        RECT 3524.420 3155.140 3528.830 3155.250 ;
        RECT 3516.160 3153.640 3528.830 3155.140 ;
        RECT 3516.160 3153.560 3528.825 3153.640 ;
        RECT 3516.160 3153.540 3528.820 3153.560 ;
        RECT 3459.540 3149.900 3463.865 3149.960 ;
        RECT 3459.540 3148.300 3471.950 3149.900 ;
        RECT 3459.540 3148.190 3463.865 3148.300 ;
        RECT 3518.450 3146.690 3522.630 3146.780 ;
        RECT 3516.000 3145.090 3522.630 3146.690 ;
        RECT 3518.450 3144.980 3522.630 3145.090 ;
        RECT 3465.540 3141.450 3469.865 3141.555 ;
        RECT 3465.540 3139.850 3471.950 3141.450 ;
        RECT 3465.540 3139.785 3469.865 3139.850 ;
        RECT 3524.415 3138.240 3528.600 3138.320 ;
        RECT 3516.000 3136.640 3528.600 3138.240 ;
        RECT 3524.415 3136.545 3528.600 3136.640 ;
        RECT 3459.570 3133.000 3463.895 3133.100 ;
        RECT 3459.570 3131.400 3471.950 3133.000 ;
        RECT 3459.570 3131.330 3463.895 3131.400 ;
        RECT 191.280 3097.380 203.560 3102.650 ;
        RECT 175.230 3089.470 187.510 3094.740 ;
        RECT 59.120 3067.280 63.315 3067.395 ;
        RECT 41.440 3065.680 63.315 3067.280 ;
        RECT 59.120 3065.590 63.315 3065.680 ;
        RECT 65.150 3063.780 69.345 3063.850 ;
        RECT 41.440 3062.180 69.500 3063.780 ;
        RECT 65.150 3062.045 69.345 3062.180 ;
        RECT 59.135 3043.250 63.345 3043.340 ;
        RECT 57.010 3041.650 63.430 3043.250 ;
        RECT 59.135 3041.540 63.345 3041.650 ;
        RECT 65.170 3034.800 69.380 3034.865 ;
        RECT 57.010 3033.200 69.390 3034.800 ;
        RECT 65.170 3033.120 69.380 3033.200 ;
        RECT 59.175 3026.350 63.385 3026.390 ;
        RECT 57.010 3024.750 63.385 3026.350 ;
        RECT 59.175 3024.645 63.385 3024.750 ;
        RECT 65.155 3017.900 69.365 3017.975 ;
        RECT 57.010 3016.300 69.390 3017.900 ;
        RECT 65.155 3016.230 69.365 3016.300 ;
        RECT 59.155 3009.450 63.365 3009.525 ;
        RECT 57.010 3007.850 63.400 3009.450 ;
        RECT 59.155 3007.780 63.365 3007.850 ;
        RECT 65.200 3001.000 69.410 3001.075 ;
        RECT 57.010 2999.400 69.410 3001.000 ;
        RECT 65.200 2999.330 69.410 2999.400 ;
        RECT 3346.930 2988.740 3352.340 2994.230 ;
        RECT 3328.400 2980.650 3333.810 2986.140 ;
        RECT 3465.680 2974.280 3469.810 2974.340 ;
        RECT 3465.680 2972.680 3487.520 2974.280 ;
        RECT 3465.680 2972.625 3469.810 2972.680 ;
        RECT 3459.625 2970.780 3463.755 2970.855 ;
        RECT 3459.460 2969.180 3487.520 2970.780 ;
        RECT 3459.625 2969.140 3463.755 2969.180 ;
        RECT 3518.470 2955.490 3522.655 2955.575 ;
        RECT 3516.160 2953.890 3522.770 2955.490 ;
        RECT 3518.470 2953.800 3522.655 2953.890 ;
        RECT 3465.520 2950.250 3469.845 2950.350 ;
        RECT 3465.520 2948.650 3471.950 2950.250 ;
        RECT 3465.520 2948.580 3469.845 2948.650 ;
        RECT 3524.475 2947.040 3528.660 2947.120 ;
        RECT 3516.160 2945.440 3528.830 2947.040 ;
        RECT 3524.475 2945.345 3528.660 2945.440 ;
        RECT 3459.535 2941.800 3463.860 2941.860 ;
        RECT 3459.535 2940.200 3471.950 2941.800 ;
        RECT 3459.535 2940.090 3463.860 2940.200 ;
        RECT 3518.445 2938.590 3522.630 2938.705 ;
        RECT 3516.160 2936.990 3522.740 2938.590 ;
        RECT 3518.445 2936.930 3522.630 2936.990 ;
        RECT 3465.635 2933.350 3469.960 2933.435 ;
        RECT 3465.635 2931.750 3471.950 2933.350 ;
        RECT 3465.635 2931.665 3469.960 2931.750 ;
        RECT 3524.420 2930.140 3528.830 2930.250 ;
        RECT 3516.160 2928.640 3528.830 2930.140 ;
        RECT 3516.160 2928.560 3528.825 2928.640 ;
        RECT 3516.160 2928.540 3528.820 2928.560 ;
        RECT 3459.540 2924.900 3463.865 2924.960 ;
        RECT 3459.540 2923.300 3471.950 2924.900 ;
        RECT 3459.540 2923.190 3463.865 2923.300 ;
        RECT 3518.450 2921.690 3522.630 2921.780 ;
        RECT 3516.000 2920.090 3522.630 2921.690 ;
        RECT 3518.450 2919.980 3522.630 2920.090 ;
        RECT 3465.540 2916.450 3469.865 2916.555 ;
        RECT 3465.540 2914.850 3471.950 2916.450 ;
        RECT 3465.540 2914.785 3469.865 2914.850 ;
        RECT 3524.415 2913.240 3528.600 2913.320 ;
        RECT 3516.000 2911.640 3528.600 2913.240 ;
        RECT 3524.415 2911.545 3528.600 2911.640 ;
        RECT 3459.570 2908.000 3463.895 2908.100 ;
        RECT 3459.570 2906.400 3471.950 2908.000 ;
        RECT 3459.570 2906.330 3463.895 2906.400 ;
        RECT 191.280 2886.680 203.560 2891.950 ;
        RECT 175.230 2878.770 187.510 2884.040 ;
        RECT 59.120 2851.280 63.315 2851.395 ;
        RECT 41.440 2849.680 63.315 2851.280 ;
        RECT 59.120 2849.590 63.315 2849.680 ;
        RECT 65.150 2847.780 69.345 2847.850 ;
        RECT 41.440 2846.180 69.500 2847.780 ;
        RECT 65.150 2846.045 69.345 2846.180 ;
        RECT 59.135 2827.250 63.345 2827.340 ;
        RECT 57.010 2825.650 63.430 2827.250 ;
        RECT 59.135 2825.540 63.345 2825.650 ;
        RECT 65.170 2818.800 69.380 2818.865 ;
        RECT 57.010 2817.200 69.390 2818.800 ;
        RECT 65.170 2817.120 69.380 2817.200 ;
        RECT 59.175 2810.350 63.385 2810.390 ;
        RECT 57.010 2808.750 63.385 2810.350 ;
        RECT 59.175 2808.645 63.385 2808.750 ;
        RECT 65.155 2801.900 69.365 2801.975 ;
        RECT 57.010 2800.300 69.390 2801.900 ;
        RECT 65.155 2800.230 69.365 2800.300 ;
        RECT 59.155 2793.450 63.365 2793.525 ;
        RECT 57.010 2791.850 63.400 2793.450 ;
        RECT 59.155 2791.780 63.365 2791.850 ;
        RECT 65.200 2785.000 69.410 2785.075 ;
        RECT 57.010 2783.400 69.410 2785.000 ;
        RECT 65.200 2783.330 69.410 2783.400 ;
        RECT 3346.930 2762.740 3352.340 2768.230 ;
        RECT 3328.400 2754.650 3333.810 2760.140 ;
        RECT 3465.680 2748.280 3469.810 2748.340 ;
        RECT 3465.680 2746.680 3487.520 2748.280 ;
        RECT 3465.680 2746.625 3469.810 2746.680 ;
        RECT 3459.625 2744.780 3463.755 2744.855 ;
        RECT 3459.460 2743.180 3487.520 2744.780 ;
        RECT 3459.625 2743.140 3463.755 2743.180 ;
        RECT 3518.470 2729.490 3522.655 2729.575 ;
        RECT 3516.160 2727.890 3522.770 2729.490 ;
        RECT 3518.470 2727.800 3522.655 2727.890 ;
        RECT 3465.520 2724.250 3469.845 2724.350 ;
        RECT 3465.520 2722.650 3471.950 2724.250 ;
        RECT 3465.520 2722.580 3469.845 2722.650 ;
        RECT 3524.475 2721.040 3528.660 2721.120 ;
        RECT 3516.160 2719.440 3528.830 2721.040 ;
        RECT 3524.475 2719.345 3528.660 2719.440 ;
        RECT 3459.535 2715.800 3463.860 2715.860 ;
        RECT 3459.535 2714.200 3471.950 2715.800 ;
        RECT 3459.535 2714.090 3463.860 2714.200 ;
        RECT 3518.445 2712.590 3522.630 2712.705 ;
        RECT 3516.160 2710.990 3522.740 2712.590 ;
        RECT 3518.445 2710.930 3522.630 2710.990 ;
        RECT 3465.635 2707.350 3469.960 2707.435 ;
        RECT 3465.635 2705.750 3471.950 2707.350 ;
        RECT 3465.635 2705.665 3469.960 2705.750 ;
        RECT 3524.420 2704.140 3528.830 2704.250 ;
        RECT 3516.160 2702.640 3528.830 2704.140 ;
        RECT 3516.160 2702.560 3528.825 2702.640 ;
        RECT 3516.160 2702.540 3528.820 2702.560 ;
        RECT 3459.540 2698.900 3463.865 2698.960 ;
        RECT 3459.540 2697.300 3471.950 2698.900 ;
        RECT 3459.540 2697.190 3463.865 2697.300 ;
        RECT 3518.450 2695.690 3522.630 2695.780 ;
        RECT 3516.000 2694.090 3522.630 2695.690 ;
        RECT 3518.450 2693.980 3522.630 2694.090 ;
        RECT 3465.540 2690.450 3469.865 2690.555 ;
        RECT 3465.540 2688.850 3471.950 2690.450 ;
        RECT 3465.540 2688.785 3469.865 2688.850 ;
        RECT 3524.415 2687.240 3528.600 2687.320 ;
        RECT 3516.000 2685.640 3528.600 2687.240 ;
        RECT 3524.415 2685.545 3528.600 2685.640 ;
        RECT 3459.570 2682.000 3463.895 2682.100 ;
        RECT 3459.570 2680.400 3471.950 2682.000 ;
        RECT 3459.570 2680.330 3463.895 2680.400 ;
        RECT 191.280 2665.380 203.560 2670.650 ;
        RECT 175.230 2657.470 187.510 2662.740 ;
        RECT 59.120 2635.280 63.315 2635.395 ;
        RECT 41.440 2633.680 63.315 2635.280 ;
        RECT 59.120 2633.590 63.315 2633.680 ;
        RECT 65.150 2631.780 69.345 2631.850 ;
        RECT 41.440 2630.180 69.500 2631.780 ;
        RECT 65.150 2630.045 69.345 2630.180 ;
        RECT 59.135 2611.250 63.345 2611.340 ;
        RECT 57.010 2609.650 63.430 2611.250 ;
        RECT 59.135 2609.540 63.345 2609.650 ;
        RECT 65.170 2602.800 69.380 2602.865 ;
        RECT 57.010 2601.200 69.390 2602.800 ;
        RECT 65.170 2601.120 69.380 2601.200 ;
        RECT 59.175 2594.350 63.385 2594.390 ;
        RECT 57.010 2592.750 63.385 2594.350 ;
        RECT 59.175 2592.645 63.385 2592.750 ;
        RECT 65.155 2585.900 69.365 2585.975 ;
        RECT 57.010 2584.300 69.390 2585.900 ;
        RECT 65.155 2584.230 69.365 2584.300 ;
        RECT 59.155 2577.450 63.365 2577.525 ;
        RECT 57.010 2575.850 63.400 2577.450 ;
        RECT 59.155 2575.780 63.365 2575.850 ;
        RECT 65.200 2569.000 69.410 2569.075 ;
        RECT 57.010 2567.400 69.410 2569.000 ;
        RECT 65.200 2567.330 69.410 2567.400 ;
        RECT 3346.930 2537.740 3352.340 2543.230 ;
        RECT 3328.400 2529.650 3333.810 2535.140 ;
        RECT 3465.680 2523.280 3469.810 2523.340 ;
        RECT 3465.680 2521.680 3487.520 2523.280 ;
        RECT 3465.680 2521.625 3469.810 2521.680 ;
        RECT 3459.625 2519.780 3463.755 2519.855 ;
        RECT 3459.460 2518.180 3487.520 2519.780 ;
        RECT 3459.625 2518.140 3463.755 2518.180 ;
        RECT 3518.470 2504.490 3522.655 2504.575 ;
        RECT 3516.160 2502.890 3522.770 2504.490 ;
        RECT 3518.470 2502.800 3522.655 2502.890 ;
        RECT 3465.520 2499.250 3469.845 2499.350 ;
        RECT 3465.520 2497.650 3471.950 2499.250 ;
        RECT 3465.520 2497.580 3469.845 2497.650 ;
        RECT 3524.475 2496.040 3528.660 2496.120 ;
        RECT 3516.160 2494.440 3528.830 2496.040 ;
        RECT 3524.475 2494.345 3528.660 2494.440 ;
        RECT 3459.535 2490.800 3463.860 2490.860 ;
        RECT 3459.535 2489.200 3471.950 2490.800 ;
        RECT 3459.535 2489.090 3463.860 2489.200 ;
        RECT 3518.445 2487.590 3522.630 2487.705 ;
        RECT 3516.160 2485.990 3522.740 2487.590 ;
        RECT 3518.445 2485.930 3522.630 2485.990 ;
        RECT 3465.635 2482.350 3469.960 2482.435 ;
        RECT 3465.635 2480.750 3471.950 2482.350 ;
        RECT 3465.635 2480.665 3469.960 2480.750 ;
        RECT 3524.420 2479.140 3528.830 2479.250 ;
        RECT 3516.160 2477.640 3528.830 2479.140 ;
        RECT 3516.160 2477.560 3528.825 2477.640 ;
        RECT 3516.160 2477.540 3528.820 2477.560 ;
        RECT 3459.540 2473.900 3463.865 2473.960 ;
        RECT 3459.540 2472.300 3471.950 2473.900 ;
        RECT 3459.540 2472.190 3463.865 2472.300 ;
        RECT 3518.450 2470.690 3522.630 2470.780 ;
        RECT 3516.000 2469.090 3522.630 2470.690 ;
        RECT 3518.450 2468.980 3522.630 2469.090 ;
        RECT 3465.540 2465.450 3469.865 2465.555 ;
        RECT 3465.540 2463.850 3471.950 2465.450 ;
        RECT 3465.540 2463.785 3469.865 2463.850 ;
        RECT 3524.415 2462.240 3528.600 2462.320 ;
        RECT 3516.000 2460.640 3528.600 2462.240 ;
        RECT 3524.415 2460.545 3528.600 2460.640 ;
        RECT 3459.570 2457.000 3463.895 2457.100 ;
        RECT 3459.570 2455.400 3471.950 2457.000 ;
        RECT 3459.570 2455.330 3463.895 2455.400 ;
        RECT 3346.930 2317.740 3352.340 2323.230 ;
        RECT 3328.400 2309.650 3333.810 2315.140 ;
        RECT 3465.680 2303.280 3469.810 2303.340 ;
        RECT 3465.680 2301.680 3487.520 2303.280 ;
        RECT 3465.680 2301.625 3469.810 2301.680 ;
        RECT 3459.625 2299.780 3463.755 2299.855 ;
        RECT 3459.460 2298.180 3487.520 2299.780 ;
        RECT 3459.625 2298.140 3463.755 2298.180 ;
        RECT 3518.470 2284.490 3522.655 2284.575 ;
        RECT 3516.160 2282.890 3522.770 2284.490 ;
        RECT 3518.470 2282.800 3522.655 2282.890 ;
        RECT 3465.520 2279.250 3469.845 2279.350 ;
        RECT 3465.520 2277.650 3471.950 2279.250 ;
        RECT 3465.520 2277.580 3469.845 2277.650 ;
        RECT 3524.475 2276.040 3528.660 2276.120 ;
        RECT 3516.160 2274.440 3528.830 2276.040 ;
        RECT 3524.475 2274.345 3528.660 2274.440 ;
        RECT 3459.535 2270.800 3463.860 2270.860 ;
        RECT 3459.535 2269.200 3471.950 2270.800 ;
        RECT 3459.535 2269.090 3463.860 2269.200 ;
        RECT 3518.445 2267.590 3522.630 2267.705 ;
        RECT 3516.160 2265.990 3522.740 2267.590 ;
        RECT 3518.445 2265.930 3522.630 2265.990 ;
        RECT 3465.635 2262.350 3469.960 2262.435 ;
        RECT 3465.635 2260.750 3471.950 2262.350 ;
        RECT 3465.635 2260.665 3469.960 2260.750 ;
        RECT 3524.420 2259.140 3528.830 2259.250 ;
        RECT 3516.160 2257.640 3528.830 2259.140 ;
        RECT 3516.160 2257.560 3528.825 2257.640 ;
        RECT 3516.160 2257.540 3528.820 2257.560 ;
        RECT 3459.540 2253.900 3463.865 2253.960 ;
        RECT 3459.540 2252.300 3471.950 2253.900 ;
        RECT 3459.540 2252.190 3463.865 2252.300 ;
        RECT 3518.450 2250.690 3522.630 2250.780 ;
        RECT 3516.000 2249.090 3522.630 2250.690 ;
        RECT 3518.450 2248.980 3522.630 2249.090 ;
        RECT 3465.540 2245.450 3469.865 2245.555 ;
        RECT 3465.540 2243.850 3471.950 2245.450 ;
        RECT 3465.540 2243.785 3469.865 2243.850 ;
        RECT 3524.415 2242.240 3528.600 2242.320 ;
        RECT 3516.000 2240.640 3528.600 2242.240 ;
        RECT 3524.415 2240.545 3528.600 2240.640 ;
        RECT 3459.570 2237.000 3463.895 2237.100 ;
        RECT 3459.570 2235.400 3471.950 2237.000 ;
        RECT 3459.570 2235.330 3463.895 2235.400 ;
        RECT 191.280 2027.380 203.560 2032.650 ;
        RECT 175.230 2019.470 187.510 2024.740 ;
        RECT 59.120 1997.280 63.315 1997.395 ;
        RECT 41.440 1995.680 63.315 1997.280 ;
        RECT 59.120 1995.590 63.315 1995.680 ;
        RECT 65.150 1993.780 69.345 1993.850 ;
        RECT 41.440 1992.180 69.500 1993.780 ;
        RECT 65.150 1992.045 69.345 1992.180 ;
        RECT 59.135 1973.250 63.345 1973.340 ;
        RECT 57.010 1971.650 63.430 1973.250 ;
        RECT 59.135 1971.540 63.345 1971.650 ;
        RECT 65.170 1964.800 69.380 1964.865 ;
        RECT 57.010 1963.200 69.390 1964.800 ;
        RECT 65.170 1963.120 69.380 1963.200 ;
        RECT 59.175 1956.350 63.385 1956.390 ;
        RECT 57.010 1954.750 63.385 1956.350 ;
        RECT 59.175 1954.645 63.385 1954.750 ;
        RECT 65.155 1947.900 69.365 1947.975 ;
        RECT 57.010 1946.300 69.390 1947.900 ;
        RECT 65.155 1946.230 69.365 1946.300 ;
        RECT 59.155 1939.450 63.365 1939.525 ;
        RECT 57.010 1937.850 63.400 1939.450 ;
        RECT 59.155 1937.780 63.365 1937.850 ;
        RECT 65.200 1931.000 69.410 1931.075 ;
        RECT 57.010 1929.400 69.410 1931.000 ;
        RECT 65.200 1929.330 69.410 1929.400 ;
        RECT 3346.930 1876.740 3352.340 1882.230 ;
        RECT 3328.400 1868.650 3333.810 1874.140 ;
        RECT 3465.680 1862.280 3469.810 1862.340 ;
        RECT 3465.680 1860.680 3487.520 1862.280 ;
        RECT 3465.680 1860.625 3469.810 1860.680 ;
        RECT 3459.625 1858.780 3463.755 1858.855 ;
        RECT 3459.460 1857.180 3487.520 1858.780 ;
        RECT 3459.625 1857.140 3463.755 1857.180 ;
        RECT 3518.470 1843.490 3522.655 1843.575 ;
        RECT 3516.160 1841.890 3522.770 1843.490 ;
        RECT 3518.470 1841.800 3522.655 1841.890 ;
        RECT 3465.520 1838.250 3469.845 1838.350 ;
        RECT 3465.520 1836.650 3471.950 1838.250 ;
        RECT 3465.520 1836.580 3469.845 1836.650 ;
        RECT 3524.475 1835.040 3528.660 1835.120 ;
        RECT 3516.160 1833.440 3528.830 1835.040 ;
        RECT 3524.475 1833.345 3528.660 1833.440 ;
        RECT 3459.535 1829.800 3463.860 1829.860 ;
        RECT 3459.535 1828.200 3471.950 1829.800 ;
        RECT 3459.535 1828.090 3463.860 1828.200 ;
        RECT 3518.445 1826.590 3522.630 1826.705 ;
        RECT 3516.160 1824.990 3522.740 1826.590 ;
        RECT 3518.445 1824.930 3522.630 1824.990 ;
        RECT 3465.635 1821.350 3469.960 1821.435 ;
        RECT 3465.635 1819.750 3471.950 1821.350 ;
        RECT 3465.635 1819.665 3469.960 1819.750 ;
        RECT 3524.420 1818.140 3528.830 1818.250 ;
        RECT 191.280 1811.380 203.560 1816.650 ;
        RECT 3516.160 1816.640 3528.830 1818.140 ;
        RECT 3516.160 1816.560 3528.825 1816.640 ;
        RECT 3516.160 1816.540 3528.820 1816.560 ;
        RECT 3459.540 1812.900 3463.865 1812.960 ;
        RECT 3459.540 1811.300 3471.950 1812.900 ;
        RECT 3459.540 1811.190 3463.865 1811.300 ;
        RECT 3518.450 1809.690 3522.630 1809.780 ;
        RECT 175.230 1803.470 187.510 1808.740 ;
        RECT 3516.000 1808.090 3522.630 1809.690 ;
        RECT 3518.450 1807.980 3522.630 1808.090 ;
        RECT 3465.540 1804.450 3469.865 1804.555 ;
        RECT 3465.540 1802.850 3471.950 1804.450 ;
        RECT 3465.540 1802.785 3469.865 1802.850 ;
        RECT 3524.415 1801.240 3528.600 1801.320 ;
        RECT 3516.000 1799.640 3528.600 1801.240 ;
        RECT 3524.415 1799.545 3528.600 1799.640 ;
        RECT 3459.570 1796.000 3463.895 1796.100 ;
        RECT 3459.570 1794.400 3471.950 1796.000 ;
        RECT 3459.570 1794.330 3463.895 1794.400 ;
        RECT 59.120 1781.280 63.315 1781.395 ;
        RECT 41.440 1779.680 63.315 1781.280 ;
        RECT 59.120 1779.590 63.315 1779.680 ;
        RECT 65.150 1777.780 69.345 1777.850 ;
        RECT 41.440 1776.180 69.500 1777.780 ;
        RECT 65.150 1776.045 69.345 1776.180 ;
        RECT 59.135 1757.250 63.345 1757.340 ;
        RECT 57.010 1755.650 63.430 1757.250 ;
        RECT 59.135 1755.540 63.345 1755.650 ;
        RECT 65.170 1748.800 69.380 1748.865 ;
        RECT 57.010 1747.200 69.390 1748.800 ;
        RECT 65.170 1747.120 69.380 1747.200 ;
        RECT 59.175 1740.350 63.385 1740.390 ;
        RECT 57.010 1738.750 63.385 1740.350 ;
        RECT 59.175 1738.645 63.385 1738.750 ;
        RECT 65.155 1731.900 69.365 1731.975 ;
        RECT 57.010 1730.300 69.390 1731.900 ;
        RECT 65.155 1730.230 69.365 1730.300 ;
        RECT 59.155 1723.450 63.365 1723.525 ;
        RECT 57.010 1721.850 63.400 1723.450 ;
        RECT 59.155 1721.780 63.365 1721.850 ;
        RECT 65.200 1715.000 69.410 1715.075 ;
        RECT 57.010 1713.400 69.410 1715.000 ;
        RECT 65.200 1713.330 69.410 1713.400 ;
        RECT 3346.930 1650.740 3352.340 1656.230 ;
        RECT 3328.400 1642.650 3333.810 1648.140 ;
        RECT 3465.680 1636.280 3469.810 1636.340 ;
        RECT 3465.680 1634.680 3487.520 1636.280 ;
        RECT 3465.680 1634.625 3469.810 1634.680 ;
        RECT 3459.625 1632.780 3463.755 1632.855 ;
        RECT 3459.460 1631.180 3487.520 1632.780 ;
        RECT 3459.625 1631.140 3463.755 1631.180 ;
        RECT 3518.470 1617.490 3522.655 1617.575 ;
        RECT 3516.160 1615.890 3522.770 1617.490 ;
        RECT 3518.470 1615.800 3522.655 1615.890 ;
        RECT 3465.520 1612.250 3469.845 1612.350 ;
        RECT 3465.520 1610.650 3471.950 1612.250 ;
        RECT 3465.520 1610.580 3469.845 1610.650 ;
        RECT 3524.475 1609.040 3528.660 1609.120 ;
        RECT 3516.160 1607.440 3528.830 1609.040 ;
        RECT 3524.475 1607.345 3528.660 1607.440 ;
        RECT 191.280 1600.380 203.560 1605.650 ;
        RECT 3459.535 1603.800 3463.860 1603.860 ;
        RECT 3459.535 1602.200 3471.950 1603.800 ;
        RECT 3459.535 1602.090 3463.860 1602.200 ;
        RECT 3518.445 1600.590 3522.630 1600.705 ;
        RECT 3516.160 1598.990 3522.740 1600.590 ;
        RECT 3518.445 1598.930 3522.630 1598.990 ;
        RECT 175.230 1592.470 187.510 1597.740 ;
        RECT 3465.635 1595.350 3469.960 1595.435 ;
        RECT 3465.635 1593.750 3471.950 1595.350 ;
        RECT 3465.635 1593.665 3469.960 1593.750 ;
        RECT 3524.420 1592.140 3528.830 1592.250 ;
        RECT 3516.160 1590.640 3528.830 1592.140 ;
        RECT 3516.160 1590.560 3528.825 1590.640 ;
        RECT 3516.160 1590.540 3528.820 1590.560 ;
        RECT 3459.540 1586.900 3463.865 1586.960 ;
        RECT 3459.540 1585.300 3471.950 1586.900 ;
        RECT 3459.540 1585.190 3463.865 1585.300 ;
        RECT 3518.450 1583.690 3522.630 1583.780 ;
        RECT 3516.000 1582.090 3522.630 1583.690 ;
        RECT 3518.450 1581.980 3522.630 1582.090 ;
        RECT 3465.540 1578.450 3469.865 1578.555 ;
        RECT 3465.540 1576.850 3471.950 1578.450 ;
        RECT 3465.540 1576.785 3469.865 1576.850 ;
        RECT 3524.415 1575.240 3528.600 1575.320 ;
        RECT 3516.000 1573.640 3528.600 1575.240 ;
        RECT 3524.415 1573.545 3528.600 1573.640 ;
        RECT 3459.570 1570.000 3463.895 1570.100 ;
        RECT 3459.570 1568.400 3471.950 1570.000 ;
        RECT 3459.570 1568.330 3463.895 1568.400 ;
        RECT 59.120 1565.280 63.315 1565.395 ;
        RECT 41.440 1563.680 63.315 1565.280 ;
        RECT 59.120 1563.590 63.315 1563.680 ;
        RECT 65.150 1561.780 69.345 1561.850 ;
        RECT 41.440 1560.180 69.500 1561.780 ;
        RECT 65.150 1560.045 69.345 1560.180 ;
        RECT 59.135 1541.250 63.345 1541.340 ;
        RECT 57.010 1539.650 63.430 1541.250 ;
        RECT 59.135 1539.540 63.345 1539.650 ;
        RECT 65.170 1532.800 69.380 1532.865 ;
        RECT 57.010 1531.200 69.390 1532.800 ;
        RECT 65.170 1531.120 69.380 1531.200 ;
        RECT 59.175 1524.350 63.385 1524.390 ;
        RECT 57.010 1522.750 63.385 1524.350 ;
        RECT 59.175 1522.645 63.385 1522.750 ;
        RECT 65.155 1515.900 69.365 1515.975 ;
        RECT 57.010 1514.300 69.390 1515.900 ;
        RECT 65.155 1514.230 69.365 1514.300 ;
        RECT 59.155 1507.450 63.365 1507.525 ;
        RECT 57.010 1505.850 63.400 1507.450 ;
        RECT 59.155 1505.780 63.365 1505.850 ;
        RECT 65.200 1499.000 69.410 1499.075 ;
        RECT 57.010 1497.400 69.410 1499.000 ;
        RECT 65.200 1497.330 69.410 1497.400 ;
        RECT 3346.930 1425.740 3352.340 1431.230 ;
        RECT 3328.400 1417.650 3333.810 1423.140 ;
        RECT 3465.680 1411.280 3469.810 1411.340 ;
        RECT 3465.680 1409.680 3487.520 1411.280 ;
        RECT 3465.680 1409.625 3469.810 1409.680 ;
        RECT 3459.625 1407.780 3463.755 1407.855 ;
        RECT 3459.460 1406.180 3487.520 1407.780 ;
        RECT 3459.625 1406.140 3463.755 1406.180 ;
        RECT 3518.470 1392.490 3522.655 1392.575 ;
        RECT 3516.160 1390.890 3522.770 1392.490 ;
        RECT 3518.470 1390.800 3522.655 1390.890 ;
        RECT 3465.520 1387.250 3469.845 1387.350 ;
        RECT 3465.520 1385.650 3471.950 1387.250 ;
        RECT 3465.520 1385.580 3469.845 1385.650 ;
        RECT 191.280 1379.380 203.560 1384.650 ;
        RECT 3524.475 1384.040 3528.660 1384.120 ;
        RECT 3516.160 1382.440 3528.830 1384.040 ;
        RECT 3524.475 1382.345 3528.660 1382.440 ;
        RECT 3459.535 1378.800 3463.860 1378.860 ;
        RECT 3459.535 1377.200 3471.950 1378.800 ;
        RECT 3459.535 1377.090 3463.860 1377.200 ;
        RECT 175.230 1371.470 187.510 1376.740 ;
        RECT 3518.445 1375.590 3522.630 1375.705 ;
        RECT 3516.160 1373.990 3522.740 1375.590 ;
        RECT 3518.445 1373.930 3522.630 1373.990 ;
        RECT 3465.635 1370.350 3469.960 1370.435 ;
        RECT 3465.635 1368.750 3471.950 1370.350 ;
        RECT 3465.635 1368.665 3469.960 1368.750 ;
        RECT 3524.420 1367.140 3528.830 1367.250 ;
        RECT 3516.160 1365.640 3528.830 1367.140 ;
        RECT 3516.160 1365.560 3528.825 1365.640 ;
        RECT 3516.160 1365.540 3528.820 1365.560 ;
        RECT 3459.540 1361.900 3463.865 1361.960 ;
        RECT 3459.540 1360.300 3471.950 1361.900 ;
        RECT 3459.540 1360.190 3463.865 1360.300 ;
        RECT 3518.450 1358.690 3522.630 1358.780 ;
        RECT 3516.000 1357.090 3522.630 1358.690 ;
        RECT 3518.450 1356.980 3522.630 1357.090 ;
        RECT 3465.540 1353.450 3469.865 1353.555 ;
        RECT 3465.540 1351.850 3471.950 1353.450 ;
        RECT 3465.540 1351.785 3469.865 1351.850 ;
        RECT 3524.415 1350.240 3528.600 1350.320 ;
        RECT 59.120 1349.280 63.315 1349.395 ;
        RECT 41.440 1347.680 63.315 1349.280 ;
        RECT 3516.000 1348.640 3528.600 1350.240 ;
        RECT 3524.415 1348.545 3528.600 1348.640 ;
        RECT 59.120 1347.590 63.315 1347.680 ;
        RECT 65.150 1345.780 69.345 1345.850 ;
        RECT 41.440 1344.180 69.500 1345.780 ;
        RECT 3459.570 1345.000 3463.895 1345.100 ;
        RECT 65.150 1344.045 69.345 1344.180 ;
        RECT 3459.570 1343.400 3471.950 1345.000 ;
        RECT 3459.570 1343.330 3463.895 1343.400 ;
        RECT 59.135 1325.250 63.345 1325.340 ;
        RECT 57.010 1323.650 63.430 1325.250 ;
        RECT 59.135 1323.540 63.345 1323.650 ;
        RECT 65.170 1316.800 69.380 1316.865 ;
        RECT 57.010 1315.200 69.390 1316.800 ;
        RECT 65.170 1315.120 69.380 1315.200 ;
        RECT 59.175 1308.350 63.385 1308.390 ;
        RECT 57.010 1306.750 63.385 1308.350 ;
        RECT 59.175 1306.645 63.385 1306.750 ;
        RECT 65.155 1299.900 69.365 1299.975 ;
        RECT 57.010 1298.300 69.390 1299.900 ;
        RECT 65.155 1298.230 69.365 1298.300 ;
        RECT 59.155 1291.450 63.365 1291.525 ;
        RECT 57.010 1289.850 63.400 1291.450 ;
        RECT 59.155 1289.780 63.365 1289.850 ;
        RECT 65.200 1283.000 69.410 1283.075 ;
        RECT 57.010 1281.400 69.410 1283.000 ;
        RECT 65.200 1281.330 69.410 1281.400 ;
        RECT 3226.020 1219.420 3285.680 1222.520 ;
        RECT 191.030 1209.940 203.700 1216.810 ;
        RECT 3230.830 1214.620 3285.680 1217.720 ;
        RECT 248.660 1209.820 276.830 1212.920 ;
        RECT 3324.310 1210.870 3336.710 1217.550 ;
        RECT 3340.310 1214.600 3352.710 1222.280 ;
        RECT 184.040 1177.390 187.530 1207.790 ;
        RECT 248.660 1205.020 272.030 1208.120 ;
        RECT 3346.930 1200.740 3352.340 1206.230 ;
        RECT 3328.400 1192.650 3333.810 1198.140 ;
        RECT 3465.680 1186.280 3469.810 1186.340 ;
        RECT 3465.680 1184.680 3487.520 1186.280 ;
        RECT 3465.680 1184.625 3469.810 1184.680 ;
        RECT 3459.625 1182.780 3463.755 1182.855 ;
        RECT 3459.460 1181.180 3487.520 1182.780 ;
        RECT 3459.625 1181.140 3463.755 1181.180 ;
        RECT 3518.470 1167.490 3522.655 1167.575 ;
        RECT 3516.160 1165.890 3522.770 1167.490 ;
        RECT 3518.470 1165.800 3522.655 1165.890 ;
        RECT 3465.520 1162.250 3469.845 1162.350 ;
        RECT 3465.520 1160.650 3471.950 1162.250 ;
        RECT 3465.520 1160.580 3469.845 1160.650 ;
        RECT 3524.475 1159.040 3528.660 1159.120 ;
        RECT 3516.160 1157.440 3528.830 1159.040 ;
        RECT 3524.475 1157.345 3528.660 1157.440 ;
        RECT 3459.535 1153.800 3463.860 1153.860 ;
        RECT 3459.535 1152.200 3471.950 1153.800 ;
        RECT 3459.535 1152.090 3463.860 1152.200 ;
        RECT 3518.445 1150.590 3522.630 1150.705 ;
        RECT 3516.160 1148.990 3522.740 1150.590 ;
        RECT 3518.445 1148.930 3522.630 1148.990 ;
        RECT 3465.635 1145.350 3469.960 1145.435 ;
        RECT 3465.635 1143.750 3471.950 1145.350 ;
        RECT 3465.635 1143.665 3469.960 1143.750 ;
        RECT 3524.420 1142.140 3528.830 1142.250 ;
        RECT 3516.160 1140.640 3528.830 1142.140 ;
        RECT 3516.160 1140.560 3528.825 1140.640 ;
        RECT 3516.160 1140.540 3528.820 1140.560 ;
        RECT 3459.540 1136.900 3463.865 1136.960 ;
        RECT 3459.540 1135.300 3471.950 1136.900 ;
        RECT 3459.540 1135.190 3463.865 1135.300 ;
        RECT 3518.450 1133.690 3522.630 1133.780 ;
        RECT 59.120 1133.280 63.315 1133.395 ;
        RECT 41.440 1131.680 63.315 1133.280 ;
        RECT 3516.000 1132.090 3522.630 1133.690 ;
        RECT 3518.450 1131.980 3522.630 1132.090 ;
        RECT 59.120 1131.590 63.315 1131.680 ;
        RECT 65.150 1129.780 69.345 1129.850 ;
        RECT 41.440 1128.180 69.500 1129.780 ;
        RECT 3465.540 1128.450 3469.865 1128.555 ;
        RECT 65.150 1128.045 69.345 1128.180 ;
        RECT 3465.540 1126.850 3471.950 1128.450 ;
        RECT 3465.540 1126.785 3469.865 1126.850 ;
        RECT 3524.415 1125.240 3528.600 1125.320 ;
        RECT 3516.000 1123.640 3528.600 1125.240 ;
        RECT 3524.415 1123.545 3528.600 1123.640 ;
        RECT 3459.570 1120.000 3463.895 1120.100 ;
        RECT 3459.570 1118.400 3471.950 1120.000 ;
        RECT 3459.570 1118.330 3463.895 1118.400 ;
        RECT 59.135 1109.250 63.345 1109.340 ;
        RECT 57.010 1107.650 63.430 1109.250 ;
        RECT 59.135 1107.540 63.345 1107.650 ;
        RECT 65.170 1100.800 69.380 1100.865 ;
        RECT 57.010 1099.200 69.390 1100.800 ;
        RECT 65.170 1099.120 69.380 1099.200 ;
        RECT 59.175 1092.350 63.385 1092.390 ;
        RECT 57.010 1090.750 63.385 1092.350 ;
        RECT 59.175 1090.645 63.385 1090.750 ;
        RECT 65.155 1083.900 69.365 1083.975 ;
        RECT 57.010 1082.300 69.390 1083.900 ;
        RECT 65.155 1082.230 69.365 1082.300 ;
        RECT 59.155 1075.450 63.365 1075.525 ;
        RECT 57.010 1073.850 63.400 1075.450 ;
        RECT 59.155 1073.780 63.365 1073.850 ;
        RECT 65.200 1067.000 69.410 1067.075 ;
        RECT 57.010 1065.400 69.410 1067.000 ;
        RECT 65.200 1065.330 69.410 1065.400 ;
        RECT 3346.930 974.740 3352.340 980.230 ;
        RECT 3328.400 966.650 3333.810 972.140 ;
        RECT 3465.680 960.280 3469.810 960.340 ;
        RECT 3465.680 958.680 3487.520 960.280 ;
        RECT 3465.680 958.625 3469.810 958.680 ;
        RECT 3459.625 956.780 3463.755 956.855 ;
        RECT 3459.460 955.180 3487.520 956.780 ;
        RECT 3459.625 955.140 3463.755 955.180 ;
        RECT 3518.470 941.490 3522.655 941.575 ;
        RECT 3516.160 939.890 3522.770 941.490 ;
        RECT 3518.470 939.800 3522.655 939.890 ;
        RECT 3465.520 936.250 3469.845 936.350 ;
        RECT 3465.520 934.650 3471.950 936.250 ;
        RECT 3465.520 934.580 3469.845 934.650 ;
        RECT 3524.475 933.040 3528.660 933.120 ;
        RECT 3516.160 931.440 3528.830 933.040 ;
        RECT 3524.475 931.345 3528.660 931.440 ;
        RECT 3459.535 927.800 3463.860 927.860 ;
        RECT 3459.535 926.200 3471.950 927.800 ;
        RECT 3459.535 926.090 3463.860 926.200 ;
        RECT 3518.445 924.590 3522.630 924.705 ;
        RECT 3516.160 922.990 3522.740 924.590 ;
        RECT 3518.445 922.930 3522.630 922.990 ;
        RECT 3465.635 919.350 3469.960 919.435 ;
        RECT 3465.635 917.750 3471.950 919.350 ;
        RECT 3465.635 917.665 3469.960 917.750 ;
        RECT 59.120 917.280 63.315 917.395 ;
        RECT 41.440 915.680 63.315 917.280 ;
        RECT 3524.420 916.140 3528.830 916.250 ;
        RECT 59.120 915.590 63.315 915.680 ;
        RECT 3516.160 914.640 3528.830 916.140 ;
        RECT 3516.160 914.560 3528.825 914.640 ;
        RECT 3516.160 914.540 3528.820 914.560 ;
        RECT 65.150 913.780 69.345 913.850 ;
        RECT 41.440 912.180 69.500 913.780 ;
        RECT 65.150 912.045 69.345 912.180 ;
        RECT 3459.540 910.900 3463.865 910.960 ;
        RECT 3459.540 909.300 3471.950 910.900 ;
        RECT 3459.540 909.190 3463.865 909.300 ;
        RECT 3518.450 907.690 3522.630 907.780 ;
        RECT 3516.000 906.090 3522.630 907.690 ;
        RECT 3518.450 905.980 3522.630 906.090 ;
        RECT 3465.540 902.450 3469.865 902.555 ;
        RECT 3465.540 900.850 3471.950 902.450 ;
        RECT 3465.540 900.785 3469.865 900.850 ;
        RECT 3524.415 899.240 3528.600 899.320 ;
        RECT 3516.000 897.640 3528.600 899.240 ;
        RECT 3524.415 897.545 3528.600 897.640 ;
        RECT 3459.570 894.000 3463.895 894.100 ;
        RECT 59.135 893.250 63.345 893.340 ;
        RECT 57.010 891.650 63.430 893.250 ;
        RECT 3459.570 892.400 3471.950 894.000 ;
        RECT 3459.570 892.330 3463.895 892.400 ;
        RECT 59.135 891.540 63.345 891.650 ;
        RECT 65.170 884.800 69.380 884.865 ;
        RECT 57.010 883.200 69.390 884.800 ;
        RECT 65.170 883.120 69.380 883.200 ;
        RECT 59.175 876.350 63.385 876.390 ;
        RECT 57.010 874.750 63.385 876.350 ;
        RECT 59.175 874.645 63.385 874.750 ;
        RECT 65.155 867.900 69.365 867.975 ;
        RECT 57.010 866.300 69.390 867.900 ;
        RECT 65.155 866.230 69.365 866.300 ;
        RECT 59.155 859.450 63.365 859.525 ;
        RECT 57.010 857.850 63.400 859.450 ;
        RECT 59.155 857.780 63.365 857.850 ;
        RECT 65.200 851.000 69.410 851.075 ;
        RECT 57.010 849.400 69.410 851.000 ;
        RECT 65.200 849.330 69.410 849.400 ;
        RECT 3346.930 749.740 3352.340 755.230 ;
        RECT 3328.400 741.650 3333.810 747.140 ;
        RECT 3465.680 735.280 3469.810 735.340 ;
        RECT 3465.680 733.680 3487.520 735.280 ;
        RECT 3465.680 733.625 3469.810 733.680 ;
        RECT 3459.625 731.780 3463.755 731.855 ;
        RECT 3459.460 730.180 3487.520 731.780 ;
        RECT 3459.625 730.140 3463.755 730.180 ;
        RECT 3518.470 716.490 3522.655 716.575 ;
        RECT 3516.160 714.890 3522.770 716.490 ;
        RECT 3518.470 714.800 3522.655 714.890 ;
        RECT 3465.520 711.250 3469.845 711.350 ;
        RECT 3465.520 709.650 3471.950 711.250 ;
        RECT 3465.520 709.580 3469.845 709.650 ;
        RECT 3524.475 708.040 3528.660 708.120 ;
        RECT 3516.160 706.440 3528.830 708.040 ;
        RECT 3524.475 706.345 3528.660 706.440 ;
        RECT 3459.535 702.800 3463.860 702.860 ;
        RECT 3459.535 701.200 3471.950 702.800 ;
        RECT 3459.535 701.090 3463.860 701.200 ;
        RECT 3518.445 699.590 3522.630 699.705 ;
        RECT 3516.160 697.990 3522.740 699.590 ;
        RECT 3518.445 697.930 3522.630 697.990 ;
        RECT 3465.635 694.350 3469.960 694.435 ;
        RECT 3465.635 692.750 3471.950 694.350 ;
        RECT 3465.635 692.665 3469.960 692.750 ;
        RECT 3524.420 691.140 3528.830 691.250 ;
        RECT 3516.160 689.640 3528.830 691.140 ;
        RECT 3516.160 689.560 3528.825 689.640 ;
        RECT 3516.160 689.540 3528.820 689.560 ;
        RECT 3459.540 685.900 3463.865 685.960 ;
        RECT 3459.540 684.300 3471.950 685.900 ;
        RECT 3459.540 684.190 3463.865 684.300 ;
        RECT 3518.450 682.690 3522.630 682.780 ;
        RECT 3516.000 681.090 3522.630 682.690 ;
        RECT 3518.450 680.980 3522.630 681.090 ;
        RECT 3465.540 677.450 3469.865 677.555 ;
        RECT 3465.540 675.850 3471.950 677.450 ;
        RECT 3465.540 675.785 3469.865 675.850 ;
        RECT 3524.415 674.240 3528.600 674.320 ;
        RECT 3516.000 672.640 3528.600 674.240 ;
        RECT 3524.415 672.545 3528.600 672.640 ;
        RECT 3459.570 669.000 3463.895 669.100 ;
        RECT 3459.570 667.400 3471.950 669.000 ;
        RECT 3459.570 667.330 3463.895 667.400 ;
        RECT 3346.930 523.740 3352.340 529.230 ;
        RECT 3328.400 515.650 3333.810 521.140 ;
        RECT 3465.680 509.280 3469.810 509.340 ;
        RECT 3465.680 507.680 3487.520 509.280 ;
        RECT 3465.680 507.625 3469.810 507.680 ;
        RECT 3459.625 505.780 3463.755 505.855 ;
        RECT 3459.460 504.180 3487.520 505.780 ;
        RECT 3459.625 504.140 3463.755 504.180 ;
        RECT 3518.470 490.490 3522.655 490.575 ;
        RECT 3516.160 488.890 3522.770 490.490 ;
        RECT 3518.470 488.800 3522.655 488.890 ;
        RECT 3465.520 485.250 3469.845 485.350 ;
        RECT 3465.520 483.650 3471.950 485.250 ;
        RECT 3465.520 483.580 3469.845 483.650 ;
        RECT 3524.475 482.040 3528.660 482.120 ;
        RECT 3516.160 480.440 3528.830 482.040 ;
        RECT 3524.475 480.345 3528.660 480.440 ;
        RECT 3459.535 476.800 3463.860 476.860 ;
        RECT 3459.535 475.200 3471.950 476.800 ;
        RECT 3459.535 475.090 3463.860 475.200 ;
        RECT 3518.445 473.590 3522.630 473.705 ;
        RECT 3516.160 471.990 3522.740 473.590 ;
        RECT 3518.445 471.930 3522.630 471.990 ;
        RECT 3465.635 468.350 3469.960 468.435 ;
        RECT 3465.635 466.750 3471.950 468.350 ;
        RECT 3465.635 466.665 3469.960 466.750 ;
        RECT 3524.420 465.140 3528.830 465.250 ;
        RECT 3516.160 463.640 3528.830 465.140 ;
        RECT 3516.160 463.560 3528.825 463.640 ;
        RECT 3516.160 463.540 3528.820 463.560 ;
        RECT 3459.540 459.900 3463.865 459.960 ;
        RECT 3459.540 458.300 3471.950 459.900 ;
        RECT 3459.540 458.190 3463.865 458.300 ;
        RECT 3518.450 456.690 3522.630 456.780 ;
        RECT 3516.000 455.090 3522.630 456.690 ;
        RECT 3518.450 454.980 3522.630 455.090 ;
        RECT 3465.540 451.450 3469.865 451.555 ;
        RECT 3465.540 449.850 3471.950 451.450 ;
        RECT 3465.540 449.785 3469.865 449.850 ;
        RECT 3524.415 448.240 3528.600 448.320 ;
        RECT 3516.000 446.640 3528.600 448.240 ;
        RECT 3524.415 446.545 3528.600 446.640 ;
        RECT 3459.570 443.000 3463.895 443.100 ;
        RECT 3459.570 441.400 3471.950 443.000 ;
        RECT 3459.570 441.330 3463.895 441.400 ;
  END
END caravel_power_routing
END LIBRARY

