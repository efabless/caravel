* NGSPICE file created from housekeeping.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtn_1 abstract view
.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

.subckt housekeeping VGND VPWR debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oeb
+ pad_flash_csb pad_flash_csb_oeb pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ieb
+ pad_flash_io0_oeb pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ieb pad_flash_io1_oeb
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out[0] pwr_ctrl_out[1]
+ pwr_ctrl_out[2] pwr_ctrl_out[3] qspi_enabled reset ser_rx ser_tx serial_clock serial_data_1
+ serial_data_2 serial_load serial_resetn spi_csb spi_enabled spi_sck spi_sdi spi_sdo
+ spi_sdoenb spimemio_flash_clk spimemio_flash_csb spimemio_flash_io0_di spimemio_flash_io0_do
+ spimemio_flash_io0_oeb spimemio_flash_io1_di spimemio_flash_io1_do spimemio_flash_io1_oeb
+ spimemio_flash_io2_di spimemio_flash_io2_do spimemio_flash_io2_oeb spimemio_flash_io3_di
+ spimemio_flash_io3_do spimemio_flash_io3_oeb sram_ro_addr[0] sram_ro_addr[1] sram_ro_addr[2]
+ sram_ro_addr[3] sram_ro_addr[4] sram_ro_addr[5] sram_ro_addr[6] sram_ro_addr[7]
+ sram_ro_clk sram_ro_csb sram_ro_data[0] sram_ro_data[10] sram_ro_data[11] sram_ro_data[12]
+ sram_ro_data[13] sram_ro_data[14] sram_ro_data[15] sram_ro_data[16] sram_ro_data[17]
+ sram_ro_data[18] sram_ro_data[19] sram_ro_data[1] sram_ro_data[20] sram_ro_data[21]
+ sram_ro_data[22] sram_ro_data[23] sram_ro_data[24] sram_ro_data[25] sram_ro_data[26]
+ sram_ro_data[27] sram_ro_data[28] sram_ro_data[29] sram_ro_data[2] sram_ro_data[30]
+ sram_ro_data[31] sram_ro_data[3] sram_ro_data[4] sram_ro_data[5] sram_ro_data[6]
+ sram_ro_data[7] sram_ro_data[8] sram_ro_data[9] trap uart_enabled user_clock usr1_vcc_pwrgood
+ usr1_vdd_pwrgood usr2_vcc_pwrgood usr2_vdd_pwrgood wb_ack_o wb_adr_i[0] wb_adr_i[10]
+ wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17]
+ wb_adr_i[18] wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23]
+ wb_adr_i[24] wb_adr_i[25] wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2]
+ wb_adr_i[30] wb_adr_i[31] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7]
+ wb_adr_i[8] wb_adr_i[9] wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11]
+ wb_dat_i[12] wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18]
+ wb_dat_i[19] wb_dat_i[1] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24]
+ wb_dat_i[25] wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30]
+ wb_dat_i[31] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8]
+ wb_dat_i[9] wb_dat_o[0] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14]
+ wb_dat_o[15] wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20]
+ wb_dat_o[21] wb_dat_o[22] wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27]
+ wb_dat_o[28] wb_dat_o[29] wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4]
+ wb_dat_o[5] wb_dat_o[6] wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0]
+ wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] wb_stb_i wb_we_i
XFILLER_39_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7963_ _9368_/Q _7960_/X _7962_/X _9320_/Q VGND VGND VPWR VPWR _7963_/X sky130_fd_sc_hd__a22o_1
XFILLER_82_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6914_ _6521_/B _6460_/B _6812_/Y _6973_/C _6514_/Y VGND VGND VPWR VPWR _6915_/C
+ sky130_fd_sc_hd__a32o_1
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7894_ _9498_/Q _9497_/Q _7902_/B VGND VGND VPWR VPWR _7904_/B sky130_fd_sc_hd__and3_1
X_6845_ _6603_/A _6828_/X _6782_/X _6844_/Y VGND VGND VPWR VPWR _6929_/B sky130_fd_sc_hd__o211a_1
XFILLER_23_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9564_ _9564_/A _5104_/Y VGND VGND VPWR VPWR mgmt_gpio_out[10] sky130_fd_sc_hd__ebufn_8
XFILLER_168_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6776_ _6668_/A _6775_/X _6440_/A _6976_/B VGND VGND VPWR VPWR _6924_/D sky130_fd_sc_hd__a2bb2o_1
X_8515_ _9461_/Q _8348_/X _8411_/X _9341_/Q _8514_/X VGND VGND VPWR VPWR _8525_/B
+ sky130_fd_sc_hd__a221o_1
X_5727_ _5727_/A _7043_/B VGND VGND VPWR VPWR _5736_/S sky130_fd_sc_hd__nand2_4
XFILLER_109_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9495_ _9520_/CLK _9495_/D fanout470/X VGND VGND VPWR VPWR _9495_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_148_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8446_ _9378_/Q _8337_/X _8384_/X _9194_/Q _8445_/X VGND VGND VPWR VPWR _8449_/C
+ sky130_fd_sc_hd__a221o_1
X_5658_ _5658_/A VGND VGND VPWR VPWR _8918_/D sky130_fd_sc_hd__clkbuf_1
X_4609_ _9151_/Q _7091_/A _5806_/A _8987_/Q VGND VGND VPWR VPWR _4609_/X sky130_fd_sc_hd__a22o_1
XFILLER_124_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8377_ _8385_/A _8377_/B VGND VGND VPWR VPWR _8378_/A sky130_fd_sc_hd__nor2_4
X_5589_ _5589_/A VGND VGND VPWR VPWR _8889_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold340 _7630_/X VGND VGND VPWR VPWR _7631_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7328_ _7328_/A VGND VGND VPWR VPWR _9250_/D sky130_fd_sc_hd__clkbuf_1
Xhold351 _7805_/X VGND VGND VPWR VPWR _7806_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 _7788_/X VGND VGND VPWR VPWR _7789_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold373 hold373/A VGND VGND VPWR VPWR hold373/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 _5461_/X VGND VGND VPWR VPWR _5462_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7259_ _7259_/A VGND VGND VPWR VPWR _9220_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold395 hold395/A VGND VGND VPWR VPWR hold395/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1040 hold1149/X VGND VGND VPWR VPWR _5854_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1051 _9106_/Q VGND VGND VPWR VPWR _6827_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 _5826_/X VGND VGND VPWR VPWR _8989_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1073 _7080_/X VGND VGND VPWR VPWR _7081_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1084 _5844_/X VGND VGND VPWR VPWR _8995_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1095 _9397_/Q VGND VGND VPWR VPWR hold241/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_202 _8304_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_213 _8346_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_224 _8854_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_235 _9212_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_246 wb_dat_i[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_257 _5174_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_268 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_279 input38/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4960_ _4960_/A _4960_/B _4960_/C _4960_/D VGND VGND VPWR VPWR _4961_/C sky130_fd_sc_hd__or4_1
XFILLER_64_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4891_ _7158_/A _4891_/B VGND VGND VPWR VPWR _7129_/A sky130_fd_sc_hd__nor2_2
XFILLER_60_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6630_ _6664_/B _6859_/B VGND VGND VPWR VPWR _6824_/A sky130_fd_sc_hd__or2_1
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6561_ _6562_/A _6562_/B VGND VGND VPWR VPWR _6561_/X sky130_fd_sc_hd__or2_1
X_8300_ _8355_/A _8392_/C _8389_/C VGND VGND VPWR VPWR _8301_/A sky130_fd_sc_hd__and3b_4
X_5512_ _5512_/A VGND VGND VPWR VPWR _8855_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9280_ _9328_/CLK _9280_/D fanout463/X VGND VGND VPWR VPWR _9280_/Q sky130_fd_sc_hd__dfstp_1
X_6492_ _6732_/B _6492_/B VGND VGND VPWR VPWR _6618_/B sky130_fd_sc_hd__nor2_2
XFILLER_8_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8231_ _9101_/Q _8275_/B VGND VGND VPWR VPWR _8231_/X sky130_fd_sc_hd__or2_1
X_5443_ _5443_/A VGND VGND VPWR VPWR _5443_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_145_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8162_ _8162_/A _8162_/B _8162_/C _8162_/D VGND VGND VPWR VPWR _8162_/X sky130_fd_sc_hd__or4_1
X_5374_ _5374_/A VGND VGND VPWR VPWR _5374_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7113_ _7113_/A _7284_/B VGND VGND VPWR VPWR _7124_/S sky130_fd_sc_hd__nand2_2
XFILLER_87_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8093_ _9212_/Q _7923_/X _7997_/X _9364_/Q _8092_/X VGND VGND VPWR VPWR _8097_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_141_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7044_ _5947_/X _9126_/Q _7054_/S VGND VGND VPWR VPWR _7044_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8995_ _9475_/CLK _8995_/D fanout481/X VGND VGND VPWR VPWR _9577_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_27_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7946_ _9496_/Q _7991_/B _8000_/B VGND VGND VPWR VPWR _7947_/A sky130_fd_sc_hd__and3_2
XFILLER_42_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7877_ _9494_/Q VGND VGND VPWR VPWR _7929_/B sky130_fd_sc_hd__inv_2
XFILLER_168_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6828_ _6828_/A _6828_/B _6635_/A VGND VGND VPWR VPWR _6828_/X sky130_fd_sc_hd__or3b_2
XFILLER_23_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6759_ _6759_/A _6759_/B _6759_/C VGND VGND VPWR VPWR _6761_/B sky130_fd_sc_hd__or3_1
X_9547_ _9550_/CLK _9547_/D _8709_/B VGND VGND VPWR VPWR _9547_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_12_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9478_ _9485_/CLK _9478_/D fanout405/X VGND VGND VPWR VPWR _9478_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_12_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8429_ _9466_/Q _8312_/X _8376_/X _9426_/Q VGND VGND VPWR VPWR _8429_/X sky130_fd_sc_hd__a22o_1
XFILLER_136_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold170 _5616_/X VGND VGND VPWR VPWR _5617_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 _7243_/X VGND VGND VPWR VPWR _7244_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 _9452_/Q VGND VGND VPWR VPWR hold192/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5090_ _9379_/Q VGND VGND VPWR VPWR _5090_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7800_ _7800_/A VGND VGND VPWR VPWR _9464_/D sky130_fd_sc_hd__clkbuf_1
X_8780_ _8831_/CLK _8780_/D _5323_/X VGND VGND VPWR VPWR _8780_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5992_ _9067_/Q _4549_/X _5994_/S VGND VGND VPWR VPWR _5993_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7731_ _7731_/A VGND VGND VPWR VPWR _9432_/D sky130_fd_sc_hd__clkbuf_1
X_4943_ input43/X _4582_/A _6055_/A _9094_/Q _4942_/X VGND VGND VPWR VPWR _4949_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7662_ _7517_/X hold935/X _7676_/S VGND VGND VPWR VPWR _7663_/A sky130_fd_sc_hd__mux2_1
X_4874_ _8909_/Q _5630_/A _7132_/A _9166_/Q VGND VGND VPWR VPWR _4874_/X sky130_fd_sc_hd__a22o_1
XFILLER_177_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6613_ _6926_/B _6597_/Y _6605_/X wire367/X VGND VGND VPWR VPWR _6613_/X sky130_fd_sc_hd__o211a_1
X_9401_ _9427_/CLK _9401_/D fanout479/X VGND VGND VPWR VPWR hold92/A sky130_fd_sc_hd__dfstp_4
X_7593_ _7430_/X hold711/X hold75/X VGND VGND VPWR VPWR _7594_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6544_ _6382_/X _6484_/X _6809_/D _6542_/X _8735_/A VGND VGND VPWR VPWR _6544_/X
+ sky130_fd_sc_hd__a221o_1
X_9332_ _9468_/CLK _9332_/D fanout466/X VGND VGND VPWR VPWR _9332_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_9_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_5_0_csclk clkbuf_3_5_0_csclk/A VGND VGND VPWR VPWR _9303_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_180_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9263_ _9325_/CLK _9263_/D fanout464/X VGND VGND VPWR VPWR _9263_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_161_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6475_ _6588_/A _6546_/A _6987_/A _6475_/D VGND VGND VPWR VPWR _6484_/A sky130_fd_sc_hd__or4_1
XFILLER_118_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8214_ _8969_/Q _7967_/X _7999_/X _8949_/Q VGND VGND VPWR VPWR _8214_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5426_ _8820_/Q _5398_/X _5435_/S VGND VGND VPWR VPWR _5426_/X sky130_fd_sc_hd__mux2_1
Xoutput220 _5257_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[21] sky130_fd_sc_hd__buf_12
X_9194_ _9194_/CLK _9194_/D fanout456/X VGND VGND VPWR VPWR _9194_/Q sky130_fd_sc_hd__dfrtp_2
Xoutput231 _5266_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[31] sky130_fd_sc_hd__buf_12
X_5235__1 _5235__1/A VGND VGND VPWR VPWR _8779_/CLK sky130_fd_sc_hd__inv_2
Xoutput242 _5243_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[7] sky130_fd_sc_hd__buf_12
XFILLER_160_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput253 _5167_/Y VGND VGND VPWR VPWR pad_flash_csb_oeb sky130_fd_sc_hd__buf_12
X_8145_ _9414_/Q _7967_/X _7999_/X _9430_/Q VGND VGND VPWR VPWR _8145_/X sky130_fd_sc_hd__a22o_1
X_5357_ _5357_/A VGND VGND VPWR VPWR _5357_/X sky130_fd_sc_hd__clkbuf_1
Xoutput264 _9120_/Q VGND VGND VPWR VPWR pll_dco_ena sky130_fd_sc_hd__buf_12
XFILLER_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput275 _8811_/Q VGND VGND VPWR VPWR pll_trim[10] sky130_fd_sc_hd__buf_12
XFILLER_160_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput286 _9136_/Q VGND VGND VPWR VPWR pll_trim[20] sky130_fd_sc_hd__buf_12
Xoutput297 _8824_/Q VGND VGND VPWR VPWR pll_trim[7] sky130_fd_sc_hd__buf_12
XFILLER_114_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8076_ _9243_/Q _7949_/X _8224_/B _9419_/Q _8075_/X VGND VGND VPWR VPWR _8082_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_141_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5288_ _5288_/A VGND VGND VPWR VPWR _9026_/D sky130_fd_sc_hd__clkbuf_1
X_7027_ _7027_/A _7139_/B VGND VGND VPWR VPWR _7030_/S sky130_fd_sc_hd__nand2_1
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8978_ _9466_/CLK _8978_/D fanout472/X VGND VGND VPWR VPWR _8978_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_82_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7929_ _9495_/Q _7929_/B VGND VGND VPWR VPWR _8000_/B sky130_fd_sc_hd__and2_2
XFILLER_70_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire369 _6612_/Y VGND VGND VPWR VPWR wire369/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout480 fanout482/X VGND VGND VPWR VPWR fanout480/X sky130_fd_sc_hd__clkbuf_2
Xfanout491 fanout495/X VGND VGND VPWR VPWR fanout491/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4590_ _4590_/A _4590_/B _4590_/C _4590_/D VGND VGND VPWR VPWR _4591_/C sky130_fd_sc_hd__or4_1
XFILLER_115_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold906 hold906/A VGND VGND VPWR VPWR hold906/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold917 hold917/A VGND VGND VPWR VPWR hold917/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold928 _9328_/Q VGND VGND VPWR VPWR hold928/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold939 hold939/A VGND VGND VPWR VPWR hold939/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6260_ _6279_/A _7001_/A VGND VGND VPWR VPWR _6851_/A sky130_fd_sc_hd__nor2_1
XFILLER_127_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5211_ _9015_/Q input77/X _5277_/B VGND VGND VPWR VPWR _5212_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6191_ _6628_/B _6891_/B VGND VGND VPWR VPWR _6609_/A sky130_fd_sc_hd__nor2_8
X_5142_ _9032_/Q VGND VGND VPWR VPWR _5271_/A sky130_fd_sc_hd__buf_2
XFILLER_96_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5073_ _5453_/C VGND VGND VPWR VPWR _7025_/B sky130_fd_sc_hd__buf_2
XFILLER_96_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8901_ _9184_/CLK _8901_/D fanout438/X VGND VGND VPWR VPWR _8901_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_65_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8832_ _9178_/CLK _8832_/D fanout493/X VGND VGND VPWR VPWR _8832_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_92_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8763_ _9034_/Q _8763_/A2 _8763_/B1 _5871_/A VGND VGND VPWR VPWR _8763_/X sky130_fd_sc_hd__a22o_1
XFILLER_52_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5975_ _5975_/A VGND VGND VPWR VPWR _9059_/D sky130_fd_sc_hd__clkbuf_1
X_4926_ input4/X _4477_/Y _5656_/A _8918_/Q _4925_/X VGND VGND VPWR VPWR _4931_/B
+ sky130_fd_sc_hd__a221o_1
X_7714_ _7714_/A VGND VGND VPWR VPWR _9424_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8694_ _8987_/Q _8292_/X _8294_/X _8882_/Q VGND VGND VPWR VPWR _8694_/X sky130_fd_sc_hd__a22o_1
X_4857_ _4857_/A1 _4483_/Y _4450_/Y _9457_/Q _4856_/X VGND VGND VPWR VPWR _4864_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_60_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7645_ _7645_/A VGND VGND VPWR VPWR _7645_/X sky130_fd_sc_hd__buf_6
XFILLER_178_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7576_ _7430_/X hold714/X hold78/X VGND VGND VPWR VPWR _7577_/A sky130_fd_sc_hd__mux2_1
X_4788_ _8935_/Q _5693_/A _7032_/A _9123_/Q _4787_/X VGND VGND VPWR VPWR _4791_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6527_ _6527_/A _6528_/B VGND VGND VPWR VPWR _6642_/B sky130_fd_sc_hd__or2_1
X_9315_ _9465_/CLK _9315_/D fanout474/X VGND VGND VPWR VPWR _9315_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_181_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9246_ _9437_/CLK _9246_/D fanout419/X VGND VGND VPWR VPWR _9246_/Q sky130_fd_sc_hd__dfrtp_1
X_6458_ _6895_/B _6830_/A _6457_/X VGND VGND VPWR VPWR _6468_/C sky130_fd_sc_hd__o21ai_1
XFILLER_133_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5409_ hold26/X _8761_/A1 _5413_/S VGND VGND VPWR VPWR hold27/A sky130_fd_sc_hd__mux2_8
X_9177_ _9464_/CLK _9177_/D fanout420/X VGND VGND VPWR VPWR _9177_/Q sky130_fd_sc_hd__dfrtp_1
X_6389_ _6973_/A _6839_/B VGND VGND VPWR VPWR _6471_/C sky130_fd_sc_hd__xnor2_1
XFILLER_161_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8128_ _9189_/Q _8010_/B _8117_/X _8127_/X _8105_/X VGND VGND VPWR VPWR _8128_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_88_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8059_ _8059_/A _8059_/B _8059_/C _8059_/D VGND VGND VPWR VPWR _8059_/X sky130_fd_sc_hd__or4_2
XFILLER_28_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5760_ _5760_/A VGND VGND VPWR VPWR _8962_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4711_ _4711_/A _4711_/B _4711_/C _4711_/D VGND VGND VPWR VPWR _4724_/B sky130_fd_sc_hd__or4_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5691_ hold516/X _5690_/X _5691_/S VGND VGND VPWR VPWR _5692_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7430_ _7645_/A VGND VGND VPWR VPWR _7430_/X sky130_fd_sc_hd__clkbuf_2
X_4642_ _4665_/A _7158_/B VGND VGND VPWR VPWR _5784_/A sky130_fd_sc_hd__nor2_8
X_7361_ _7361_/A VGND VGND VPWR VPWR _9265_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4573_ _4573_/A _4573_/B _4573_/C _4573_/D VGND VGND VPWR VPWR _4591_/A sky130_fd_sc_hd__or4_1
XFILLER_116_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap400 _4402_/B VGND VGND VPWR VPWR _4476_/A sky130_fd_sc_hd__buf_4
XFILLER_162_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold703 _9479_/Q VGND VGND VPWR VPWR hold703/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6312_ _6312_/A _6312_/B VGND VGND VPWR VPWR _6788_/B sky130_fd_sc_hd__or2_1
Xhold714 _9362_/Q VGND VGND VPWR VPWR hold714/X sky130_fd_sc_hd__dlygate4sd3_1
X_9100_ _9442_/CLK _9100_/D fanout437/X VGND VGND VPWR VPWR _9100_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7292_ _7292_/A VGND VGND VPWR VPWR _9235_/D sky130_fd_sc_hd__clkbuf_1
Xhold725 hold725/A VGND VGND VPWR VPWR hold725/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 _7636_/X VGND VGND VPWR VPWR _7637_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 _7549_/X VGND VGND VPWR VPWR _7550_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 hold758/A VGND VGND VPWR VPWR _7055_/A sky130_fd_sc_hd__dlygate4sd3_1
X_9031_ _9551_/CLK _9031_/D _8709_/B VGND VGND VPWR VPWR _9031_/Q sky130_fd_sc_hd__dfrtp_1
Xhold769 _9234_/Q VGND VGND VPWR VPWR hold769/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6243_ _6243_/A _6716_/B VGND VGND VPWR VPWR _6744_/A sky130_fd_sc_hd__or2b_2
XFILLER_89_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6174_ _6297_/A _6297_/B _6156_/B VGND VGND VPWR VPWR _6345_/A sky130_fd_sc_hd__nor3b_4
X_5125_ _5120_/X _6312_/A _5125_/C _5125_/D VGND VGND VPWR VPWR _8705_/B sky130_fd_sc_hd__and4bb_2
XFILLER_111_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5056_ _5056_/A VGND VGND VPWR VPWR _8786_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8815_ _9487_/CLK _8815_/D fanout411/X VGND VGND VPWR VPWR _8815_/Q sky130_fd_sc_hd__dfstp_2
Xclkbuf_1_0_1_wb_clk_i clkbuf_1_0_1_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_52_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8746_ _8746_/A VGND VGND VPWR VPWR _9544_/D sky130_fd_sc_hd__clkbuf_1
X_5958_ _5653_/X hold356/X _5958_/S VGND VGND VPWR VPWR _5958_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4909_ _4909_/A _4909_/B _4909_/C _4909_/D VGND VGND VPWR VPWR _4922_/C sky130_fd_sc_hd__or4_1
XFILLER_178_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8677_ _8851_/Q _8400_/B _8663_/X _8676_/X _8627_/S VGND VGND VPWR VPWR _8677_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_139_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5889_ _9558_/A hold34/X _5898_/S VGND VGND VPWR VPWR _5889_/X sky130_fd_sc_hd__mux2_1
X_7628_ _7430_/X hold408/X _7638_/S VGND VGND VPWR VPWR _7628_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7559_ _7430_/X hold723/X hold99/A VGND VGND VPWR VPWR _7560_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_2_2_0_csclk clkbuf_2_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_5_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_134_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9229_ _9469_/CLK _9229_/D fanout458/X VGND VGND VPWR VPWR _9229_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold30 hold30/A VGND VGND VPWR VPWR hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A VGND VGND VPWR VPWR hold41/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold52 hold52/A VGND VGND VPWR VPWR hold52/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold63 hold63/A VGND VGND VPWR VPWR hold63/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold74 hold74/A VGND VGND VPWR VPWR hold74/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold85 hold85/A VGND VGND VPWR VPWR hold85/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 hold96/A VGND VGND VPWR VPWR hold96/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_5 _5911_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6930_ _6628_/A _6473_/Y _6710_/C _6867_/B VGND VGND VPWR VPWR _6989_/A sky130_fd_sc_hd__a211o_1
XFILLER_81_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6861_ _6861_/A _6946_/C _6964_/C _6861_/D VGND VGND VPWR VPWR _6864_/B sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_6_csclk _9359_/CLK VGND VGND VPWR VPWR _9367_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_62_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8600_ _8600_/A _8600_/B _8600_/C _8600_/D VGND VGND VPWR VPWR _8601_/D sky130_fd_sc_hd__or4_1
XFILLER_179_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5812_ hold606/X _5683_/X _5816_/S VGND VGND VPWR VPWR _5813_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9580_ _9580_/A _5088_/Y VGND VGND VPWR VPWR mgmt_gpio_out[26] sky130_fd_sc_hd__ebufn_8
X_6792_ _6792_/A _7001_/B VGND VGND VPWR VPWR _6806_/B sky130_fd_sc_hd__nor2_1
XFILLER_34_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_0_0_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR clkbuf_2_1_0_mgmt_gpio_in[4]/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_179_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8531_ _9374_/Q _8682_/B VGND VGND VPWR VPWR _8531_/X sky130_fd_sc_hd__and2_1
X_5743_ _5647_/X hold811/X _5747_/S VGND VGND VPWR VPWR _5744_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8462_ _9443_/Q _8301_/A _8356_/C _9483_/Q VGND VGND VPWR VPWR _8462_/X sky130_fd_sc_hd__a22o_1
X_5674_ _5650_/X hold395/X _5676_/S VGND VGND VPWR VPWR _5675_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4625_ _4635_/A _4891_/B VGND VGND VPWR VPWR _5656_/A sky130_fd_sc_hd__nor2_4
X_7413_ _7233_/X hold787/X _7423_/S VGND VGND VPWR VPWR _7414_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8393_ _9216_/Q _8391_/X _8411_/A _9336_/Q VGND VGND VPWR VPWR _8393_/X sky130_fd_sc_hd__a22o_1
XFILLER_175_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold500 hold500/A VGND VGND VPWR VPWR hold500/X sky130_fd_sc_hd__dlygate4sd3_1
X_7344_ _7233_/X hold781/X _7354_/S VGND VGND VPWR VPWR _7345_/A sky130_fd_sc_hd__mux2_1
X_4556_ _4758_/A _4794_/B VGND VGND VPWR VPWR _7043_/A sky130_fd_sc_hd__nor2_4
Xhold511 _7786_/X VGND VGND VPWR VPWR _7787_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold522 hold522/A VGND VGND VPWR VPWR hold522/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 _9279_/Q VGND VGND VPWR VPWR hold533/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold544 _9049_/Q VGND VGND VPWR VPWR hold544/X sky130_fd_sc_hd__dlygate4sd3_1
X_7275_ _7239_/X hold167/X _7282_/S VGND VGND VPWR VPWR _7275_/X sky130_fd_sc_hd__mux2_1
Xhold555 _6010_/X VGND VGND VPWR VPWR _6011_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold566 hold566/A VGND VGND VPWR VPWR hold566/X sky130_fd_sc_hd__dlygate4sd3_1
X_4487_ _9455_/Q _7764_/A _4483_/Y _4487_/B2 _4486_/X VGND VGND VPWR VPWR _4495_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold577 _8925_/Q VGND VGND VPWR VPWR hold577/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 hold588/A VGND VGND VPWR VPWR hold588/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9014_ _9181_/CLK _9014_/D fanout488/X VGND VGND VPWR VPWR _9559_/A sky130_fd_sc_hd__dfrtp_1
X_6226_ _6437_/A _6716_/A _6416_/A VGND VGND VPWR VPWR _6510_/A sky130_fd_sc_hd__nor3_4
Xhold599 _7534_/X VGND VGND VPWR VPWR _7535_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6157_ _6228_/A _6249_/A VGND VGND VPWR VPWR _6158_/B sky130_fd_sc_hd__or2_2
Xhold1200 _7142_/X VGND VGND VPWR VPWR hold803/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1211 _9359_/Q VGND VGND VPWR VPWR hold841/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1222 _9430_/Q VGND VGND VPWR VPWR hold196/A sky130_fd_sc_hd__dlygate4sd3_1
X_5108_ _9235_/Q VGND VGND VPWR VPWR _5108_/Y sky130_fd_sc_hd__inv_2
Xhold1233 _9096_/Q VGND VGND VPWR VPWR hold600/A sky130_fd_sc_hd__dlygate4sd3_1
X_6088_ _6182_/A _6088_/B _6093_/B VGND VGND VPWR VPWR _6089_/B sky130_fd_sc_hd__and3_1
Xhold1244 _5302_/X VGND VGND VPWR VPWR _5303_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1255 _9079_/Q VGND VGND VPWR VPWR hold884/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1266 _8923_/Q VGND VGND VPWR VPWR hold847/A sky130_fd_sc_hd__dlygate4sd3_1
X_5039_ _5068_/B _5039_/B VGND VGND VPWR VPWR _5127_/A sky130_fd_sc_hd__nand2_1
XFILLER_45_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1277 _8868_/Q VGND VGND VPWR VPWR hold906/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_406 hold27/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8729_ _5287_/A _8729_/A2 _8729_/B1 _5275_/A _8728_/X VGND VGND VPWR VPWR _8729_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_185_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput120 sram_ro_data[5] VGND VGND VPWR VPWR _4589_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput131 wb_adr_i[0] VGND VGND VPWR VPWR _6317_/A sky130_fd_sc_hd__clkbuf_4
Xinput142 wb_adr_i[1] VGND VGND VPWR VPWR _6167_/A sky130_fd_sc_hd__clkbuf_2
Xinput153 wb_adr_i[2] VGND VGND VPWR VPWR _6167_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xinput164 wb_dat_i[0] VGND VGND VPWR VPWR _8728_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput175 wb_dat_i[1] VGND VGND VPWR VPWR _8740_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput186 wb_dat_i[2] VGND VGND VPWR VPWR _8744_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput197 wb_sel_i[0] VGND VGND VPWR VPWR _8734_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4410_ _9287_/Q _7391_/A _7339_/A _9263_/Q VGND VGND VPWR VPWR _4410_/X sky130_fd_sc_hd__a22o_2
XFILLER_145_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5390_ _8809_/Q _5387_/X _5416_/S VGND VGND VPWR VPWR _5390_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7060_ _9133_/Q _5809_/X _7072_/S VGND VGND VPWR VPWR _7060_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6011_ _6011_/A VGND VGND VPWR VPWR _9075_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7962_ _7962_/A VGND VGND VPWR VPWR _7962_/X sky130_fd_sc_hd__buf_6
X_6913_ _6396_/B _6445_/Y _6523_/X _6905_/A _6433_/B VGND VGND VPWR VPWR _6997_/C
+ sky130_fd_sc_hd__a2111o_1
X_7893_ _7920_/B _8375_/A _8342_/B _7875_/X _7893_/B2 VGND VGND VPWR VPWR _9498_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_63_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6844_ _6844_/A _6844_/B VGND VGND VPWR VPWR _6844_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9563_ _9563_/A _5105_/Y VGND VGND VPWR VPWR mgmt_gpio_out[9] sky130_fd_sc_hd__ebufn_2
X_6775_ _6779_/A _6775_/B _6775_/C VGND VGND VPWR VPWR _6775_/X sky130_fd_sc_hd__or3_1
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8514_ _9221_/Q _8391_/X _8367_/X _9477_/Q _8513_/X VGND VGND VPWR VPWR _8514_/X
+ sky130_fd_sc_hd__a221o_2
X_5726_ hold20/X VGND VGND VPWR VPWR _7043_/B sky130_fd_sc_hd__buf_12
X_9494_ _9520_/CLK _9494_/D fanout469/X VGND VGND VPWR VPWR _9494_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_109_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8445_ _9434_/Q _7908_/X _8335_/X _9274_/Q VGND VGND VPWR VPWR _8445_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5657_ hold930/X _5505_/X _5665_/S VGND VGND VPWR VPWR _5658_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4608_ _4665_/A _4891_/B VGND VGND VPWR VPWR _5806_/A sky130_fd_sc_hd__nor2_2
X_5588_ hold749/X _5587_/X _5594_/S VGND VGND VPWR VPWR _5589_/A sky130_fd_sc_hd__mux2_1
X_8376_ _8376_/A VGND VGND VPWR VPWR _8376_/X sky130_fd_sc_hd__buf_6
Xhold330 _9189_/Q VGND VGND VPWR VPWR hold330/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4539_ _4539_/A VGND VGND VPWR VPWR _4539_/X sky130_fd_sc_hd__clkbuf_4
Xhold341 _7041_/X VGND VGND VPWR VPWR _7042_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7327_ hold720/X _6048_/X _7337_/S VGND VGND VPWR VPWR _7327_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold352 _9196_/Q VGND VGND VPWR VPWR hold352/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold363 _9106_/Q VGND VGND VPWR VPWR hold363/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 _9179_/Q VGND VGND VPWR VPWR hold374/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 _7070_/X VGND VGND VPWR VPWR _7071_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7258_ _7239_/X hold165/X _7264_/S VGND VGND VPWR VPWR _7258_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold396 _8936_/Q VGND VGND VPWR VPWR hold396/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6209_ _6790_/B _6799_/A VGND VGND VPWR VPWR _6209_/X sky130_fd_sc_hd__or2_1
X_7189_ _7189_/A VGND VGND VPWR VPWR _9189_/D sky130_fd_sc_hd__clkbuf_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1030 _8784_/Q VGND VGND VPWR VPWR _5059_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1041 hold1186/X VGND VGND VPWR VPWR _5893_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1052 _9544_/Q VGND VGND VPWR VPWR _8745_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1063 _5822_/X VGND VGND VPWR VPWR _5823_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1074 _7081_/X VGND VGND VPWR VPWR _9142_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1085 _7613_/X VGND VGND VPWR VPWR _7614_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1096 _8908_/Q VGND VGND VPWR VPWR hold849/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_203 _8360_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_214 _8701_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_225 _8854_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_236 _9212_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_247 wb_dat_i[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_258 _5174_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_269 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_71_csclk _9090_/CLK VGND VGND VPWR VPWR _9203_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4890_ _7111_/B VGND VGND VPWR VPWR _4890_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_86_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _9383_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_80_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6560_ _6560_/A _6560_/B VGND VGND VPWR VPWR _6960_/A sky130_fd_sc_hd__or2_1
XFILLER_13_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5511_ hold601/X _5395_/X _5515_/S VGND VGND VPWR VPWR _5511_/X sky130_fd_sc_hd__mux2_1
X_6491_ _6790_/B _6651_/A VGND VGND VPWR VPWR _6925_/A sky130_fd_sc_hd__nor2_1
XFILLER_8_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5442_ _7011_/A _7013_/B VGND VGND VPWR VPWR _5443_/A sky130_fd_sc_hd__and2_1
X_8230_ _8970_/Q _7967_/X _7990_/X _8870_/Q _8229_/X VGND VGND VPWR VPWR _8238_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5373_ _5375_/A _5378_/B VGND VGND VPWR VPWR _5374_/A sky130_fd_sc_hd__and2_1
X_8161_ _9223_/Q _7927_/X _8023_/B _9311_/Q _8160_/X VGND VGND VPWR VPWR _8162_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_172_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_24_csclk _9303_/CLK VGND VGND VPWR VPWR _9305_/CLK sky130_fd_sc_hd__clkbuf_16
X_7112_ _9156_/Q _4944_/Y _7139_/B _7111_/X VGND VGND VPWR VPWR _7112_/X sky130_fd_sc_hd__o211a_1
XFILLER_99_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8092_ _9324_/Q _7962_/X _7988_/X _9436_/Q VGND VGND VPWR VPWR _8092_/X sky130_fd_sc_hd__a22o_1
X_7043_ _7043_/A _7043_/B VGND VGND VPWR VPWR _7054_/S sky130_fd_sc_hd__nand2_2
XFILLER_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_39_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _9178_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_55_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_1_0_csclk clkbuf_3_1_0_csclk/A VGND VGND VPWR VPWR _9359_/CLK sky130_fd_sc_hd__clkbuf_8
X_8994_ _9468_/CLK _8994_/D fanout477/X VGND VGND VPWR VPWR _9576_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_82_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7945_ _9200_/Q _7938_/X _7940_/X _9248_/Q _7944_/X VGND VGND VPWR VPWR _7965_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7876_ _7920_/B _7991_/B _7989_/B _7876_/B1 _7875_/X VGND VGND VPWR VPWR _9493_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_179_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6827_ _6753_/Y _6786_/Y _6826_/X _6908_/A _6827_/B2 VGND VGND VPWR VPWR _9106_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_51_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9546_ _9551_/CLK _9546_/D fanout500/X VGND VGND VPWR VPWR _9546_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_10_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6758_ _6758_/A _6758_/B _6758_/C _6834_/A VGND VGND VPWR VPWR _6761_/A sky130_fd_sc_hd__or4b_1
XFILLER_149_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5709_ hold663/X _5683_/X _5713_/S VGND VGND VPWR VPWR _5710_/A sky130_fd_sc_hd__mux2_1
XFILLER_176_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9477_ _9477_/CLK _9477_/D fanout406/X VGND VGND VPWR VPWR _9477_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6689_ _6421_/A _6441_/B _6609_/B _6481_/A VGND VGND VPWR VPWR _6689_/X sky130_fd_sc_hd__o211a_1
XFILLER_109_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8428_ _8428_/A VGND VGND VPWR VPWR _9521_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8359_ _8363_/A _8359_/B VGND VGND VPWR VPWR _8379_/A sky130_fd_sc_hd__nor2_2
XFILLER_163_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold160 _6075_/X VGND VGND VPWR VPWR _6076_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold171 _8937_/Q VGND VGND VPWR VPWR hold171/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 _9177_/Q VGND VGND VPWR VPWR hold182/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold193 _7773_/X VGND VGND VPWR VPWR _7774_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5991_ _5991_/A VGND VGND VPWR VPWR _9066_/D sky130_fd_sc_hd__clkbuf_1
X_7730_ _5387_/X hold900/X hold86/X VGND VGND VPWR VPWR _7731_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4942_ _9368_/Q _7588_/A _5948_/A _9048_/Q VGND VGND VPWR VPWR _4942_/X sky130_fd_sc_hd__a22o_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7661_ _7661_/A _7695_/B VGND VGND VPWR VPWR _7676_/S sky130_fd_sc_hd__nand2_8
X_4873_ _4873_/A _4873_/B _4873_/C _4873_/D VGND VGND VPWR VPWR _4884_/C sky130_fd_sc_hd__or4_1
XFILLER_178_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9400_ _9416_/CLK _9400_/D fanout425/X VGND VGND VPWR VPWR _9400_/Q sky130_fd_sc_hd__dfstp_1
X_6612_ _6228_/Y _6973_/B _6607_/Y _6608_/Y _6611_/Y VGND VGND VPWR VPWR _6612_/Y
+ sky130_fd_sc_hd__a2111oi_1
X_7592_ _7592_/A VGND VGND VPWR VPWR _9369_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9331_ _9419_/CLK _9331_/D fanout491/X VGND VGND VPWR VPWR _9331_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6543_ _6543_/A _6543_/B VGND VGND VPWR VPWR _8735_/A sky130_fd_sc_hd__nor2_8
XFILLER_146_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9262_ _9325_/CLK _9262_/D fanout460/X VGND VGND VPWR VPWR _9262_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_173_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6474_ _6481_/A _6404_/Y _6469_/X _6473_/Y VGND VGND VPWR VPWR _6475_/D sky130_fd_sc_hd__a211o_1
X_8213_ _9075_/Q _8034_/X _8210_/X _8212_/X VGND VGND VPWR VPWR _8216_/C sky130_fd_sc_hd__a211o_1
XFILLER_146_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5425_ _5425_/A VGND VGND VPWR VPWR _8819_/D sky130_fd_sc_hd__clkbuf_1
Xoutput210 _5248_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[12] sky130_fd_sc_hd__buf_12
XFILLER_133_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput221 _5258_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[22] sky130_fd_sc_hd__buf_12
X_9193_ _9195_/CLK _9193_/D fanout467/X VGND VGND VPWR VPWR _9193_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput232 _5267_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[32] sky130_fd_sc_hd__buf_12
Xoutput243 _5244_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[8] sky130_fd_sc_hd__buf_12
XFILLER_133_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5356_ _5375_/A _5356_/B VGND VGND VPWR VPWR _5357_/A sky130_fd_sc_hd__and2_1
Xoutput254 _5178_/X VGND VGND VPWR VPWR pad_flash_io0_do sky130_fd_sc_hd__buf_12
X_8144_ _9238_/Q _8034_/X _8141_/X _8143_/X VGND VGND VPWR VPWR _8149_/B sky130_fd_sc_hd__a211o_1
Xoutput265 _9121_/Q VGND VGND VPWR VPWR pll_div[0] sky130_fd_sc_hd__buf_12
Xoutput276 _8812_/Q VGND VGND VPWR VPWR pll_trim[11] sky130_fd_sc_hd__buf_12
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput287 _9137_/Q VGND VGND VPWR VPWR pll_trim[21] sky130_fd_sc_hd__buf_12
Xoutput298 _8809_/Q VGND VGND VPWR VPWR pll_trim[8] sky130_fd_sc_hd__buf_12
X_5287_ _5287_/A _5287_/B VGND VGND VPWR VPWR _5288_/A sky130_fd_sc_hd__and2_1
X_8075_ _9315_/Q _8008_/B _7979_/A _9227_/Q _7984_/X VGND VGND VPWR VPWR _8075_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7026_ _7026_/A VGND VGND VPWR VPWR _7026_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_75_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8977_ _9087_/CLK _8977_/D fanout447/X VGND VGND VPWR VPWR _8977_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_82_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7928_ _9496_/Q VGND VGND VPWR VPWR _7998_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_169_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7859_ _9488_/Q _9489_/Q _7858_/Y VGND VGND VPWR VPWR _7860_/B sky130_fd_sc_hd__a21o_1
XFILLER_168_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9529_ _9529_/CLK _9529_/D fanout448/X VGND VGND VPWR VPWR _9529_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout470 fanout497/X VGND VGND VPWR VPWR fanout470/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout481 fanout482/X VGND VGND VPWR VPWR fanout481/X sky130_fd_sc_hd__clkbuf_4
XFILLER_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout492 fanout495/X VGND VGND VPWR VPWR fanout492/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold907 _7092_/X VGND VGND VPWR VPWR _7093_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold918 hold918/A VGND VGND VPWR VPWR hold918/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold929 _9344_/Q VGND VGND VPWR VPWR hold929/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5210_ _5210_/A VGND VGND VPWR VPWR _9562_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_89_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6190_ _6190_/A VGND VGND VPWR VPWR _6624_/B sky130_fd_sc_hd__buf_2
X_5141_ _5135_/X _5139_/Y _5155_/B _7919_/A3 VGND VGND VPWR VPWR _8999_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_96_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5072_ _7158_/C VGND VGND VPWR VPWR _5453_/C sky130_fd_sc_hd__buf_4
XFILLER_96_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8900_ _9442_/CLK _8900_/D fanout438/X VGND VGND VPWR VPWR _8900_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_56_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8831_ _8831_/CLK _8831_/D _5451_/X VGND VGND VPWR VPWR _8831_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8762_ _8762_/A VGND VGND VPWR VPWR _9548_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5974_ _9059_/Q _4549_/X _5976_/S VGND VGND VPWR VPWR _5975_/A sky130_fd_sc_hd__mux2_1
X_7713_ _5387_/X hold888/X hold95/X VGND VGND VPWR VPWR _7714_/A sky130_fd_sc_hd__mux2_1
X_4925_ _9352_/Q _4427_/Y _6043_/A _9089_/Q VGND VGND VPWR VPWR _4925_/X sky130_fd_sc_hd__a22o_1
X_8693_ _9078_/Q _8322_/X _8333_/X _8867_/Q _8692_/X VGND VGND VPWR VPWR _8700_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7644_ _7644_/A VGND VGND VPWR VPWR _9393_/D sky130_fd_sc_hd__clkbuf_1
X_4856_ _9201_/Q _7211_/A _5573_/A _8884_/Q VGND VGND VPWR VPWR _4856_/X sky130_fd_sc_hd__a22o_2
XFILLER_178_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7575_ _7575_/A VGND VGND VPWR VPWR _9361_/D sky130_fd_sc_hd__clkbuf_1
X_4787_ _9482_/Q _4898_/A2 _4500_/Y input13/X VGND VGND VPWR VPWR _4787_/X sky130_fd_sc_hd__a22o_1
X_9314_ _9452_/CLK _9314_/D fanout429/X VGND VGND VPWR VPWR _9314_/Q sky130_fd_sc_hd__dfrtp_4
X_6526_ _6906_/B _6926_/A VGND VGND VPWR VPWR _6917_/B sky130_fd_sc_hd__or2_1
XFILLER_119_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9245_ _9477_/CLK _9245_/D fanout406/X VGND VGND VPWR VPWR _9245_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6457_ _6514_/A _6524_/C VGND VGND VPWR VPWR _6457_/X sky130_fd_sc_hd__or2_1
XFILLER_173_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5408_ _5408_/A VGND VGND VPWR VPWR _8814_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9176_ _9464_/CLK _9176_/D fanout420/X VGND VGND VPWR VPWR _9176_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6388_ _6794_/A _6175_/A _6633_/A _6387_/Y VGND VGND VPWR VPWR _6667_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8127_ _8127_/A _8127_/B _8127_/C _8127_/D VGND VGND VPWR VPWR _8127_/X sky130_fd_sc_hd__or4_1
XFILLER_87_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5339_ _5353_/A _5356_/B VGND VGND VPWR VPWR _5340_/A sky130_fd_sc_hd__and2_1
XFILLER_75_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8058_ _9354_/Q _8020_/A _7990_/A _9274_/Q _8057_/X VGND VGND VPWR VPWR _8059_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_102_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7009_ _7009_/A _7009_/B _7009_/C _7008_/X VGND VGND VPWR VPWR _7010_/A sky130_fd_sc_hd__or4b_1
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _9307_/Q _7446_/A _7781_/A _9459_/Q _4709_/X VGND VGND VPWR VPWR _4711_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_30_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5690_ _5690_/A VGND VGND VPWR VPWR _5690_/X sky130_fd_sc_hd__buf_4
XFILLER_175_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4641_ _4667_/A _7126_/B VGND VGND VPWR VPWR _5948_/A sky130_fd_sc_hd__nor2_4
XFILLER_147_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4572_ _9317_/Q _7463_/A _7091_/A _9152_/Q _4571_/X VGND VGND VPWR VPWR _4573_/D
+ sky130_fd_sc_hd__a221o_1
X_7360_ _7359_/X hold144/X _7372_/S VGND VGND VPWR VPWR _7360_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap401 _5051_/C VGND VGND VPWR VPWR _5045_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_116_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold704 _7830_/X VGND VGND VPWR VPWR _7831_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6311_ _6402_/A _6311_/B VGND VGND VPWR VPWR _6715_/B sky130_fd_sc_hd__nor2_4
Xhold715 hold715/A VGND VGND VPWR VPWR hold715/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 _7218_/X VGND VGND VPWR VPWR _7219_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7291_ _7236_/X _9235_/Q _7300_/S VGND VGND VPWR VPWR _7291_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold737 hold737/A VGND VGND VPWR VPWR hold737/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold748 _7096_/X VGND VGND VPWR VPWR _7097_/A sky130_fd_sc_hd__dlygate4sd3_1
X_9030_ _9551_/CLK _9030_/D fanout499/X VGND VGND VPWR VPWR _9030_/Q sky130_fd_sc_hd__dfrtp_4
Xhold759 _9310_/Q VGND VGND VPWR VPWR hold759/X sky130_fd_sc_hd__dlygate4sd3_1
X_6242_ _6227_/Y _6194_/B _6144_/A _6158_/B VGND VGND VPWR VPWR _6250_/B sky130_fd_sc_hd__o22a_1
X_6173_ _6415_/A _6317_/B _6318_/A VGND VGND VPWR VPWR _6297_/B sky130_fd_sc_hd__and3_1
X_5124_ input150/X input151/X _5124_/C _5124_/D VGND VGND VPWR VPWR _5125_/D sky130_fd_sc_hd__and4bb_1
XFILLER_85_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5055_ _5057_/A1 _5055_/A1 _5065_/S VGND VGND VPWR VPWR _5056_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8814_ _9487_/CLK _8814_/D fanout411/X VGND VGND VPWR VPWR _8814_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_111_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8745_ _8744_/X _8745_/A1 _8765_/S VGND VGND VPWR VPWR _8746_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5957_ _5957_/A VGND VGND VPWR VPWR _9051_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4908_ _9147_/Q _7091_/A _6066_/A _9099_/Q _4907_/X VGND VGND VPWR VPWR _4909_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_139_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8676_ _8701_/A _8676_/B _8676_/C VGND VGND VPWR VPWR _8676_/X sky130_fd_sc_hd__or3_1
X_5888_ _9180_/Q hold24/X _5897_/S VGND VGND VPWR VPWR hold34/A sky130_fd_sc_hd__mux2_1
XFILLER_139_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7627_ hold91/X VGND VGND VPWR VPWR _9385_/D sky130_fd_sc_hd__clkbuf_1
X_4839_ _9465_/Q _7798_/A _7266_/A _9225_/Q VGND VGND VPWR VPWR _4839_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7558_ _7558_/A VGND VGND VPWR VPWR _9353_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6509_ _6967_/B _6926_/B _6895_/A VGND VGND VPWR VPWR _6509_/X sky130_fd_sc_hd__a21o_1
XFILLER_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7489_ _7489_/A VGND VGND VPWR VPWR _9323_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9228_ _9452_/CLK _9228_/D fanout415/X VGND VGND VPWR VPWR _9228_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9159_ _9161_/CLK _9159_/D fanout440/X VGND VGND VPWR VPWR _9159_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_121_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold20 hold20/A VGND VGND VPWR VPWR hold20/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold31 hold31/A VGND VGND VPWR VPWR hold31/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold42 hold42/A VGND VGND VPWR VPWR hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A VGND VGND VPWR VPWR hold53/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold64 hold64/A VGND VGND VPWR VPWR hold64/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold75 hold75/A VGND VGND VPWR VPWR hold75/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold86 hold86/A VGND VGND VPWR VPWR hold86/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A VGND VGND VPWR VPWR hold97/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_6 _9075_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6860_ _6876_/B _6860_/B VGND VGND VPWR VPWR _6861_/D sky130_fd_sc_hd__and2b_1
XFILLER_62_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5811_ _5811_/A VGND VGND VPWR VPWR _8984_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6791_ _6791_/A VGND VGND VPWR VPWR _7001_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_50_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8530_ _9422_/Q _8402_/A _8378_/A _9358_/Q _8529_/X VGND VGND VPWR VPWR _8537_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5742_ _5742_/A VGND VGND VPWR VPWR _8954_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8461_ _9411_/Q _8506_/B _8456_/X _8458_/X _8460_/X VGND VGND VPWR VPWR _8461_/X
+ sky130_fd_sc_hd__a2111o_1
X_5673_ _5673_/A VGND VGND VPWR VPWR _8925_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7412_ _7412_/A VGND VGND VPWR VPWR _9289_/D sky130_fd_sc_hd__clkbuf_1
X_4624_ _8821_/Q _5418_/A _5296_/A _8776_/Q _4623_/X VGND VGND VPWR VPWR _4633_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_163_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8392_ _8392_/A _8398_/A _8392_/C VGND VGND VPWR VPWR _8411_/A sky130_fd_sc_hd__and3_4
XFILLER_135_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold501 _8910_/Q VGND VGND VPWR VPWR hold501/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7343_ _7343_/A VGND VGND VPWR VPWR _9257_/D sky130_fd_sc_hd__clkbuf_1
X_4555_ _4555_/A _4555_/B VGND VGND VPWR VPWR _4794_/B sky130_fd_sc_hd__nand2_8
Xhold512 _9101_/Q VGND VGND VPWR VPWR hold512/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 _5906_/X VGND VGND VPWR VPWR _5907_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 _7389_/X VGND VGND VPWR VPWR _7390_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold545 _5952_/X VGND VGND VPWR VPWR _5953_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 _9100_/Q VGND VGND VPWR VPWR hold556/X sky130_fd_sc_hd__dlygate4sd3_1
X_7274_ _7274_/A VGND VGND VPWR VPWR _9227_/D sky130_fd_sc_hd__clkbuf_1
X_4486_ _9407_/Q _7661_/A _4485_/Y _9375_/Q VGND VGND VPWR VPWR _4486_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold567 _9183_/Q VGND VGND VPWR VPWR hold567/X sky130_fd_sc_hd__dlygate4sd3_1
X_9013_ _9181_/CLK _9013_/D fanout487/X VGND VGND VPWR VPWR _9558_/A sky130_fd_sc_hd__dfrtp_1
Xhold578 _8935_/Q VGND VGND VPWR VPWR hold578/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold589 _7120_/X VGND VGND VPWR VPWR _7121_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6225_ _6635_/A _6628_/B VGND VGND VPWR VPWR _6897_/A sky130_fd_sc_hd__nor2_4
XFILLER_131_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6156_ _6739_/B _6156_/B VGND VGND VPWR VPWR _6249_/A sky130_fd_sc_hd__nand2_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1201 _8892_/Q VGND VGND VPWR VPWR hold804/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1212 _9322_/Q VGND VGND VPWR VPWR hold722/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1223 _9164_/Q VGND VGND VPWR VPWR hold916/A sky130_fd_sc_hd__dlygate4sd3_1
X_5107_ _9243_/Q VGND VGND VPWR VPWR _5107_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1234 _8978_/Q VGND VGND VPWR VPWR hold882/A sky130_fd_sc_hd__dlygate4sd3_1
X_6087_ _6437_/A _6175_/A _6095_/B VGND VGND VPWR VPWR _6093_/B sky130_fd_sc_hd__and3_1
XFILLER_111_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1245 _8949_/Q VGND VGND VPWR VPWR hold455/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1256 _8775_/Q VGND VGND VPWR VPWR hold397/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1267 _9428_/Q VGND VGND VPWR VPWR hold354/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1278 _8879_/Q VGND VGND VPWR VPWR hold459/A sky130_fd_sc_hd__dlygate4sd3_1
X_5038_ _5035_/B _8806_/Q _5021_/A _4550_/S _5039_/B VGND VGND VPWR VPWR _5051_/C
+ sky130_fd_sc_hd__a2111oi_2
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6989_ _6989_/A _6989_/B _6989_/C VGND VGND VPWR VPWR _7008_/A sky130_fd_sc_hd__or3_1
XFILLER_53_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8728_ _5271_/A _8728_/A2 _8728_/B1 _8727_/Y VGND VGND VPWR VPWR _8728_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8659_ _8916_/Q _8298_/X _8370_/X _9087_/Q VGND VGND VPWR VPWR _8659_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput110 sram_ro_data[25] VGND VGND VPWR VPWR _4857_/A1 sky130_fd_sc_hd__buf_2
XFILLER_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput121 sram_ro_data[6] VGND VGND VPWR VPWR _4514_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_163_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput132 wb_adr_i[10] VGND VGND VPWR VPWR _6080_/D sky130_fd_sc_hd__clkbuf_1
Xinput143 wb_adr_i[20] VGND VGND VPWR VPWR _5121_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput154 wb_adr_i[30] VGND VGND VPWR VPWR input154/X sky130_fd_sc_hd__clkbuf_1
Xinput165 wb_dat_i[10] VGND VGND VPWR VPWR _8743_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput176 wb_dat_i[20] VGND VGND VPWR VPWR _8752_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput187 wb_dat_i[30] VGND VGND VPWR VPWR _8760_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput198 wb_sel_i[1] VGND VGND VPWR VPWR _8769_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6010_ _5951_/X hold554/X _6019_/S VGND VGND VPWR VPWR _6010_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7961_ _9496_/Q _7984_/C _7992_/C VGND VGND VPWR VPWR _7962_/A sky130_fd_sc_hd__and3_2
X_6912_ _6912_/A VGND VGND VPWR VPWR _9107_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7892_ _9498_/Q _9497_/Q VGND VGND VPWR VPWR _8342_/B sky130_fd_sc_hd__nor2b_2
XFILLER_23_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6843_ _6354_/B _6761_/B _6843_/C _6843_/D VGND VGND VPWR VPWR _7006_/C sky130_fd_sc_hd__and4bb_1
X_9562_ _9562_/A _5106_/Y VGND VGND VPWR VPWR mgmt_gpio_out[8] sky130_fd_sc_hd__ebufn_8
X_6774_ _6230_/X _6811_/B _6672_/C _6660_/A _6422_/B VGND VGND VPWR VPWR _6987_/D
+ sky130_fd_sc_hd__a32o_1
X_8513_ _9445_/Q _8398_/B _8344_/X _9485_/Q VGND VGND VPWR VPWR _8513_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5725_ _5725_/A VGND VGND VPWR VPWR _8947_/D sky130_fd_sc_hd__clkbuf_1
X_9493_ _9520_/CLK _9493_/D fanout469/X VGND VGND VPWR VPWR _9493_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_148_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8444_ _9226_/Q _8388_/X _8379_/X _9202_/Q _8443_/X VGND VGND VPWR VPWR _8449_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5656_ _5656_/A _5715_/B VGND VGND VPWR VPWR _5665_/S sky130_fd_sc_hd__and2_2
XFILLER_108_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4607_ _4635_/A _7126_/B VGND VGND VPWR VPWR _5795_/A sky130_fd_sc_hd__nor2_8
X_8375_ _8375_/A _8389_/A _8398_/A VGND VGND VPWR VPWR _8376_/A sky130_fd_sc_hd__and3_4
XFILLER_163_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5587_ _5951_/A VGND VGND VPWR VPWR _5587_/X sky130_fd_sc_hd__buf_4
Xhold320 _9486_/Q VGND VGND VPWR VPWR hold320/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 _7188_/X VGND VGND VPWR VPWR _7189_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7326_ _7326_/A VGND VGND VPWR VPWR _9249_/D sky130_fd_sc_hd__clkbuf_1
X_4538_ _9532_/Q _9161_/Q _9162_/Q VGND VGND VPWR VPWR _4539_/A sky130_fd_sc_hd__mux2_1
Xhold342 _7526_/X VGND VGND VPWR VPWR _7527_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold353 _7203_/X VGND VGND VPWR VPWR _7204_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold364 _7771_/X VGND VGND VPWR VPWR _7772_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold375 _7166_/X VGND VGND VPWR VPWR _7167_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7257_ _7257_/A VGND VGND VPWR VPWR _9219_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold386 hold386/A VGND VGND VPWR VPWR hold386/X sky130_fd_sc_hd__dlygate4sd3_1
X_4469_ _4475_/A hold64/A VGND VGND VPWR VPWR _4470_/A sky130_fd_sc_hd__or2_1
Xhold397 hold397/A VGND VGND VPWR VPWR hold397/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6208_ _6329_/B VGND VGND VPWR VPWR _6799_/A sky130_fd_sc_hd__buf_2
X_7188_ hold330/X _5465_/A _7192_/S VGND VGND VPWR VPWR _7188_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6139_ _6334_/B _6858_/B VGND VGND VPWR VPWR _6546_/A sky130_fd_sc_hd__nor2_1
Xhold1020 _9530_/Q VGND VGND VPWR VPWR _8653_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1031 _9030_/Q VGND VGND VPWR VPWR _6543_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1042 _5883_/X VGND VGND VPWR VPWR _5884_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1053 _9542_/Q VGND VGND VPWR VPWR _8737_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1064 _5823_/X VGND VGND VPWR VPWR _8988_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1075 _5850_/X VGND VGND VPWR VPWR _5851_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1086 _7471_/X VGND VGND VPWR VPWR _7472_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_204 _8360_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1097 _9380_/Q VGND VGND VPWR VPWR hold310/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_215 _8388_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_226 _9363_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_237 _9070_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_248 wb_dat_i[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_259 _5174_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_5_csclk _9359_/CLK VGND VGND VPWR VPWR _9461_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_123_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5510_ _5510_/A VGND VGND VPWR VPWR _8854_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6490_ _6535_/A _6862_/B VGND VGND VPWR VPWR _6966_/B sky130_fd_sc_hd__nor2_1
XFILLER_9_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5441_ _5441_/A VGND VGND VPWR VPWR _8826_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8160_ _9399_/Q _7977_/X _8159_/X _8008_/B VGND VGND VPWR VPWR _8160_/X sky130_fd_sc_hd__a22o_1
X_5372_ _5372_/A VGND VGND VPWR VPWR _5372_/X sky130_fd_sc_hd__clkbuf_1
X_7111_ _7111_/A _7111_/B _7126_/C VGND VGND VPWR VPWR _7111_/X sky130_fd_sc_hd__or3_1
XFILLER_153_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8091_ _9252_/Q _7940_/X _7969_/X _9292_/Q _8090_/X VGND VGND VPWR VPWR _8097_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_141_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7042_ _7042_/A VGND VGND VPWR VPWR _9125_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8993_ _9370_/CLK _8993_/D fanout477/X VGND VGND VPWR VPWR _9575_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_27_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7944_ _9352_/Q _8020_/A _8034_/A _9232_/Q VGND VGND VPWR VPWR _7944_/X sky130_fd_sc_hd__a22o_1
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7875_ _8996_/Q _7902_/B VGND VGND VPWR VPWR _7875_/X sky130_fd_sc_hd__or2_1
XFILLER_179_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6826_ _6809_/C _6807_/X _6808_/X _6825_/X VGND VGND VPWR VPWR _6826_/X sky130_fd_sc_hd__a31o_1
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9545_ _9550_/CLK _9545_/D fanout500/X VGND VGND VPWR VPWR _9545_/Q sky130_fd_sc_hd__dfrtp_1
X_6757_ _6799_/A _6874_/A _6781_/B _6514_/A _6756_/X VGND VGND VPWR VPWR _6834_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5708_ _5708_/A VGND VGND VPWR VPWR _8939_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9476_ _9476_/CLK _9476_/D fanout414/X VGND VGND VPWR VPWR _9476_/Q sky130_fd_sc_hd__dfrtp_1
X_6688_ _6345_/X _6673_/B _6421_/A _6445_/Y VGND VGND VPWR VPWR _6700_/C sky130_fd_sc_hd__a22o_1
XFILLER_164_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8427_ _8427_/A0 _8426_/X _8653_/S VGND VGND VPWR VPWR _8428_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5639_ _5639_/A VGND VGND VPWR VPWR _8911_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8358_ _8358_/A _8358_/B _8358_/C _8370_/A VGND VGND VPWR VPWR _8361_/C sky130_fd_sc_hd__or4_1
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold150 _5560_/X VGND VGND VPWR VPWR _5561_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7309_ _7233_/X hold560/X _7319_/S VGND VGND VPWR VPWR _7309_/X sky130_fd_sc_hd__mux2_1
Xhold161 _9345_/Q VGND VGND VPWR VPWR hold161/X sky130_fd_sc_hd__dlygate4sd3_1
X_8289_ _8356_/A VGND VGND VPWR VPWR _8289_/X sky130_fd_sc_hd__buf_6
Xhold172 _5702_/X VGND VGND VPWR VPWR _5703_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 _7162_/X VGND VGND VPWR VPWR _7163_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold194 _9470_/Q VGND VGND VPWR VPWR hold194/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5990_ _9066_/Q _4591_/X _5994_/S VGND VGND VPWR VPWR _5991_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4941_ _5281_/A _4811_/A _4734_/Y _4941_/B2 _4940_/X VGND VGND VPWR VPWR _4949_/A
+ sky130_fd_sc_hd__a221o_1
X_7660_ _7660_/A VGND VGND VPWR VPWR _9399_/D sky130_fd_sc_hd__clkbuf_1
X_4872_ hold88/A _7695_/A _7481_/A _9321_/Q _4871_/X VGND VGND VPWR VPWR _4873_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_177_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6611_ _6609_/Y _6610_/X _6967_/A VGND VGND VPWR VPWR _6611_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_32_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7591_ _7556_/X _7591_/A1 hold75/X VGND VGND VPWR VPWR _7592_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9330_ _9370_/CLK _9330_/D fanout477/X VGND VGND VPWR VPWR _9330_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6542_ _6664_/B _6867_/A _6754_/C _6542_/D VGND VGND VPWR VPWR _6542_/X sky130_fd_sc_hd__or4_1
XFILLER_20_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9261_ _9325_/CLK _9261_/D fanout460/X VGND VGND VPWR VPWR _9261_/Q sky130_fd_sc_hd__dfrtp_4
X_6473_ _6589_/C _6828_/A _6665_/B VGND VGND VPWR VPWR _6473_/Y sky130_fd_sc_hd__nor3_1
X_8212_ _9080_/Q _7949_/X _7973_/X _8854_/Q _8211_/X VGND VGND VPWR VPWR _8212_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_145_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5424_ _8819_/Q _5395_/X _5435_/S VGND VGND VPWR VPWR _5424_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9192_ _9272_/CLK _9192_/D fanout422/X VGND VGND VPWR VPWR _9192_/Q sky130_fd_sc_hd__dfstp_1
Xoutput211 _5249_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[13] sky130_fd_sc_hd__buf_12
Xoutput222 _5259_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[23] sky130_fd_sc_hd__buf_12
Xoutput233 _5268_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[33] sky130_fd_sc_hd__buf_12
X_8143_ _9246_/Q _7949_/X _7973_/X _9198_/Q _8142_/X VGND VGND VPWR VPWR _8143_/X
+ sky130_fd_sc_hd__a221o_1
Xoutput244 _5245_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[9] sky130_fd_sc_hd__buf_12
X_5355_ _7025_/A VGND VGND VPWR VPWR _5375_/A sky130_fd_sc_hd__clkbuf_2
Xoutput255 _5173_/A VGND VGND VPWR VPWR pad_flash_io0_ieb sky130_fd_sc_hd__buf_12
XFILLER_99_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput266 _9122_/Q VGND VGND VPWR VPWR pll_div[1] sky130_fd_sc_hd__buf_12
Xoutput277 _8813_/Q VGND VGND VPWR VPWR pll_trim[12] sky130_fd_sc_hd__buf_12
Xoutput288 _9138_/Q VGND VGND VPWR VPWR pll_trim[22] sky130_fd_sc_hd__buf_12
Xoutput299 _8810_/Q VGND VGND VPWR VPWR pll_trim[9] sky130_fd_sc_hd__buf_12
XFILLER_101_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8074_ _9251_/Q _7940_/X _8001_/X _9267_/Q _8073_/X VGND VGND VPWR VPWR _8082_/A
+ sky130_fd_sc_hd__a221o_1
X_5286_ _5286_/A VGND VGND VPWR VPWR _5286_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7025_ _7025_/A _7025_/B VGND VGND VPWR VPWR _7026_/A sky130_fd_sc_hd__and2_1
XFILLER_101_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8976_ _9092_/CLK _8976_/D fanout451/X VGND VGND VPWR VPWR _8976_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_43_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7927_ _7927_/A VGND VGND VPWR VPWR _7927_/X sky130_fd_sc_hd__buf_8
XFILLER_24_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7858_ _8997_/Q _8999_/Q VGND VGND VPWR VPWR _7858_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6809_ _6754_/B _6867_/A _6809_/C _6809_/D VGND VGND VPWR VPWR _6907_/B sky130_fd_sc_hd__and4bb_1
XFILLER_168_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7789_ _7789_/A VGND VGND VPWR VPWR _9459_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9528_ _9532_/CLK _9528_/D fanout448/X VGND VGND VPWR VPWR _9528_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9459_ _9459_/CLK _9459_/D fanout491/X VGND VGND VPWR VPWR _9459_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_70_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _9089_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_109_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_85_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _9462_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout460 fanout461/X VGND VGND VPWR VPWR fanout460/X sky130_fd_sc_hd__clkbuf_4
XFILLER_93_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout471 fanout496/X VGND VGND VPWR VPWR fanout471/X sky130_fd_sc_hd__buf_4
XFILLER_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout482 fanout483/X VGND VGND VPWR VPWR fanout482/X sky130_fd_sc_hd__buf_2
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout493 fanout494/X VGND VGND VPWR VPWR fanout493/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_23_csclk _9210_/CLK VGND VGND VPWR VPWR _9290_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_14_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_38_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _9006_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_183_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold908 _9192_/Q VGND VGND VPWR VPWR hold908/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_127_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold919 _9408_/Q VGND VGND VPWR VPWR hold919/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5140_ _9488_/Q _9490_/Q _9491_/Q _9489_/Q VGND VGND VPWR VPWR _5155_/B sky130_fd_sc_hd__or4b_1
XFILLER_123_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5071_ _9211_/Q _9164_/Q _5071_/C VGND VGND VPWR VPWR _7158_/C sky130_fd_sc_hd__nor3_1
XFILLER_96_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8830_ _8831_/CLK _8830_/D _5449_/X VGND VGND VPWR VPWR hold94/A sky130_fd_sc_hd__dfrtp_4
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8761_ _8760_/X _8761_/A1 _8765_/S VGND VGND VPWR VPWR _8762_/A sky130_fd_sc_hd__mux2_1
X_5973_ _5973_/A VGND VGND VPWR VPWR _9058_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7712_ _7712_/A hold21/A VGND VGND VPWR VPWR hold95/A sky130_fd_sc_hd__nand2_8
X_4924_ _8809_/Q _5388_/A _7032_/A _9121_/Q _4923_/X VGND VGND VPWR VPWR _4931_/A
+ sky130_fd_sc_hd__a221o_1
X_8692_ _8877_/Q _8316_/X _8327_/X _9093_/Q VGND VGND VPWR VPWR _8692_/X sky130_fd_sc_hd__a22o_1
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7643_ _7556_/X _7643_/A1 hold84/X VGND VGND VPWR VPWR _7644_/A sky130_fd_sc_hd__mux2_1
X_4855_ _9281_/Q _7391_/A _5727_/A _8949_/Q _4854_/X VGND VGND VPWR VPWR _4884_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_138_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7574_ _7556_/X _7574_/A1 hold78/X VGND VGND VPWR VPWR _7575_/A sky130_fd_sc_hd__mux2_1
X_4786_ _9386_/Q _4445_/Y _4734_/Y _4786_/B2 _4785_/X VGND VGND VPWR VPWR _4791_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9313_ _9449_/CLK _9313_/D fanout474/X VGND VGND VPWR VPWR _9313_/Q sky130_fd_sc_hd__dfstp_2
X_6525_ _6794_/A _6409_/B _6904_/C VGND VGND VPWR VPWR _6540_/C sky130_fd_sc_hd__o21a_1
X_9244_ _9413_/CLK _9244_/D fanout459/X VGND VGND VPWR VPWR _9244_/Q sky130_fd_sc_hd__dfrtp_2
X_6456_ _6895_/B _6466_/A _6514_/A VGND VGND VPWR VPWR _6468_/B sky130_fd_sc_hd__a21oi_1
XFILLER_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5407_ _8814_/Q _5465_/A _5416_/S VGND VGND VPWR VPWR _5407_/X sky130_fd_sc_hd__mux2_1
X_9175_ _9468_/CLK _9175_/D fanout466/X VGND VGND VPWR VPWR _9175_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6387_ _6973_/A _6839_/B _6721_/A VGND VGND VPWR VPWR _6387_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_88_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8126_ _9309_/Q _8023_/B _7977_/X _9397_/Q _8125_/X VGND VGND VPWR VPWR _8127_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5338_ _5338_/A VGND VGND VPWR VPWR _5338_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_125_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8057_ _9402_/Q _7931_/A _7933_/A _9338_/Q VGND VGND VPWR VPWR _8057_/X sky130_fd_sc_hd__a22o_1
XFILLER_102_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5269_ _9459_/Q VGND VGND VPWR VPWR _5269_/Y sky130_fd_sc_hd__inv_2
X_7008_ _7008_/A _7008_/B _6982_/X VGND VGND VPWR VPWR _7008_/X sky130_fd_sc_hd__or3b_1
XFILLER_141_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8959_ _9088_/CLK _8959_/D fanout454/X VGND VGND VPWR VPWR _8959_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_188_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4640_ _4667_/A _4685_/B VGND VGND VPWR VPWR _5518_/A sky130_fd_sc_hd__nor2_8
XFILLER_30_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4571_ input8/X _4406_/Y _5418_/A _8822_/Q _4570_/X VGND VGND VPWR VPWR _4571_/X
+ sky130_fd_sc_hd__a221o_1
Xmax_cap402 _4550_/S VGND VGND VPWR VPWR _4886_/S sky130_fd_sc_hd__clkbuf_2
X_6310_ _6795_/A _6507_/A _6314_/C VGND VGND VPWR VPWR _6362_/C sky130_fd_sc_hd__and3_1
XFILLER_190_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold705 hold705/A VGND VGND VPWR VPWR _7134_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7290_ _7290_/A VGND VGND VPWR VPWR _9234_/D sky130_fd_sc_hd__clkbuf_1
Xhold716 _9215_/Q VGND VGND VPWR VPWR hold716/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold727 hold727/A VGND VGND VPWR VPWR hold727/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold738 _9487_/Q VGND VGND VPWR VPWR hold738/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold749 hold749/A VGND VGND VPWR VPWR hold749/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6241_ _6279_/A _6241_/B VGND VGND VPWR VPWR _6568_/A sky130_fd_sc_hd__nor2_1
XFILLER_171_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6172_ _6317_/B _6318_/A _6415_/A VGND VGND VPWR VPWR _6297_/A sky130_fd_sc_hd__a21oi_2
XFILLER_130_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5123_ input155/X input154/X _5123_/C _5123_/D VGND VGND VPWR VPWR _5125_/C sky130_fd_sc_hd__and4bb_1
XFILLER_85_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5054_ _5054_/A VGND VGND VPWR VPWR _8787_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8813_ _9484_/CLK _8813_/D fanout428/X VGND VGND VPWR VPWR _8813_/Q sky130_fd_sc_hd__dfrtp_2
X_8744_ _5271_/A _8744_/A2 _8744_/B1 _8727_/Y _8743_/X VGND VGND VPWR VPWR _8744_/X
+ sky130_fd_sc_hd__a221o_1
X_5956_ _5650_/X hold674/X _5958_/S VGND VGND VPWR VPWR _5956_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4907_ _9312_/Q _7463_/A _5573_/A _8883_/Q VGND VGND VPWR VPWR _4907_/X sky130_fd_sc_hd__a22o_1
XFILLER_33_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8675_ _8675_/A _8675_/B _8675_/C _8675_/D VGND VGND VPWR VPWR _8676_/C sky130_fd_sc_hd__or4_1
X_5887_ _5887_/A VGND VGND VPWR VPWR _9012_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4838_ _9249_/Q _7321_/A _5540_/A _8869_/Q _4837_/X VGND VGND VPWR VPWR _4841_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7626_ _7556_/X hold90/X _7638_/S VGND VGND VPWR VPWR hold91/A sky130_fd_sc_hd__mux2_1
XFILLER_138_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7557_ _7556_/X _9353_/Q hold99/X VGND VGND VPWR VPWR _7557_/X sky130_fd_sc_hd__mux2_1
X_4769_ _9370_/Q _7588_/A _7211_/A _9202_/Q _4768_/X VGND VGND VPWR VPWR _4772_/C
+ sky130_fd_sc_hd__a221o_1
X_6508_ _6508_/A _6508_/B VGND VGND VPWR VPWR _6508_/Y sky130_fd_sc_hd__nand2_1
XFILLER_106_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7488_ _7433_/X _9323_/Q _7497_/S VGND VGND VPWR VPWR _7488_/X sky130_fd_sc_hd__mux2_1
X_9227_ _9227_/CLK _9227_/D fanout467/X VGND VGND VPWR VPWR _9227_/Q sky130_fd_sc_hd__dfrtp_4
X_6439_ _6518_/A _6862_/A VGND VGND VPWR VPWR _6462_/B sky130_fd_sc_hd__nor2_4
XFILLER_162_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9158_ _9162_/CLK _9158_/D fanout440/X VGND VGND VPWR VPWR _9158_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8109_ _9205_/Q _7938_/X _7960_/X _9373_/Q VGND VGND VPWR VPWR _8109_/X sky130_fd_sc_hd__a22o_1
XFILLER_121_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold10 hold10/A VGND VGND VPWR VPWR hold10/X sky130_fd_sc_hd__dlygate4sd3_1
X_9089_ _9089_/CLK _9089_/D fanout434/X VGND VGND VPWR VPWR _9089_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_29_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold21 hold21/A VGND VGND VPWR VPWR hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A VGND VGND VPWR VPWR hold32/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold43 hold43/A VGND VGND VPWR VPWR hold43/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold54 hold54/A VGND VGND VPWR VPWR hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A VGND VGND VPWR VPWR hold65/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold76 hold76/A VGND VGND VPWR VPWR hold7/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold87/A VGND VGND VPWR VPWR hold87/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold98 hold98/A VGND VGND VPWR VPWR hold98/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_7 _9077_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5810_ hold526/X _5809_/X _5816_/S VGND VGND VPWR VPWR _5811_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6790_ _6790_/A _6790_/B _6790_/C VGND VGND VPWR VPWR _6791_/A sky130_fd_sc_hd__and3_1
XFILLER_34_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5741_ _5633_/X hold850/X _5747_/S VGND VGND VPWR VPWR _5742_/A sky130_fd_sc_hd__mux2_1
XFILLER_187_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8460_ _9315_/Q _8372_/X _8369_/X _9323_/Q _8459_/X VGND VGND VPWR VPWR _8460_/X
+ sky130_fd_sc_hd__a221o_1
X_5672_ _5647_/X hold577/X _5676_/S VGND VGND VPWR VPWR _5673_/A sky130_fd_sc_hd__mux2_1
X_7411_ _7359_/X hold389/X _7423_/S VGND VGND VPWR VPWR _7412_/A sky130_fd_sc_hd__mux2_1
X_4623_ _9388_/Q _4445_/Y _5762_/A _8967_/Q VGND VGND VPWR VPWR _4623_/X sky130_fd_sc_hd__a22o_1
X_8391_ _8391_/A VGND VGND VPWR VPWR _8391_/X sky130_fd_sc_hd__buf_4
XFILLER_129_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7342_ _7147_/X hold119/X _7354_/S VGND VGND VPWR VPWR _7342_/X sky130_fd_sc_hd__mux2_1
X_4554_ _9373_/Q _4485_/Y _7623_/A _9389_/Q _4553_/X VGND VGND VPWR VPWR _4573_/A
+ sky130_fd_sc_hd__a221o_1
Xhold502 _5636_/X VGND VGND VPWR VPWR _5637_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 _6071_/X VGND VGND VPWR VPWR _6072_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold524 _5907_/X VGND VGND VPWR VPWR _9019_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold535 _8900_/Q VGND VGND VPWR VPWR hold535/X sky130_fd_sc_hd__dlygate4sd3_1
X_7273_ _7236_/X _9227_/Q _7282_/S VGND VGND VPWR VPWR _7273_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4485_ _4674_/A _5474_/B VGND VGND VPWR VPWR _4485_/Y sky130_fd_sc_hd__nor2_4
Xhold546 hold546/A VGND VGND VPWR VPWR hold546/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold557 _9544_/Q VGND VGND VPWR VPWR hold557/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9012_ _9181_/CLK _9012_/D fanout488/X VGND VGND VPWR VPWR _9557_/A sky130_fd_sc_hd__dfrtp_4
Xhold568 _7174_/X VGND VGND VPWR VPWR _7175_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold579 _9050_/Q VGND VGND VPWR VPWR hold579/X sky130_fd_sc_hd__dlygate4sd3_1
X_6224_ _6249_/A VGND VGND VPWR VPWR _6967_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6155_ _6151_/Y _6152_/X _6392_/A VGND VGND VPWR VPWR _6156_/B sky130_fd_sc_hd__a21oi_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1202 _7140_/X VGND VGND VPWR VPWR hold867/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _9251_/Q VGND VGND VPWR VPWR _5106_/Y sky130_fd_sc_hd__inv_2
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1213 _5886_/X VGND VGND VPWR VPWR hold200/A sky130_fd_sc_hd__dlygate4sd3_1
X_6086_ _6891_/A _6317_/A _6167_/B _6167_/C VGND VGND VPWR VPWR _6095_/B sky130_fd_sc_hd__o211a_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1224 _8903_/Q VGND VGND VPWR VPWR hold923/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1235 _8904_/Q VGND VGND VPWR VPWR hold525/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1246 _7087_/X VGND VGND VPWR VPWR hold802/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1257 _8869_/Q VGND VGND VPWR VPWR hold532/A sky130_fd_sc_hd__dlygate4sd3_1
X_5037_ _5037_/A VGND VGND VPWR VPWR _8791_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1268 _8926_/Q VGND VGND VPWR VPWR hold395/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1279 _9330_/Q VGND VGND VPWR VPWR hold719/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6988_ _6988_/A _6988_/B _6988_/C VGND VGND VPWR VPWR _6989_/C sky130_fd_sc_hd__or3_1
XFILLER_25_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8727_ _9033_/Q _9032_/Q _9034_/Q VGND VGND VPWR VPWR _8727_/Y sky130_fd_sc_hd__nor3_4
X_5939_ _9044_/Q _8719_/A1 _5945_/S VGND VGND VPWR VPWR _5940_/A sky130_fd_sc_hd__mux2_2
XFILLER_139_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8658_ _8966_/Q _8346_/X _8386_/X _8936_/Q _8657_/X VGND VGND VPWR VPWR _8663_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_178_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7609_ hold114/X _5951_/A _7621_/S VGND VGND VPWR VPWR _7610_/A sky130_fd_sc_hd__mux2_1
X_8589_ _8928_/Q _8398_/B _8344_/X _8893_/Q VGND VGND VPWR VPWR _8589_/X sky130_fd_sc_hd__a22o_1
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput100 sram_ro_data[16] VGND VGND VPWR VPWR _4918_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput111 sram_ro_data[26] VGND VGND VPWR VPWR _4780_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_76_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput122 sram_ro_data[7] VGND VGND VPWR VPWR _4446_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput133 wb_adr_i[11] VGND VGND VPWR VPWR _6080_/C sky130_fd_sc_hd__clkbuf_1
Xinput144 wb_adr_i[21] VGND VGND VPWR VPWR _6192_/A sky130_fd_sc_hd__clkbuf_2
Xinput155 wb_adr_i[31] VGND VGND VPWR VPWR input155/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput166 wb_dat_i[11] VGND VGND VPWR VPWR _8747_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput177 wb_dat_i[21] VGND VGND VPWR VPWR _8756_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput188 wb_dat_i[31] VGND VGND VPWR VPWR _8763_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput199 wb_sel_i[2] VGND VGND VPWR VPWR _8732_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_76_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7960_ _7960_/A VGND VGND VPWR VPWR _7960_/X sky130_fd_sc_hd__buf_8
XFILLER_54_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6911_ _6911_/A _6911_/B _6911_/C VGND VGND VPWR VPWR _6912_/A sky130_fd_sc_hd__or3_1
XFILLER_82_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7891_ _7891_/A VGND VGND VPWR VPWR _9497_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6842_ _6882_/B _6842_/B VGND VGND VPWR VPWR _6843_/D sky130_fd_sc_hd__nor2_1
XFILLER_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9561_ _9561_/A _5107_/Y VGND VGND VPWR VPWR mgmt_gpio_out[7] sky130_fd_sc_hd__ebufn_8
X_6773_ _6481_/A _6768_/A _6693_/Y _6772_/Y VGND VGND VPWR VPWR _6983_/A sky130_fd_sc_hd__a31o_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5724_ hold485/X _5690_/X _5724_/S VGND VGND VPWR VPWR _5725_/A sky130_fd_sc_hd__mux2_1
X_8512_ _8512_/A _8512_/B _8512_/C _8512_/D VGND VGND VPWR VPWR _8512_/X sky130_fd_sc_hd__or4_1
X_9492_ _9520_/CLK _9492_/D fanout469/X VGND VGND VPWR VPWR _9492_/Q sky130_fd_sc_hd__dfrtp_4
X_8443_ _9386_/Q _8292_/X _8294_/X _9290_/Q VGND VGND VPWR VPWR _8443_/X sky130_fd_sc_hd__a22o_1
X_5655_ _5655_/A VGND VGND VPWR VPWR _8917_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4606_ _4656_/A _4891_/B VGND VGND VPWR VPWR _5618_/A sky130_fd_sc_hd__nor2_8
XFILLER_148_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8374_ _9472_/Q _8367_/X _8369_/X _9320_/Q _8373_/X VGND VGND VPWR VPWR _8396_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_191_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5586_ _5586_/A VGND VGND VPWR VPWR _8888_/D sky130_fd_sc_hd__clkbuf_1
Xhold310 hold310/A VGND VGND VPWR VPWR hold310/X sky130_fd_sc_hd__dlygate4sd3_1
X_7325_ hold108/X _5951_/A _7337_/S VGND VGND VPWR VPWR _7326_/A sky130_fd_sc_hd__mux2_1
Xhold321 _7845_/X VGND VGND VPWR VPWR _7846_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4537_ _7126_/A _7126_/B VGND VGND VPWR VPWR _7113_/A sky130_fd_sc_hd__nor2_8
XFILLER_190_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold332 _9317_/Q VGND VGND VPWR VPWR hold332/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold343 _7561_/X VGND VGND VPWR VPWR _7562_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold354 hold354/A VGND VGND VPWR VPWR hold354/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 _7506_/X VGND VGND VPWR VPWR _7507_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7256_ _7236_/X _9219_/Q _7264_/S VGND VGND VPWR VPWR _7256_/X sky130_fd_sc_hd__mux2_1
X_4468_ hold10/X _4468_/B VGND VGND VPWR VPWR _4475_/A sky130_fd_sc_hd__nand2_1
XFILLER_132_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold376 _7702_/X VGND VGND VPWR VPWR _7703_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 hold387/A VGND VGND VPWR VPWR hold387/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 hold398/A VGND VGND VPWR VPWR hold398/X sky130_fd_sc_hd__dlygate4sd3_1
X_6207_ _6262_/A _6558_/B VGND VGND VPWR VPWR _6329_/B sky130_fd_sc_hd__or2_1
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7187_ _7187_/A VGND VGND VPWR VPWR _9188_/D sky130_fd_sc_hd__clkbuf_1
X_4399_ _9154_/Q _7091_/A _7228_/A _9215_/Q _4398_/X VGND VGND VPWR VPWR _4431_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_58_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6138_ _6341_/A VGND VGND VPWR VPWR _6334_/B sky130_fd_sc_hd__clkbuf_4
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1010 _9493_/Q VGND VGND VPWR VPWR _7876_/B1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 _9502_/Q VGND VGND VPWR VPWR _7910_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1032 _9032_/Q VGND VGND VPWR VPWR _5871_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1043 _9361_/Q VGND VGND VPWR VPWR _7574_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_6069_ hold556/X _5809_/X _6075_/S VGND VGND VPWR VPWR _6070_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1054 _8786_/Q VGND VGND VPWR VPWR hold26/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1065 _5840_/X VGND VGND VPWR VPWR _5841_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1076 _5851_/X VGND VGND VPWR VPWR _9001_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1087 _7578_/X VGND VGND VPWR VPWR _7579_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_205 _8360_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1098 _7615_/X VGND VGND VPWR VPWR _7616_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_216 _8657_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_227 _8964_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_238 _9240_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_249 wb_dat_i[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5440_ _5301_/X _8826_/Q _5440_/S VGND VGND VPWR VPWR _5440_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5371_ _5375_/A _5378_/B VGND VGND VPWR VPWR _5372_/A sky130_fd_sc_hd__and2_1
XFILLER_114_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7110_ _7110_/A VGND VGND VPWR VPWR _7110_/X sky130_fd_sc_hd__clkbuf_1
X_8090_ _9284_/Q _7953_/B _8003_/X _9300_/Q VGND VGND VPWR VPWR _8090_/X sky130_fd_sc_hd__a22o_1
XFILLER_153_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7041_ _6018_/X _9125_/Q _7041_/S VGND VGND VPWR VPWR _7041_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8992_ _9427_/CLK _8992_/D fanout478/X VGND VGND VPWR VPWR _9574_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_103_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7943_ _8275_/B _7996_/B _8002_/B VGND VGND VPWR VPWR _8034_/A sky130_fd_sc_hd__and3_4
XFILLER_36_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7874_ _9493_/Q _9492_/Q VGND VGND VPWR VPWR _7989_/B sky130_fd_sc_hd__and2_4
XFILLER_23_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A VGND VGND VPWR VPWR _9551_/CLK sky130_fd_sc_hd__clkbuf_8
X_6825_ _6907_/B _6824_/X _8735_/A VGND VGND VPWR VPWR _6825_/X sky130_fd_sc_hd__a21o_1
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9544_ _9550_/CLK _9544_/D fanout500/X VGND VGND VPWR VPWR _9544_/Q sky130_fd_sc_hd__dfrtp_1
X_6756_ _6799_/A _6779_/A _6895_/B _6514_/A VGND VGND VPWR VPWR _6756_/X sky130_fd_sc_hd__o22a_1
XFILLER_149_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5707_ hold583/X _5587_/X _5713_/S VGND VGND VPWR VPWR _5708_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9475_ _9475_/CLK _9475_/D fanout482/X VGND VGND VPWR VPWR _9475_/Q sky130_fd_sc_hd__dfrtp_4
X_6687_ _6441_/B _6445_/Y _6937_/A VGND VGND VPWR VPWR _6700_/B sky130_fd_sc_hd__a21o_1
XFILLER_163_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8426_ _9520_/Q _8425_/X _8627_/S VGND VGND VPWR VPWR _8426_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5638_ _5311_/X hold672/X _5640_/S VGND VGND VPWR VPWR _5638_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5569_ hold410/X _5398_/X _5571_/S VGND VGND VPWR VPWR _5570_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8357_ _8357_/A _8357_/B _8389_/C VGND VGND VPWR VPWR _8370_/A sky130_fd_sc_hd__and3_2
XFILLER_128_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold140 _6019_/X VGND VGND VPWR VPWR _6020_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 _9157_/Q VGND VGND VPWR VPWR hold151/X sky130_fd_sc_hd__dlygate4sd3_1
X_7308_ _7308_/A VGND VGND VPWR VPWR _9241_/D sky130_fd_sc_hd__clkbuf_1
Xhold162 _8917_/Q VGND VGND VPWR VPWR hold162/X sky130_fd_sc_hd__dlygate4sd3_1
X_8288_ _8392_/A _8357_/A _8392_/C VGND VGND VPWR VPWR _8356_/A sky130_fd_sc_hd__and3_2
Xhold173 _8982_/Q VGND VGND VPWR VPWR hold173/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold184 _9460_/Q VGND VGND VPWR VPWR hold184/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 _7811_/X VGND VGND VPWR VPWR _7812_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7239_ hold24/X VGND VGND VPWR VPWR _7239_/X sky130_fd_sc_hd__buf_6
XFILLER_104_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4940_ _9448_/Q _7764_/A _4406_/Y input34/X VGND VGND VPWR VPWR _4940_/X sky130_fd_sc_hd__a22o_1
XFILLER_91_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4871_ input21/X _4460_/Y _4734_/Y _4871_/B2 VGND VGND VPWR VPWR _4871_/X sky130_fd_sc_hd__a22o_1
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6610_ _6610_/A _6610_/B VGND VGND VPWR VPWR _6610_/X sky130_fd_sc_hd__or2_1
XFILLER_177_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7590_ _7590_/A VGND VGND VPWR VPWR _9368_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6541_ _6978_/A _6541_/B VGND VGND VPWR VPWR _6542_/D sky130_fd_sc_hd__nand2_1
XFILLER_193_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9260_ _9328_/CLK _9260_/D fanout463/X VGND VGND VPWR VPWR _9260_/Q sky130_fd_sc_hd__dfrtp_1
X_6472_ _6668_/A _6477_/A VGND VGND VPWR VPWR _6665_/B sky130_fd_sc_hd__or2_1
XFILLER_118_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5423_ _5423_/A VGND VGND VPWR VPWR _8818_/D sky130_fd_sc_hd__clkbuf_1
X_8211_ _9090_/Q _7958_/X _8224_/B _8959_/Q VGND VGND VPWR VPWR _8211_/X sky130_fd_sc_hd__a22o_1
X_9191_ _9486_/CLK _9191_/D fanout416/X VGND VGND VPWR VPWR _9191_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_145_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput212 _5250_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[14] sky130_fd_sc_hd__buf_12
Xoutput223 _5260_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[24] sky130_fd_sc_hd__buf_12
Xoutput234 _5269_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[34] sky130_fd_sc_hd__buf_12
X_5354_ _5354_/A VGND VGND VPWR VPWR _5354_/X sky130_fd_sc_hd__clkbuf_1
X_8142_ _9262_/Q _7958_/X _8224_/B _9422_/Q VGND VGND VPWR VPWR _8142_/X sky130_fd_sc_hd__a22o_1
Xoutput245 _5218_/X VGND VGND VPWR VPWR mgmt_gpio_out[0] sky130_fd_sc_hd__buf_12
Xoutput256 _5173_/Y VGND VGND VPWR VPWR pad_flash_io0_oeb sky130_fd_sc_hd__buf_12
Xoutput267 _9123_/Q VGND VGND VPWR VPWR pll_div[2] sky130_fd_sc_hd__buf_12
Xoutput278 _8814_/Q VGND VGND VPWR VPWR pll_trim[13] sky130_fd_sc_hd__buf_12
X_8073_ _9283_/Q _7953_/B _8003_/X _9299_/Q VGND VGND VPWR VPWR _8073_/X sky130_fd_sc_hd__a22o_1
Xoutput289 _9139_/Q VGND VGND VPWR VPWR pll_trim[23] sky130_fd_sc_hd__buf_12
X_5285_ _9169_/Q _5285_/B VGND VGND VPWR VPWR _5286_/A sky130_fd_sc_hd__and2_1
X_7024_ _7024_/A VGND VGND VPWR VPWR _7024_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8975_ _9243_/CLK _8975_/D fanout469/X VGND VGND VPWR VPWR _8975_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_55_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7926_ _8206_/B _7991_/B _7996_/B VGND VGND VPWR VPWR _7927_/A sky130_fd_sc_hd__and3_2
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7857_ _7863_/D VGND VGND VPWR VPWR _7857_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_4_csclk _9359_/CLK VGND VGND VPWR VPWR _9464_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6808_ _6248_/A _6479_/A _6891_/B _6377_/X VGND VGND VPWR VPWR _6808_/X sky130_fd_sc_hd__o31a_1
XFILLER_23_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7788_ _7648_/X _9459_/Q _7796_/S VGND VGND VPWR VPWR _7788_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9527_ _9529_/CLK _9527_/D fanout448/X VGND VGND VPWR VPWR _9527_/Q sky130_fd_sc_hd__dfrtp_1
X_6739_ _6739_/A _6739_/B VGND VGND VPWR VPWR _6739_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9458_ _9474_/CLK _9458_/D fanout427/X VGND VGND VPWR VPWR _9458_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8409_ _9313_/Q _8372_/X _8369_/X _9321_/Q _8408_/X VGND VGND VPWR VPWR _8409_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_124_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9389_ _9469_/CLK _9389_/D fanout458/X VGND VGND VPWR VPWR _9389_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_152_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout450 fanout456/X VGND VGND VPWR VPWR fanout450/X sky130_fd_sc_hd__buf_4
Xfanout461 fanout462/X VGND VGND VPWR VPWR fanout461/X sky130_fd_sc_hd__buf_4
XFILLER_171_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout472 fanout496/X VGND VGND VPWR VPWR fanout472/X sky130_fd_sc_hd__buf_2
XFILLER_59_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout483 fanout496/X VGND VGND VPWR VPWR fanout483/X sky130_fd_sc_hd__clkbuf_2
XFILLER_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout494 fanout495/X VGND VGND VPWR VPWR fanout494/X sky130_fd_sc_hd__buf_2
XFILLER_74_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold909 _7109_/X VGND VGND VPWR VPWR _7110_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5070_ _5070_/A VGND VGND VPWR VPWR _5330_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_96_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8760_ _5287_/A _8760_/A2 _8760_/B1 _8727_/Y _8759_/X VGND VGND VPWR VPWR _8760_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_18_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5972_ _9058_/Q _4591_/X _5976_/S VGND VGND VPWR VPWR _5973_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7711_ _7711_/A VGND VGND VPWR VPWR _9423_/D sky130_fd_sc_hd__clkbuf_1
X_4923_ _8893_/Q _5596_/A _5762_/A _8963_/Q VGND VGND VPWR VPWR _4923_/X sky130_fd_sc_hd__a22o_1
XFILLER_52_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8691_ _8912_/Q _8348_/X _8411_/X _8927_/Q _8690_/X VGND VGND VPWR VPWR _8701_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7642_ _7642_/A VGND VGND VPWR VPWR _9392_/D sky130_fd_sc_hd__clkbuf_1
X_4854_ _9185_/Q _7176_/A _5678_/A _8929_/Q VGND VGND VPWR VPWR _4854_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4785_ _8920_/Q _5656_/A _7077_/A _9143_/Q VGND VGND VPWR VPWR _4785_/X sky130_fd_sc_hd__a22o_1
X_7573_ _7573_/A VGND VGND VPWR VPWR _9360_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9312_ _9416_/CLK _9312_/D fanout461/X VGND VGND VPWR VPWR _9312_/Q sky130_fd_sc_hd__dfstp_1
X_6524_ _6906_/C _6524_/B _6524_/C VGND VGND VPWR VPWR _6904_/C sky130_fd_sc_hd__or3_1
XFILLER_109_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9243_ _9243_/CLK _9243_/D fanout469/X VGND VGND VPWR VPWR _9243_/Q sky130_fd_sc_hd__dfrtp_4
X_6455_ _6455_/A _6643_/A _6455_/C _6455_/D VGND VGND VPWR VPWR _6468_/A sky130_fd_sc_hd__or4_1
X_5406_ hold15/X VGND VGND VPWR VPWR _5465_/A sky130_fd_sc_hd__buf_4
X_9174_ _9468_/CLK _9174_/D fanout466/X VGND VGND VPWR VPWR _9174_/Q sky130_fd_sc_hd__dfrtp_1
X_6386_ _6716_/A _6672_/B VGND VGND VPWR VPWR _6691_/A sky130_fd_sc_hd__xnor2_1
XFILLER_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8125_ _9213_/Q _7923_/X _7973_/X _9197_/Q VGND VGND VPWR VPWR _8125_/X sky130_fd_sc_hd__a22o_1
X_5337_ _5353_/A _5356_/B VGND VGND VPWR VPWR _5338_/A sky130_fd_sc_hd__and2_1
XFILLER_125_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8056_ _9202_/Q _7938_/A _8077_/A _9346_/Q _8055_/X VGND VGND VPWR VPWR _8059_/C
+ sky130_fd_sc_hd__a221o_1
X_5268_ _9451_/Q VGND VGND VPWR VPWR _5268_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7007_ _6929_/Y _7007_/B _7007_/C VGND VGND VPWR VPWR _7008_/B sky130_fd_sc_hd__and3b_1
X_5199_ _9170_/Q input80/X _5279_/B VGND VGND VPWR VPWR _5200_/A sky130_fd_sc_hd__mux2_4
XFILLER_56_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8958_ _9162_/CLK _8958_/D fanout436/X VGND VGND VPWR VPWR _8958_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_43_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7909_ _7909_/A _7909_/B VGND VGND VPWR VPWR _7909_/Y sky130_fd_sc_hd__nor2_1
X_8889_ _9051_/CLK _8889_/D fanout453/X VGND VGND VPWR VPWR _8889_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4570_ _9357_/Q _7553_/A _7284_/A _9237_/Q VGND VGND VPWR VPWR _4570_/X sky130_fd_sc_hd__a22o_2
XFILLER_156_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap403 hold17/X VGND VGND VPWR VPWR hold18/A sky130_fd_sc_hd__buf_2
XFILLER_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold706 hold706/A VGND VGND VPWR VPWR hold706/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold717 _7247_/X VGND VGND VPWR VPWR _7248_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold728 hold728/A VGND VGND VPWR VPWR hold728/X sky130_fd_sc_hd__dlygate4sd3_1
X_6240_ _6266_/A _6241_/B VGND VGND VPWR VPWR _6857_/B sky130_fd_sc_hd__nor2_1
Xhold739 _7847_/X VGND VGND VPWR VPWR _7848_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6171_ _6504_/A VGND VGND VPWR VPWR _6415_/A sky130_fd_sc_hd__clkinv_2
XFILLER_131_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5122_ _6192_/A _6504_/A _6504_/B _6504_/C VGND VGND VPWR VPWR _6312_/A sky130_fd_sc_hd__a211o_2
XFILLER_69_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5053_ _5055_/A1 hold4/X _5065_/S VGND VGND VPWR VPWR _5054_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8812_ _9474_/CLK _8812_/D fanout427/X VGND VGND VPWR VPWR _8812_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_65_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8743_ _5287_/A _8743_/A2 _8743_/B1 _5275_/A VGND VGND VPWR VPWR _8743_/X sky130_fd_sc_hd__a22o_1
X_5955_ _5955_/A VGND VGND VPWR VPWR _9050_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4906_ _9432_/Q _4906_/A2 _6007_/A _9074_/Q _4905_/X VGND VGND VPWR VPWR _4909_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8674_ _8775_/Q _8304_/X _8324_/X _9082_/Q _8673_/X VGND VGND VPWR VPWR _8675_/D
+ sky130_fd_sc_hd__a221o_1
X_5886_ _9557_/A hold199/X _5898_/S VGND VGND VPWR VPWR _5886_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_84_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _9456_/CLK sky130_fd_sc_hd__clkbuf_16
X_7625_ _7625_/A VGND VGND VPWR VPWR _9384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4837_ _8919_/Q _5656_/A _5296_/A _8773_/Q VGND VGND VPWR VPWR _4837_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7556_ hold37/X VGND VGND VPWR VPWR _7556_/X sky130_fd_sc_hd__clkbuf_2
X_4768_ _9418_/Q _7695_/A _7712_/A _9426_/Q VGND VGND VPWR VPWR _4768_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6507_ _6507_/A _6510_/A VGND VGND VPWR VPWR _6508_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4699_ _8861_/Q _5518_/A _6055_/A _9097_/Q _4698_/X VGND VGND VPWR VPWR _4702_/C
+ sky130_fd_sc_hd__a221o_1
X_7487_ _7487_/A VGND VGND VPWR VPWR _9322_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9226_ _9466_/CLK _9226_/D fanout472/X VGND VGND VPWR VPWR _9226_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_162_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6438_ _6438_/A VGND VGND VPWR VPWR _6862_/A sky130_fd_sc_hd__buf_4
XFILLER_106_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9157_ _9162_/CLK _9157_/D fanout440/X VGND VGND VPWR VPWR _9157_/Q sky130_fd_sc_hd__dfrtp_4
X_6369_ _6402_/A _6955_/B _6364_/X _6955_/A _6664_/B VGND VGND VPWR VPWR _6369_/X
+ sky130_fd_sc_hd__a2111o_1
X_8108_ hold989/X _8017_/X _8106_/X _8107_/X VGND VGND VPWR VPWR _9511_/D sky130_fd_sc_hd__o22a_1
XFILLER_29_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9088_ _9088_/CLK _9088_/D fanout455/X VGND VGND VPWR VPWR _9088_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_102_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold11 hold11/A VGND VGND VPWR VPWR hold11/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 hold94/X VGND VGND VPWR VPWR hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A VGND VGND VPWR VPWR hold33/X sky130_fd_sc_hd__buf_12
XFILLER_48_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8039_ _9185_/Q _8010_/B _8027_/X _8037_/X _8627_/S VGND VGND VPWR VPWR _8039_/X
+ sky130_fd_sc_hd__o221a_1
Xhold44 hold44/A VGND VGND VPWR VPWR hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A VGND VGND VPWR VPWR hold55/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold66 hold66/A VGND VGND VPWR VPWR hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold7/X VGND VGND VPWR VPWR hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A VGND VGND VPWR VPWR hold88/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A VGND VGND VPWR VPWR hold99/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_37_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _9172_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] VGND VGND VPWR VPWR clkbuf_0_mgmt_gpio_in[4]/X
+ sky130_fd_sc_hd__clkbuf_16
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_8 _9129_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5740_ _5740_/A VGND VGND VPWR VPWR _8953_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5671_ _5671_/A VGND VGND VPWR VPWR _8924_/D sky130_fd_sc_hd__clkbuf_1
X_7410_ _7410_/A VGND VGND VPWR VPWR _9288_/D sky130_fd_sc_hd__clkbuf_1
X_4622_ _4665_/A _5453_/B VGND VGND VPWR VPWR _5762_/A sky130_fd_sc_hd__nor2_4
X_8390_ _8657_/B VGND VGND VPWR VPWR _8506_/B sky130_fd_sc_hd__buf_6
XFILLER_128_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4553_ _9485_/Q _7832_/A _7249_/A _9221_/Q VGND VGND VPWR VPWR _4553_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7341_ _7341_/A VGND VGND VPWR VPWR _9256_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold503 _9442_/Q VGND VGND VPWR VPWR hold503/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 _8774_/Q VGND VGND VPWR VPWR hold514/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 hold525/A VGND VGND VPWR VPWR hold525/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4484_ _4858_/B _4675_/B VGND VGND VPWR VPWR _4484_/Y sky130_fd_sc_hd__nor2_4
Xhold536 _5612_/X VGND VGND VPWR VPWR _5613_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7272_ _7272_/A VGND VGND VPWR VPWR _9226_/D sky130_fd_sc_hd__clkbuf_1
Xhold547 _9083_/Q VGND VGND VPWR VPWR hold547/X sky130_fd_sc_hd__dlygate4sd3_1
X_9011_ _9181_/CLK _9011_/D fanout487/X VGND VGND VPWR VPWR _9556_/A sky130_fd_sc_hd__dfrtp_4
Xhold558 _5304_/X VGND VGND VPWR VPWR hold12/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 _8960_/Q VGND VGND VPWR VPWR hold569/X sky130_fd_sc_hd__dlygate4sd3_1
X_6223_ _6790_/A _6266_/A _6881_/A VGND VGND VPWR VPWR _6257_/A sky130_fd_sc_hd__a21oi_1
XFILLER_116_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6154_ _6151_/Y _6153_/Y _6312_/A VGND VGND VPWR VPWR _6392_/A sky130_fd_sc_hd__o21a_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1203 _9484_/Q VGND VGND VPWR VPWR hold573/A sky130_fd_sc_hd__dlygate4sd3_1
X_5105_ _9259_/Q VGND VGND VPWR VPWR _5105_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6085_ _6167_/A VGND VGND VPWR VPWR _6891_/A sky130_fd_sc_hd__buf_4
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1214 _9374_/Q VGND VGND VPWR VPWR hold727/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1225 _9468_/Q VGND VGND VPWR VPWR hold350/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1236 _8853_/Q VGND VGND VPWR VPWR hold917/A sky130_fd_sc_hd__dlygate4sd3_1
X_5036_ _8791_/Q _5067_/B _5036_/S VGND VGND VPWR VPWR _5037_/A sky130_fd_sc_hd__mux2_1
Xhold1247 _9318_/Q VGND VGND VPWR VPWR hold398/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1258 _7084_/X VGND VGND VPWR VPWR hold66/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 _8907_/Q VGND VGND VPWR VPWR hold622/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6987_ _6987_/A _6987_/B _6987_/C _6987_/D VGND VGND VPWR VPWR _6988_/C sky130_fd_sc_hd__or4_1
XFILLER_80_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8726_ _8726_/A VGND VGND VPWR VPWR _9541_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5938_ _5938_/A VGND VGND VPWR VPWR _9043_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8657_ _8971_/Q _8657_/B VGND VGND VPWR VPWR _8657_/X sky130_fd_sc_hd__and2_1
X_5869_ _5869_/A VGND VGND VPWR VPWR _5869_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7608_ _7608_/A VGND VGND VPWR VPWR _9376_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8588_ _8588_/A _8588_/B _8588_/C _8588_/D VGND VGND VPWR VPWR _8588_/X sky130_fd_sc_hd__or4_1
XFILLER_147_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7539_ _7359_/X hold161/X _7551_/S VGND VGND VPWR VPWR _7540_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9209_ _9219_/CLK _9209_/D fanout467/X VGND VGND VPWR VPWR _9209_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_122_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput101 sram_ro_data[17] VGND VGND VPWR VPWR _4880_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput112 sram_ro_data[27] VGND VGND VPWR VPWR _4695_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_103_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput123 sram_ro_data[8] VGND VGND VPWR VPWR _4904_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_76_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput134 wb_adr_i[12] VGND VGND VPWR VPWR _6079_/B sky130_fd_sc_hd__clkbuf_1
Xinput145 wb_adr_i[22] VGND VGND VPWR VPWR _6504_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_103_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput156 wb_adr_i[3] VGND VGND VPWR VPWR _6167_/B sky130_fd_sc_hd__clkbuf_4
Xinput167 wb_dat_i[12] VGND VGND VPWR VPWR _8751_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput178 wb_dat_i[22] VGND VGND VPWR VPWR _8759_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput189 wb_dat_i[3] VGND VGND VPWR VPWR _8748_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_721 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6910_ hold62/A _8735_/A _6942_/A _6886_/X _6909_/X VGND VGND VPWR VPWR _6911_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_47_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7890_ _7875_/X _7920_/B _9497_/Q VGND VGND VPWR VPWR _7891_/A sky130_fd_sc_hd__mux2_1
X_6841_ _6924_/C _6770_/B _6841_/C _6841_/D VGND VGND VPWR VPWR _6846_/B sky130_fd_sc_hd__and4bb_1
XFILLER_23_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9560_ _9560_/A _5108_/Y VGND VGND VPWR VPWR mgmt_gpio_out[6] sky130_fd_sc_hd__ebufn_8
XFILLER_50_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6772_ _6772_/A _6772_/B VGND VGND VPWR VPWR _6772_/Y sky130_fd_sc_hd__nor2_1
X_8511_ _9317_/Q _8372_/X _8369_/X _9325_/Q _8510_/X VGND VGND VPWR VPWR _8512_/D
+ sky130_fd_sc_hd__a221o_1
X_5723_ _5723_/A VGND VGND VPWR VPWR _8946_/D sky130_fd_sc_hd__clkbuf_1
X_9491_ _9532_/CLK _9491_/D fanout441/X VGND VGND VPWR VPWR _9491_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8442_ _9234_/Q _8322_/X _8333_/X _9266_/Q _8441_/X VGND VGND VPWR VPWR _8449_/A
+ sky130_fd_sc_hd__a221o_1
X_5654_ _5653_/X hold162/X _5654_/S VGND VGND VPWR VPWR _5654_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4605_ _9308_/Q _7446_/A _7113_/A _9157_/Q _4604_/X VGND VGND VPWR VPWR _4617_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_176_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8373_ _9248_/Q _8370_/X _8372_/X _9312_/Q VGND VGND VPWR VPWR _8373_/X sky130_fd_sc_hd__a22o_1
XFILLER_175_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5585_ hold939/X _5505_/X _5594_/S VGND VGND VPWR VPWR _5586_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold300 _7777_/X VGND VGND VPWR VPWR _7778_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7324_ _7324_/A VGND VGND VPWR VPWR _9248_/D sky130_fd_sc_hd__clkbuf_1
Xhold311 _9301_/Q VGND VGND VPWR VPWR hold311/X sky130_fd_sc_hd__dlygate4sd3_1
X_4536_ _4555_/A _4536_/B VGND VGND VPWR VPWR _7126_/B sky130_fd_sc_hd__nand2_8
Xhold322 _9190_/Q VGND VGND VPWR VPWR hold322/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold333 _7475_/X VGND VGND VPWR VPWR _7476_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold344 _7052_/X VGND VGND VPWR VPWR _7053_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold355 hold355/A VGND VGND VPWR VPWR _7435_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7255_ _7255_/A VGND VGND VPWR VPWR _9218_/D sky130_fd_sc_hd__clkbuf_1
Xhold366 hold366/A VGND VGND VPWR VPWR hold366/X sky130_fd_sc_hd__dlygate4sd3_1
X_4467_ _4492_/A hold33/X VGND VGND VPWR VPWR _7815_/A sky130_fd_sc_hd__nor2_8
Xhold377 _5433_/X VGND VGND VPWR VPWR _5434_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold388 _8916_/Q VGND VGND VPWR VPWR hold388/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold399 hold399/A VGND VGND VPWR VPWR hold399/X sky130_fd_sc_hd__dlygate4sd3_1
X_6206_ _6232_/B _6309_/A VGND VGND VPWR VPWR _6558_/B sky130_fd_sc_hd__or2_2
X_7186_ hold345/X _5690_/A _7192_/S VGND VGND VPWR VPWR _7187_/A sky130_fd_sc_hd__mux2_1
X_4398_ _9399_/Q _7640_/A _7463_/A _9319_/Q VGND VGND VPWR VPWR _4398_/X sky130_fd_sc_hd__a22o_1
XFILLER_98_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1000 _8788_/Q VGND VGND VPWR VPWR _5050_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6137_ _6794_/A _6811_/A VGND VGND VPWR VPWR _6341_/A sky130_fd_sc_hd__nand2_2
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1011 _9491_/Q VGND VGND VPWR VPWR _7868_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1022 _8807_/Q VGND VGND VPWR VPWR _4970_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1033 _5868_/X VGND VGND VPWR VPWR _5869_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1044 _9393_/Q VGND VGND VPWR VPWR _7643_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_6068_ _6068_/A VGND VGND VPWR VPWR _9099_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1055 _8801_/Q VGND VGND VPWR VPWR _5000_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 _5841_/X VGND VGND VPWR VPWR _8994_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1077 _5837_/X VGND VGND VPWR VPWR _5838_/A sky130_fd_sc_hd__dlygate4sd3_1
X_5019_ _5019_/A VGND VGND VPWR VPWR _5019_/Y sky130_fd_sc_hd__inv_2
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1088 _7649_/X VGND VGND VPWR VPWR _7650_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1099 _8942_/Q VGND VGND VPWR VPWR hold616/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_206 _8310_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_217 _8657_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_228 _9394_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_239 _8797_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8709_ _9026_/Q _8709_/B VGND VGND VPWR VPWR _8710_/A sky130_fd_sc_hd__and2_1
XFILLER_9_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5370_ _5370_/A VGND VGND VPWR VPWR _5370_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7040_ _7040_/A VGND VGND VPWR VPWR _9124_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8991_ _9006_/CLK _8991_/D fanout494/X VGND VGND VPWR VPWR _9573_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_27_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7942_ _7998_/A _7996_/B _7992_/C VGND VGND VPWR VPWR _8020_/A sky130_fd_sc_hd__and3_2
XFILLER_36_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7873_ _9493_/Q _9492_/Q VGND VGND VPWR VPWR _7991_/B sky130_fd_sc_hd__nor2_8
XFILLER_51_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6824_ _6824_/A _6824_/B _6824_/C _6824_/D VGND VGND VPWR VPWR _6824_/X sky130_fd_sc_hd__or4_1
XFILLER_50_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9543_ _9551_/CLK _9543_/D fanout500/X VGND VGND VPWR VPWR hold68/A sky130_fd_sc_hd__dfrtp_1
X_6755_ _6895_/B _6781_/B _6830_/A VGND VGND VPWR VPWR _6758_/C sky130_fd_sc_hd__a21oi_1
XFILLER_50_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5706_ _5706_/A VGND VGND VPWR VPWR _8938_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9474_ _9474_/CLK _9474_/D fanout429/X VGND VGND VPWR VPWR _9474_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6686_ _6345_/X _6230_/X _6844_/B VGND VGND VPWR VPWR _6700_/A sky130_fd_sc_hd__a21o_1
X_8425_ _8404_/X _8410_/X _8424_/X _8400_/B _9185_/Q VGND VGND VPWR VPWR _8425_/X
+ sky130_fd_sc_hd__o32a_1
X_5637_ _5637_/A VGND VGND VPWR VPWR _8910_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8356_ _8356_/A _8356_/B _8356_/C _8367_/A VGND VGND VPWR VPWR _8361_/B sky130_fd_sc_hd__or4_1
X_5568_ _5568_/A VGND VGND VPWR VPWR _8880_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold130 _5782_/X VGND VGND VPWR VPWR _5783_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7307_ _7147_/X hold268/X _7319_/S VGND VGND VPWR VPWR _7307_/X sky130_fd_sc_hd__mux2_1
Xhold141 _8872_/Q VGND VGND VPWR VPWR hold141/X sky130_fd_sc_hd__dlygate4sd3_1
X_4519_ _8815_/Q _5388_/A _7228_/A _9214_/Q VGND VGND VPWR VPWR _4519_/X sky130_fd_sc_hd__a22o_1
XFILLER_105_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold152 _7114_/X VGND VGND VPWR VPWR _7115_/A sky130_fd_sc_hd__dlygate4sd3_1
X_8287_ _9500_/Q _9499_/Q VGND VGND VPWR VPWR _8392_/C sky130_fd_sc_hd__nor2_4
X_5499_ _5499_/A VGND VGND VPWR VPWR _8850_/D sky130_fd_sc_hd__clkbuf_1
Xhold163 _5654_/X VGND VGND VPWR VPWR _5655_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold174 _5804_/X VGND VGND VPWR VPWR _5805_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _7790_/X VGND VGND VPWR VPWR _7791_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7238_ _7238_/A VGND VGND VPWR VPWR _9211_/D sky130_fd_sc_hd__clkbuf_1
Xhold196 hold196/A VGND VGND VPWR VPWR hold196/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7169_ _7169_/A VGND VGND VPWR VPWR _7169_/X sky130_fd_sc_hd__clkbuf_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4870_ input44/X _4582_/A _5738_/A _8954_/Q _4869_/X VGND VGND VPWR VPWR _4873_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6540_ _6517_/X _6523_/X _6540_/C _6540_/D VGND VGND VPWR VPWR _6541_/B sky130_fd_sc_hd__and4bb_1
XFILLER_185_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6471_ _6721_/A _6775_/B _6471_/C VGND VGND VPWR VPWR _6477_/A sky130_fd_sc_hd__or3_1
XFILLER_173_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8210_ _9070_/Q _7979_/X _7993_/X _8984_/Q VGND VGND VPWR VPWR _8210_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5422_ _8818_/Q _5392_/X _5435_/S VGND VGND VPWR VPWR _5422_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9190_ _9288_/CLK _9190_/D fanout425/X VGND VGND VPWR VPWR _9190_/Q sky130_fd_sc_hd__dfrtp_4
Xoutput213 _5251_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[15] sky130_fd_sc_hd__buf_12
Xoutput224 _5261_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[25] sky130_fd_sc_hd__buf_12
X_8141_ _9230_/Q _7979_/X _7993_/X _9390_/Q VGND VGND VPWR VPWR _8141_/X sky130_fd_sc_hd__a22o_1
Xoutput235 _5198_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[35] sky130_fd_sc_hd__buf_12
X_5353_ _5353_/A _5356_/B VGND VGND VPWR VPWR _5354_/A sky130_fd_sc_hd__and2_1
Xoutput246 _5216_/X VGND VGND VPWR VPWR mgmt_gpio_out[1] sky130_fd_sc_hd__buf_12
Xoutput257 _9553_/X VGND VGND VPWR VPWR pad_flash_io1_do sky130_fd_sc_hd__buf_12
Xoutput268 _9124_/Q VGND VGND VPWR VPWR pll_div[3] sky130_fd_sc_hd__buf_12
Xoutput279 _8815_/Q VGND VGND VPWR VPWR pll_trim[14] sky130_fd_sc_hd__buf_12
XFILLER_87_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8072_ _8072_/A _8072_/B _8072_/C _8072_/D VGND VGND VPWR VPWR _8072_/X sky130_fd_sc_hd__or4_2
X_5284_ _5284_/A VGND VGND VPWR VPWR _5284_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7023_ _7025_/A _7025_/B VGND VGND VPWR VPWR _7024_/A sky130_fd_sc_hd__and2_1
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8974_ _9243_/CLK _8974_/D fanout469/X VGND VGND VPWR VPWR _8974_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_55_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7925_ _9495_/Q _7929_/B VGND VGND VPWR VPWR _7996_/B sky130_fd_sc_hd__nor2_4
XFILLER_24_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7856_ _7856_/A VGND VGND VPWR VPWR _9488_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6807_ _6807_/A _6807_/B _6939_/A VGND VGND VPWR VPWR _6807_/X sky130_fd_sc_hd__or3b_1
XFILLER_11_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7787_ _7787_/A VGND VGND VPWR VPWR _9458_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4999_ hold39/A _5040_/B _4997_/Y _4998_/X VGND VGND VPWR VPWR _4999_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9526_ _9529_/CLK _9526_/D fanout447/X VGND VGND VPWR VPWR _9526_/Q sky130_fd_sc_hd__dfrtp_1
X_6738_ _6738_/A _6867_/A _6964_/A VGND VGND VPWR VPWR _6741_/C sky130_fd_sc_hd__or3_1
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9457_ _9473_/CLK _9457_/D fanout430/X VGND VGND VPWR VPWR _9457_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_164_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6669_ _6779_/A _6764_/B VGND VGND VPWR VPWR _6924_/B sky130_fd_sc_hd__nor2_1
XFILLER_136_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8408_ _9297_/Q _8314_/X _8331_/X hold92/A VGND VGND VPWR VPWR _8408_/X sky130_fd_sc_hd__a22o_1
X_9388_ _9468_/CLK _9388_/D fanout466/X VGND VGND VPWR VPWR _9388_/Q sky130_fd_sc_hd__dfrtp_4
X_8339_ _9400_/Q _8331_/X _8333_/X _9264_/Q _8338_/X VGND VGND VPWR VPWR _8351_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_155_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout440 fanout441/X VGND VGND VPWR VPWR fanout440/X sky130_fd_sc_hd__clkbuf_4
XFILLER_48_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout451 fanout453/X VGND VGND VPWR VPWR fanout451/X sky130_fd_sc_hd__buf_4
Xfanout462 fanout498/X VGND VGND VPWR VPWR fanout462/X sky130_fd_sc_hd__clkbuf_4
XFILLER_120_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout473 fanout474/X VGND VGND VPWR VPWR fanout473/X sky130_fd_sc_hd__clkbuf_4
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout484 fanout496/X VGND VGND VPWR VPWR fanout484/X sky130_fd_sc_hd__buf_4
XFILLER_59_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout495 fanout496/X VGND VGND VPWR VPWR fanout495/X sky130_fd_sc_hd__clkbuf_2
XFILLER_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5971_ _5971_/A VGND VGND VPWR VPWR _9057_/D sky130_fd_sc_hd__buf_1
X_7710_ _5415_/X hold643/X _7710_/S VGND VGND VPWR VPWR _7710_/X sky130_fd_sc_hd__mux2_1
X_4922_ _4922_/A _4922_/B _4922_/C _4922_/D VGND VGND VPWR VPWR _4961_/A sky130_fd_sc_hd__or4_1
XFILLER_52_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8690_ _8932_/Q _8398_/B _8344_/X _8897_/Q _8689_/X VGND VGND VPWR VPWR _8690_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_45_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7641_ _7517_/X hold924/X hold84/X VGND VGND VPWR VPWR _7642_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4853_ _4853_/A _4853_/B _4853_/C _4853_/D VGND VGND VPWR VPWR _4885_/B sky130_fd_sc_hd__or4_1
XFILLER_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7572_ _7517_/X hold904/X hold78/X VGND VGND VPWR VPWR _7573_/A sky130_fd_sc_hd__mux2_1
X_4784_ _9402_/Q _7661_/A _5540_/A _8870_/Q _4783_/X VGND VGND VPWR VPWR _4791_/A
+ sky130_fd_sc_hd__a221o_4
X_9311_ _9398_/CLK _9311_/D _5070_/A VGND VGND VPWR VPWR _9311_/Q sky130_fd_sc_hd__dfrtp_2
Xclkbuf_opt_2_0_csclk _8954_/CLK VGND VGND VPWR VPWR clkbuf_opt_2_0_csclk/X sky130_fd_sc_hd__clkbuf_16
X_6523_ _6897_/A _6518_/Y _6857_/C _6657_/B VGND VGND VPWR VPWR _6523_/X sky130_fd_sc_hd__a211o_1
XFILLER_158_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9242_ _9474_/CLK _9242_/D fanout429/X VGND VGND VPWR VPWR _9242_/Q sky130_fd_sc_hd__dfrtp_4
X_6454_ _6759_/B _6844_/A _6657_/A _6648_/A VGND VGND VPWR VPWR _6455_/D sky130_fd_sc_hd__or4b_1
XFILLER_174_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5405_ hold14/X _5405_/A1 _5413_/S VGND VGND VPWR VPWR _5405_/X sky130_fd_sc_hd__mux2_8
X_9173_ _9173_/CLK _9173_/D fanout459/X VGND VGND VPWR VPWR _9173_/Q sky130_fd_sc_hd__dfrtp_1
X_6385_ _6672_/B _6384_/X VGND VGND VPWR VPWR _6470_/A sky130_fd_sc_hd__or2b_1
XFILLER_161_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8124_ _9237_/Q _8034_/X _8224_/B _9421_/Q _8123_/X VGND VGND VPWR VPWR _8127_/C
+ sky130_fd_sc_hd__a221o_1
X_5336_ _5453_/C VGND VGND VPWR VPWR _5356_/B sky130_fd_sc_hd__buf_4
XFILLER_142_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8055_ _9410_/Q _7967_/A _8068_/B _9426_/Q VGND VGND VPWR VPWR _8055_/X sky130_fd_sc_hd__a22o_1
XFILLER_141_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5267_ _9443_/Q VGND VGND VPWR VPWR _5267_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7006_ _7002_/B _7006_/B _7006_/C _7006_/D VGND VGND VPWR VPWR _7007_/C sky130_fd_sc_hd__and4b_1
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5198_ _5198_/A VGND VGND VPWR VPWR _5198_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8957_ _9241_/CLK _8957_/D fanout450/X VGND VGND VPWR VPWR _8957_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_43_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7908_ _7908_/A VGND VGND VPWR VPWR _7908_/X sky130_fd_sc_hd__clkbuf_16
X_8888_ _9051_/CLK _8888_/D fanout444/X VGND VGND VPWR VPWR _8888_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_70_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7839_ _5398_/X _9483_/Q _7847_/S VGND VGND VPWR VPWR _7839_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9509_ _9520_/CLK _9509_/D fanout454/X VGND VGND VPWR VPWR _9509_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold707 _9036_/Q VGND VGND VPWR VPWR hold707/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold718 hold718/A VGND VGND VPWR VPWR hold718/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold729 _5416_/X VGND VGND VPWR VPWR _5417_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6170_ _6182_/A _6170_/B _6170_/C _6170_/D VGND VGND VPWR VPWR _6318_/A sky130_fd_sc_hd__and4_1
Xclkbuf_leaf_3_csclk _9359_/CLK VGND VGND VPWR VPWR _9471_/CLK sky130_fd_sc_hd__clkbuf_16
X_5121_ _5121_/A VGND VGND VPWR VPWR _6504_/A sky130_fd_sc_hd__buf_4
XFILLER_97_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5052_ _5021_/A _5045_/B _5050_/X _5051_/X VGND VGND VPWR VPWR _8788_/D sky130_fd_sc_hd__a211o_1
XFILLER_57_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8811_ _9476_/CLK _8811_/D fanout427/X VGND VGND VPWR VPWR _8811_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_53_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8742_ _8742_/A VGND VGND VPWR VPWR _9543_/D sky130_fd_sc_hd__clkbuf_1
X_5954_ _5647_/X hold579/X _5958_/S VGND VGND VPWR VPWR _5954_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4905_ _8903_/Q _5618_/A _5918_/A _9035_/Q VGND VGND VPWR VPWR _4905_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8673_ _9051_/Q _8289_/X _8341_/X _8891_/Q VGND VGND VPWR VPWR _8673_/X sky130_fd_sc_hd__a22o_1
X_5885_ _9179_/Q _7648_/A _5897_/S VGND VGND VPWR VPWR _5885_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7624_ _7517_/X hold887/X _7638_/S VGND VGND VPWR VPWR _7625_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4836_ _9449_/Q _4836_/A2 _5506_/A _8854_/Q _4835_/X VGND VGND VPWR VPWR _4841_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7555_ _7555_/A VGND VGND VPWR VPWR _9352_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4767_ _9338_/Q _7519_/A _7356_/A _9266_/Q _4766_/X VGND VGND VPWR VPWR _4772_/B
+ sky130_fd_sc_hd__a221o_1
X_6506_ _6655_/C _6508_/B VGND VGND VPWR VPWR _6506_/Y sky130_fd_sc_hd__nor2_1
XFILLER_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7486_ _7430_/X hold722/X _7497_/S VGND VGND VPWR VPWR _7487_/A sky130_fd_sc_hd__mux2_1
X_4698_ _5071_/C _4811_/A _4416_/Y _9203_/Q VGND VGND VPWR VPWR _4698_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9225_ _9465_/CLK _9225_/D fanout471/X VGND VGND VPWR VPWR _9225_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_161_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6437_ _6437_/A _6716_/A _6850_/A VGND VGND VPWR VPWR _6438_/A sky130_fd_sc_hd__or3_1
XFILLER_105_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9156_ _9452_/CLK _9156_/D fanout415/X VGND VGND VPWR VPWR _9156_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6368_ _6479_/A _6895_/B VGND VGND VPWR VPWR _6664_/B sky130_fd_sc_hd__nor2_1
XFILLER_96_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8107_ _5139_/A hold974/X _8013_/X VGND VGND VPWR VPWR _8107_/X sky130_fd_sc_hd__a21o_1
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5319_ _5319_/A VGND VGND VPWR VPWR _5319_/X sky130_fd_sc_hd__clkbuf_1
X_9087_ _9087_/CLK _9087_/D fanout447/X VGND VGND VPWR VPWR _9087_/Q sky130_fd_sc_hd__dfrtp_2
X_6299_ _6345_/B _6547_/B VGND VGND VPWR VPWR _6365_/B sky130_fd_sc_hd__nand2_1
Xhold12 hold12/A VGND VGND VPWR VPWR hold12/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold23 hold23/A VGND VGND VPWR VPWR hold23/X sky130_fd_sc_hd__dlygate4sd3_1
X_8038_ _8652_/S VGND VGND VPWR VPWR _8627_/S sky130_fd_sc_hd__buf_6
XFILLER_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold34 hold34/A VGND VGND VPWR VPWR hold34/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold45 hold45/A VGND VGND VPWR VPWR hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A VGND VGND VPWR VPWR hold56/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold67 hold67/A VGND VGND VPWR VPWR hold67/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold78 hold78/A VGND VGND VPWR VPWR hold78/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold89 hold89/A VGND VGND VPWR VPWR hold89/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_9 _9141_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5670_ _5633_/X hold444/X _5676_/S VGND VGND VPWR VPWR _5671_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4621_ _4635_/A _4794_/B VGND VGND VPWR VPWR _5296_/A sky130_fd_sc_hd__nor2_8
XFILLER_175_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7340_ _7302_/X hold926/X _7354_/S VGND VGND VPWR VPWR _7341_/A sky130_fd_sc_hd__mux2_1
X_4552_ _4552_/A VGND VGND VPWR VPWR _9117_/D sky130_fd_sc_hd__clkbuf_1
Xhold504 _7752_/X VGND VGND VPWR VPWR _7753_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold515 _5307_/X VGND VGND VPWR VPWR _5308_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7271_ _7233_/X hold764/X _7282_/S VGND VGND VPWR VPWR _7272_/A sky130_fd_sc_hd__mux2_1
Xhold526 hold526/A VGND VGND VPWR VPWR hold526/X sky130_fd_sc_hd__dlygate4sd3_1
X_4483_ _4492_/A _7126_/A VGND VGND VPWR VPWR _4483_/Y sky130_fd_sc_hd__nor2_8
Xhold537 _9481_/Q VGND VGND VPWR VPWR hold537/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold548 _6030_/X VGND VGND VPWR VPWR _6031_/A sky130_fd_sc_hd__dlygate4sd3_1
X_9010_ _9464_/CLK _9010_/D fanout420/X VGND VGND VPWR VPWR _9010_/Q sky130_fd_sc_hd__dfrtp_1
Xhold559 _6013_/X VGND VGND VPWR VPWR _6014_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6222_ _6222_/A VGND VGND VPWR VPWR _6881_/A sky130_fd_sc_hd__buf_2
XFILLER_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6153_ _6504_/B _6504_/C VGND VGND VPWR VPWR _6153_/Y sky130_fd_sc_hd__nand2_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5104_ _9267_/Q VGND VGND VPWR VPWR _5104_/Y sky130_fd_sc_hd__inv_2
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ _6084_/A VGND VGND VPWR VPWR _6175_/A sky130_fd_sc_hd__clkbuf_2
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1204 _8948_/Q VGND VGND VPWR VPWR hold831/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1215 _8977_/Q VGND VGND VPWR VPWR hold641/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1226 _9084_/Q VGND VGND VPWR VPWR hold898/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1237 _8964_/Q VGND VGND VPWR VPWR hold553/A sky130_fd_sc_hd__dlygate4sd3_1
X_5035_ _8808_/Q _5035_/B _5068_/B _8827_/Q VGND VGND VPWR VPWR _5036_/S sky130_fd_sc_hd__and4b_1
Xhold1248 _9303_/Q VGND VGND VPWR VPWR hold848/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1259 _8973_/Q VGND VGND VPWR VPWR hold915/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6986_ _6420_/B _6828_/A _6241_/B _6841_/C _6985_/X VGND VGND VPWR VPWR _7007_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5937_ _9043_/Q _4752_/X _5945_/S VGND VGND VPWR VPWR _5938_/A sky130_fd_sc_hd__mux2_1
X_8725_ _9541_/Q _4507_/X _8725_/S VGND VGND VPWR VPWR _8726_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8656_ _8961_/Q _8402_/X _8378_/X _8946_/Q _8655_/X VGND VGND VPWR VPWR _8663_/A
+ sky130_fd_sc_hd__a221o_1
X_5868_ _9007_/Q _5867_/X _5868_/S VGND VGND VPWR VPWR _5868_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7607_ hold878/X _5761_/A _7621_/S VGND VGND VPWR VPWR _7607_/X sky130_fd_sc_hd__mux2_1
X_4819_ _4818_/X hold961/X _4964_/B VGND VGND VPWR VPWR _4819_/X sky130_fd_sc_hd__mux2_1
X_8587_ _9099_/Q _8372_/X _8369_/X _8903_/Q _8586_/X VGND VGND VPWR VPWR _8588_/D
+ sky130_fd_sc_hd__a221o_1
X_5799_ _5799_/A VGND VGND VPWR VPWR _8979_/D sky130_fd_sc_hd__clkbuf_1
X_7538_ _7538_/A VGND VGND VPWR VPWR _9344_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7469_ hold566/X _6048_/X _7479_/S VGND VGND VPWR VPWR _7470_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9208_ _9398_/CLK _9208_/D _5332_/A VGND VGND VPWR VPWR _9208_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_134_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9139_ _9480_/CLK _9139_/D fanout412/X VGND VGND VPWR VPWR _9139_/Q sky130_fd_sc_hd__dfstp_1
Xinput102 sram_ro_data[18] VGND VGND VPWR VPWR _4759_/A1 sky130_fd_sc_hd__buf_2
Xinput113 sram_ro_data[28] VGND VGND VPWR VPWR _4616_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput124 sram_ro_data[9] VGND VGND VPWR VPWR _4821_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput135 wb_adr_i[13] VGND VGND VPWR VPWR _6079_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput146 wb_adr_i[23] VGND VGND VPWR VPWR _6504_/B sky130_fd_sc_hd__clkbuf_1
Xinput157 wb_adr_i[4] VGND VGND VPWR VPWR _6181_/A sky130_fd_sc_hd__buf_4
Xinput168 wb_dat_i[13] VGND VGND VPWR VPWR _8755_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput179 wb_dat_i[23] VGND VGND VPWR VPWR _8764_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_17_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_83_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _9485_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_79_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6840_ _6334_/B _6658_/A _6839_/Y _6665_/B VGND VGND VPWR VPWR _6841_/D sky130_fd_sc_hd__o22a_1
XFILLER_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6771_ _6422_/B _6521_/B _6460_/B _6704_/A _6330_/Y VGND VGND VPWR VPWR _6922_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8510_ _9301_/Q _8314_/X _8331_/X _9405_/Q VGND VGND VPWR VPWR _8510_/X sky130_fd_sc_hd__a22o_1
X_5722_ hold678/X _5687_/X _5724_/S VGND VGND VPWR VPWR _5723_/A sky130_fd_sc_hd__mux2_1
X_9490_ _9531_/CLK _9490_/D fanout441/X VGND VGND VPWR VPWR _9490_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_21_csclk _9210_/CLK VGND VGND VPWR VPWR _9276_/CLK sky130_fd_sc_hd__clkbuf_16
X_8441_ _9282_/Q _8316_/X _8327_/X _9258_/Q VGND VGND VPWR VPWR _8441_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5653_ hold24/X VGND VGND VPWR VPWR _5653_/X sky130_fd_sc_hd__buf_4
XFILLER_175_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4604_ _9356_/Q _4427_/Y _5506_/A _8857_/Q VGND VGND VPWR VPWR _4604_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8372_ _8372_/A VGND VGND VPWR VPWR _8372_/X sky130_fd_sc_hd__buf_6
XFILLER_163_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5584_ _5584_/A _5715_/B VGND VGND VPWR VPWR _5594_/S sky130_fd_sc_hd__and2_2
XFILLER_117_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_36_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _9419_/CLK sky130_fd_sc_hd__clkbuf_16
X_7323_ hold840/X _7126_/C _7337_/S VGND VGND VPWR VPWR _7324_/A sky130_fd_sc_hd__mux2_1
X_4535_ _9398_/Q _7640_/A _4531_/Y _4532_/X _4534_/X VGND VGND VPWR VPWR _4549_/C
+ sky130_fd_sc_hd__a2111o_1
Xhold301 _9325_/Q VGND VGND VPWR VPWR hold301/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 _7440_/X VGND VGND VPWR VPWR _7441_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 _7190_/X VGND VGND VPWR VPWR _7191_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 hold334/A VGND VGND VPWR VPWR hold334/X sky130_fd_sc_hd__dlygate4sd3_1
X_7254_ _7233_/X hold570/X _7264_/S VGND VGND VPWR VPWR _7254_/X sky130_fd_sc_hd__mux2_1
Xhold345 hold345/A VGND VGND VPWR VPWR hold345/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4466_ _4499_/A _7158_/B VGND VGND VPWR VPWR _5418_/A sky130_fd_sc_hd__nor2_8
Xhold356 _9052_/Q VGND VGND VPWR VPWR hold356/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold367 _8843_/Q VGND VGND VPWR VPWR hold367/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold378 hold378/A VGND VGND VPWR VPWR _7840_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 _9289_/Q VGND VGND VPWR VPWR hold389/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6205_ _6178_/A _6178_/B _6232_/C VGND VGND VPWR VPWR _6309_/A sky130_fd_sc_hd__a21bo_1
X_7185_ _7185_/A VGND VGND VPWR VPWR _9187_/D sky130_fd_sc_hd__clkbuf_1
X_4397_ _4656_/A _4748_/B VGND VGND VPWR VPWR _7463_/A sky130_fd_sc_hd__nor2_8
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6136_ _6248_/A _6420_/B VGND VGND VPWR VPWR _6811_/A sky130_fd_sc_hd__nor2_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1001 _9529_/Q VGND VGND VPWR VPWR _8628_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1012 _8792_/Q VGND VGND VPWR VPWR _5032_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1023 _9500_/Q VGND VGND VPWR VPWR _7901_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_6067_ hold894/X _5761_/X _6075_/S VGND VGND VPWR VPWR _6068_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1034 _5869_/X VGND VGND VPWR VPWR _9007_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1045 _9369_/Q VGND VGND VPWR VPWR _7591_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1056 hold76/A VGND VGND VPWR VPWR _5009_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 _5880_/X VGND VGND VPWR VPWR _5881_/A sky130_fd_sc_hd__dlygate4sd3_1
X_5018_ _5018_/A VGND VGND VPWR VPWR _8797_/D sky130_fd_sc_hd__clkbuf_1
Xhold1078 _5838_/X VGND VGND VPWR VPWR _8993_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1089 _7595_/X VGND VGND VPWR VPWR _7596_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_207 _8312_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_218 _8506_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_229 _9424_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6969_ _6969_/A _6969_/B _6969_/C _6968_/X VGND VGND VPWR VPWR _6970_/D sky130_fd_sc_hd__or4b_1
X_8708_ _9533_/Q _8705_/Y _8706_/Y _8707_/X VGND VGND VPWR VPWR _9533_/D sky130_fd_sc_hd__a31o_1
XFILLER_179_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8639_ _8860_/Q _8391_/X _8367_/X _9096_/Q _8638_/X VGND VGND VPWR VPWR _8639_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_167_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold890 hold890/A VGND VGND VPWR VPWR hold890/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8990_ _9006_/CLK _8990_/D fanout494/X VGND VGND VPWR VPWR _9572_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_55_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7941_ _9493_/Q _9492_/Q VGND VGND VPWR VPWR _7992_/C sky130_fd_sc_hd__and2b_4
X_7872_ _7902_/B VGND VGND VPWR VPWR _7920_/B sky130_fd_sc_hd__inv_2
XFILLER_36_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6823_ _6812_/Y _6813_/X _6817_/Y _6821_/X _6822_/X VGND VGND VPWR VPWR _6824_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_51_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6754_ _6754_/A _6754_/B _6754_/C _6382_/X VGND VGND VPWR VPWR _6931_/A sky130_fd_sc_hd__or4b_4
X_9542_ _9550_/CLK _9542_/D fanout499/X VGND VGND VPWR VPWR _9542_/Q sky130_fd_sc_hd__dfrtp_1
X_5705_ hold903/X _5505_/X _5713_/S VGND VGND VPWR VPWR _5706_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9473_ _9473_/CLK _9473_/D fanout431/X VGND VGND VPWR VPWR _9473_/Q sky130_fd_sc_hd__dfstp_1
X_6685_ _6967_/B _6926_/A VGND VGND VPWR VPWR _6844_/B sky130_fd_sc_hd__nor2_1
XFILLER_176_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5636_ _5306_/X hold501/X _5640_/S VGND VGND VPWR VPWR _5636_/X sky130_fd_sc_hd__mux2_1
X_8424_ _8701_/A _8424_/B _8424_/C VGND VGND VPWR VPWR _8424_/X sky130_fd_sc_hd__or3_1
XFILLER_163_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8355_ _8355_/A _8385_/B VGND VGND VPWR VPWR _8367_/A sky130_fd_sc_hd__nor2_4
XFILLER_191_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5567_ hold788/X _5395_/X _5571_/S VGND VGND VPWR VPWR _5568_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7306_ _7306_/A VGND VGND VPWR VPWR _9240_/D sky130_fd_sc_hd__clkbuf_1
Xhold120 _7342_/X VGND VGND VPWR VPWR _7343_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4518_ input59/X _5901_/A _4409_/Y _9262_/Q _4517_/X VGND VGND VPWR VPWR _4521_/C
+ sky130_fd_sc_hd__a221o_1
Xhold131 _8776_/Q VGND VGND VPWR VPWR hold131/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8286_ _9501_/Q _9502_/Q VGND VGND VPWR VPWR _8357_/A sky130_fd_sc_hd__nor2_2
Xhold142 _5549_/X VGND VGND VPWR VPWR _5550_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 _5910_/X VGND VGND VPWR VPWR _5911_/A sky130_fd_sc_hd__dlygate4sd3_1
X_5498_ hold592/X _5395_/X _5502_/S VGND VGND VPWR VPWR _5498_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold164 _7066_/X VGND VGND VPWR VPWR _7067_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 _9441_/Q VGND VGND VPWR VPWR hold175/X sky130_fd_sc_hd__dlygate4sd3_1
X_7237_ _7236_/X _9211_/Q _7247_/S VGND VGND VPWR VPWR _7237_/X sky130_fd_sc_hd__mux2_1
Xhold186 _8862_/Q VGND VGND VPWR VPWR hold186/X sky130_fd_sc_hd__dlygate4sd3_1
X_4449_ _4492_/B _5474_/B VGND VGND VPWR VPWR _4449_/Y sky130_fd_sc_hd__nor2_8
XFILLER_132_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold197 _9545_/Q VGND VGND VPWR VPWR hold197/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7168_ _6018_/X _9180_/Q _7174_/S VGND VGND VPWR VPWR _7168_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6119_ _6192_/A _6312_/A VGND VGND VPWR VPWR _6415_/B sky130_fd_sc_hd__nor2_2
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7099_ _7099_/A VGND VGND VPWR VPWR _9150_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6470_ _6470_/A _6691_/A VGND VGND VPWR VPWR _6775_/B sky130_fd_sc_hd__nand2_1
XFILLER_71_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5421_ _5421_/A VGND VGND VPWR VPWR _8817_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput203 _5282_/X VGND VGND VPWR VPWR debug_in sky130_fd_sc_hd__buf_12
X_8140_ _8140_/A _8140_/B _8140_/C _8140_/D VGND VGND VPWR VPWR _8149_/A sky130_fd_sc_hd__or4_1
XFILLER_160_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5352_ _5352_/A VGND VGND VPWR VPWR _5352_/X sky130_fd_sc_hd__clkbuf_1
Xoutput214 _5252_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[16] sky130_fd_sc_hd__buf_12
Xoutput225 _5185_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[26] sky130_fd_sc_hd__buf_12
Xoutput236 _5195_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[36] sky130_fd_sc_hd__buf_12
Xoutput247 _5204_/X VGND VGND VPWR VPWR mgmt_gpio_out[35] sky130_fd_sc_hd__buf_12
XFILLER_114_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput258 _5176_/Y VGND VGND VPWR VPWR pad_flash_io1_ieb sky130_fd_sc_hd__buf_12
X_8071_ _9331_/Q _7981_/X _7993_/X _9387_/Q _8070_/X VGND VGND VPWR VPWR _8072_/D
+ sky130_fd_sc_hd__a221o_1
Xoutput269 _9125_/Q VGND VGND VPWR VPWR pll_div[4] sky130_fd_sc_hd__buf_12
X_5283_ _9168_/Q _5283_/B VGND VGND VPWR VPWR _5284_/A sky130_fd_sc_hd__and2_1
XFILLER_87_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7022_ _7022_/A VGND VGND VPWR VPWR _7022_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_102_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8973_ _9087_/CLK _8973_/D fanout447/X VGND VGND VPWR VPWR _8973_/Q sky130_fd_sc_hd__dfrtp_4
X_7924_ _8181_/B VGND VGND VPWR VPWR _8206_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_70_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7855_ _7865_/A _7855_/B _7855_/C VGND VGND VPWR VPWR _7856_/A sky130_fd_sc_hd__and3_1
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6806_ _6867_/B _6806_/B _6806_/C _6806_/D VGND VGND VPWR VPWR _6807_/B sky130_fd_sc_hd__or4_1
XFILLER_169_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4998_ _8801_/Q _5002_/B VGND VGND VPWR VPWR _4998_/X sky130_fd_sc_hd__or2_1
X_7786_ _7645_/X hold510/X _7796_/S VGND VGND VPWR VPWR _7786_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9525_ _9529_/CLK _9525_/D fanout451/X VGND VGND VPWR VPWR _9525_/Q sky130_fd_sc_hd__dfrtp_1
X_6737_ _6228_/Y _6860_/B _6608_/Y VGND VGND VPWR VPWR _6856_/B sky130_fd_sc_hd__a21o_1
XFILLER_137_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9456_ _9456_/CLK _9456_/D fanout404/X VGND VGND VPWR VPWR _9456_/Q sky130_fd_sc_hd__dfstp_2
X_6668_ _6668_/A _6775_/B _6695_/A VGND VGND VPWR VPWR _6764_/B sky130_fd_sc_hd__or3_1
XFILLER_192_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5619_ hold923/X _5505_/X _5627_/S VGND VGND VPWR VPWR _5620_/A sky130_fd_sc_hd__mux2_1
X_8407_ _9449_/Q _8310_/X _8381_/X _9361_/Q _8406_/X VGND VGND VPWR VPWR _8407_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_191_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9387_ _9475_/CLK _9387_/D fanout482/X VGND VGND VPWR VPWR _9387_/Q sky130_fd_sc_hd__dfrtp_4
X_6599_ _6419_/A _6597_/A _6597_/B _6340_/Y _6507_/A VGND VGND VPWR VPWR _6851_/C
+ sky130_fd_sc_hd__a32o_1
XFILLER_3_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8338_ _9272_/Q _8335_/X _8337_/X _9376_/Q VGND VGND VPWR VPWR _8338_/X sky130_fd_sc_hd__a22o_1
XFILLER_117_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8269_ _8982_/Q _7931_/X _8268_/X VGND VGND VPWR VPWR _8272_/C sky130_fd_sc_hd__a21o_1
XFILLER_48_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout430 fanout432/X VGND VGND VPWR VPWR fanout430/X sky130_fd_sc_hd__clkbuf_4
Xfanout441 fanout449/X VGND VGND VPWR VPWR fanout441/X sky130_fd_sc_hd__buf_4
Xfanout452 fanout453/X VGND VGND VPWR VPWR fanout452/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout463 fanout464/X VGND VGND VPWR VPWR fanout463/X sky130_fd_sc_hd__clkbuf_4
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout474 fanout496/X VGND VGND VPWR VPWR fanout474/X sky130_fd_sc_hd__clkbuf_4
XFILLER_74_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout485 fanout496/X VGND VGND VPWR VPWR fanout485/X sky130_fd_sc_hd__buf_2
XFILLER_19_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout496 fanout497/X VGND VGND VPWR VPWR fanout496/X sky130_fd_sc_hd__clkbuf_4
XFILLER_19_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5970_ _9057_/Q _8719_/A1 _5976_/S VGND VGND VPWR VPWR _5971_/A sky130_fd_sc_hd__mux2_2
XFILLER_80_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4921_ _4921_/A _4921_/B _4921_/C _4921_/D VGND VGND VPWR VPWR _4922_/D sky130_fd_sc_hd__or4_1
XFILLER_33_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4852_ _4852_/A _4852_/B _4852_/C _4852_/D VGND VGND VPWR VPWR _4853_/D sky130_fd_sc_hd__or4_1
X_7640_ _7640_/A _7695_/B VGND VGND VPWR VPWR hold84/A sky130_fd_sc_hd__nand2_8
XFILLER_33_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_390 _9490_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7571_ _7571_/A _7695_/B VGND VGND VPWR VPWR hold78/A sky130_fd_sc_hd__nand2_8
XFILLER_20_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4783_ _8975_/Q _5784_/A _5642_/A _8915_/Q VGND VGND VPWR VPWR _4783_/X sky130_fd_sc_hd__a22o_1
X_9310_ _9398_/CLK _9310_/D fanout419/X VGND VGND VPWR VPWR _9310_/Q sky130_fd_sc_hd__dfrtp_2
X_6522_ _6926_/B _6528_/B VGND VGND VPWR VPWR _6657_/B sky130_fd_sc_hd__nor2_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9241_ _9241_/CLK _9241_/D fanout467/X VGND VGND VPWR VPWR _9241_/Q sky130_fd_sc_hd__dfstp_1
X_6453_ _6535_/A _6453_/B VGND VGND VPWR VPWR _6648_/A sky130_fd_sc_hd__or2_1
XFILLER_109_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5404_ _5404_/A VGND VGND VPWR VPWR _8813_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9172_ _9172_/CLK _9172_/D fanout494/X VGND VGND VPWR VPWR _9588_/A sky130_fd_sc_hd__dfrtp_1
X_6384_ _6317_/A _6175_/A _6633_/A _6437_/A VGND VGND VPWR VPWR _6384_/X sky130_fd_sc_hd__a31o_1
X_8123_ _9325_/Q _7962_/X _8003_/X _9301_/Q VGND VGND VPWR VPWR _8123_/X sky130_fd_sc_hd__a22o_1
X_5335_ _5335_/A VGND VGND VPWR VPWR _5335_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8054_ _9234_/Q _8034_/A _8052_/X _8053_/X VGND VGND VPWR VPWR _8059_/B sky130_fd_sc_hd__a211o_1
XFILLER_87_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5266_ _9435_/Q VGND VGND VPWR VPWR _5266_/Y sky130_fd_sc_hd__inv_2
X_7005_ _6331_/Y _6566_/B _6455_/A _6643_/A VGND VGND VPWR VPWR _7006_/D sky130_fd_sc_hd__a211oi_1
X_5197_ _5196_/Y input82/X _5279_/B VGND VGND VPWR VPWR _5198_/A sky130_fd_sc_hd__mux2_8
XFILLER_110_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8956_ _9091_/CLK _8956_/D fanout455/X VGND VGND VPWR VPWR _8956_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7907_ _8392_/A _8389_/A _8336_/A VGND VGND VPWR VPWR _7908_/A sky130_fd_sc_hd__and3_2
XFILLER_34_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8887_ _9449_/CLK _8887_/D fanout473/X VGND VGND VPWR VPWR _8887_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_169_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7838_ _7838_/A VGND VGND VPWR VPWR _9482_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7769_ _7645_/X hold488/X _7779_/S VGND VGND VPWR VPWR _7769_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__1160_ clkbuf_0__1160_/X VGND VGND VPWR VPWR _8719_/A1 sky130_fd_sc_hd__clkbuf_16
X_9508_ _9520_/CLK _9508_/D fanout454/X VGND VGND VPWR VPWR _9508_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9439_ _9477_/CLK _9439_/D fanout409/X VGND VGND VPWR VPWR _9439_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_165_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold708 _5921_/X VGND VGND VPWR VPWR _5922_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold719 hold719/A VGND VGND VPWR VPWR hold719/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5120_ _5120_/A _5120_/B _5120_/C _5120_/D VGND VGND VPWR VPWR _5120_/X sky130_fd_sc_hd__or4_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5051_ _5067_/B _5068_/C _5051_/C VGND VGND VPWR VPWR _5051_/X sky130_fd_sc_hd__and3_1
XFILLER_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8810_ _9484_/CLK _8810_/D fanout427/X VGND VGND VPWR VPWR _8810_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_92_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8741_ _8740_/X hold68/X _8765_/S VGND VGND VPWR VPWR _8742_/A sky130_fd_sc_hd__mux2_1
X_5953_ _5953_/A VGND VGND VPWR VPWR _9049_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4904_ _4904_/A1 _4488_/Y _7623_/A _9384_/Q _4903_/X VGND VGND VPWR VPWR _4909_/B
+ sky130_fd_sc_hd__a221o_1
X_5884_ _5884_/A VGND VGND VPWR VPWR _9011_/D sky130_fd_sc_hd__clkbuf_1
X_8672_ _8976_/Q _8337_/X _8384_/X _8856_/Q _8671_/X VGND VGND VPWR VPWR _8675_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7623_ _7623_/A _7695_/B VGND VGND VPWR VPWR _7638_/S sky130_fd_sc_hd__nand2_8
X_4835_ _9273_/Q _4938_/A2 _7228_/A _9209_/Q VGND VGND VPWR VPWR _4835_/X sky130_fd_sc_hd__a22o_1
X_7554_ _7517_/X hold889/X hold99/A VGND VGND VPWR VPWR _7555_/A sky130_fd_sc_hd__mux2_1
X_4766_ _9282_/Q _7391_/A _5795_/A _8980_/Q VGND VGND VPWR VPWR _4766_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6505_ _6524_/B _6524_/C VGND VGND VPWR VPWR _6508_/B sky130_fd_sc_hd__or2_1
XFILLER_147_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7485_ _7485_/A VGND VGND VPWR VPWR _9321_/D sky130_fd_sc_hd__clkbuf_1
X_4697_ _9235_/Q _7284_/A _5750_/A _8961_/Q _4696_/X VGND VGND VPWR VPWR _4702_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_107_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9224_ _9272_/CLK _9224_/D fanout419/X VGND VGND VPWR VPWR _9224_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_162_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6436_ _6482_/A _6815_/B VGND VGND VPWR VPWR _6436_/Y sky130_fd_sc_hd__nand2_1
XFILLER_146_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9155_ _9462_/CLK _9155_/D fanout408/X VGND VGND VPWR VPWR _9155_/Q sky130_fd_sc_hd__dfrtp_1
X_6367_ _6495_/B VGND VGND VPWR VPWR _6895_/B sky130_fd_sc_hd__buf_4
X_5318_ _5330_/A _5334_/B VGND VGND VPWR VPWR _5319_/A sky130_fd_sc_hd__and2_1
X_8106_ _9188_/Q _8010_/B _8104_/X _8105_/X VGND VGND VPWR VPWR _8106_/X sky130_fd_sc_hd__o211a_1
X_6298_ _6739_/A _6558_/C _6788_/A VGND VGND VPWR VPWR _6376_/A sky130_fd_sc_hd__nor3b_1
X_9086_ _9088_/CLK _9086_/D fanout455/X VGND VGND VPWR VPWR _9086_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold13 hold13/A VGND VGND VPWR VPWR hold13/X sky130_fd_sc_hd__dlygate4sd3_1
X_8037_ _8037_/A _8037_/B _8037_/C _8037_/D VGND VGND VPWR VPWR _8037_/X sky130_fd_sc_hd__or4_2
X_5249_ _9291_/Q VGND VGND VPWR VPWR _5249_/Y sky130_fd_sc_hd__inv_2
Xhold24 hold24/A VGND VGND VPWR VPWR hold24/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold35 hold85/X VGND VGND VPWR VPWR hold35/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold46 hold46/A VGND VGND VPWR VPWR hold46/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold57 hold57/A VGND VGND VPWR VPWR hold57/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold68 hold68/A VGND VGND VPWR VPWR hold68/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A VGND VGND VPWR VPWR hold79/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8939_ _9161_/CLK _8939_/D fanout445/X VGND VGND VPWR VPWR _8939_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_71_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4620_ _9468_/Q _7798_/A _4502_/Y _4620_/B2 _4619_/X VGND VGND VPWR VPWR _4633_/A
+ sky130_fd_sc_hd__a221o_1
X_4551_ _4550_/X hold963/X _4964_/B VGND VGND VPWR VPWR _4551_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold505 hold505/A VGND VGND VPWR VPWR hold505/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7270_ _7270_/A VGND VGND VPWR VPWR _9225_/D sky130_fd_sc_hd__clkbuf_1
X_4482_ _7158_/A _4861_/A VGND VGND VPWR VPWR _7764_/A sky130_fd_sc_hd__nor2_8
Xhold516 hold516/A VGND VGND VPWR VPWR hold516/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold527 _9247_/Q VGND VGND VPWR VPWR hold527/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 _8945_/Q VGND VGND VPWR VPWR hold538/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6221_ _6562_/A _6558_/B VGND VGND VPWR VPWR _6222_/A sky130_fd_sc_hd__or2_1
Xhold549 _7062_/X VGND VGND VPWR VPWR _7063_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6152_ _6192_/A _6504_/A VGND VGND VPWR VPWR _6152_/X sky130_fd_sc_hd__or2_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _9275_/Q VGND VGND VPWR VPWR _5103_/Y sky130_fd_sc_hd__inv_2
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _6181_/A _6181_/B VGND VGND VPWR VPWR _6084_/A sky130_fd_sc_hd__and2_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1205 _9396_/Q VGND VGND VPWR VPWR hold366/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 _8894_/Q VGND VGND VPWR VPWR hold522/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _8807_/Q VGND VGND VPWR VPWR _5035_/B sky130_fd_sc_hd__inv_2
Xhold1227 _9226_/Q VGND VGND VPWR VPWR hold764/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1238 _9306_/Q VGND VGND VPWR VPWR hold706/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 _7054_/X VGND VGND VPWR VPWR hold758/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6985_ _6524_/C _6772_/B _6983_/Y _6984_/X VGND VGND VPWR VPWR _6985_/X sky130_fd_sc_hd__o211a_1
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8724_ _8724_/A VGND VGND VPWR VPWR _9540_/D sky130_fd_sc_hd__clkbuf_1
X_5936_ _5936_/A VGND VGND VPWR VPWR _9042_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8655_ _8901_/Q _8312_/X _8376_/X _8951_/Q VGND VGND VPWR VPWR _8655_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5867_ hold469/X hold5/X _5867_/S VGND VGND VPWR VPWR _5867_/X sky130_fd_sc_hd__mux2_1
X_7606_ hold54/X VGND VGND VPWR VPWR _7621_/S sky130_fd_sc_hd__buf_6
X_4818_ _9112_/Q _4817_/X _4886_/S VGND VGND VPWR VPWR _4818_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8586_ _8883_/Q _8314_/X _8331_/X _8978_/Q VGND VGND VPWR VPWR _8586_/X sky130_fd_sc_hd__a22o_1
X_5798_ _5633_/X hold454/X _5804_/S VGND VGND VPWR VPWR _5799_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7537_ _7517_/X hold929/X _7551_/S VGND VGND VPWR VPWR _7538_/A sky130_fd_sc_hd__mux2_1
X_4749_ _9475_/Q _7815_/A _7077_/A _9144_/Q VGND VGND VPWR VPWR _4749_/X sky130_fd_sc_hd__a22o_2
XFILLER_147_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7468_ _7468_/A VGND VGND VPWR VPWR _9313_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9207_ _9437_/CLK _9207_/D fanout419/X VGND VGND VPWR VPWR _9207_/Q sky130_fd_sc_hd__dfrtp_1
X_6419_ _6419_/A _6503_/A VGND VGND VPWR VPWR _6900_/A sky130_fd_sc_hd__nand2_4
XFILLER_134_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7399_ _7399_/A VGND VGND VPWR VPWR _9283_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9138_ _9480_/CLK _9138_/D fanout412/X VGND VGND VPWR VPWR _9138_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_1_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput103 sram_ro_data[19] VGND VGND VPWR VPWR _4704_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_163_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput114 sram_ro_data[29] VGND VGND VPWR VPWR _4575_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9069_ _9069_/CLK _9069_/D fanout434/X VGND VGND VPWR VPWR _9069_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput125 trap VGND VGND VPWR VPWR _5228_/A1 sky130_fd_sc_hd__buf_4
Xinput136 wb_adr_i[14] VGND VGND VPWR VPWR _6079_/D sky130_fd_sc_hd__clkbuf_1
Xinput147 wb_adr_i[24] VGND VGND VPWR VPWR _5118_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_56_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput158 wb_adr_i[5] VGND VGND VPWR VPWR _6181_/B sky130_fd_sc_hd__buf_2
XFILLER_48_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput169 wb_dat_i[14] VGND VGND VPWR VPWR _8759_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_2_csclk _9359_/CLK VGND VGND VPWR VPWR _9463_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6770_ _6838_/A _6770_/B _6770_/C _7006_/B VGND VGND VPWR VPWR _6784_/A sky130_fd_sc_hd__or4b_1
XFILLER_22_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5721_ _5721_/A VGND VGND VPWR VPWR _8945_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8440_ _9458_/Q _8348_/X _8411_/X _9338_/Q _8439_/X VGND VGND VPWR VPWR _8450_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_175_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5652_ _5652_/A VGND VGND VPWR VPWR _8916_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4603_ _4758_/A _4891_/B VGND VGND VPWR VPWR _5506_/A sky130_fd_sc_hd__nor2_4
XFILLER_129_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8371_ _8398_/A _8392_/C _8389_/C VGND VGND VPWR VPWR _8372_/A sky130_fd_sc_hd__and3_4
X_5583_ _5583_/A VGND VGND VPWR VPWR _8887_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7322_ _7322_/A VGND VGND VPWR VPWR _7337_/S sky130_fd_sc_hd__buf_8
X_4534_ _9294_/Q _7408_/A _7176_/A _9190_/Q _4533_/X VGND VGND VPWR VPWR _4534_/X
+ sky130_fd_sc_hd__a221o_1
Xhold302 _7492_/X VGND VGND VPWR VPWR _7493_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold313 _5411_/X VGND VGND VPWR VPWR _5412_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold324 _9462_/Q VGND VGND VPWR VPWR hold324/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 hold335/A VGND VGND VPWR VPWR hold335/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 _7822_/X VGND VGND VPWR VPWR _7823_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4465_ _4465_/A _4465_/B VGND VGND VPWR VPWR _7158_/B sky130_fd_sc_hd__nand2_8
X_7253_ _7253_/A VGND VGND VPWR VPWR _9217_/D sky130_fd_sc_hd__clkbuf_1
Xhold357 _5958_/X VGND VGND VPWR VPWR _5959_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold368 _5482_/X VGND VGND VPWR VPWR _5483_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6204_ _6297_/A _6297_/B _6156_/B VGND VGND VPWR VPWR _6232_/B sky130_fd_sc_hd__or3b_2
Xhold379 _9446_/Q VGND VGND VPWR VPWR hold379/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7184_ _9187_/Q hold46/X _7192_/S VGND VGND VPWR VPWR _7184_/X sky130_fd_sc_hd__mux2_1
X_4396_ _4396_/A _4465_/A VGND VGND VPWR VPWR _4748_/B sky130_fd_sc_hd__nand2_8
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6135_ _6167_/C _6167_/B VGND VGND VPWR VPWR _6420_/B sky130_fd_sc_hd__nand2b_4
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1002 _9521_/Q VGND VGND VPWR VPWR _8427_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1013 _9498_/Q VGND VGND VPWR VPWR _7893_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1024 _8793_/Q VGND VGND VPWR VPWR _5029_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6066_ _6066_/A _7132_/B VGND VGND VPWR VPWR _6075_/S sky130_fd_sc_hd__and2_2
XFILLER_100_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1035 _9549_/Q VGND VGND VPWR VPWR _5413_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1046 _9425_/Q VGND VGND VPWR VPWR _7715_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1057 _9545_/Q VGND VGND VPWR VPWR _8749_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5017_ hold994/X _8797_/Q _5017_/S VGND VGND VPWR VPWR _5018_/A sky130_fd_sc_hd__mux2_1
Xhold1068 _5881_/X VGND VGND VPWR VPWR _9010_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 _5834_/X VGND VGND VPWR VPWR _5835_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_54_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_208 _8402_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_219 _8400_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6968_ _6744_/A _6728_/B _6790_/B _6736_/A _6241_/B VGND VGND VPWR VPWR _6968_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_41_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8707_ _8706_/A _8705_/B _9031_/D VGND VGND VPWR VPWR _8707_/X sky130_fd_sc_hd__o21a_1
X_5919_ _5629_/X hold890/X _5927_/S VGND VGND VPWR VPWR _5920_/A sky130_fd_sc_hd__mux2_1
X_6899_ _6830_/Y _6812_/Y _6898_/Y _6636_/Y VGND VGND VPWR VPWR _6915_/B sky130_fd_sc_hd__a211o_1
XFILLER_139_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8638_ _8930_/Q _8301_/A _8356_/C _8895_/Q VGND VGND VPWR VPWR _8638_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8569_ _9391_/Q _8292_/X _8294_/X _9295_/Q VGND VGND VPWR VPWR _8569_/X sky130_fd_sc_hd__a22o_1
XFILLER_154_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold880 _8968_/Q VGND VGND VPWR VPWR hold880/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 hold891/A VGND VGND VPWR VPWR hold891/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7940_ _7940_/A VGND VGND VPWR VPWR _7940_/X sky130_fd_sc_hd__buf_8
XFILLER_103_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7871_ _7871_/A VGND VGND VPWR VPWR _9492_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6822_ _6822_/A _6822_/B VGND VGND VPWR VPWR _6822_/X sky130_fd_sc_hd__or2_1
XFILLER_168_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9541_ _9541_/CLK _9541_/D VGND VGND VPWR VPWR _9541_/Q sky130_fd_sc_hd__dfxtp_1
X_6753_ _6865_/B _6753_/B VGND VGND VPWR VPWR _6753_/Y sky130_fd_sc_hd__nor2_1
XFILLER_148_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5704_ _5704_/A _5715_/B VGND VGND VPWR VPWR _5713_/S sky130_fd_sc_hd__and2_2
XFILLER_148_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9472_ _9476_/CLK _9472_/D fanout414/X VGND VGND VPWR VPWR _9472_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_148_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6684_ _6340_/Y _6673_/B _6897_/B _6518_/Y VGND VGND VPWR VPWR _6759_/C sky130_fd_sc_hd__a22o_1
X_8423_ _8423_/A _8423_/B _8423_/C _8423_/D VGND VGND VPWR VPWR _8424_/C sky130_fd_sc_hd__or4_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5635_ _5635_/A VGND VGND VPWR VPWR _8909_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8354_ _8354_/A _8354_/B _8354_/C _8391_/A VGND VGND VPWR VPWR _8361_/A sky130_fd_sc_hd__or4_1
X_5566_ _5566_/A VGND VGND VPWR VPWR _8879_/D sky130_fd_sc_hd__clkbuf_1
Xhold110 _8836_/Q VGND VGND VPWR VPWR hold110/X sky130_fd_sc_hd__dlygate4sd3_1
X_7305_ _7302_/X hold920/X _7319_/S VGND VGND VPWR VPWR _7306_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold121 _8927_/Q VGND VGND VPWR VPWR hold121/X sky130_fd_sc_hd__dlygate4sd3_1
X_4517_ _9446_/Q _7746_/A _7729_/A _9438_/Q VGND VGND VPWR VPWR _4517_/X sky130_fd_sc_hd__a22o_1
Xhold132 _5316_/X VGND VGND VPWR VPWR _5317_/A sky130_fd_sc_hd__dlygate4sd3_1
X_5497_ _5497_/A VGND VGND VPWR VPWR _8849_/D sky130_fd_sc_hd__clkbuf_1
X_8285_ _9519_/Q _8017_/X _8284_/X VGND VGND VPWR VPWR _8285_/X sky130_fd_sc_hd__o21a_1
Xhold143 _9281_/Q VGND VGND VPWR VPWR hold143/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 _5911_/X VGND VGND VPWR VPWR _9021_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 _9220_/Q VGND VGND VPWR VPWR hold165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 _9461_/Q VGND VGND VPWR VPWR hold176/X sky130_fd_sc_hd__dlygate4sd3_1
X_7236_ _7648_/A VGND VGND VPWR VPWR _7236_/X sky130_fd_sc_hd__clkbuf_4
X_4448_ hold60/X _4858_/B VGND VGND VPWR VPWR _7374_/A sky130_fd_sc_hd__nor2_8
Xhold187 _5527_/X VGND VGND VPWR VPWR _5528_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold198 _5309_/X VGND VGND VPWR VPWR hold45/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4379_ hold51/X hold82/X VGND VGND VPWR VPWR _4432_/B sky130_fd_sc_hd__or2b_1
XFILLER_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7167_ _7167_/A VGND VGND VPWR VPWR _9179_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6118_ _6118_/A VGND VGND VPWR VPWR _6748_/B sky130_fd_sc_hd__clkbuf_4
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7098_ _6015_/X _9150_/Q _7106_/S VGND VGND VPWR VPWR _7098_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6049_ hold753/X _6048_/X _6053_/S VGND VGND VPWR VPWR _6050_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_82_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _9477_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_139_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_csclk _9210_/CLK VGND VGND VPWR VPWR _9436_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_76_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_35_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _9005_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5420_ _8817_/Q _5387_/X _5435_/S VGND VGND VPWR VPWR _5420_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5351_ _5353_/A _5356_/B VGND VGND VPWR VPWR _5352_/A sky130_fd_sc_hd__and2_1
Xoutput204 _9156_/Q VGND VGND VPWR VPWR irq[0] sky130_fd_sc_hd__buf_12
XFILLER_154_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput215 _5253_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[17] sky130_fd_sc_hd__buf_12
Xoutput226 _5262_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[27] sky130_fd_sc_hd__buf_12
Xoutput237 _5192_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[37] sky130_fd_sc_hd__buf_12
XFILLER_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput248 _5189_/X VGND VGND VPWR VPWR mgmt_gpio_out[36] sky130_fd_sc_hd__buf_12
XFILLER_5_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput259 _5176_/A VGND VGND VPWR VPWR pad_flash_io1_oeb sky130_fd_sc_hd__buf_12
X_5282_ _5282_/A VGND VGND VPWR VPWR _5282_/X sky130_fd_sc_hd__clkbuf_1
X_8070_ _9379_/Q _7947_/X _7990_/A _9275_/Q VGND VGND VPWR VPWR _8070_/X sky130_fd_sc_hd__a22o_1
XFILLER_4_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7021_ _7025_/A _7025_/B VGND VGND VPWR VPWR _7022_/A sky130_fd_sc_hd__and2_1
XFILLER_99_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8972_ _9427_/CLK _8972_/D fanout478/X VGND VGND VPWR VPWR _8972_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_55_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7923_ _7923_/A VGND VGND VPWR VPWR _7923_/X sky130_fd_sc_hd__buf_8
XFILLER_70_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7854_ _9488_/Q _7863_/D VGND VGND VPWR VPWR _7855_/C sky130_fd_sc_hd__or2_1
XFILLER_23_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6805_ _6870_/A _6959_/D _6805_/C VGND VGND VPWR VPWR _6806_/D sky130_fd_sc_hd__or3_1
XFILLER_169_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7785_ _7785_/A VGND VGND VPWR VPWR _9457_/D sky130_fd_sc_hd__clkbuf_1
X_4997_ _5040_/B _4997_/B VGND VGND VPWR VPWR _4997_/Y sky130_fd_sc_hd__nor2_1
X_9524_ _9529_/CLK _9524_/D fanout451/X VGND VGND VPWR VPWR _9524_/Q sky130_fd_sc_hd__dfrtp_1
X_6736_ _6736_/A _6736_/B VGND VGND VPWR VPWR _6860_/B sky130_fd_sc_hd__nand2_1
XFILLER_176_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9455_ _9471_/CLK _9455_/D fanout421/X VGND VGND VPWR VPWR _9455_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6667_ _6667_/A _6692_/B VGND VGND VPWR VPWR _6695_/A sky130_fd_sc_hd__or2_1
X_8406_ _9329_/Q _8298_/X _8370_/X _9249_/Q VGND VGND VPWR VPWR _8406_/X sky130_fd_sc_hd__a22o_1
X_5618_ _5618_/A _5715_/B VGND VGND VPWR VPWR _5627_/S sky130_fd_sc_hd__and2_2
X_9386_ _9467_/CLK _9386_/D fanout476/X VGND VGND VPWR VPWR _9386_/Q sky130_fd_sc_hd__dfrtp_4
X_6598_ _6852_/A _6597_/Y _6272_/D VGND VGND VPWR VPWR _6853_/C sky130_fd_sc_hd__o21ai_1
XFILLER_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8337_ _8337_/A VGND VGND VPWR VPWR _8337_/X sky130_fd_sc_hd__buf_8
XFILLER_145_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5549_ _5315_/X hold141/X _5549_/S VGND VGND VPWR VPWR _5549_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8268_ _9093_/Q _7958_/X _8001_/X _8867_/Q VGND VGND VPWR VPWR _8268_/X sky130_fd_sc_hd__a22o_1
XFILLER_155_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7219_ _7219_/A VGND VGND VPWR VPWR _9203_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout420 fanout424/X VGND VGND VPWR VPWR fanout420/X sky130_fd_sc_hd__clkbuf_4
Xfanout431 fanout432/X VGND VGND VPWR VPWR fanout431/X sky130_fd_sc_hd__clkbuf_2
X_8199_ _8924_/Q _7933_/X _8020_/X _8944_/Q _8198_/X VGND VGND VPWR VPWR _8216_/A
+ sky130_fd_sc_hd__a221o_1
Xfanout442 fanout449/X VGND VGND VPWR VPWR fanout442/X sky130_fd_sc_hd__clkbuf_2
Xfanout453 fanout456/X VGND VGND VPWR VPWR fanout453/X sky130_fd_sc_hd__clkbuf_4
Xfanout464 fanout498/X VGND VGND VPWR VPWR fanout464/X sky130_fd_sc_hd__clkbuf_4
XFILLER_59_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout475 fanout483/X VGND VGND VPWR VPWR fanout475/X sky130_fd_sc_hd__clkbuf_4
Xfanout486 fanout488/X VGND VGND VPWR VPWR fanout486/X sky130_fd_sc_hd__clkbuf_4
XFILLER_171_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout497 fanout498/X VGND VGND VPWR VPWR fanout497/X sky130_fd_sc_hd__clkbuf_4
XFILLER_100_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A VGND VGND VPWR VPWR _5226_/A1 sky130_fd_sc_hd__buf_12
XFILLER_69_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4920_ _9232_/Q _4428_/Y _5493_/A _8848_/Q _4919_/X VGND VGND VPWR VPWR _4921_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_33_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4851_ _8959_/Q _5750_/A _5642_/A _8914_/Q _4850_/X VGND VGND VPWR VPWR _4852_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_380 _4857_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_391 _7321_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7570_ _7570_/A VGND VGND VPWR VPWR _9359_/D sky130_fd_sc_hd__clkbuf_1
X_4782_ _4782_/A _4782_/B _4782_/C VGND VGND VPWR VPWR _4817_/A sky130_fd_sc_hd__or3_1
X_6521_ _6609_/A _6521_/B VGND VGND VPWR VPWR _6528_/B sky130_fd_sc_hd__nand2_1
XFILLER_158_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9240_ _9461_/CLK _9240_/D fanout420/X VGND VGND VPWR VPWR _9240_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_158_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6452_ _6967_/B _6453_/B VGND VGND VPWR VPWR _6657_/A sky130_fd_sc_hd__nor2_1
XFILLER_146_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5403_ _8813_/Q _5402_/X _5416_/S VGND VGND VPWR VPWR _5403_/X sky130_fd_sc_hd__mux2_1
X_9171_ _9173_/CLK _9171_/D fanout459/X VGND VGND VPWR VPWR _9171_/Q sky130_fd_sc_hd__dfrtp_1
X_6383_ _6891_/B _6828_/A VGND VGND VPWR VPWR _6673_/B sky130_fd_sc_hd__nor2_4
XFILLER_161_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8122_ _9261_/Q _7958_/X _7969_/X _9293_/Q _8121_/X VGND VGND VPWR VPWR _8127_/B
+ sky130_fd_sc_hd__a221o_1
X_5334_ _5353_/A _5334_/B VGND VGND VPWR VPWR _5335_/A sky130_fd_sc_hd__and2_1
XFILLER_0_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8053_ _9258_/Q _7958_/A _7971_/A _9418_/Q VGND VGND VPWR VPWR _8053_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5265_ _9427_/Q VGND VGND VPWR VPWR _5265_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7004_ _7004_/A _7004_/B _7004_/C VGND VGND VPWR VPWR _7009_/C sky130_fd_sc_hd__and3_1
X_5196_ _9467_/Q VGND VGND VPWR VPWR _5196_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8955_ _8955_/CLK _8955_/D fanout455/X VGND VGND VPWR VPWR _8955_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_55_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7906_ _9502_/Q _9501_/Q VGND VGND VPWR VPWR _8336_/A sky130_fd_sc_hd__and2b_1
XFILLER_70_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8886_ _9283_/CLK _8886_/D fanout484/X VGND VGND VPWR VPWR _8886_/Q sky130_fd_sc_hd__dfrtp_4
X_7837_ _5395_/X hold633/X _7847_/S VGND VGND VPWR VPWR _7837_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7768_ _7768_/A VGND VGND VPWR VPWR _9449_/D sky130_fd_sc_hd__clkbuf_1
X_9507_ _9531_/CLK _9507_/D fanout454/X VGND VGND VPWR VPWR _9507_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6719_ _6967_/A VGND VGND VPWR VPWR _6719_/Y sky130_fd_sc_hd__inv_2
XFILLER_177_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7699_ hold89/X VGND VGND VPWR VPWR _9417_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9438_ _9477_/CLK _9438_/D fanout409/X VGND VGND VPWR VPWR _9438_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9369_ _9475_/CLK _9369_/D fanout481/X VGND VGND VPWR VPWR _9369_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_117_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold709 _7050_/X VGND VGND VPWR VPWR _7051_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5050_ _5050_/A _5050_/B VGND VGND VPWR VPWR _5050_/X sky130_fd_sc_hd__and2_1
XFILLER_97_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8740_ _5271_/A _8740_/A2 _8740_/B1 _8727_/Y _8739_/X VGND VGND VPWR VPWR _8740_/X
+ sky130_fd_sc_hd__a221o_1
X_5952_ _5951_/X hold544/X _5958_/S VGND VGND VPWR VPWR _5952_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4903_ _8938_/Q _5704_/A _5296_/A _8772_/Q VGND VGND VPWR VPWR _4903_/X sky130_fd_sc_hd__a22o_1
X_8671_ _8941_/Q _7908_/X _8335_/X _8871_/Q VGND VGND VPWR VPWR _8671_/X sky130_fd_sc_hd__a22o_1
X_5883_ _9556_/A hold13/X _5898_/S VGND VGND VPWR VPWR _5883_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7622_ _7622_/A VGND VGND VPWR VPWR _9383_/D sky130_fd_sc_hd__clkbuf_1
X_4834_ _4834_/A1 _4444_/Y _4449_/Y _9241_/Q _4833_/X VGND VGND VPWR VPWR _4841_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_60_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7553_ _7553_/A _7695_/B VGND VGND VPWR VPWR hold99/A sky130_fd_sc_hd__nand2_8
X_4765_ input22/X _4460_/Y _7815_/A _9474_/Q _4764_/X VGND VGND VPWR VPWR _4772_/A
+ sky130_fd_sc_hd__a221o_4
XFILLER_193_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6504_ _6504_/A _6504_/B _6504_/C _6192_/A VGND VGND VPWR VPWR _6655_/C sky130_fd_sc_hd__or4b_4
XFILLER_146_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7484_ _7359_/X hold125/X _7497_/S VGND VGND VPWR VPWR _7484_/X sky130_fd_sc_hd__mux2_1
X_4696_ _9211_/Q _7228_/A _5948_/A _9051_/Q VGND VGND VPWR VPWR _4696_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9223_ _9485_/CLK _9223_/D fanout406/X VGND VGND VPWR VPWR _9223_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_107_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6435_ _6435_/A _6830_/A VGND VGND VPWR VPWR _6643_/A sky130_fd_sc_hd__nor2_1
XFILLER_162_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9154_ _9456_/CLK _9154_/D fanout406/X VGND VGND VPWR VPWR _9154_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_161_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6366_ _6440_/A _6420_/B VGND VGND VPWR VPWR _6495_/B sky130_fd_sc_hd__or2_2
XFILLER_161_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8105_ _8652_/S VGND VGND VPWR VPWR _8105_/X sky130_fd_sc_hd__buf_4
XFILLER_114_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5317_ _5317_/A VGND VGND VPWR VPWR _8776_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9085_ _9088_/CLK _9085_/D fanout455/X VGND VGND VPWR VPWR _9085_/Q sky130_fd_sc_hd__dfrtp_2
X_6297_ _6297_/A _6297_/B VGND VGND VPWR VPWR _6788_/A sky130_fd_sc_hd__or2_1
XFILLER_0_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8036_ _9233_/Q _8034_/X _7993_/X hold90/A _8035_/X VGND VGND VPWR VPWR _8037_/D
+ sky130_fd_sc_hd__a221o_1
Xhold14 hold14/A VGND VGND VPWR VPWR hold14/X sky130_fd_sc_hd__dlygate4sd3_1
X_5248_ _9283_/Q VGND VGND VPWR VPWR _5248_/Y sky130_fd_sc_hd__inv_2
Xhold25 hold25/A VGND VGND VPWR VPWR hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A VGND VGND VPWR VPWR hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A VGND VGND VPWR VPWR hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 hold58/A VGND VGND VPWR VPWR hold58/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold69 hold69/A VGND VGND VPWR VPWR hold69/X sky130_fd_sc_hd__dlygate4sd3_1
X_5179_ _8795_/Q _5179_/B VGND VGND VPWR VPWR _5180_/A sky130_fd_sc_hd__and2b_1
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8938_ _9089_/CLK _8938_/D fanout433/X VGND VGND VPWR VPWR _8938_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8869_ _9181_/CLK _8869_/D fanout486/X VGND VGND VPWR VPWR _8869_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4550_ _9116_/Q _4549_/X _4550_/S VGND VGND VPWR VPWR _4550_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold506 _8842_/Q VGND VGND VPWR VPWR hold506/X sky130_fd_sc_hd__dlygate4sd3_1
X_4481_ _9439_/Q _7729_/A _4477_/Y input33/X _4480_/X VGND VGND VPWR VPWR _4495_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold517 _9465_/Q VGND VGND VPWR VPWR hold517/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold528 _7319_/X VGND VGND VPWR VPWR _7320_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6220_ _6344_/A _6344_/B VGND VGND VPWR VPWR _6562_/A sky130_fd_sc_hd__nand2_4
Xhold539 _5720_/X VGND VGND VPWR VPWR _5721_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6151_ _6192_/A _6504_/A VGND VGND VPWR VPWR _6151_/Y sky130_fd_sc_hd__nand2_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _9283_/Q VGND VGND VPWR VPWR _5102_/Y sky130_fd_sc_hd__inv_2
X_6082_ _6169_/A VGND VGND VPWR VPWR _6437_/A sky130_fd_sc_hd__clkbuf_4
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1206 _8848_/Q VGND VGND VPWR VPWR hold940/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1217 _8963_/Q VGND VGND VPWR VPWR hold892/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5033_ _5067_/B _5068_/C _4550_/S _5032_/X VGND VGND VPWR VPWR _8792_/D sky130_fd_sc_hd__a31o_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1228 _8924_/Q VGND VGND VPWR VPWR hold444/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1239 _8889_/Q VGND VGND VPWR VPWR hold749/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6984_ _6764_/A _6781_/C _6779_/C _6453_/B _6967_/B VGND VGND VPWR VPWR _6984_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_25_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8723_ _9540_/Q _4549_/X _8725_/S VGND VGND VPWR VPWR _8724_/A sky130_fd_sc_hd__mux2_1
X_5935_ _9042_/Q _4817_/X _5945_/S VGND VGND VPWR VPWR _5936_/A sky130_fd_sc_hd__mux2_1
X_8654_ _8654_/A VGND VGND VPWR VPWR _9530_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5866_ _5866_/A VGND VGND VPWR VPWR _5866_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_178_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7605_ _7605_/A hold19/X VGND VGND VPWR VPWR hold54/A sky130_fd_sc_hd__and2_1
XFILLER_166_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4817_ _4817_/A _4817_/B _4817_/C _4817_/D VGND VGND VPWR VPWR _4817_/X sky130_fd_sc_hd__or4_4
X_8585_ _8918_/Q _8310_/X _8381_/X _8953_/Q _8584_/X VGND VGND VPWR VPWR _8588_/C
+ sky130_fd_sc_hd__a221o_1
X_5797_ _5797_/A VGND VGND VPWR VPWR _8978_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7536_ _7536_/A _7695_/B VGND VGND VPWR VPWR _7551_/S sky130_fd_sc_hd__nand2_8
X_4748_ _7158_/A _4748_/B VGND VGND VPWR VPWR _7077_/A sky130_fd_sc_hd__nor2_4
XFILLER_5_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7467_ hold109/X _5951_/A _7479_/S VGND VGND VPWR VPWR _7468_/A sky130_fd_sc_hd__mux2_1
X_4679_ _9292_/Q _7408_/A _6066_/A _9103_/Q VGND VGND VPWR VPWR _4679_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9206_ _9437_/CLK _9206_/D fanout409/X VGND VGND VPWR VPWR _9206_/Q sky130_fd_sc_hd__dfrtp_1
X_6418_ _6495_/B _6435_/A _6449_/B VGND VGND VPWR VPWR _6433_/B sky130_fd_sc_hd__a21oi_1
XFILLER_162_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7398_ _7236_/X _9283_/Q _7406_/S VGND VGND VPWR VPWR _7398_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9137_ _9480_/CLK _9137_/D fanout412/X VGND VGND VPWR VPWR _9137_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_1_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6349_ _6215_/A _6281_/A _6973_/B _6510_/A _6345_/A VGND VGND VPWR VPWR _6349_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_1_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput104 sram_ro_data[1] VGND VGND VPWR VPWR _4834_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9068_ _9110_/CLK _9068_/D VGND VGND VPWR VPWR _9068_/Q sky130_fd_sc_hd__dfxtp_1
Xinput115 sram_ro_data[2] VGND VGND VPWR VPWR _4793_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput126 uart_enabled VGND VGND VPWR VPWR _5277_/B sky130_fd_sc_hd__clkbuf_1
Xinput137 wb_adr_i[15] VGND VGND VPWR VPWR _6079_/C sky130_fd_sc_hd__clkbuf_1
Xinput148 wb_adr_i[25] VGND VGND VPWR VPWR input148/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8019_ _9329_/Q _7981_/X _7997_/X _9361_/Q _8018_/X VGND VGND VPWR VPWR _8027_/A
+ sky130_fd_sc_hd__a221o_1
Xinput159 wb_adr_i[6] VGND VGND VPWR VPWR _6169_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_56_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5720_ hold538/X _5683_/X _5724_/S VGND VGND VPWR VPWR _5720_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5651_ _5650_/X hold388/X _5654_/S VGND VGND VPWR VPWR _5652_/A sky130_fd_sc_hd__mux2_1
X_4602_ _9412_/Q _4438_/Y _5727_/A _8952_/Q _4601_/X VGND VGND VPWR VPWR _4690_/A
+ sky130_fd_sc_hd__a221o_1
X_8370_ _8370_/A VGND VGND VPWR VPWR _8370_/X sky130_fd_sc_hd__buf_6
XFILLER_175_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5582_ _5315_/X hold157/X _5582_/S VGND VGND VPWR VPWR _5582_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7321_ _7321_/A hold19/X VGND VGND VPWR VPWR _7322_/A sky130_fd_sc_hd__and2_1
X_4533_ _9302_/Q _4457_/Y _7284_/A _9238_/Q VGND VGND VPWR VPWR _4533_/X sky130_fd_sc_hd__a22o_1
Xhold303 _9324_/Q VGND VGND VPWR VPWR hold303/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold314 _9260_/Q VGND VGND VPWR VPWR hold314/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold325 _7794_/X VGND VGND VPWR VPWR _7795_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7252_ _7147_/X hold242/X _7264_/S VGND VGND VPWR VPWR _7252_/X sky130_fd_sc_hd__mux2_1
X_4464_ hold33/X _4878_/A VGND VGND VPWR VPWR _7832_/A sky130_fd_sc_hd__nor2_4
Xhold336 hold336/A VGND VGND VPWR VPWR hold336/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 _7488_/X VGND VGND VPWR VPWR _7489_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 _9254_/Q VGND VGND VPWR VPWR hold358/X sky130_fd_sc_hd__dlygate4sd3_1
X_6203_ _6716_/A _6344_/A VGND VGND VPWR VPWR _6262_/A sky130_fd_sc_hd__or2_2
Xhold369 _5430_/X VGND VGND VPWR VPWR _5431_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7183_ _7183_/A VGND VGND VPWR VPWR _9186_/D sky130_fd_sc_hd__clkbuf_1
X_4395_ hold64/X VGND VGND VPWR VPWR _4465_/A sky130_fd_sc_hd__inv_4
XFILLER_131_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6134_ _6479_/A _6764_/A VGND VGND VPWR VPWR _6778_/A sky130_fd_sc_hd__nor2_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1003 _8808_/Q VGND VGND VPWR VPWR _4969_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _6065_/A VGND VGND VPWR VPWR _9098_/D sky130_fd_sc_hd__clkbuf_1
Xhold1014 _9526_/Q VGND VGND VPWR VPWR _8553_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1025 _9489_/Q VGND VGND VPWR VPWR _7861_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1036 _5413_/X VGND VGND VPWR VPWR hold5/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 _9547_/Q VGND VGND VPWR VPWR _5405_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1058 _9547_/Q VGND VGND VPWR VPWR _8757_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5016_ _5068_/C _5016_/B VGND VGND VPWR VPWR _5017_/S sky130_fd_sc_hd__nand2_1
Xhold1069 _5862_/X VGND VGND VPWR VPWR _5863_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_209 _8333_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6967_ _6967_/A _6967_/B _6967_/C VGND VGND VPWR VPWR _6969_/B sky130_fd_sc_hd__nor3_1
XFILLER_41_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5918_ _5918_/A _7043_/B VGND VGND VPWR VPWR _5927_/S sky130_fd_sc_hd__nand2_4
X_8706_ _8706_/A _8706_/B VGND VGND VPWR VPWR _8706_/Y sky130_fd_sc_hd__nand2_1
X_6898_ _6898_/A _6900_/B VGND VGND VPWR VPWR _6898_/Y sky130_fd_sc_hd__nor2_1
X_8637_ _8970_/Q _8506_/B _8632_/X _8634_/X _8636_/X VGND VGND VPWR VPWR _8637_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_166_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5849_ _8841_/Q hold37/X _5867_/S VGND VGND VPWR VPWR hold38/A sky130_fd_sc_hd__mux2_1
XFILLER_22_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8568_ _9239_/Q _8322_/X _8333_/X _9271_/Q _8567_/X VGND VGND VPWR VPWR _8575_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7519_ _7519_/A _7695_/B VGND VGND VPWR VPWR _7534_/S sky130_fd_sc_hd__nand2_8
X_8499_ _8499_/A _8499_/B _8499_/C _8499_/D VGND VGND VPWR VPWR _8500_/C sky130_fd_sc_hd__or4_2
XFILLER_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold870 hold870/A VGND VGND VPWR VPWR hold870/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold881 hold881/A VGND VGND VPWR VPWR hold881/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold892 hold892/A VGND VGND VPWR VPWR hold892/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7870_ _7902_/B _7869_/Y _9492_/Q VGND VGND VPWR VPWR _7871_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6821_ _6462_/B _6812_/Y _6819_/Y _6820_/Y VGND VGND VPWR VPWR _6821_/X sky130_fd_sc_hd__a211o_1
XFILLER_35_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9540_ _9541_/CLK _9540_/D VGND VGND VPWR VPWR _9540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6752_ _6752_/A _6752_/B VGND VGND VPWR VPWR _6753_/B sky130_fd_sc_hd__nor2_1
XFILLER_50_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5703_ _5703_/A VGND VGND VPWR VPWR _8937_/D sky130_fd_sc_hd__clkbuf_1
X_9471_ _9471_/CLK _9471_/D fanout421/X VGND VGND VPWR VPWR _9471_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6683_ _6419_/A _6897_/B _6503_/A _6355_/C VGND VGND VPWR VPWR _6703_/B sky130_fd_sc_hd__a31o_1
XFILLER_176_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8422_ _9209_/Q _8289_/X _8341_/X _9305_/Q _8421_/X VGND VGND VPWR VPWR _8423_/D
+ sky130_fd_sc_hd__a221o_1
X_5634_ _5633_/X hold728/X _5640_/S VGND VGND VPWR VPWR _5635_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8353_ _8363_/A _8385_/B VGND VGND VPWR VPWR _8391_/A sky130_fd_sc_hd__nor2_4
X_5565_ hold459/X _5392_/X _5571_/S VGND VGND VPWR VPWR _5566_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold100 _7557_/X VGND VGND VPWR VPWR _7558_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7304_ _7304_/A _7499_/B VGND VGND VPWR VPWR _7319_/S sky130_fd_sc_hd__nand2_8
Xhold111 _5463_/X VGND VGND VPWR VPWR _5464_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4516_ _4516_/A1 _4483_/Y _7211_/A _9206_/Q _4515_/X VGND VGND VPWR VPWR _4521_/B
+ sky130_fd_sc_hd__a221o_1
X_8284_ _5130_/A _9518_/Q _8013_/A _8283_/X VGND VGND VPWR VPWR _8284_/X sky130_fd_sc_hd__a211o_1
Xhold122 _5676_/X VGND VGND VPWR VPWR _5677_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5496_ hold477/X _5392_/X _5502_/S VGND VGND VPWR VPWR _5496_/X sky130_fd_sc_hd__mux2_1
Xhold133 _9297_/Q VGND VGND VPWR VPWR hold133/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold144 _9265_/Q VGND VGND VPWR VPWR hold144/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold155 _9098_/Q VGND VGND VPWR VPWR hold155/X sky130_fd_sc_hd__dlygate4sd3_1
X_7235_ _7235_/A VGND VGND VPWR VPWR _9210_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4447_ hold33/X _4858_/B VGND VGND VPWR VPWR _4447_/Y sky130_fd_sc_hd__nor2_1
Xhold166 _7258_/X VGND VGND VPWR VPWR _7259_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 _7792_/X VGND VGND VPWR VPWR _7793_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 _9422_/Q VGND VGND VPWR VPWR hold188/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold199 _5885_/X VGND VGND VPWR VPWR hold199/X sky130_fd_sc_hd__dlygate4sd3_1
X_7166_ _6015_/X hold374/X _7174_/S VGND VGND VPWR VPWR _7166_/X sky130_fd_sc_hd__mux2_1
X_4378_ _4402_/B _4425_/B VGND VGND VPWR VPWR _4858_/B sky130_fd_sc_hd__nand2_8
Xclkbuf_leaf_1_csclk _9359_/CLK VGND VGND VPWR VPWR _9398_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6117_ _6628_/A _6589_/C _6628_/B VGND VGND VPWR VPWR _6118_/A sky130_fd_sc_hd__or3_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7097_ _7097_/A VGND VGND VPWR VPWR _9149_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6048_ _7645_/A VGND VGND VPWR VPWR _6048_/X sky130_fd_sc_hd__buf_8
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7999_ _8068_/B VGND VGND VPWR VPWR _7999_/X sky130_fd_sc_hd__buf_6
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_0_0_mgmt_gpio_in[4] clkbuf_2_1_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _8831_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_150_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5350_ _5350_/A VGND VGND VPWR VPWR _5350_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_173_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput205 _5284_/X VGND VGND VPWR VPWR irq[1] sky130_fd_sc_hd__buf_12
Xoutput216 _5254_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[18] sky130_fd_sc_hd__buf_12
Xoutput227 _5263_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[28] sky130_fd_sc_hd__buf_12
Xoutput238 _5238_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[3] sky130_fd_sc_hd__buf_12
Xoutput249 _5187_/X VGND VGND VPWR VPWR mgmt_gpio_out[37] sky130_fd_sc_hd__buf_12
X_5281_ _5281_/A input1/X VGND VGND VPWR VPWR _5282_/A sky130_fd_sc_hd__and2_1
X_7020_ _7020_/A VGND VGND VPWR VPWR _7020_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8971_ _9419_/CLK _8971_/D fanout491/X VGND VGND VPWR VPWR _8971_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_95_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7922_ _8181_/B _7989_/B _7984_/C VGND VGND VPWR VPWR _7923_/A sky130_fd_sc_hd__and3_2
XFILLER_48_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7853_ _9488_/Q _7863_/D VGND VGND VPWR VPWR _7855_/B sky130_fd_sc_hd__nand2_1
XFILLER_130_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6804_ _6957_/A _6872_/D _6803_/X VGND VGND VPWR VPWR _6805_/C sky130_fd_sc_hd__or3b_1
X_7784_ _5392_/X hold476/X _7796_/S VGND VGND VPWR VPWR _7785_/A sky130_fd_sc_hd__mux2_1
X_4996_ _4996_/A VGND VGND VPWR VPWR _8802_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9523_ _9529_/CLK _9523_/D fanout451/X VGND VGND VPWR VPWR _9523_/Q sky130_fd_sc_hd__dfrtp_1
X_6735_ _6863_/D _6966_/D _6851_/D _6735_/D VGND VGND VPWR VPWR _6751_/A sky130_fd_sc_hd__or4_1
XFILLER_149_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9454_ _9462_/CLK _9454_/D fanout408/X VGND VGND VPWR VPWR _9454_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6666_ _6973_/A _6666_/B VGND VGND VPWR VPWR _6692_/B sky130_fd_sc_hd__xnor2_1
XFILLER_164_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5617_ _5617_/A VGND VGND VPWR VPWR _8902_/D sky130_fd_sc_hd__clkbuf_1
X_8405_ _9369_/Q _8346_/X _8386_/X _9345_/Q VGND VGND VPWR VPWR _8405_/X sky130_fd_sc_hd__a22o_1
X_9385_ _9427_/CLK _9385_/D fanout479/X VGND VGND VPWR VPWR hold90/A sky130_fd_sc_hd__dfstp_2
XFILLER_191_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6597_ _6597_/A _6597_/B VGND VGND VPWR VPWR _6597_/Y sky130_fd_sc_hd__nand2_2
XFILLER_152_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8336_ _8336_/A _8357_/B _8389_/C VGND VGND VPWR VPWR _8337_/A sky130_fd_sc_hd__and3_2
X_5548_ _5548_/A VGND VGND VPWR VPWR _8871_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8267_ _8862_/Q _7927_/X _8023_/B _8892_/Q _8266_/X VGND VGND VPWR VPWR _8272_/B
+ sky130_fd_sc_hd__a221o_1
X_5479_ _5479_/A VGND VGND VPWR VPWR _8841_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7218_ _6015_/X _9203_/Q _7226_/S VGND VGND VPWR VPWR _7218_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout410 fanout457/X VGND VGND VPWR VPWR fanout410/X sky130_fd_sc_hd__buf_2
X_8198_ _8979_/Q _7931_/X _7990_/X _8869_/Q VGND VGND VPWR VPWR _8198_/X sky130_fd_sc_hd__a22o_1
Xfanout421 fanout424/X VGND VGND VPWR VPWR fanout421/X sky130_fd_sc_hd__clkbuf_4
XFILLER_132_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout432 fanout435/X VGND VGND VPWR VPWR fanout432/X sky130_fd_sc_hd__buf_4
Xfanout443 fanout449/X VGND VGND VPWR VPWR fanout443/X sky130_fd_sc_hd__clkbuf_4
Xfanout454 fanout455/X VGND VGND VPWR VPWR fanout454/X sky130_fd_sc_hd__clkbuf_4
X_7149_ _7149_/A VGND VGND VPWR VPWR _7149_/X sky130_fd_sc_hd__clkbuf_1
Xfanout465 fanout498/X VGND VGND VPWR VPWR fanout465/X sky130_fd_sc_hd__clkbuf_4
Xfanout476 fanout483/X VGND VGND VPWR VPWR fanout476/X sky130_fd_sc_hd__clkbuf_4
XFILLER_101_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout487 fanout488/X VGND VGND VPWR VPWR fanout487/X sky130_fd_sc_hd__clkbuf_2
Xfanout498 input75/X VGND VGND VPWR VPWR fanout498/X sky130_fd_sc_hd__buf_4
XFILLER_74_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4850_ _8818_/Q _5418_/A _6055_/A _9095_/Q VGND VGND VPWR VPWR _4850_/X sky130_fd_sc_hd__a22o_2
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_370 _8796_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_381 _4562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_392 _5468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4781_ _4781_/A _4781_/B _4781_/C _4781_/D VGND VGND VPWR VPWR _4782_/C sky130_fd_sc_hd__or4_1
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6520_ _6520_/A _6967_/C VGND VGND VPWR VPWR _6857_/C sky130_fd_sc_hd__nor2_1
XFILLER_118_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6451_ _6926_/B _6453_/B VGND VGND VPWR VPWR _6844_/A sky130_fd_sc_hd__nor2_1
X_5402_ _5690_/A VGND VGND VPWR VPWR _5402_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_146_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9170_ _9464_/CLK _9170_/D fanout420/X VGND VGND VPWR VPWR _9170_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6382_ _6393_/A _6668_/A _9033_/Q VGND VGND VPWR VPWR _6382_/X sky130_fd_sc_hd__o21a_1
XFILLER_133_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8121_ _9357_/Q _8020_/X _8008_/B _8120_/X VGND VGND VPWR VPWR _8121_/X sky130_fd_sc_hd__a22o_1
X_5333_ _7025_/A VGND VGND VPWR VPWR _5353_/A sky130_fd_sc_hd__buf_4
XFILLER_114_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8052_ _9242_/Q _7949_/A _7973_/A _9194_/Q VGND VGND VPWR VPWR _8052_/X sky130_fd_sc_hd__a22o_1
XFILLER_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5264_ _9419_/Q VGND VGND VPWR VPWR _5264_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7003_ _7003_/A _7003_/B _7003_/C _7003_/D VGND VGND VPWR VPWR _7004_/C sky130_fd_sc_hd__or4_1
XFILLER_87_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5195_ _5195_/A VGND VGND VPWR VPWR _5195_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_81_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _9486_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8954_ _8954_/CLK _8954_/D fanout469/X VGND VGND VPWR VPWR _8954_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_43_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7905_ _7898_/Y _7903_/Y _7909_/B VGND VGND VPWR VPWR _9501_/D sky130_fd_sc_hd__a21oi_1
X_8885_ _9283_/CLK _8885_/D fanout484/X VGND VGND VPWR VPWR _8885_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7836_ _7836_/A VGND VGND VPWR VPWR _9481_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4979_ _5021_/A _4979_/B VGND VGND VPWR VPWR _5014_/S sky130_fd_sc_hd__nand2_4
XFILLER_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7767_ _5392_/X hold499/X _7779_/S VGND VGND VPWR VPWR _7768_/A sky130_fd_sc_hd__mux2_1
X_9506_ _9529_/CLK _9506_/D fanout442/X VGND VGND VPWR VPWR _9506_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_7_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6718_ _6623_/Y _6717_/Y _6618_/B _7002_/A VGND VGND VPWR VPWR _6853_/D sky130_fd_sc_hd__a211o_1
XFILLER_137_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7698_ _7556_/X hold88/X _7710_/S VGND VGND VPWR VPWR hold89/A sky130_fd_sc_hd__mux2_1
XFILLER_192_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9437_ _9437_/CLK _9437_/D fanout410/X VGND VGND VPWR VPWR _9437_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6649_ _6811_/B _6811_/C VGND VGND VPWR VPWR _6658_/A sky130_fd_sc_hd__nand2_1
XFILLER_50_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9368_ _9416_/CLK _9368_/D fanout425/X VGND VGND VPWR VPWR _9368_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_152_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_34_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _9283_/CLK sky130_fd_sc_hd__clkbuf_16
X_8319_ _9501_/Q _9502_/Q VGND VGND VPWR VPWR _8320_/A sky130_fd_sc_hd__or2_1
XFILLER_105_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9299_ _9459_/CLK _9299_/D fanout479/X VGND VGND VPWR VPWR _9299_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_105_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_49_csclk _8954_/CLK VGND VGND VPWR VPWR _9241_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_115_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5951_ _5951_/A VGND VGND VPWR VPWR _5951_/X sky130_fd_sc_hd__buf_4
XFILLER_18_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4902_ _9248_/Q _7321_/A _5540_/A _8868_/Q _4901_/X VGND VGND VPWR VPWR _4909_/A
+ sky130_fd_sc_hd__a221o_1
X_8670_ _9072_/Q _8388_/X _8379_/X _9038_/Q _8669_/X VGND VGND VPWR VPWR _8675_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5882_ _9178_/Q hold12/X _5897_/S VGND VGND VPWR VPWR hold13/A sky130_fd_sc_hd__mux2_1
X_7621_ hold224/X _7514_/A _7621_/S VGND VGND VPWR VPWR _7622_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4833_ _8864_/Q _5529_/A _5773_/A _8969_/Q VGND VGND VPWR VPWR _4833_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7552_ _7552_/A VGND VGND VPWR VPWR _9351_/D sky130_fd_sc_hd__clkbuf_1
X_4764_ input5/X _4406_/Y _5678_/A _8930_/Q VGND VGND VPWR VPWR _4764_/X sky130_fd_sc_hd__a22o_1
X_6503_ _6503_/A VGND VGND VPWR VPWR _6521_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_147_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7483_ _7483_/A VGND VGND VPWR VPWR _9320_/D sky130_fd_sc_hd__clkbuf_1
X_4695_ _4695_/A1 _4483_/Y _7605_/A _9379_/Q _4694_/X VGND VGND VPWR VPWR _4702_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9222_ _9477_/CLK _9222_/D fanout409/X VGND VGND VPWR VPWR _9222_/Q sky130_fd_sc_hd__dfrtp_2
X_6434_ _6900_/A _6524_/C VGND VGND VPWR VPWR _6455_/A sky130_fd_sc_hd__nor2_1
XFILLER_161_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9153_ _9456_/CLK _9153_/D fanout407/X VGND VGND VPWR VPWR _9153_/Q sky130_fd_sc_hd__dfrtp_4
X_6365_ _6790_/B _6365_/B VGND VGND VPWR VPWR _6955_/A sky130_fd_sc_hd__nor2_1
XFILLER_115_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8104_ _8104_/A _8104_/B _8104_/C _8104_/D VGND VGND VPWR VPWR _8104_/X sky130_fd_sc_hd__or4_4
X_5316_ _5315_/X hold131/X _5316_/S VGND VGND VPWR VPWR _5316_/X sky130_fd_sc_hd__mux2_1
X_9084_ _9084_/CLK _9084_/D fanout447/X VGND VGND VPWR VPWR _9084_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_115_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6296_ _6479_/A _6790_/A VGND VGND VPWR VPWR _6585_/B sky130_fd_sc_hd__nor2_1
XFILLER_114_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8035_ _9225_/Q _7979_/X _8003_/X _9297_/Q VGND VGND VPWR VPWR _8035_/X sky130_fd_sc_hd__a22o_1
X_5247_ _9275_/Q VGND VGND VPWR VPWR _5247_/Y sky130_fd_sc_hd__inv_2
Xhold15 hold15/A VGND VGND VPWR VPWR hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 hold26/A VGND VGND VPWR VPWR hold26/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold37 hold69/X VGND VGND VPWR VPWR hold37/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold48 hold48/A VGND VGND VPWR VPWR hold48/X sky130_fd_sc_hd__dlygate4sd3_1
X_5178_ _5178_/A VGND VGND VPWR VPWR _5178_/X sky130_fd_sc_hd__clkbuf_1
Xhold59 hold59/A VGND VGND VPWR VPWR hold59/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8937_ _9465_/CLK _8937_/D fanout472/X VGND VGND VPWR VPWR _8937_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8868_ _9466_/CLK _8868_/D fanout471/X VGND VGND VPWR VPWR _8868_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7819_ _7819_/A VGND VGND VPWR VPWR _9473_/D sky130_fd_sc_hd__clkbuf_1
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8799_ _5168_/A1 _8799_/D _5366_/X VGND VGND VPWR VPWR hold8/A sky130_fd_sc_hd__dfrtp_2
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4480_ _9351_/Q _7536_/A _4811_/A _5283_/B VGND VGND VPWR VPWR _4480_/X sky130_fd_sc_hd__a22o_1
XFILLER_128_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold507 _5480_/X VGND VGND VPWR VPWR _5481_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 _8841_/Q VGND VGND VPWR VPWR hold518/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold529 hold529/A VGND VGND VPWR VPWR hold529/X sky130_fd_sc_hd__dlygate4sd3_1
X_6150_ _6150_/A VGND VGND VPWR VPWR _6895_/A sky130_fd_sc_hd__buf_4
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _9291_/Q VGND VGND VPWR VPWR _5101_/Y sky130_fd_sc_hd__inv_2
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6081_ _6170_/B _6170_/C _6170_/D VGND VGND VPWR VPWR _6088_/B sky130_fd_sc_hd__and3_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__1160_ _4690_/X VGND VGND VPWR VPWR clkbuf_0__1160_/X sky130_fd_sc_hd__clkbuf_16
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1207 _9090_/Q VGND VGND VPWR VPWR hold866/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5032_ _5021_/A _4964_/A _5032_/B1 VGND VGND VPWR VPWR _5032_/X sky130_fd_sc_hd__o21a_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1218 _8962_/Q VGND VGND VPWR VPWR hold642/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1229 _9382_/Q VGND VGND VPWR VPWR hold386/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_93_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6983_ _6983_/A VGND VGND VPWR VPWR _6983_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8722_ _8722_/A VGND VGND VPWR VPWR _9539_/D sky130_fd_sc_hd__clkbuf_1
X_5934_ _5934_/A VGND VGND VPWR VPWR _9041_/D sky130_fd_sc_hd__clkbuf_1
X_8653_ _8653_/A0 _8652_/X _8653_/S VGND VGND VPWR VPWR _8654_/A sky130_fd_sc_hd__mux2_1
X_5865_ _9006_/Q hold28/X _5868_/S VGND VGND VPWR VPWR _5865_/X sky130_fd_sc_hd__mux2_1
X_4816_ _4816_/A _4816_/B _4816_/C _4816_/D VGND VGND VPWR VPWR _4817_/D sky130_fd_sc_hd__or4_1
X_7604_ _7604_/A VGND VGND VPWR VPWR _9375_/D sky130_fd_sc_hd__clkbuf_1
X_8584_ _8913_/Q _8298_/X _8370_/X _9084_/Q VGND VGND VPWR VPWR _8584_/X sky130_fd_sc_hd__a22o_1
X_5796_ _5629_/X hold882/X _5804_/S VGND VGND VPWR VPWR _5797_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7535_ _7535_/A VGND VGND VPWR VPWR _9343_/D sky130_fd_sc_hd__clkbuf_1
X_4747_ _9267_/Q _4458_/Y _5618_/A _8906_/Q _4746_/X VGND VGND VPWR VPWR _4751_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_107_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7466_ _7466_/A VGND VGND VPWR VPWR _9312_/D sky130_fd_sc_hd__clkbuf_1
X_4678_ hold60/X _7158_/B VGND VGND VPWR VPWR _6066_/A sky130_fd_sc_hd__nor2_8
XFILLER_134_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9205_ _9461_/CLK _9205_/D fanout423/X VGND VGND VPWR VPWR _9205_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6417_ _6518_/A _6527_/A VGND VGND VPWR VPWR _6449_/B sky130_fd_sc_hd__or2_4
X_7397_ _7397_/A VGND VGND VPWR VPWR _9282_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9136_ _9476_/CLK _9136_/D fanout414/X VGND VGND VPWR VPWR _9136_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_162_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6348_ _6635_/A _6440_/A VGND VGND VPWR VPWR _6973_/B sky130_fd_sc_hd__nor2_8
XFILLER_49_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9067_ _9110_/CLK _9067_/D VGND VGND VPWR VPWR _9067_/Q sky130_fd_sc_hd__dfxtp_1
Xinput105 sram_ro_data[20] VGND VGND VPWR VPWR _4620_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_102_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6279_ _6279_/A VGND VGND VPWR VPWR _6281_/A sky130_fd_sc_hd__clkinv_2
Xinput116 sram_ro_data[30] VGND VGND VPWR VPWR _4516_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput127 usr1_vcc_pwrgood VGND VGND VPWR VPWR _4736_/B2 sky130_fd_sc_hd__clkbuf_2
Xinput138 wb_adr_i[16] VGND VGND VPWR VPWR _6078_/B sky130_fd_sc_hd__clkbuf_1
X_8018_ hold92/A _7931_/A _7999_/X _9425_/Q VGND VGND VPWR VPWR _8018_/X sky130_fd_sc_hd__a22o_1
Xinput149 wb_adr_i[26] VGND VGND VPWR VPWR _5124_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5650_ _7648_/A VGND VGND VPWR VPWR _5650_/X sky130_fd_sc_hd__buf_4
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4601_ _4601_/A1 _4444_/Y _4598_/X _4600_/X VGND VGND VPWR VPWR _4601_/X sky130_fd_sc_hd__a211o_1
X_5581_ _5581_/A VGND VGND VPWR VPWR _8886_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7320_ _7320_/A VGND VGND VPWR VPWR _9247_/D sky130_fd_sc_hd__clkbuf_1
X_4532_ _9486_/Q _7832_/A _4455_/Y _9326_/Q VGND VGND VPWR VPWR _4532_/X sky130_fd_sc_hd__a22o_1
XFILLER_184_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold304 _7490_/X VGND VGND VPWR VPWR _7491_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7251_ _7251_/A VGND VGND VPWR VPWR _9216_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold315 _7348_/X VGND VGND VPWR VPWR _7349_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4463_ _4463_/A _4463_/B _4463_/C _4463_/D VGND VGND VPWR VPWR _4506_/B sky130_fd_sc_hd__or4_1
XFILLER_144_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold326 hold326/A VGND VGND VPWR VPWR hold326/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 hold337/A VGND VGND VPWR VPWR hold337/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 _7453_/X VGND VGND VPWR VPWR _7454_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6202_ _6790_/B _6800_/A VGND VGND VPWR VPWR _6591_/A sky130_fd_sc_hd__or2_1
Xhold359 _7335_/X VGND VGND VPWR VPWR _7336_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7182_ hold743/X _6048_/X _7192_/S VGND VGND VPWR VPWR _7182_/X sky130_fd_sc_hd__mux2_1
X_4394_ hold63/X hold41/X VGND VGND VPWR VPWR hold64/A sky130_fd_sc_hd__nand2_1
XFILLER_98_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6133_ _6402_/A _6839_/A VGND VGND VPWR VPWR _6764_/A sky130_fd_sc_hd__nand2_4
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1004 _9504_/Q VGND VGND VPWR VPWR _7914_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_6064_ _6018_/X hold155/X _6064_/S VGND VGND VPWR VPWR _6064_/X sky130_fd_sc_hd__mux2_1
Xhold1015 _9033_/Q VGND VGND VPWR VPWR _5871_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1026 _9031_/Q VGND VGND VPWR VPWR _8706_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5015_ _5015_/A VGND VGND VPWR VPWR _8798_/D sky130_fd_sc_hd__clkbuf_1
Xhold1037 hold1199/X VGND VGND VPWR VPWR _5899_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1048 _5405_/X VGND VGND VPWR VPWR hold15/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 _5828_/X VGND VGND VPWR VPWR _5829_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6966_ _6966_/A _6966_/B _6966_/C _6966_/D VGND VGND VPWR VPWR _6994_/C sky130_fd_sc_hd__or4_1
X_8705_ _8705_/A _8705_/B VGND VGND VPWR VPWR _8705_/Y sky130_fd_sc_hd__nand2_1
X_5917_ _5917_/A VGND VGND VPWR VPWR _5917_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6897_ _6897_/A _6897_/B VGND VGND VPWR VPWR _6900_/B sky130_fd_sc_hd__nor2_1
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8636_ _9101_/Q _8372_/A _8369_/A _8905_/Q _8635_/X VGND VGND VPWR VPWR _8636_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5848_ _5848_/A VGND VGND VPWR VPWR _9000_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8567_ _9287_/Q _8316_/X _8327_/X _9263_/Q VGND VGND VPWR VPWR _8567_/X sky130_fd_sc_hd__a22o_2
XFILLER_166_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5779_ _5779_/A VGND VGND VPWR VPWR _8970_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7518_ hold20/A VGND VGND VPWR VPWR _7695_/B sky130_fd_sc_hd__buf_12
X_8498_ _9212_/Q _8289_/X _8341_/X _9308_/Q _8497_/X VGND VGND VPWR VPWR _8499_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7449_ _7359_/X hold394/X _7461_/S VGND VGND VPWR VPWR _7450_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold860 _5420_/X VGND VGND VPWR VPWR _5421_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 _9216_/Q VGND VGND VPWR VPWR hold871/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 hold882/A VGND VGND VPWR VPWR hold882/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold893 _9232_/Q VGND VGND VPWR VPWR hold893/X sky130_fd_sc_hd__dlygate4sd3_1
X_9119_ _9456_/CLK _9119_/D fanout404/X VGND VGND VPWR VPWR _9119_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6820_ _6894_/B _6895_/B VGND VGND VPWR VPWR _6820_/Y sky130_fd_sc_hd__nor2_1
X_6751_ _6751_/A _6751_/B _6946_/B _6751_/D VGND VGND VPWR VPWR _6752_/B sky130_fd_sc_hd__or4_1
XFILLER_50_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_1_0_wb_clk_i rebuffer3/X VGND VGND VPWR VPWR clkbuf_1_1_1_wb_clk_i/A sky130_fd_sc_hd__buf_8
X_5702_ _5653_/X hold171/X _5702_/S VGND VGND VPWR VPWR _5702_/X sky130_fd_sc_hd__mux2_1
X_9470_ _9471_/CLK _9470_/D fanout421/X VGND VGND VPWR VPWR _9470_/Q sky130_fd_sc_hd__dfrtp_2
X_6682_ _6897_/B _6503_/A _6429_/B _6758_/B VGND VGND VPWR VPWR _6703_/A sky130_fd_sc_hd__a31o_1
XFILLER_149_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8421_ _9393_/Q _8304_/A _8354_/C _9241_/Q VGND VGND VPWR VPWR _8421_/X sky130_fd_sc_hd__a22o_1
X_5633_ _5951_/A VGND VGND VPWR VPWR _5633_/X sky130_fd_sc_hd__buf_4
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5564_ _5564_/A VGND VGND VPWR VPWR _8878_/D sky130_fd_sc_hd__clkbuf_1
X_8352_ _8352_/A _8389_/C VGND VGND VPWR VPWR _8385_/B sky130_fd_sc_hd__nand2_2
XFILLER_176_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4515_ _9350_/Q _7536_/A _7091_/A _9153_/Q VGND VGND VPWR VPWR _4515_/X sky130_fd_sc_hd__a22o_1
Xhold101 _5895_/X VGND VGND VPWR VPWR _5896_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7303_ hold20/X VGND VGND VPWR VPWR _7499_/B sky130_fd_sc_hd__buf_12
XFILLER_117_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold112 _9546_/Q VGND VGND VPWR VPWR hold112/X sky130_fd_sc_hd__dlygate4sd3_1
X_8283_ _8852_/Q _8009_/A _8272_/X _8282_/X _8627_/S VGND VGND VPWR VPWR _8283_/X
+ sky130_fd_sc_hd__o221a_1
X_5495_ _5495_/A VGND VGND VPWR VPWR _8848_/D sky130_fd_sc_hd__clkbuf_1
Xhold123 _8952_/Q VGND VGND VPWR VPWR hold123/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold134 _9225_/Q VGND VGND VPWR VPWR hold134/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 _7360_/X VGND VGND VPWR VPWR _7361_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold156 _6064_/X VGND VGND VPWR VPWR _6065_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4446_ _4446_/A1 _4444_/Y _7623_/A _9391_/Q VGND VGND VPWR VPWR _4463_/A sky130_fd_sc_hd__a22o_1
X_7234_ _7233_/X hold865/X _7247_/S VGND VGND VPWR VPWR _7235_/A sky130_fd_sc_hd__mux2_1
Xhold167 _9228_/Q VGND VGND VPWR VPWR hold167/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 _9437_/Q VGND VGND VPWR VPWR hold178/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 _7708_/X VGND VGND VPWR VPWR _7709_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7165_ _7165_/A VGND VGND VPWR VPWR _9178_/D sky130_fd_sc_hd__clkbuf_1
X_4377_ hold10/X _4468_/B VGND VGND VPWR VPWR _4425_/B sky130_fd_sc_hd__nor2_8
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116_ _6248_/A _6794_/A VGND VGND VPWR VPWR _6628_/B sky130_fd_sc_hd__nand2_8
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7096_ _6012_/X _9149_/Q _7106_/S VGND VGND VPWR VPWR _7096_/X sky130_fd_sc_hd__mux2_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6047_ _6047_/A VGND VGND VPWR VPWR _9090_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7998_ _7998_/A _8002_/B _8002_/C VGND VGND VPWR VPWR _8068_/B sky130_fd_sc_hd__and3_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6949_ _6739_/Y _6721_/X _6732_/Y _6924_/C _6469_/B VGND VGND VPWR VPWR _6950_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_186_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8619_ _9070_/Q _8388_/A _8379_/A _9036_/Q _8618_/X VGND VGND VPWR VPWR _8624_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_10_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold690 _7127_/X VGND VGND VPWR VPWR _9163_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput206 _5286_/X VGND VGND VPWR VPWR irq[2] sky130_fd_sc_hd__buf_12
Xoutput217 _5255_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[19] sky130_fd_sc_hd__buf_12
XFILLER_126_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput228 _5264_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[29] sky130_fd_sc_hd__buf_12
XFILLER_154_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput239 _5240_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[4] sky130_fd_sc_hd__buf_12
X_5280_ _5280_/A VGND VGND VPWR VPWR _5280_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8970_ _9419_/CLK _8970_/D fanout492/X VGND VGND VPWR VPWR _8970_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7921_ _9495_/Q _9494_/Q VGND VGND VPWR VPWR _7984_/C sky130_fd_sc_hd__nor2_4
XFILLER_82_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7852_ _8997_/Q _8999_/Q _8998_/Q _7851_/Y VGND VGND VPWR VPWR _7863_/D sky130_fd_sc_hd__o31a_1
XFILLER_51_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6803_ _6603_/A _6881_/A _6871_/B _7001_/A _7001_/B VGND VGND VPWR VPWR _6803_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7783_ _7783_/A VGND VGND VPWR VPWR _9456_/D sky130_fd_sc_hd__clkbuf_1
X_4995_ _4994_/X hold80/A _5014_/S VGND VGND VPWR VPWR _4996_/A sky130_fd_sc_hd__mux2_1
X_9522_ _9529_/CLK _9522_/D fanout451/X VGND VGND VPWR VPWR _9522_/Q sky130_fd_sc_hd__dfrtp_1
X_6734_ _6715_/B _6673_/A _6195_/B _6597_/A _6733_/X VGND VGND VPWR VPWR _6735_/D
+ sky130_fd_sc_hd__a221o_1
X_9453_ _9453_/CLK _9453_/D fanout461/X VGND VGND VPWR VPWR _9453_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6665_ _6790_/C _6665_/B VGND VGND VPWR VPWR _6710_/C sky130_fd_sc_hd__nor2_1
XFILLER_177_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8404_ hold88/A _8402_/X _8378_/X _9353_/Q _8403_/X VGND VGND VPWR VPWR _8404_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_164_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5616_ _5315_/X hold169/X _5616_/S VGND VGND VPWR VPWR _5616_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9384_ _9471_/CLK _9384_/D _5070_/A VGND VGND VPWR VPWR _9384_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_176_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6596_ _6850_/B _6596_/B VGND VGND VPWR VPWR _6852_/A sky130_fd_sc_hd__or2_1
XFILLER_164_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8335_ _8358_/C VGND VGND VPWR VPWR _8335_/X sky130_fd_sc_hd__buf_8
X_5547_ _5311_/X hold387/X _5549_/S VGND VGND VPWR VPWR _5548_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8266_ _8927_/Q _7933_/A _7999_/X _8952_/Q VGND VGND VPWR VPWR _8266_/X sky130_fd_sc_hd__a22o_1
X_5478_ _5301_/X hold518/X _5490_/S VGND VGND VPWR VPWR _5478_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4429_ _9359_/Q _7553_/A _7284_/A _9239_/Q VGND VGND VPWR VPWR _4429_/X sky130_fd_sc_hd__a22o_1
X_7217_ _7217_/A VGND VGND VPWR VPWR _9202_/D sky130_fd_sc_hd__clkbuf_1
Xfanout411 fanout413/X VGND VGND VPWR VPWR fanout411/X sky130_fd_sc_hd__clkbuf_4
X_8197_ _8197_/A VGND VGND VPWR VPWR _9515_/D sky130_fd_sc_hd__clkbuf_1
Xfanout422 fanout424/X VGND VGND VPWR VPWR fanout422/X sky130_fd_sc_hd__clkbuf_4
Xfanout433 fanout434/X VGND VGND VPWR VPWR fanout433/X sky130_fd_sc_hd__clkbuf_4
XFILLER_132_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout444 fanout449/X VGND VGND VPWR VPWR fanout444/X sky130_fd_sc_hd__clkbuf_4
X_7148_ _7147_/X _9171_/Q _7156_/S VGND VGND VPWR VPWR _7148_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout455 fanout456/X VGND VGND VPWR VPWR fanout455/X sky130_fd_sc_hd__clkbuf_4
Xfanout466 fanout498/X VGND VGND VPWR VPWR fanout466/X sky130_fd_sc_hd__buf_2
XFILLER_48_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout477 fanout483/X VGND VGND VPWR VPWR fanout477/X sky130_fd_sc_hd__clkbuf_4
XFILLER_48_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7079_ _7079_/A VGND VGND VPWR VPWR _9141_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout488 fanout496/X VGND VGND VPWR VPWR fanout488/X sky130_fd_sc_hd__buf_2
Xfanout499 _8709_/B VGND VGND VPWR VPWR fanout499/X sky130_fd_sc_hd__clkbuf_4
XFILLER_74_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_360 _7969_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_371 _9168_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_382 _9147_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_393 _5471_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4780_ _9226_/Q _4454_/Y _4483_/Y _4780_/B2 _4779_/X VGND VGND VPWR VPWR _4781_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_0_csclk _9359_/CLK VGND VGND VPWR VPWR _9437_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6450_ _6973_/B _6597_/B VGND VGND VPWR VPWR _6453_/B sky130_fd_sc_hd__nand2_1
XFILLER_118_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5401_ hold24/X VGND VGND VPWR VPWR _5690_/A sky130_fd_sc_hd__buf_6
X_6381_ _6415_/B _6391_/B VGND VGND VPWR VPWR _6668_/A sky130_fd_sc_hd__nand2_1
XFILLER_161_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5332_ _5332_/A VGND VGND VPWR VPWR _7025_/A sky130_fd_sc_hd__clkbuf_2
X_8120_ _9317_/Q _8275_/B VGND VGND VPWR VPWR _8120_/X sky130_fd_sc_hd__or2_1
X_8051_ _9226_/Q _7979_/X _7993_/X _9386_/Q VGND VGND VPWR VPWR _8059_/A sky130_fd_sc_hd__a22o_1
X_5263_ _9411_/Q VGND VGND VPWR VPWR _5263_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7002_ _7002_/A _7002_/B _7002_/C _7002_/D VGND VGND VPWR VPWR _7003_/D sky130_fd_sc_hd__or4_1
X_5194_ _5193_/Y input90/X _5194_/S VGND VGND VPWR VPWR _5195_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8953_ _9241_/CLK _8953_/D fanout450/X VGND VGND VPWR VPWR _8953_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7904_ _9501_/Q _7904_/B _8389_/A VGND VGND VPWR VPWR _7909_/B sky130_fd_sc_hd__and3_1
XFILLER_71_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8884_ _9283_/CLK _8884_/D fanout484/X VGND VGND VPWR VPWR _8884_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_36_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7835_ _5392_/X hold537/X _7847_/S VGND VGND VPWR VPWR _7836_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7766_ _7766_/A VGND VGND VPWR VPWR _9448_/D sky130_fd_sc_hd__clkbuf_1
X_4978_ _8829_/Q _5016_/B _5127_/B _5040_/B VGND VGND VPWR VPWR _4979_/B sky130_fd_sc_hd__a31o_1
X_9505_ _9529_/CLK _9505_/D fanout442/X VGND VGND VPWR VPWR _9505_/Q sky130_fd_sc_hd__dfrtp_1
X_6717_ _6725_/B VGND VGND VPWR VPWR _6717_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7697_ _7697_/A VGND VGND VPWR VPWR _9416_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9436_ _9436_/CLK _9436_/D fanout462/X VGND VGND VPWR VPWR _9436_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6648_ _6648_/A _6729_/B VGND VGND VPWR VPWR _6661_/B sky130_fd_sc_hd__nand2_1
XFILLER_165_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9367_ _9367_/CLK _9367_/D fanout422/X VGND VGND VPWR VPWR _9367_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6579_ _6315_/Y _6551_/Y _6578_/X _6869_/A _6869_/D VGND VGND VPWR VPWR _6579_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_117_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8318_ _9448_/Q _8310_/X _8312_/X _9464_/Q _8317_/X VGND VGND VPWR VPWR _8351_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_164_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9298_ _9467_/CLK _9298_/D fanout475/X VGND VGND VPWR VPWR _9298_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8249_ _8891_/Q _8023_/B _8246_/X _8248_/X VGND VGND VPWR VPWR _8250_/C sky130_fd_sc_hd__a211o_1
XFILLER_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5950_ _5950_/A VGND VGND VPWR VPWR _9048_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4901_ _9328_/Q _4459_/Y _7228_/A _9208_/Q VGND VGND VPWR VPWR _4901_/X sky130_fd_sc_hd__a22o_1
XFILLER_45_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5881_ _5881_/A VGND VGND VPWR VPWR _5881_/X sky130_fd_sc_hd__clkbuf_1
X_7620_ _7620_/A VGND VGND VPWR VPWR _9382_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4832_ _9337_/Q _4414_/Y _5562_/A _8879_/Q _4831_/X VGND VGND VPWR VPWR _4853_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA_190 _7997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7551_ _7514_/X hold595/X _7551_/S VGND VGND VPWR VPWR _7551_/X sky130_fd_sc_hd__mux2_1
X_4763_ _4763_/A _4763_/B _4763_/C _4763_/D VGND VGND VPWR VPWR _4782_/A sky130_fd_sc_hd__or4_1
XFILLER_147_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6502_ _6966_/B _6502_/B _6726_/B _6501_/X VGND VGND VPWR VPWR _6517_/A sky130_fd_sc_hd__or4b_1
XFILLER_159_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4694_ _9243_/Q _4449_/Y _6066_/A hold71/A VGND VGND VPWR VPWR _4694_/X sky130_fd_sc_hd__a22o_1
X_7482_ _7302_/X hold927/X _7497_/S VGND VGND VPWR VPWR _7483_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9221_ _9477_/CLK _9221_/D fanout406/X VGND VGND VPWR VPWR _9221_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6433_ _6922_/A _6433_/B _6433_/C _6432_/X VGND VGND VPWR VPWR _6469_/C sky130_fd_sc_hd__or4b_1
XFILLER_20_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9152_ _9456_/CLK _9152_/D fanout404/X VGND VGND VPWR VPWR _9152_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_161_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6364_ _6364_/A _6948_/B _6364_/C _6363_/X VGND VGND VPWR VPWR _6364_/X sky130_fd_sc_hd__or4b_1
XFILLER_115_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8103_ _9204_/Q _7938_/X _8077_/X _9348_/Q _8102_/X VGND VGND VPWR VPWR _8104_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5315_ hold24/X VGND VGND VPWR VPWR _5315_/X sky130_fd_sc_hd__buf_6
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9083_ _9162_/CLK _9083_/D fanout441/X VGND VGND VPWR VPWR _9083_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_88_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6295_ _6479_/A _6873_/B VGND VGND VPWR VPWR _6867_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8034_ _8034_/A VGND VGND VPWR VPWR _8034_/X sky130_fd_sc_hd__buf_6
XFILLER_102_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5246_ _9267_/Q VGND VGND VPWR VPWR _5246_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold16 hold16/A VGND VGND VPWR VPWR hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A VGND VGND VPWR VPWR hold27/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold38 hold38/A VGND VGND VPWR VPWR hold38/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 hold49/A VGND VGND VPWR VPWR hold49/X sky130_fd_sc_hd__dlygate4sd3_1
X_5177_ input85/X _5067_/B _8795_/Q VGND VGND VPWR VPWR _5178_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8936_ _9005_/CLK _8936_/D fanout490/X VGND VGND VPWR VPWR _8936_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_37_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8867_ _9467_/CLK _8867_/D fanout471/X VGND VGND VPWR VPWR _8867_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7818_ _5392_/X hold475/X _7830_/S VGND VGND VPWR VPWR _7819_/A sky130_fd_sc_hd__mux2_1
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8798_ _8831_/CLK _8798_/D _5364_/X VGND VGND VPWR VPWR hold76/A sky130_fd_sc_hd__dfrtp_4
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7749_ _7749_/A VGND VGND VPWR VPWR _9440_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9419_ _9419_/CLK _9419_/D fanout491/X VGND VGND VPWR VPWR _9419_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_80_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _9487_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_190_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold508 _8860_/Q VGND VGND VPWR VPWR hold508/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold519 _5478_/X VGND VGND VPWR VPWR _5479_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_124_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5100_ _9299_/Q VGND VGND VPWR VPWR _5100_/Y sky130_fd_sc_hd__inv_2
X_6080_ _6080_/A _6080_/B _6080_/C _6080_/D VGND VGND VPWR VPWR _6170_/D sky130_fd_sc_hd__and4_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _5031_/A _5031_/B VGND VGND VPWR VPWR _8793_/D sky130_fd_sc_hd__nor2_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1208 _9373_/Q VGND VGND VPWR VPWR hold227/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1219 _7133_/X VGND VGND VPWR VPWR hold705/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6982_ _6761_/C _6982_/B _6982_/C _6982_/D VGND VGND VPWR VPWR _6982_/X sky130_fd_sc_hd__and4b_1
XFILLER_80_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8721_ _9539_/Q _4591_/X _8725_/S VGND VGND VPWR VPWR _8722_/A sky130_fd_sc_hd__mux2_1
X_5933_ _9041_/Q _4885_/X _5945_/S VGND VGND VPWR VPWR _5934_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_33_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _9449_/CLK sky130_fd_sc_hd__clkbuf_16
X_8652_ _9529_/Q _8651_/X _8652_/S VGND VGND VPWR VPWR _8652_/X sky130_fd_sc_hd__mux2_1
X_5864_ _8846_/Q hold27/X _5867_/S VGND VGND VPWR VPWR hold28/A sky130_fd_sc_hd__mux2_1
XFILLER_21_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7603_ _7514_/X hold584/X hold75/X VGND VGND VPWR VPWR _7603_/X sky130_fd_sc_hd__mux2_1
X_4815_ _9466_/Q _7798_/A _7553_/A _9354_/Q _4814_/X VGND VGND VPWR VPWR _4816_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_166_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8583_ _8963_/Q _8346_/X _8386_/X _8933_/Q _8582_/X VGND VGND VPWR VPWR _8588_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_193_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5795_ _5795_/A _7043_/B VGND VGND VPWR VPWR _5804_/S sky130_fd_sc_hd__nand2_4
X_7534_ _7514_/X hold598/X _7534_/S VGND VGND VPWR VPWR _7534_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_48_csclk _8954_/CLK VGND VGND VPWR VPWR _9227_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_119_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4746_ _9355_/Q _7553_/A _5667_/A _8926_/Q VGND VGND VPWR VPWR _4746_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7465_ hold852/X _7126_/C _7479_/S VGND VGND VPWR VPWR _7466_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4677_ _9284_/Q _7391_/A _7463_/A _9316_/Q _4676_/X VGND VGND VPWR VPWR _4688_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9204_ _9392_/CLK _9204_/D fanout425/X VGND VGND VPWR VPWR _9204_/Q sky130_fd_sc_hd__dfrtp_4
X_6416_ _6416_/A _6818_/A VGND VGND VPWR VPWR _6527_/A sky130_fd_sc_hd__or2_2
XFILLER_134_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7396_ _7233_/X hold771/X _7406_/S VGND VGND VPWR VPWR _7397_/A sky130_fd_sc_hd__mux2_1
X_9135_ _9473_/CLK _9135_/D fanout430/X VGND VGND VPWR VPWR _9135_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_150_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6347_ _6547_/A _6197_/B _6230_/C _6345_/A _6345_/C VGND VGND VPWR VPWR _6347_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9066_ _9110_/CLK _9066_/D VGND VGND VPWR VPWR _9066_/Q sky130_fd_sc_hd__dfxtp_1
X_6278_ _6311_/B _6799_/A _6209_/X _6275_/X _6277_/Y VGND VGND VPWR VPWR _6278_/X
+ sky130_fd_sc_hd__o2111a_1
Xinput106 sram_ro_data[21] VGND VGND VPWR VPWR _4579_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput117 sram_ro_data[31] VGND VGND VPWR VPWR _4487_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput128 usr1_vdd_pwrgood VGND VGND VPWR VPWR _4871_/B2 sky130_fd_sc_hd__clkbuf_2
X_8017_ _8196_/S VGND VGND VPWR VPWR _8017_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_48_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput139 wb_adr_i[17] VGND VGND VPWR VPWR _6078_/A sky130_fd_sc_hd__clkbuf_1
X_5229_ _5229_/A VGND VGND VPWR VPWR _9567_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_57_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8919_ _9051_/CLK _8919_/D fanout444/X VGND VGND VPWR VPWR _8919_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_90 _5468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__buf_8
XFILLER_67_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4600_ _5285_/B _4436_/A _4500_/Y input16/X _4599_/X VGND VGND VPWR VPWR _4600_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_175_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5580_ _5311_/X hold423/X _5582_/S VGND VGND VPWR VPWR _5581_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4531_ _4670_/B _7111_/B VGND VGND VPWR VPWR _4531_/Y sky130_fd_sc_hd__nor2_4
XFILLER_144_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold305 _9381_/Q VGND VGND VPWR VPWR hold305/X sky130_fd_sc_hd__dlygate4sd3_1
X_7250_ _7128_/X hold871/X _7264_/S VGND VGND VPWR VPWR _7251_/A sky130_fd_sc_hd__mux2_1
Xhold316 _9193_/Q VGND VGND VPWR VPWR hold316/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4462_ _9303_/Q _7425_/A _7356_/A _9271_/Q _4461_/X VGND VGND VPWR VPWR _4463_/D
+ sky130_fd_sc_hd__a221o_1
Xhold327 _7100_/X VGND VGND VPWR VPWR _7101_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 _5407_/X VGND VGND VPWR VPWR _5408_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold349 _7543_/X VGND VGND VPWR VPWR _7544_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6201_ _6266_/A VGND VGND VPWR VPWR _6790_/B sky130_fd_sc_hd__buf_4
XFILLER_144_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4393_ hold60/X VGND VGND VPWR VPWR _4656_/A sky130_fd_sc_hd__buf_12
X_7181_ _7181_/A VGND VGND VPWR VPWR _9185_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6132_ _6167_/B _6828_/A VGND VGND VPWR VPWR _6839_/A sky130_fd_sc_hd__nor2_8
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6063_ _6063_/A VGND VGND VPWR VPWR _9097_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1005 _9515_/Q VGND VGND VPWR VPWR _8196_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1016 _8763_/X VGND VGND VPWR VPWR _8764_/C1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1027 _9548_/Q VGND VGND VPWR VPWR _8761_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5014_ _5013_/X hold76/A _5014_/S VGND VGND VPWR VPWR _5015_/A sky130_fd_sc_hd__mux2_1
Xhold1038 hold1115/X VGND VGND VPWR VPWR _5860_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 _9030_/Q VGND VGND VPWR VPWR _5126_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6965_ _6965_/A _6965_/B _6965_/C VGND VGND VPWR VPWR _6965_/Y sky130_fd_sc_hd__nor3_1
XFILLER_41_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8704_ _9532_/Q _8196_/S _8702_/X _8703_/X VGND VGND VPWR VPWR _8704_/X sky130_fd_sc_hd__o22a_1
X_5916_ _5471_/X _9585_/A _5916_/S VGND VGND VPWR VPWR _5916_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6896_ _6514_/Y _6812_/Y _6973_/C _6462_/B _6644_/X VGND VGND VPWR VPWR _6972_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8635_ _8885_/Q _8354_/B _8331_/A _8980_/Q VGND VGND VPWR VPWR _8635_/X sky130_fd_sc_hd__a22o_1
X_5847_ _9000_/Q _5845_/X _5868_/S VGND VGND VPWR VPWR _5847_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8566_ _9463_/Q _8348_/X _8411_/X _9343_/Q _8565_/X VGND VGND VPWR VPWR _8576_/C
+ sky130_fd_sc_hd__a221o_1
X_5778_ _5647_/X hold615/X _5782_/S VGND VGND VPWR VPWR _5779_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7517_ _7517_/A VGND VGND VPWR VPWR _7517_/X sky130_fd_sc_hd__clkbuf_4
X_4729_ _9419_/Q _7695_/A _5493_/A _8851_/Q _4728_/X VGND VGND VPWR VPWR _4731_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_175_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8497_ _9396_/Q _8304_/X _8324_/X _9244_/Q VGND VGND VPWR VPWR _8497_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7448_ _7448_/A VGND VGND VPWR VPWR _9304_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold850 hold850/A VGND VGND VPWR VPWR hold850/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold861 _7058_/X VGND VGND VPWR VPWR _7059_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7379_ _7233_/X hold782/X _7389_/S VGND VGND VPWR VPWR _7380_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold872 hold872/A VGND VGND VPWR VPWR hold872/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 hold883/A VGND VGND VPWR VPWR hold883/X sky130_fd_sc_hd__dlygate4sd3_1
X_9118_ _5235__1/A _9118_/D _7026_/X VGND VGND VPWR VPWR _9118_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_107_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold894 hold894/A VGND VGND VPWR VPWR hold894/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9049_ _9184_/CLK _9049_/D fanout443/X VGND VGND VPWR VPWR _9049_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6750_ _6969_/A _6857_/D _6859_/C _6861_/A VGND VGND VPWR VPWR _6751_/D sky130_fd_sc_hd__or4_1
XFILLER_50_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5701_ _5701_/A VGND VGND VPWR VPWR _8936_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6681_ _6802_/A _6779_/A VGND VGND VPWR VPWR _6758_/B sky130_fd_sc_hd__nor2_1
XFILLER_188_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8420_ _9377_/Q _8337_/X _8384_/X _9193_/Q _8419_/X VGND VGND VPWR VPWR _8423_/C
+ sky130_fd_sc_hd__a221o_1
X_5632_ _5632_/A VGND VGND VPWR VPWR _8908_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8351_ _8351_/A _8351_/B _8351_/C _8351_/D VGND VGND VPWR VPWR _8397_/B sky130_fd_sc_hd__or4_1
X_5563_ hold932/X _5505_/X _5571_/S VGND VGND VPWR VPWR _5564_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7302_ _7517_/A VGND VGND VPWR VPWR _7302_/X sky130_fd_sc_hd__buf_4
X_4514_ _4514_/A1 _4444_/Y _7356_/A _9270_/Q _4513_/X VGND VGND VPWR VPWR _4521_/A
+ sky130_fd_sc_hd__a221o_1
X_8282_ _8282_/A _8282_/B _8282_/C _8282_/D VGND VGND VPWR VPWR _8282_/X sky130_fd_sc_hd__or4_1
Xhold102 _5896_/X VGND VGND VPWR VPWR _9015_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5494_ hold940/X _5387_/X _5502_/S VGND VGND VPWR VPWR _5495_/A sky130_fd_sc_hd__mux2_1
Xhold113 _5538_/X VGND VGND VPWR VPWR _5539_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 _5736_/X VGND VGND VPWR VPWR _5737_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold135 _9201_/Q VGND VGND VPWR VPWR hold135/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7233_ _7645_/A VGND VGND VPWR VPWR _7233_/X sky130_fd_sc_hd__buf_4
X_4445_ _4861_/A _4635_/A VGND VGND VPWR VPWR _4445_/Y sky130_fd_sc_hd__nor2_4
Xhold146 _7148_/X VGND VGND VPWR VPWR _7149_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 _8887_/Q VGND VGND VPWR VPWR hold157/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 _7275_/X VGND VGND VPWR VPWR _7276_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 _7740_/X VGND VGND VPWR VPWR _7741_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7164_ _6012_/X hold486/X _7174_/S VGND VGND VPWR VPWR _7164_/X sky130_fd_sc_hd__mux2_1
X_4376_ _4758_/A _4685_/B VGND VGND VPWR VPWR _7091_/A sky130_fd_sc_hd__nor2_8
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6115_ _6317_/A VGND VGND VPWR VPWR _6794_/A sky130_fd_sc_hd__buf_4
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7095_ _7095_/A VGND VGND VPWR VPWR _9148_/D sky130_fd_sc_hd__clkbuf_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ hold866/X _5809_/X _6053_/S VGND VGND VPWR VPWR _6047_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7997_ _7997_/A VGND VGND VPWR VPWR _7997_/X sky130_fd_sc_hd__buf_8
XFILLER_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6948_ _6948_/A _6948_/B _6947_/X VGND VGND VPWR VPWR _6964_/D sky130_fd_sc_hd__or3b_1
XFILLER_41_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6879_ _6227_/Y _6510_/Y _6508_/A _6610_/X _6232_/B VGND VGND VPWR VPWR _6879_/X
+ sky130_fd_sc_hd__a41o_1
X_8618_ _8984_/Q _8292_/A _8358_/A _8879_/Q VGND VGND VPWR VPWR _8618_/X sky130_fd_sc_hd__a22o_1
XFILLER_167_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8549_ _8549_/A _8549_/B _8549_/C _8549_/D VGND VGND VPWR VPWR _8550_/D sky130_fd_sc_hd__or4_1
XFILLER_108_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold680 _7222_/X VGND VGND VPWR VPWR _7223_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold691 _9263_/Q VGND VGND VPWR VPWR hold691/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput207 _5223_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[0] sky130_fd_sc_hd__buf_12
XFILLER_154_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput218 _5221_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[1] sky130_fd_sc_hd__buf_12
XFILLER_99_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput229 _5239_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[2] sky130_fd_sc_hd__buf_12
XFILLER_5_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7920_ _8997_/Q _7920_/B VGND VGND VPWR VPWR _7920_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7851_ _8997_/Q _7911_/B VGND VGND VPWR VPWR _7851_/Y sky130_fd_sc_hd__nand2_1
XFILLER_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6802_ _6802_/A _7001_/B VGND VGND VPWR VPWR _6872_/D sky130_fd_sc_hd__nor2_1
XFILLER_24_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7782_ _5387_/X hold936/X _7796_/S VGND VGND VPWR VPWR _7783_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4994_ hold50/A _4360_/Y _4997_/B VGND VGND VPWR VPWR _4994_/X sky130_fd_sc_hd__mux2_1
XFILLER_168_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9521_ _9529_/CLK _9521_/D fanout451/X VGND VGND VPWR VPWR _9521_/Q sky130_fd_sc_hd__dfrtp_1
X_6733_ _6623_/Y _6732_/Y _6959_/A VGND VGND VPWR VPWR _6733_/X sky130_fd_sc_hd__a21o_1
XFILLER_149_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9452_ _9452_/CLK _9452_/D fanout416/X VGND VGND VPWR VPWR _9452_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_177_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6664_ _6778_/A _6664_/B VGND VGND VPWR VPWR _6964_/A sky130_fd_sc_hd__or2_2
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8403_ _9465_/Q _8312_/X _8376_/X _9425_/Q VGND VGND VPWR VPWR _8403_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5615_ _5615_/A VGND VGND VPWR VPWR _8901_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9383_ _9383_/CLK _9383_/D fanout409/X VGND VGND VPWR VPWR _9383_/Q sky130_fd_sc_hd__dfrtp_2
X_6595_ _6597_/A _6503_/A _6413_/B _6217_/B _6507_/A VGND VGND VPWR VPWR _6944_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_192_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8334_ _8392_/A _8357_/A _8357_/B VGND VGND VPWR VPWR _8358_/C sky130_fd_sc_hd__and3_2
XFILLER_129_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5546_ _5546_/A VGND VGND VPWR VPWR _8870_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8265_ _8942_/Q _7988_/X _7990_/X _8872_/Q _8264_/X VGND VGND VPWR VPWR _8272_/A
+ sky130_fd_sc_hd__a221o_1
X_5477_ _5477_/A VGND VGND VPWR VPWR _8840_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7216_ _6012_/X hold779/X _7226_/S VGND VGND VPWR VPWR _7216_/X sky130_fd_sc_hd__mux2_1
X_4428_ _7111_/A _4492_/B VGND VGND VPWR VPWR _4428_/Y sky130_fd_sc_hd__nor2_2
X_8196_ _8196_/A0 _8195_/X _8196_/S VGND VGND VPWR VPWR _8197_/A sky130_fd_sc_hd__mux2_1
Xfanout412 fanout413/X VGND VGND VPWR VPWR fanout412/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout423 fanout424/X VGND VGND VPWR VPWR fanout423/X sky130_fd_sc_hd__clkbuf_4
XFILLER_160_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout434 fanout435/X VGND VGND VPWR VPWR fanout434/X sky130_fd_sc_hd__buf_2
XFILLER_86_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7147_ hold37/X VGND VGND VPWR VPWR _7147_/X sky130_fd_sc_hd__clkbuf_8
Xfanout445 fanout446/X VGND VGND VPWR VPWR fanout445/X sky130_fd_sc_hd__clkbuf_4
X_4359_ hold81/X hold774/X hold73/X VGND VGND VPWR VPWR hold82/A sky130_fd_sc_hd__mux2_1
XFILLER_86_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout456 fanout457/X VGND VGND VPWR VPWR fanout456/X sky130_fd_sc_hd__buf_4
Xfanout467 fanout497/X VGND VGND VPWR VPWR fanout467/X sky130_fd_sc_hd__buf_4
Xfanout478 fanout483/X VGND VGND VPWR VPWR fanout478/X sky130_fd_sc_hd__buf_2
X_7078_ _9141_/Q _5761_/X hold65/X VGND VGND VPWR VPWR _7078_/X sky130_fd_sc_hd__mux2_1
Xfanout489 fanout495/X VGND VGND VPWR VPWR fanout489/X sky130_fd_sc_hd__clkbuf_4
XFILLER_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6029_ _6029_/A VGND VGND VPWR VPWR _9082_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_350 _7264_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_361 _7999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_372 wb_dat_i[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_383 _7695_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_394 _5951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5400_ _5400_/A VGND VGND VPWR VPWR _8812_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6380_ _6504_/A _6380_/B VGND VGND VPWR VPWR _6391_/B sky130_fd_sc_hd__xnor2_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5331_ _5331_/A VGND VGND VPWR VPWR _5331_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_126_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8050_ _8050_/A _8050_/B _8050_/C _8050_/D VGND VGND VPWR VPWR _8050_/X sky130_fd_sc_hd__or4_1
X_5262_ _9403_/Q VGND VGND VPWR VPWR _5262_/Y sky130_fd_sc_hd__inv_2
X_7001_ _7001_/A _7001_/B VGND VGND VPWR VPWR _7002_/D sky130_fd_sc_hd__nor2_1
XFILLER_114_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5193_ _9475_/Q VGND VGND VPWR VPWR _5193_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8952_ _9467_/CLK _8952_/D fanout476/X VGND VGND VPWR VPWR _8952_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_83_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7903_ _7903_/A _7909_/A VGND VGND VPWR VPWR _7903_/Y sky130_fd_sc_hd__nor2_1
X_8883_ _9449_/CLK _8883_/D fanout473/X VGND VGND VPWR VPWR _8883_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_70_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_4_0_csclk clkbuf_3_5_0_csclk/A VGND VGND VPWR VPWR _9210_/CLK sky130_fd_sc_hd__clkbuf_8
X_7834_ _7834_/A VGND VGND VPWR VPWR _9480_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7765_ _5387_/X hold826/X _7779_/S VGND VGND VPWR VPWR _7766_/A sky130_fd_sc_hd__mux2_1
X_4977_ _8788_/Q _4977_/B VGND VGND VPWR VPWR _5127_/B sky130_fd_sc_hd__nand2_1
X_9504_ _9529_/CLK _9504_/D fanout441/X VGND VGND VPWR VPWR _9504_/Q sky130_fd_sc_hd__dfrtp_1
X_6716_ _6716_/A _6716_/B _6742_/B VGND VGND VPWR VPWR _6725_/B sky130_fd_sc_hd__or3_2
X_7696_ _7517_/X hold902/X _7710_/S VGND VGND VPWR VPWR _7697_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9435_ _9475_/CLK _9435_/D fanout491/X VGND VGND VPWR VPWR _9435_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6647_ _6736_/B _6781_/B _6900_/A VGND VGND VPWR VPWR _6661_/A sky130_fd_sc_hd__a21oi_1
XFILLER_165_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9366_ _9367_/CLK _9366_/D fanout422/X VGND VGND VPWR VPWR _9366_/Q sky130_fd_sc_hd__dfrtp_2
X_6578_ _6328_/Y _6551_/Y _6935_/B _6577_/X VGND VGND VPWR VPWR _6578_/X sky130_fd_sc_hd__a211o_1
XFILLER_166_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8317_ _9296_/Q _8314_/X _8316_/X _9280_/Q VGND VGND VPWR VPWR _8317_/X sky130_fd_sc_hd__a22o_1
X_5529_ _5529_/A _5693_/B VGND VGND VPWR VPWR _5538_/S sky130_fd_sc_hd__nand2_4
X_9297_ _9459_/CLK _9297_/D fanout479/X VGND VGND VPWR VPWR _9297_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_59_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8248_ _8966_/Q _7960_/X _7988_/X _8941_/Q _8247_/X VGND VGND VPWR VPWR _8248_/X
+ sky130_fd_sc_hd__a221o_1
X_8179_ _8903_/Q _7962_/A _7988_/A _8938_/Q VGND VGND VPWR VPWR _8179_/X sky130_fd_sc_hd__a22o_1
XFILLER_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4900_ _8888_/Q _5584_/A _4897_/X _4899_/X VGND VGND VPWR VPWR _4922_/B sky130_fd_sc_hd__a211o_1
X_5880_ _9010_/Q hold70/X _5898_/S VGND VGND VPWR VPWR _5880_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4831_ _9305_/Q _7446_/A _7139_/A _9169_/Q VGND VGND VPWR VPWR _4831_/X sky130_fd_sc_hd__a22o_1
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_180 _7973_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_191 _7997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7550_ _7550_/A VGND VGND VPWR VPWR _9350_/D sky130_fd_sc_hd__clkbuf_1
X_4762_ input37/X _4436_/A _6021_/A _9081_/Q _4761_/X VGND VGND VPWR VPWR _4763_/D
+ sky130_fd_sc_hd__a221o_1
X_6501_ _6748_/B _6514_/A _6830_/A _6967_/C VGND VGND VPWR VPWR _6501_/X sky130_fd_sc_hd__o22a_1
XFILLER_147_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7481_ _7481_/A _7499_/B VGND VGND VPWR VPWR _7497_/S sky130_fd_sc_hd__nand2_8
X_4693_ _4693_/A VGND VGND VPWR VPWR _9115_/D sky130_fd_sc_hd__buf_1
X_9220_ _9452_/CLK _9220_/D fanout415/X VGND VGND VPWR VPWR _9220_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_174_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6432_ _6772_/A _6425_/X _6843_/C _6431_/X VGND VGND VPWR VPWR _6432_/X sky130_fd_sc_hd__o211a_1
XFILLER_174_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9151_ _9456_/CLK _9151_/D fanout404/X VGND VGND VPWR VPWR _9151_/Q sky130_fd_sc_hd__dfrtp_4
X_6363_ _6790_/B _6906_/C _6524_/B _6736_/A _6858_/B VGND VGND VPWR VPWR _6363_/X
+ sky130_fd_sc_hd__o32a_1
X_8102_ _9412_/Q _7967_/X _7999_/X _9428_/Q VGND VGND VPWR VPWR _8102_/X sky130_fd_sc_hd__a22o_1
X_5314_ hold23/X hold112/X _5413_/S VGND VGND VPWR VPWR hold24/A sky130_fd_sc_hd__mux2_8
X_9082_ _9162_/CLK _9082_/D fanout439/X VGND VGND VPWR VPWR _9082_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_115_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6294_ _6610_/A VGND VGND VPWR VPWR _6873_/B sky130_fd_sc_hd__buf_4
XFILLER_88_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8033_ _9201_/Q _7938_/X _7949_/X _9241_/Q _8032_/X VGND VGND VPWR VPWR _8037_/C
+ sky130_fd_sc_hd__a221o_1
X_5245_ _9259_/Q VGND VGND VPWR VPWR _5245_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold17 hold17/A VGND VGND VPWR VPWR hold17/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold28 hold28/A VGND VGND VPWR VPWR hold28/X sky130_fd_sc_hd__dlygate4sd3_1
X_5176_ _5176_/A VGND VGND VPWR VPWR _5176_/Y sky130_fd_sc_hd__inv_2
Xhold39 hold39/A VGND VGND VPWR VPWR hold39/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8935_ _9005_/CLK _8935_/D fanout490/X VGND VGND VPWR VPWR _8935_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_43_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8866_ _9251_/CLK _8866_/D fanout485/X VGND VGND VPWR VPWR _8866_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A VGND VGND VPWR VPWR _9541_/CLK sky130_fd_sc_hd__clkbuf_8
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7817_ _7817_/A VGND VGND VPWR VPWR _9472_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8797_ _5168_/A1 _8797_/D _5362_/X VGND VGND VPWR VPWR _8797_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7748_ hold873/X _5761_/A _7762_/S VGND VGND VPWR VPWR _7748_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7679_ _7517_/X hold919/X _7693_/S VGND VGND VPWR VPWR _7680_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9418_ _9466_/CLK _9418_/D fanout475/X VGND VGND VPWR VPWR _9418_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_180_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9349_ _9421_/CLK _9349_/D fanout461/X VGND VGND VPWR VPWR _9349_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold509 _5523_/X VGND VGND VPWR VPWR _5524_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_167_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5030_ _5021_/A _5016_/B _5021_/X VGND VGND VPWR VPWR _5031_/B sky130_fd_sc_hd__a21oi_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1209 _5847_/X VGND VGND VPWR VPWR hold877/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6981_ _6624_/B _6828_/X _6862_/A _6926_/A _6648_/A VGND VGND VPWR VPWR _6982_/D
+ sky130_fd_sc_hd__o221a_1
X_5932_ _5932_/A VGND VGND VPWR VPWR _9040_/D sky130_fd_sc_hd__clkbuf_1
X_8720_ _8720_/A VGND VGND VPWR VPWR _9538_/D sky130_fd_sc_hd__buf_1
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8651_ _8631_/X _8637_/X _8650_/X _8399_/A _8850_/Q VGND VGND VPWR VPWR _8651_/X
+ sky130_fd_sc_hd__o32a_1
X_5863_ _5863_/A VGND VGND VPWR VPWR _5863_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7602_ _7602_/A VGND VGND VPWR VPWR _9374_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4814_ _8880_/Q _5562_/A _5573_/A _8885_/Q VGND VGND VPWR VPWR _4814_/X sky130_fd_sc_hd__a22o_1
X_8582_ _8968_/Q _8657_/B VGND VGND VPWR VPWR _8582_/X sky130_fd_sc_hd__and2_1
X_5794_ _5794_/A VGND VGND VPWR VPWR _8977_/D sky130_fd_sc_hd__clkbuf_1
X_7533_ _7533_/A VGND VGND VPWR VPWR _9342_/D sky130_fd_sc_hd__clkbuf_1
X_4745_ _9347_/Q _7536_/A _7176_/A _9187_/Q _4744_/X VGND VGND VPWR VPWR _4751_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_193_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7464_ hold61/X VGND VGND VPWR VPWR _7479_/S sky130_fd_sc_hd__buf_6
XFILLER_174_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4676_ _8927_/Q _5667_/A _5704_/A _8942_/Q VGND VGND VPWR VPWR _4676_/X sky130_fd_sc_hd__a22o_2
XFILLER_107_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6415_ _6415_/A _6415_/B VGND VGND VPWR VPWR _6518_/A sky130_fd_sc_hd__nand2_4
X_9203_ _9203_/CLK _9203_/D fanout434/X VGND VGND VPWR VPWR _9203_/Q sky130_fd_sc_hd__dfrtp_4
X_7395_ _7395_/A VGND VGND VPWR VPWR _9281_/D sky130_fd_sc_hd__clkbuf_1
X_9134_ _9476_/CLK _9134_/D fanout414/X VGND VGND VPWR VPWR _9134_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_150_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6346_ _6345_/A _6345_/C _6547_/A _6420_/B VGND VGND VPWR VPWR _6346_/X sky130_fd_sc_hd__a31o_1
XFILLER_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9065_ _9110_/CLK _9065_/D VGND VGND VPWR VPWR _9065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6277_ _6869_/A VGND VGND VPWR VPWR _6277_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput107 sram_ro_data[22] VGND VGND VPWR VPWR _4529_/A1 sky130_fd_sc_hd__clkbuf_1
X_8016_ _8653_/S VGND VGND VPWR VPWR _8196_/S sky130_fd_sc_hd__clkbuf_4
Xinput118 sram_ro_data[3] VGND VGND VPWR VPWR _4739_/A1 sky130_fd_sc_hd__clkbuf_2
X_5228_ _9005_/Q _5228_/A1 _9167_/Q VGND VGND VPWR VPWR _5229_/A sky130_fd_sc_hd__mux2_1
Xinput129 usr2_vcc_pwrgood VGND VGND VPWR VPWR _4786_/B2 sky130_fd_sc_hd__clkbuf_4
X_5159_ _8997_/Q VGND VGND VPWR VPWR _8652_/S sky130_fd_sc_hd__inv_2
XFILLER_56_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8918_ _9089_/CLK _8918_/D fanout434/X VGND VGND VPWR VPWR _8918_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_112_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_1_0_csclk clkbuf_2_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_3_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8849_ _9084_/CLK _8849_/D fanout447/X VGND VGND VPWR VPWR _8849_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_80 _5311_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 _5761_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4530_ _4530_/A _4530_/B _4530_/C _4530_/D VGND VGND VPWR VPWR _4549_/B sky130_fd_sc_hd__or4_1
XFILLER_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4461_ _9335_/Q _7499_/A _4460_/Y input28/X VGND VGND VPWR VPWR _4461_/X sky130_fd_sc_hd__a22o_1
Xhold306 _7617_/X VGND VGND VPWR VPWR _7618_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 _7197_/X VGND VGND VPWR VPWR _7198_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 _8912_/Q VGND VGND VPWR VPWR hold328/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 _7068_/X VGND VGND VPWR VPWR _7069_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6200_ _6248_/A _6794_/A _6635_/A VGND VGND VPWR VPWR _6266_/A sky130_fd_sc_hd__or3_4
X_7180_ hold574/X _5809_/X _7192_/S VGND VGND VPWR VPWR _7181_/A sky130_fd_sc_hd__mux2_1
X_4392_ hold59/X VGND VGND VPWR VPWR hold60/A sky130_fd_sc_hd__buf_8
XFILLER_98_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6131_ _6858_/B VGND VGND VPWR VPWR _6589_/D sky130_fd_sc_hd__inv_2
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _6015_/X hold490/X _6064_/S VGND VGND VPWR VPWR _6063_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1006 _9523_/Q VGND VGND VPWR VPWR _8477_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1017 _8765_/X VGND VGND VPWR VPWR _8766_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _5010_/A _5067_/B _5040_/B VGND VGND VPWR VPWR _5013_/X sky130_fd_sc_hd__mux2_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1028 _8786_/Q VGND VGND VPWR VPWR _5055_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1039 hold1161/X VGND VGND VPWR VPWR _5890_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6964_ _6964_/A _6964_/B _6964_/C _6964_/D VGND VGND VPWR VPWR _6965_/C sky130_fd_sc_hd__or4_1
XFILLER_41_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8703_ _5130_/A hold970/X _8013_/A VGND VGND VPWR VPWR _8703_/X sky130_fd_sc_hd__a21o_1
XFILLER_179_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5915_ _5915_/A VGND VGND VPWR VPWR _5915_/X sky130_fd_sc_hd__clkbuf_1
X_6895_ _6895_/A _6895_/B VGND VGND VPWR VPWR _6973_/C sky130_fd_sc_hd__nand2_2
XFILLER_22_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5846_ _5474_/B _5453_/C _5819_/X _5867_/S hold21/A VGND VGND VPWR VPWR _5868_/S
+ sky130_fd_sc_hd__o221a_4
X_8634_ _8920_/Q _8310_/X _8381_/X _8955_/Q _8633_/X VGND VGND VPWR VPWR _8634_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8565_ _9447_/Q _8398_/B _8344_/X _9487_/Q _8564_/X VGND VGND VPWR VPWR _8565_/X
+ sky130_fd_sc_hd__a221o_1
X_5777_ _5777_/A VGND VGND VPWR VPWR _8969_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7516_ _7516_/A VGND VGND VPWR VPWR _9335_/D sky130_fd_sc_hd__clkbuf_1
X_4728_ input46/X _4582_/A _7266_/A _9227_/Q VGND VGND VPWR VPWR _4728_/X sky130_fd_sc_hd__a22o_1
XFILLER_175_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8496_ _9380_/Q _8337_/X _8384_/X _9196_/Q _8495_/X VGND VGND VPWR VPWR _8499_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_175_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7447_ _7302_/X hold876/X _7461_/S VGND VGND VPWR VPWR _7448_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4659_ _7158_/A _7126_/B VGND VGND VPWR VPWR _5607_/A sky130_fd_sc_hd__nor2_4
XFILLER_107_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold840 _9248_/Q VGND VGND VPWR VPWR hold840/X sky130_fd_sc_hd__dlygate4sd3_1
X_7378_ _7378_/A VGND VGND VPWR VPWR _9273_/D sky130_fd_sc_hd__clkbuf_1
Xhold851 hold851/A VGND VGND VPWR VPWR hold851/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 hold862/A VGND VGND VPWR VPWR hold862/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold873 _9440_/Q VGND VGND VPWR VPWR hold873/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold884 hold884/A VGND VGND VPWR VPWR hold884/X sky130_fd_sc_hd__dlygate4sd3_1
X_9117_ _5235__1/A _9117_/D _7024_/X VGND VGND VPWR VPWR _9117_/Q sky130_fd_sc_hd__dfrtn_1
X_6329_ _6334_/B _6329_/B VGND VGND VPWR VPWR _6935_/A sky130_fd_sc_hd__nor2_1
XFILLER_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold895 hold895/A VGND VGND VPWR VPWR hold895/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9048_ _9069_/CLK _9048_/D fanout429/X VGND VGND VPWR VPWR _9048_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_49_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_32_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _9459_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_164_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_47_csclk _8954_/CLK VGND VGND VPWR VPWR _9219_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_48_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5700_ _5650_/X hold396/X _5702_/S VGND VGND VPWR VPWR _5701_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6680_ _6503_/A _6441_/B _6429_/B _6872_/B VGND VGND VPWR VPWR _6704_/C sky130_fd_sc_hd__a31o_1
XFILLER_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5631_ _5629_/X hold849/X _5640_/S VGND VGND VPWR VPWR _5632_/A sky130_fd_sc_hd__mux2_1
X_8350_ _9304_/Q _8341_/X _8344_/X _9480_/Q _8349_/X VGND VGND VPWR VPWR _8351_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_191_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5562_ _5562_/A _5715_/B VGND VGND VPWR VPWR _5571_/S sky130_fd_sc_hd__and2_2
XFILLER_163_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7301_ _7301_/A VGND VGND VPWR VPWR _9239_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4513_ _9222_/Q _7249_/A _7815_/A _9478_/Q VGND VGND VPWR VPWR _4513_/X sky130_fd_sc_hd__a22o_1
X_8281_ _8882_/Q _7969_/X _8077_/X _8937_/Q _8280_/X VGND VGND VPWR VPWR _8282_/D
+ sky130_fd_sc_hd__a221o_1
X_5493_ _5493_/A _5715_/B VGND VGND VPWR VPWR _5502_/S sky130_fd_sc_hd__and2_2
Xhold103 _9551_/Q VGND VGND VPWR VPWR _5292_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold114 _9377_/Q VGND VGND VPWR VPWR hold114/X sky130_fd_sc_hd__dlygate4sd3_1
X_7232_ _7232_/A VGND VGND VPWR VPWR _9209_/D sky130_fd_sc_hd__clkbuf_1
Xhold125 _9321_/Q VGND VGND VPWR VPWR hold125/X sky130_fd_sc_hd__dlygate4sd3_1
X_4444_ _7126_/A _4956_/A VGND VGND VPWR VPWR _4444_/Y sky130_fd_sc_hd__nor2_8
XFILLER_144_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold136 _7214_/X VGND VGND VPWR VPWR _7215_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 _7149_/X VGND VGND VPWR VPWR _9171_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold158 _5582_/X VGND VGND VPWR VPWR _5583_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold169 _8902_/Q VGND VGND VPWR VPWR hold169/X sky130_fd_sc_hd__dlygate4sd3_1
X_7163_ _7163_/A VGND VGND VPWR VPWR _9177_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4375_ _4476_/A _4555_/B VGND VGND VPWR VPWR _4685_/B sky130_fd_sc_hd__nand2_8
XFILLER_113_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6114_ _6167_/A VGND VGND VPWR VPWR _6248_/A sky130_fd_sc_hd__clkinv_4
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7094_ _5951_/X _9148_/Q _7106_/S VGND VGND VPWR VPWR _7094_/X sky130_fd_sc_hd__mux2_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _6045_/A VGND VGND VPWR VPWR _9089_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7996_ _7998_/A _7996_/B _8002_/B VGND VGND VPWR VPWR _7997_/A sky130_fd_sc_hd__and3_2
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6947_ _6736_/A _6732_/B _6736_/B _6876_/B VGND VGND VPWR VPWR _6947_/X sky130_fd_sc_hd__a31o_1
XFILLER_41_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6878_ _6957_/A _6956_/C _6878_/C VGND VGND VPWR VPWR _6880_/C sky130_fd_sc_hd__or3_1
X_8617_ _9075_/Q _8356_/B _8364_/B _8864_/Q _8616_/X VGND VGND VPWR VPWR _8624_/A
+ sky130_fd_sc_hd__a221o_1
X_5829_ _5829_/A VGND VGND VPWR VPWR _5829_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8548_ _9214_/Q _8289_/X _8341_/X _9310_/Q _8547_/X VGND VGND VPWR VPWR _8549_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_185_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8479_ _9468_/Q _8312_/X _8376_/X _9428_/Q VGND VGND VPWR VPWR _8479_/X sky130_fd_sc_hd__a22o_1
XFILLER_123_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold670 _9223_/Q VGND VGND VPWR VPWR hold670/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold681 _9182_/Q VGND VGND VPWR VPWR hold681/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 _7354_/X VGND VGND VPWR VPWR _7355_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput208 _5246_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[10] sky130_fd_sc_hd__buf_12
Xoutput219 _5256_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[20] sky130_fd_sc_hd__buf_12
XFILLER_126_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7850_ _8999_/Q _7850_/B _8015_/B VGND VGND VPWR VPWR _7865_/A sky130_fd_sc_hd__or3_1
XFILLER_36_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6801_ _6906_/A _6435_/A _6858_/B VGND VGND VPWR VPWR _6957_/A sky130_fd_sc_hd__a21oi_2
X_4993_ _4993_/A VGND VGND VPWR VPWR _8803_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7781_ _7781_/A hold21/A VGND VGND VPWR VPWR _7796_/S sky130_fd_sc_hd__nand2_8
X_9520_ _9520_/CLK _9520_/D fanout454/X VGND VGND VPWR VPWR _9520_/Q sky130_fd_sc_hd__dfrtp_1
X_6732_ _6732_/A _6732_/B VGND VGND VPWR VPWR _6732_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9451_ _9459_/CLK _9451_/D fanout480/X VGND VGND VPWR VPWR _9451_/Q sky130_fd_sc_hd__dfrtp_4
X_6663_ _6824_/A _6662_/X _6809_/D VGND VGND VPWR VPWR _6663_/X sky130_fd_sc_hd__o21a_1
XFILLER_149_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5614_ _5311_/X hold399/X _5616_/S VGND VGND VPWR VPWR _5615_/A sky130_fd_sc_hd__mux2_1
X_8402_ _8402_/A VGND VGND VPWR VPWR _8402_/X sky130_fd_sc_hd__buf_8
X_9382_ _9383_/CLK _9382_/D fanout409/X VGND VGND VPWR VPWR _9382_/Q sky130_fd_sc_hd__dfrtp_4
X_6594_ _6873_/B _6871_/B _6530_/D VGND VGND VPWR VPWR _6619_/A sky130_fd_sc_hd__o21ai_1
XFILLER_117_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8333_ _8364_/B VGND VGND VPWR VPWR _8333_/X sky130_fd_sc_hd__buf_8
X_5545_ _5306_/X hold491/X _5549_/S VGND VGND VPWR VPWR _5545_/X sky130_fd_sc_hd__mux2_1
X_8264_ _9073_/Q _7979_/A _7993_/A _8987_/Q VGND VGND VPWR VPWR _8264_/X sky130_fd_sc_hd__a22o_1
XFILLER_105_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_0_0_csclk clkbuf_3_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_0_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_145_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5476_ _5291_/X hold838/X _5490_/S VGND VGND VPWR VPWR _5476_/X sky130_fd_sc_hd__mux2_1
X_4427_ _4878_/A _4665_/A VGND VGND VPWR VPWR _4427_/Y sky130_fd_sc_hd__nor2_4
XFILLER_132_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7215_ _7215_/A VGND VGND VPWR VPWR _9201_/D sky130_fd_sc_hd__clkbuf_1
X_8195_ _8997_/Q _9514_/Q _8193_/X _8194_/X VGND VGND VPWR VPWR _8195_/X sky130_fd_sc_hd__a22o_1
XFILLER_160_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout413 fanout416/X VGND VGND VPWR VPWR fanout413/X sky130_fd_sc_hd__buf_2
X_7146_ _7146_/A VGND VGND VPWR VPWR _7146_/X sky130_fd_sc_hd__clkbuf_1
X_4358_ hold80/X hold22/X _4991_/A VGND VGND VPWR VPWR hold81/A sky130_fd_sc_hd__a21bo_1
Xfanout424 fanout426/X VGND VGND VPWR VPWR fanout424/X sky130_fd_sc_hd__clkbuf_2
Xfanout435 fanout457/X VGND VGND VPWR VPWR fanout435/X sky130_fd_sc_hd__buf_2
Xfanout446 fanout448/X VGND VGND VPWR VPWR fanout446/X sky130_fd_sc_hd__clkbuf_4
XFILLER_48_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout457 input75/X VGND VGND VPWR VPWR fanout457/X sky130_fd_sc_hd__buf_4
XFILLER_86_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout468 fanout497/X VGND VGND VPWR VPWR fanout468/X sky130_fd_sc_hd__buf_2
X_7077_ _7077_/A hold20/X VGND VGND VPWR VPWR hold65/A sky130_fd_sc_hd__and2_1
XFILLER_171_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout479 fanout482/X VGND VGND VPWR VPWR fanout479/X sky130_fd_sc_hd__clkbuf_4
XFILLER_86_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6028_ hold411/X _5687_/X _6030_/S VGND VGND VPWR VPWR _6028_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7979_ _7979_/A VGND VGND VPWR VPWR _7979_/X sky130_fd_sc_hd__buf_6
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_340 _5471_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_351 _7302_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_362 _8003_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_373 wb_dat_i[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_384 fanout457/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_395 _5951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5330_ _5330_/A _5334_/B VGND VGND VPWR VPWR _5331_/A sky130_fd_sc_hd__and2_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5261_ _9387_/Q VGND VGND VPWR VPWR _5261_/Y sky130_fd_sc_hd__inv_2
X_7000_ _7000_/A _7000_/B _7000_/C VGND VGND VPWR VPWR _7004_/B sky130_fd_sc_hd__nor3_1
X_5192_ _5192_/A VGND VGND VPWR VPWR _5192_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8951_ _9005_/CLK _8951_/D fanout489/X VGND VGND VPWR VPWR _8951_/Q sky130_fd_sc_hd__dfrtp_4
X_7902_ _7902_/A _7902_/B VGND VGND VPWR VPWR _7909_/A sky130_fd_sc_hd__nor2_1
X_8882_ _9089_/CLK _8882_/D fanout433/X VGND VGND VPWR VPWR _8882_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7833_ _5387_/X hold859/X _7847_/S VGND VGND VPWR VPWR _7834_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7764_ _7764_/A hold21/A VGND VGND VPWR VPWR _7779_/S sky130_fd_sc_hd__nand2_8
X_4976_ _8790_/Q _8789_/Q VGND VGND VPWR VPWR _4977_/B sky130_fd_sc_hd__nor2_1
X_9503_ _9532_/CLK _9503_/D fanout441/X VGND VGND VPWR VPWR _9503_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_189_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6715_ _6897_/A _6715_/B VGND VGND VPWR VPWR _6742_/B sky130_fd_sc_hd__nor2_1
XFILLER_20_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7695_ _7695_/A _7695_/B VGND VGND VPWR VPWR _7710_/S sky130_fd_sc_hd__nand2_8
XFILLER_149_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9434_ _9434_/CLK _9434_/D fanout450/X VGND VGND VPWR VPWR _9434_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_177_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6646_ _6646_/A _6987_/C _6977_/B _6646_/D VGND VGND VPWR VPWR _6646_/X sky130_fd_sc_hd__or4_1
XFILLER_177_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9365_ _9453_/CLK _9365_/D fanout461/X VGND VGND VPWR VPWR _9365_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6577_ _6217_/B _6551_/Y _6872_/C _6576_/X VGND VGND VPWR VPWR _6577_/X sky130_fd_sc_hd__a211o_1
XFILLER_164_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8316_ _8358_/B VGND VGND VPWR VPWR _8316_/X sky130_fd_sc_hd__buf_6
X_5528_ _5528_/A VGND VGND VPWR VPWR _8862_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9296_ _9328_/CLK _9296_/D fanout463/X VGND VGND VPWR VPWR _9296_/Q sky130_fd_sc_hd__dfstp_2
X_5459_ _5306_/X hold456/X _5472_/S VGND VGND VPWR VPWR _5459_/X sky130_fd_sc_hd__mux2_1
X_8247_ _8881_/Q _7969_/X _7981_/X _8916_/Q VGND VGND VPWR VPWR _8247_/X sky130_fd_sc_hd__a22o_1
XFILLER_79_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8178_ _9084_/Q _7940_/A _7969_/A _8878_/Q _8177_/X VGND VGND VPWR VPWR _8184_/B
+ sky130_fd_sc_hd__a221o_1
X_7129_ _7129_/A _7139_/B VGND VGND VPWR VPWR _7130_/S sky130_fd_sc_hd__nand2_1
XFILLER_87_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4830_ _7126_/A _5474_/B VGND VGND VPWR VPWR _7139_/A sky130_fd_sc_hd__nor2_4
XFILLER_61_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_170 _7960_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_181 _7977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_192 _7997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4761_ _9234_/Q _7284_/A _5296_/A _8774_/Q VGND VGND VPWR VPWR _4761_/X sky130_fd_sc_hd__a22o_1
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6500_ _6500_/A VGND VGND VPWR VPWR _6967_/C sky130_fd_sc_hd__buf_4
X_7480_ _7480_/A VGND VGND VPWR VPWR _9319_/D sky130_fd_sc_hd__clkbuf_1
X_4692_ _4691_/X _9115_/Q _4964_/B VGND VGND VPWR VPWR _4693_/A sky130_fd_sc_hd__mux2_2
XFILLER_174_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6431_ _6635_/B _6874_/A _6524_/C _6830_/A VGND VGND VPWR VPWR _6431_/X sky130_fd_sc_hd__o22a_1
XFILLER_146_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9150_ _9456_/CLK _9150_/D fanout407/X VGND VGND VPWR VPWR _9150_/Q sky130_fd_sc_hd__dfrtp_4
X_6362_ _6588_/B _6708_/B _6362_/C _6362_/D VGND VGND VPWR VPWR _6364_/C sky130_fd_sc_hd__or4_1
X_5313_ _5313_/A VGND VGND VPWR VPWR _8775_/D sky130_fd_sc_hd__clkbuf_1
X_8101_ _9236_/Q _8034_/X _8098_/X _8100_/X VGND VGND VPWR VPWR _8104_/C sky130_fd_sc_hd__a211o_1
X_6293_ _6754_/A _6754_/B _6585_/A _6291_/X _6292_/X VGND VGND VPWR VPWR _6293_/X
+ sky130_fd_sc_hd__o41a_1
X_9081_ _9161_/CLK _9081_/D fanout441/X VGND VGND VPWR VPWR _9081_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_142_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5244_ _9251_/Q VGND VGND VPWR VPWR _5244_/Y sky130_fd_sc_hd__inv_2
X_8032_ _9209_/Q _7923_/X _7988_/X _9433_/Q VGND VGND VPWR VPWR _8032_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold18 hold18/A VGND VGND VPWR VPWR hold18/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 hold29/A VGND VGND VPWR VPWR hold29/X sky130_fd_sc_hd__dlygate4sd3_1
X_5175_ _5175_/A VGND VGND VPWR VPWR _5176_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_130_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8934_ _9005_/CLK _8934_/D fanout490/X VGND VGND VPWR VPWR _8934_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_45_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8865_ _9005_/CLK _8865_/D fanout489/X VGND VGND VPWR VPWR _8865_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_52_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7816_ _5387_/X hold842/X _7830_/S VGND VGND VPWR VPWR _7817_/A sky130_fd_sc_hd__mux2_1
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8796_ _8831_/CLK _8796_/D _5360_/X VGND VGND VPWR VPWR _8796_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7747_ _7747_/A VGND VGND VPWR VPWR _7762_/S sky130_fd_sc_hd__buf_6
X_4959_ _4959_/A _4959_/B VGND VGND VPWR VPWR _4960_/D sky130_fd_sc_hd__or2_1
XFILLER_61_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7678_ _7678_/A _7695_/B VGND VGND VPWR VPWR _7693_/S sky130_fd_sc_hd__nand2_8
XFILLER_177_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9417_ _9459_/CLK _9417_/D fanout479/X VGND VGND VPWR VPWR hold88/A sky130_fd_sc_hd__dfstp_1
X_6629_ _6714_/B _6865_/A _6629_/C _6628_/X VGND VGND VPWR VPWR _6629_/X sky130_fd_sc_hd__or4b_1
XFILLER_20_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9348_ _9370_/CLK _9348_/D fanout466/X VGND VGND VPWR VPWR _9348_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9279_ _9471_/CLK _9279_/D _5070_/A VGND VGND VPWR VPWR _9279_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_79_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6980_ _9109_/Q _8735_/A _6965_/Y _6970_/X _6979_/X VGND VGND VPWR VPWR _6980_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5931_ _9040_/Q _4961_/X _5945_/S VGND VGND VPWR VPWR _5932_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8650_ _8650_/A _8650_/B _8650_/C VGND VGND VPWR VPWR _8650_/X sky130_fd_sc_hd__or3_1
XFILLER_179_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5862_ _9005_/Q hold16/X _5868_/S VGND VGND VPWR VPWR _5862_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7601_ _7494_/X hold727/X hold75/X VGND VGND VPWR VPWR _7602_/A sky130_fd_sc_hd__mux2_1
X_4813_ _5012_/A _5897_/S _5506_/A _8855_/Q _4812_/X VGND VGND VPWR VPWR _4816_/C
+ sky130_fd_sc_hd__a221o_1
X_8581_ _8958_/Q _8402_/X _8378_/X _8943_/Q _8580_/X VGND VGND VPWR VPWR _8588_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_33_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5793_ hold641/X _5690_/X _5793_/S VGND VGND VPWR VPWR _5794_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7532_ _7494_/X hold730/X _7534_/S VGND VGND VPWR VPWR _7532_/X sky130_fd_sc_hd__mux2_1
X_4744_ _9275_/Q _4938_/A2 _5562_/A _8881_/Q VGND VGND VPWR VPWR _4744_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4675_ _5453_/B _4675_/B VGND VGND VPWR VPWR _5704_/A sky130_fd_sc_hd__nor2_4
X_7463_ _7463_/A hold19/X VGND VGND VPWR VPWR hold61/A sky130_fd_sc_hd__and2_1
XFILLER_162_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9202_ _9328_/CLK _9202_/D fanout463/X VGND VGND VPWR VPWR _9202_/Q sky130_fd_sc_hd__dfrtp_2
X_6414_ _6435_/A _6514_/A VGND VGND VPWR VPWR _6922_/A sky130_fd_sc_hd__nor2_1
XFILLER_174_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7394_ _7359_/X hold143/X _7406_/S VGND VGND VPWR VPWR _7395_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9133_ _9484_/CLK _9133_/D fanout428/X VGND VGND VPWR VPWR _9133_/Q sky130_fd_sc_hd__dfstp_1
X_6345_ _6345_/A _6345_/B _6345_/C VGND VGND VPWR VPWR _6345_/X sky130_fd_sc_hd__and3_2
XFILLER_88_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9064_ _9110_/CLK _9064_/D VGND VGND VPWR VPWR _9064_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6276_ _6736_/A _6800_/A VGND VGND VPWR VPWR _6869_/A sky130_fd_sc_hd__nor2_1
XFILLER_115_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8015_ _8015_/A _8015_/B VGND VGND VPWR VPWR _8653_/S sky130_fd_sc_hd__nor2_2
Xinput108 sram_ro_data[23] VGND VGND VPWR VPWR _4503_/B2 sky130_fd_sc_hd__clkbuf_1
X_5227_ _5227_/A VGND VGND VPWR VPWR _9568_/A sky130_fd_sc_hd__buf_1
Xinput119 sram_ro_data[4] VGND VGND VPWR VPWR _4601_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5158_ _8998_/Q VGND VGND VPWR VPWR _7902_/B sky130_fd_sc_hd__buf_4
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5089_ _9387_/Q VGND VGND VPWR VPWR _5089_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8917_ _9449_/CLK _8917_/D fanout474/X VGND VGND VPWR VPWR _8917_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_71_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8848_ _8852_/CLK _8848_/D fanout443/X VGND VGND VPWR VPWR _8848_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8779_ _8779_/CLK _8779_/D _5076_/X VGND VGND VPWR VPWR _8779_/Q sky130_fd_sc_hd__dfstp_1
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_70 _5223_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_81 _5311_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_92 _5761_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4460_ _4858_/B _4499_/A VGND VGND VPWR VPWR _4460_/Y sky130_fd_sc_hd__nor2_8
Xhold307 _9244_/Q VGND VGND VPWR VPWR hold307/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold318 _9276_/Q VGND VGND VPWR VPWR hold318/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 _5640_/X VGND VGND VPWR VPWR _5641_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4391_ hold58/X _4391_/B VGND VGND VPWR VPWR hold59/A sky130_fd_sc_hd__or2_1
XFILLER_98_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6130_ _6130_/A VGND VGND VPWR VPWR _6858_/B sky130_fd_sc_hd__buf_4
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _6061_/A VGND VGND VPWR VPWR _9096_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5012_ _5012_/A VGND VGND VPWR VPWR _5067_/B sky130_fd_sc_hd__buf_8
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1007 _9509_/Q VGND VGND VPWR VPWR _8062_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1018 _9501_/Q VGND VGND VPWR VPWR _7903_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 hold36/A VGND VGND VPWR VPWR _5065_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6963_ _6906_/A _6736_/B _6858_/B VGND VGND VPWR VPWR _6964_/B sky130_fd_sc_hd__a21oi_1
X_8702_ _8852_/Q _8400_/B _8701_/X _8105_/X VGND VGND VPWR VPWR _8702_/X sky130_fd_sc_hd__o211a_1
X_5914_ _5468_/X _9584_/A _5916_/S VGND VGND VPWR VPWR _5914_/X sky130_fd_sc_hd__mux2_1
X_6894_ _6894_/A _6894_/B VGND VGND VPWR VPWR _6902_/A sky130_fd_sc_hd__nor2_1
X_8633_ _8915_/Q _8298_/A _8370_/A _9086_/Q VGND VGND VPWR VPWR _8633_/X sky130_fd_sc_hd__a22o_1
X_5845_ hold838/X _7517_/A _5867_/S VGND VGND VPWR VPWR _5845_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8564_ _9223_/Q _8391_/X _8367_/X _9479_/Q VGND VGND VPWR VPWR _8564_/X sky130_fd_sc_hd__a22o_1
X_5776_ _5633_/X hold458/X _5782_/S VGND VGND VPWR VPWR _5777_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7515_ _7514_/X hold636/X _7515_/S VGND VGND VPWR VPWR _7515_/X sky130_fd_sc_hd__mux2_1
X_4727_ input95/X _4488_/Y _5296_/A _8775_/Q VGND VGND VPWR VPWR _4731_/B sky130_fd_sc_hd__a22o_1
X_8495_ _9436_/Q _7908_/X _8335_/X _9276_/Q VGND VGND VPWR VPWR _8495_/X sky130_fd_sc_hd__a22o_1
XFILLER_135_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7446_ _7446_/A _7499_/B VGND VGND VPWR VPWR _7461_/S sky130_fd_sc_hd__nand2_8
X_4658_ _9364_/Q _7571_/A _7043_/A _9130_/Q _4657_/X VGND VGND VPWR VPWR _4673_/A
+ sky130_fd_sc_hd__a221o_1
Xinput90 spimemio_flash_io2_oeb VGND VGND VPWR VPWR input90/X sky130_fd_sc_hd__clkbuf_2
Xhold830 _8913_/Q VGND VGND VPWR VPWR hold830/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 hold841/A VGND VGND VPWR VPWR hold841/X sky130_fd_sc_hd__dlygate4sd3_1
X_7377_ _7359_/X hold393/X _7389_/S VGND VGND VPWR VPWR _7378_/A sky130_fd_sc_hd__mux2_1
X_4589_ _4589_/A1 _4444_/Y _5388_/A _8814_/Q _4588_/X VGND VGND VPWR VPWR _4590_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold852 _9312_/Q VGND VGND VPWR VPWR hold852/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold863 _7033_/X VGND VGND VPWR VPWR _7034_/A sky130_fd_sc_hd__dlygate4sd3_1
X_9116_ _5235__1/A _9116_/D _7022_/X VGND VGND VPWR VPWR _9116_/Q sky130_fd_sc_hd__dfrtn_1
Xhold874 _7748_/X VGND VGND VPWR VPWR _7749_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6328_ _6329_/B VGND VGND VPWR VPWR _6328_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold885 _7044_/X VGND VGND VPWR VPWR _7045_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold896 _5877_/X VGND VGND VPWR VPWR _5878_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9047_ _9541_/CLK _9047_/D VGND VGND VPWR VPWR _9047_/Q sky130_fd_sc_hd__dfxtp_1
X_6259_ _6338_/A VGND VGND VPWR VPWR _7001_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_131_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5630_ _5630_/A _5693_/B VGND VGND VPWR VPWR _5640_/S sky130_fd_sc_hd__nand2_4
XFILLER_85_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5561_ _5561_/A VGND VGND VPWR VPWR _8877_/D sky130_fd_sc_hd__clkbuf_1
X_7300_ _7299_/X hold562/X _7300_/S VGND VGND VPWR VPWR _7300_/X sky130_fd_sc_hd__mux2_1
X_4512_ _4512_/A VGND VGND VPWR VPWR _9118_/D sky130_fd_sc_hd__clkbuf_1
X_5492_ hold20/A VGND VGND VPWR VPWR _5715_/B sky130_fd_sc_hd__buf_2
X_8280_ _9052_/Q _7923_/X _7953_/B _8877_/Q VGND VGND VPWR VPWR _8280_/X sky130_fd_sc_hd__a22o_1
Xhold104 _5292_/X VGND VGND VPWR VPWR hold104/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 _9233_/Q VGND VGND VPWR VPWR hold115/X sky130_fd_sc_hd__dlygate4sd3_1
X_7231_ _7147_/X hold295/X _7247_/S VGND VGND VPWR VPWR _7231_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold126 _7484_/X VGND VGND VPWR VPWR _7485_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4443_ _4489_/A _4465_/B VGND VGND VPWR VPWR _4956_/A sky130_fd_sc_hd__nand2_8
Xhold137 _8844_/Q VGND VGND VPWR VPWR hold137/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold148 _9337_/Q VGND VGND VPWR VPWR hold148/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold159 _9103_/Q VGND VGND VPWR VPWR hold159/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4374_ hold10/X _4468_/B VGND VGND VPWR VPWR _4465_/B sky130_fd_sc_hd__nor2b_4
X_7162_ _7147_/X hold182/X _7174_/S VGND VGND VPWR VPWR _7162_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6113_ _6402_/A VGND VGND VPWR VPWR _6589_/C sky130_fd_sc_hd__inv_2
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7093_ _7093_/A VGND VGND VPWR VPWR _9147_/D sky130_fd_sc_hd__clkbuf_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ hold883/X _5761_/X _6053_/S VGND VGND VPWR VPWR _6045_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7995_ _9432_/Q _7988_/X _7990_/X _9272_/Q _7994_/X VGND VGND VPWR VPWR _8006_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_26_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6946_ _6946_/A _6946_/B _6946_/C _6945_/X VGND VGND VPWR VPWR _6951_/B sky130_fd_sc_hd__or4b_1
XFILLER_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6877_ _6955_/A _6955_/B _6955_/C _6955_/D VGND VGND VPWR VPWR _6878_/C sky130_fd_sc_hd__or4_1
X_8616_ _8874_/Q _8358_/B _8364_/A _9090_/Q VGND VGND VPWR VPWR _8616_/X sky130_fd_sc_hd__a22o_1
X_5828_ _9572_/A _5827_/X hold43/X VGND VGND VPWR VPWR _5828_/X sky130_fd_sc_hd__mux2_1
XFILLER_167_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8547_ _9398_/Q _8304_/X _8324_/X _9246_/Q VGND VGND VPWR VPWR _8547_/X sky130_fd_sc_hd__a22o_1
X_5759_ hold642/X _5690_/X _5759_/S VGND VGND VPWR VPWR _5760_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8478_ _8478_/A VGND VGND VPWR VPWR _9523_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7429_ _7429_/A VGND VGND VPWR VPWR _9297_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold660 _5912_/X VGND VGND VPWR VPWR _5913_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 _7264_/X VGND VGND VPWR VPWR _7265_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold682 _7172_/X VGND VGND VPWR VPWR _7173_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 _7256_/X VGND VGND VPWR VPWR _7257_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput209 _5247_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[11] sky130_fd_sc_hd__buf_12
XFILLER_126_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6800_ _6800_/A _7001_/B VGND VGND VPWR VPWR _6959_/D sky130_fd_sc_hd__nor2_1
XFILLER_91_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7780_ _7780_/A VGND VGND VPWR VPWR _9455_/D sky130_fd_sc_hd__clkbuf_1
X_4992_ _4991_/Y hold55/A _5014_/S VGND VGND VPWR VPWR _4993_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6731_ _6725_/A _6730_/X _6616_/D VGND VGND VPWR VPWR _6851_/D sky130_fd_sc_hd__o21bai_1
XFILLER_189_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9450_ _9474_/CLK _9450_/D fanout427/X VGND VGND VPWR VPWR _9450_/Q sky130_fd_sc_hd__dfrtp_4
X_6662_ _6521_/B _6634_/Y _6646_/X _6661_/X VGND VGND VPWR VPWR _6662_/X sky130_fd_sc_hd__a211o_1
XFILLER_176_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8401_ _7920_/Y _8397_/X _8400_/X _8013_/X hold946/X VGND VGND VPWR VPWR _9520_/D
+ sky130_fd_sc_hd__a32o_1
X_5613_ _5613_/A VGND VGND VPWR VPWR _8900_/D sky130_fd_sc_hd__clkbuf_1
X_9381_ _9421_/CLK _9381_/D fanout461/X VGND VGND VPWR VPWR _9381_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6593_ _6736_/B _6531_/X _6209_/X VGND VGND VPWR VPWR _6863_/C sky130_fd_sc_hd__o21ai_1
XFILLER_176_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8332_ _8375_/A _8357_/A _8357_/B VGND VGND VPWR VPWR _8364_/B sky130_fd_sc_hd__and3_2
X_5544_ _5544_/A VGND VGND VPWR VPWR _8869_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8263_ hold985/X _8196_/S _8261_/X _8262_/X VGND VGND VPWR VPWR _8263_/X sky130_fd_sc_hd__o22a_1
XFILLER_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5475_ _5475_/A VGND VGND VPWR VPWR _5490_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_145_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7214_ _7147_/X hold135/X _7226_/S VGND VGND VPWR VPWR _7214_/X sky130_fd_sc_hd__mux2_1
X_4426_ _4674_/A VGND VGND VPWR VPWR _4665_/A sky130_fd_sc_hd__buf_12
XFILLER_160_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8194_ _8848_/Q _8009_/A _8652_/S VGND VGND VPWR VPWR _8194_/X sky130_fd_sc_hd__o21a_1
XFILLER_132_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout414 fanout415/X VGND VGND VPWR VPWR fanout414/X sky130_fd_sc_hd__clkbuf_4
X_7145_ _7128_/X _9170_/Q _7156_/S VGND VGND VPWR VPWR _7145_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4357_ hold55/X _5021_/B VGND VGND VPWR VPWR _4991_/A sky130_fd_sc_hd__nand2_1
Xfanout425 fanout426/X VGND VGND VPWR VPWR fanout425/X sky130_fd_sc_hd__buf_4
XFILLER_113_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout436 fanout439/X VGND VGND VPWR VPWR fanout436/X sky130_fd_sc_hd__clkbuf_4
XFILLER_98_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout447 fanout448/X VGND VGND VPWR VPWR fanout447/X sky130_fd_sc_hd__clkbuf_4
Xfanout458 fanout459/X VGND VGND VPWR VPWR fanout458/X sky130_fd_sc_hd__clkbuf_4
X_7076_ _7076_/A VGND VGND VPWR VPWR _9140_/D sky130_fd_sc_hd__clkbuf_1
Xfanout469 fanout497/X VGND VGND VPWR VPWR fanout469/X sky130_fd_sc_hd__buf_4
XFILLER_100_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6027_ _6027_/A VGND VGND VPWR VPWR _9081_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7978_ _8181_/B _7996_/B _7992_/C VGND VGND VPWR VPWR _7979_/A sky130_fd_sc_hd__and3_2
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6929_ _6770_/C _6929_/B _6929_/C VGND VGND VPWR VPWR _6929_/Y sky130_fd_sc_hd__nand3b_1
Xclkbuf_leaf_31_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _9475_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_168_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9579_ _9579_/A _5089_/Y VGND VGND VPWR VPWR mgmt_gpio_out[25] sky130_fd_sc_hd__ebufn_8
XFILLER_183_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_46_csclk _8954_/CLK VGND VGND VPWR VPWR _9195_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_136_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold490 _9097_/Q VGND VGND VPWR VPWR hold490/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_0_0_wb_clk_i rebuffer3/A VGND VGND VPWR VPWR clkbuf_1_0_1_wb_clk_i/A sky130_fd_sc_hd__clkbuf_8
XFILLER_2_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1190 _9404_/Q VGND VGND VPWR VPWR hold373/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_330 _5187_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_341 _5761_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_352 _7302_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_363 _8346_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_374 input96/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_385 fanout457/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_396 _5951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5260_ _9379_/Q VGND VGND VPWR VPWR _5260_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5191_ _5190_/Y input92/X _5194_/S VGND VGND VPWR VPWR _5192_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8950_ _9419_/CLK _8950_/D fanout489/X VGND VGND VPWR VPWR _8950_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_49_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7901_ _7901_/A1 _7887_/B _7898_/Y _7900_/X VGND VGND VPWR VPWR _9500_/D sky130_fd_sc_hd__a31o_1
X_8881_ _9084_/CLK _8881_/D fanout444/X VGND VGND VPWR VPWR _8881_/Q sky130_fd_sc_hd__dfrtp_4
X_7832_ _7832_/A hold21/A VGND VGND VPWR VPWR _7847_/S sky130_fd_sc_hd__nand2_8
X_7763_ _7763_/A VGND VGND VPWR VPWR _9447_/D sky130_fd_sc_hd__clkbuf_1
X_4975_ _4975_/A VGND VGND VPWR VPWR _5016_/B sky130_fd_sc_hd__clkbuf_2
X_9502_ _9520_/CLK _9502_/D fanout470/X VGND VGND VPWR VPWR _9502_/Q sky130_fd_sc_hd__dfrtp_2
X_6714_ _6754_/A _6714_/B _6292_/X VGND VGND VPWR VPWR _6865_/B sky130_fd_sc_hd__or3b_2
XFILLER_149_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7694_ _7694_/A VGND VGND VPWR VPWR _9415_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9433_ _9475_/CLK _9433_/D fanout481/X VGND VGND VPWR VPWR _9433_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_20_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6645_ _6660_/B _6641_/X _6642_/Y _6997_/A _6644_/X VGND VGND VPWR VPWR _6646_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_109_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9364_ _9468_/CLK _9364_/D fanout466/X VGND VGND VPWR VPWR _9364_/Q sky130_fd_sc_hd__dfrtp_4
X_6576_ _6857_/A _6576_/B _6576_/C _6576_/D VGND VGND VPWR VPWR _6576_/X sky130_fd_sc_hd__or4_1
XFILLER_166_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8315_ _8389_/A _8357_/A _8389_/C VGND VGND VPWR VPWR _8358_/B sky130_fd_sc_hd__and3_2
XFILLER_192_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5527_ _5315_/X hold186/X _5527_/S VGND VGND VPWR VPWR _5527_/X sky130_fd_sc_hd__mux2_1
X_9295_ _9398_/CLK _9295_/D _5070_/A VGND VGND VPWR VPWR _9295_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_145_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8246_ _8976_/Q _7947_/X _7997_/X _8956_/Q VGND VGND VPWR VPWR _8246_/X sky130_fd_sc_hd__a22o_1
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5458_ _5458_/A VGND VGND VPWR VPWR _8833_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4409_ _4656_/A _4861_/A VGND VGND VPWR VPWR _4409_/Y sky130_fd_sc_hd__nor2_2
XFILLER_132_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8177_ _8873_/Q _7952_/A _8003_/A _8883_/Q VGND VGND VPWR VPWR _8177_/X sky130_fd_sc_hd__a22o_1
X_5389_ _5389_/A VGND VGND VPWR VPWR _5416_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_120_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7128_ _7517_/A VGND VGND VPWR VPWR _7128_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7059_ _7059_/A VGND VGND VPWR VPWR _9132_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_160 _7949_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_171 _7960_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_182 _7979_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_193 _8001_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4760_ _9314_/Q _7463_/A _7043_/A _9128_/Q VGND VGND VPWR VPWR _4763_/C sky130_fd_sc_hd__a22o_2
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4691_ _9114_/Q _5988_/A1 _4886_/S VGND VGND VPWR VPWR _4691_/X sky130_fd_sc_hd__mux2_2
XFILLER_119_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6430_ _6492_/B VGND VGND VPWR VPWR _6830_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_146_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6361_ _6673_/A _6839_/A _6314_/X _6360_/X VGND VGND VPWR VPWR _6362_/D sky130_fd_sc_hd__a211o_1
XFILLER_174_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8100_ _9244_/Q _7949_/X _7973_/X _9196_/Q _8099_/X VGND VGND VPWR VPWR _8100_/X
+ sky130_fd_sc_hd__a221o_1
X_5312_ _5311_/X hold397/X _5316_/S VGND VGND VPWR VPWR _5313_/A sky130_fd_sc_hd__mux2_1
X_9080_ _9162_/CLK _9080_/D fanout440/X VGND VGND VPWR VPWR _9080_/Q sky130_fd_sc_hd__dfrtp_4
X_6292_ _6479_/A _6895_/A _9034_/Q VGND VGND VPWR VPWR _6292_/X sky130_fd_sc_hd__o21a_1
X_8031_ _9281_/Q _7953_/B _7969_/X _9289_/Q _8030_/X VGND VGND VPWR VPWR _8037_/B
+ sky130_fd_sc_hd__a221o_1
X_5243_ _9243_/Q VGND VGND VPWR VPWR _5243_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold19 hold19/A VGND VGND VPWR VPWR hold19/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5174_ _8794_/Q _5174_/B VGND VGND VPWR VPWR _5175_/A sky130_fd_sc_hd__or2_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8933_ _9467_/CLK _8933_/D fanout476/X VGND VGND VPWR VPWR _8933_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8864_ _9005_/CLK _8864_/D fanout484/X VGND VGND VPWR VPWR _8864_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_52_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7815_ _7815_/A hold21/A VGND VGND VPWR VPWR _7830_/S sky130_fd_sc_hd__nand2_8
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8795_ _5168_/A1 _8795_/D _5357_/X VGND VGND VPWR VPWR _8795_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7746_ _7746_/A hold19/X VGND VGND VPWR VPWR _7747_/A sky130_fd_sc_hd__and2_1
X_4958_ _9304_/Q _7446_/A _5506_/A _8853_/Q _4957_/X VGND VGND VPWR VPWR _4959_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_184_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7677_ _7677_/A VGND VGND VPWR VPWR _9407_/D sky130_fd_sc_hd__clkbuf_1
X_4889_ _5474_/B VGND VGND VPWR VPWR _4889_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9416_ _9416_/CLK _9416_/D fanout426/X VGND VGND VPWR VPWR _9416_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6628_ _6628_/A _6628_/B _6858_/B VGND VGND VPWR VPWR _6628_/X sky130_fd_sc_hd__or3_1
XFILLER_137_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9347_ _9427_/CLK _9347_/D fanout478/X VGND VGND VPWR VPWR _9347_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_153_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6559_ _6559_/A VGND VGND VPWR VPWR _6560_/B sky130_fd_sc_hd__inv_2
XFILLER_193_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9278_ _9398_/CLK _9278_/D fanout426/X VGND VGND VPWR VPWR _9278_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_105_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8229_ _9050_/Q _7923_/X _8020_/X _8945_/Q VGND VGND VPWR VPWR _8229_/X sky130_fd_sc_hd__a22o_1
XFILLER_121_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5930_ _5930_/A VGND VGND VPWR VPWR _5945_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_19_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5861_ _8845_/Q hold15/X _5867_/S VGND VGND VPWR VPWR hold16/A sky130_fd_sc_hd__mux2_1
X_7600_ _7600_/A VGND VGND VPWR VPWR _9373_/D sky130_fd_sc_hd__clkbuf_1
X_4812_ input94/X _4488_/Y _4449_/Y _9242_/Q VGND VGND VPWR VPWR _4812_/X sky130_fd_sc_hd__a22o_1
X_8580_ _8898_/Q _8312_/X _8376_/X _8948_/Q VGND VGND VPWR VPWR _8580_/X sky130_fd_sc_hd__a22o_1
X_5792_ _5792_/A VGND VGND VPWR VPWR _8976_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7531_ _7531_/A VGND VGND VPWR VPWR _9341_/D sky130_fd_sc_hd__clkbuf_1
X_4743_ _8820_/Q _5418_/A _5607_/A _8901_/Q _4742_/X VGND VGND VPWR VPWR _4751_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7462_ _7462_/A VGND VGND VPWR VPWR _9311_/D sky130_fd_sc_hd__clkbuf_1
X_4674_ _4674_/A _7126_/B VGND VGND VPWR VPWR _5667_/A sky130_fd_sc_hd__nor2_8
XFILLER_119_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9201_ _9483_/CLK _9201_/D fanout473/X VGND VGND VPWR VPWR _9201_/Q sky130_fd_sc_hd__dfstp_1
X_6413_ _6503_/A _6413_/B VGND VGND VPWR VPWR _6514_/A sky130_fd_sc_hd__nand2_4
XFILLER_135_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7393_ _7393_/A VGND VGND VPWR VPWR _9280_/D sky130_fd_sc_hd__clkbuf_1
X_9132_ _9474_/CLK _9132_/D fanout427/X VGND VGND VPWR VPWR _9132_/Q sky130_fd_sc_hd__dfstp_1
X_6344_ _6344_/A _6344_/B VGND VGND VPWR VPWR _6345_/C sky130_fd_sc_hd__and2_1
XFILLER_115_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9063_ _9110_/CLK _9063_/D VGND VGND VPWR VPWR _9063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6275_ _6311_/B _6871_/B _6217_/Y _6272_/X _6274_/X VGND VGND VPWR VPWR _6275_/X
+ sky130_fd_sc_hd__o2111a_1
X_8014_ _7920_/Y _8007_/X _8010_/X _8013_/X hold953/X VGND VGND VPWR VPWR _9507_/D
+ sky130_fd_sc_hd__a32o_1
Xinput109 sram_ro_data[24] VGND VGND VPWR VPWR _4951_/B2 sky130_fd_sc_hd__clkbuf_2
X_5226_ _9006_/Q _5226_/A1 _9165_/Q VGND VGND VPWR VPWR _5227_/A sky130_fd_sc_hd__mux2_4
XFILLER_102_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5157_ hold999/X _5068_/C _5016_/B _5019_/A VGND VGND VPWR VPWR _8831_/D sky130_fd_sc_hd__a31o_1
XFILLER_29_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5088_ _9395_/Q VGND VGND VPWR VPWR _5088_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8916_ _9005_/CLK _8916_/D fanout490/X VGND VGND VPWR VPWR _8916_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_71_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8847_ _9172_/CLK _8847_/D fanout491/X VGND VGND VPWR VPWR _8847_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8778_ _8831_/CLK _8778_/D _5321_/X VGND VGND VPWR VPWR _8778_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7729_ _7729_/A hold21/A VGND VGND VPWR VPWR hold86/A sky130_fd_sc_hd__nand2_8
XFILLER_8_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_60 _4949_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_71 _5231_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_82 _5387_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_93 _5629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold308 _7313_/X VGND VGND VPWR VPWR _7314_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold319 _7383_/X VGND VGND VPWR VPWR _7384_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4390_ hold82/A hold51/X VGND VGND VPWR VPWR _4391_/B sky130_fd_sc_hd__nand2_1
XFILLER_125_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _6012_/X hold600/X _6064_/S VGND VGND VPWR VPWR _6061_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1008 _8829_/Q VGND VGND VPWR VPWR _5128_/B2 sky130_fd_sc_hd__dlygate4sd3_1
X_5011_ _5011_/A _5011_/B VGND VGND VPWR VPWR _8799_/D sky130_fd_sc_hd__xnor2_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1019 _8999_/Q VGND VGND VPWR VPWR _7919_/A3 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6962_ _7000_/A _7000_/B _7000_/C _7003_/C VGND VGND VPWR VPWR _6962_/X sky130_fd_sc_hd__or4_1
XFILLER_53_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8701_ _8701_/A _8701_/B _8701_/C _8701_/D VGND VGND VPWR VPWR _8701_/X sky130_fd_sc_hd__or4_1
X_5913_ _5913_/A VGND VGND VPWR VPWR _5913_/X sky130_fd_sc_hd__clkbuf_1
X_6893_ _6890_/X _6892_/X _6887_/B VGND VGND VPWR VPWR _6905_/A sky130_fd_sc_hd__a21oi_1
X_8632_ _8965_/Q _8346_/X _8386_/A _8935_/Q VGND VGND VPWR VPWR _8632_/X sky130_fd_sc_hd__a22o_1
X_5844_ _5844_/A VGND VGND VPWR VPWR _5844_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_179_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8563_ _8563_/A _8563_/B _8563_/C _8563_/D VGND VGND VPWR VPWR _8576_/B sky130_fd_sc_hd__or4_1
X_5775_ _5775_/A VGND VGND VPWR VPWR _8968_/D sky130_fd_sc_hd__clkbuf_1
X_7514_ _7514_/A VGND VGND VPWR VPWR _7514_/X sky130_fd_sc_hd__clkbuf_4
X_4726_ input23/X _4460_/Y _4500_/Y input14/X _4725_/X VGND VGND VPWR VPWR _4731_/A
+ sky130_fd_sc_hd__a221o_1
X_8494_ _9228_/Q _8388_/X _8379_/X _9204_/Q _8493_/X VGND VGND VPWR VPWR _8499_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_181_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7445_ _7445_/A VGND VGND VPWR VPWR _9303_/D sky130_fd_sc_hd__clkbuf_1
X_4657_ _9212_/Q _7228_/A _5584_/A _8892_/Q VGND VGND VPWR VPWR _4657_/X sky130_fd_sc_hd__a22o_1
Xhold820 hold820/A VGND VGND VPWR VPWR hold820/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput80 spi_sck VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput91 spimemio_flash_io3_do VGND VGND VPWR VPWR input91/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7376_ _7376_/A VGND VGND VPWR VPWR _9272_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4588_ _9397_/Q _7640_/A _4436_/A input40/X VGND VGND VPWR VPWR _4588_/X sky130_fd_sc_hd__a22o_1
Xhold831 hold831/A VGND VGND VPWR VPWR hold831/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 _9472_/Q VGND VGND VPWR VPWR hold842/X sky130_fd_sc_hd__dlygate4sd3_1
X_9115_ _5235__1/A _9115_/D _7020_/X VGND VGND VPWR VPWR _9115_/Q sky130_fd_sc_hd__dfrtn_1
Xhold853 _9272_/Q VGND VGND VPWR VPWR hold853/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold864 _7089_/X VGND VGND VPWR VPWR _7090_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6327_ _6799_/A _6874_/A VGND VGND VPWR VPWR _6869_/D sky130_fd_sc_hd__nor2_1
Xhold875 hold875/A VGND VGND VPWR VPWR _7079_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold886 _5902_/X VGND VGND VPWR VPWR _5903_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold897 _5878_/X VGND VGND VPWR VPWR _9009_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9046_ _9541_/CLK _9046_/D VGND VGND VPWR VPWR _9046_/Q sky130_fd_sc_hd__dfxtp_1
X_6258_ _6262_/A _6562_/B VGND VGND VPWR VPWR _6338_/A sky130_fd_sc_hd__or2_1
XFILLER_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5209_ _9000_/Q _5071_/C _8797_/Q VGND VGND VPWR VPWR _5210_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6189_ _6556_/B _6558_/C VGND VGND VPWR VPWR _6190_/A sky130_fd_sc_hd__or2_1
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5560_ _5315_/X hold149/X _5560_/S VGND VGND VPWR VPWR _5560_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4511_ _4509_/X hold984/X _4964_/B VGND VGND VPWR VPWR _4512_/A sky130_fd_sc_hd__mux2_1
X_5491_ _5491_/A VGND VGND VPWR VPWR _8847_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7230_ _7230_/A VGND VGND VPWR VPWR _9208_/D sky130_fd_sc_hd__clkbuf_1
Xhold105 _5452_/Y VGND VGND VPWR VPWR _7158_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4442_ _4758_/A VGND VGND VPWR VPWR _7126_/A sky130_fd_sc_hd__buf_12
Xhold116 _7287_/X VGND VGND VPWR VPWR _7288_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold127 _9329_/Q VGND VGND VPWR VPWR hold127/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 _5484_/X VGND VGND VPWR VPWR _5485_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 _8877_/Q VGND VGND VPWR VPWR hold149/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7161_ _7161_/A VGND VGND VPWR VPWR _9176_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4373_ _4372_/X hold35/X hold74/X VGND VGND VPWR VPWR _4468_/B sky130_fd_sc_hd__mux2_4
XFILLER_125_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6112_ _6167_/B VGND VGND VPWR VPWR _6628_/A sky130_fd_sc_hd__clkbuf_4
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7092_ _5947_/X _9147_/Q _7106_/S VGND VGND VPWR VPWR _7092_/X sky130_fd_sc_hd__mux2_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ _6043_/A _7132_/B VGND VGND VPWR VPWR _6053_/S sky130_fd_sc_hd__and2_4
XFILLER_140_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7994_ _9344_/Q _8077_/A _7993_/X _9384_/Q VGND VGND VPWR VPWR _7994_/X sky130_fd_sc_hd__a22o_1
XFILLER_81_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6945_ _6881_/A _6736_/A _6748_/B _6449_/B VGND VGND VPWR VPWR _6945_/X sky130_fd_sc_hd__o22a_1
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_22_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6876_ _6906_/A _6876_/B VGND VGND VPWR VPWR _6956_/C sky130_fd_sc_hd__nor2_1
X_5827_ hold456/X _7645_/A _5842_/S VGND VGND VPWR VPWR _5827_/X sky130_fd_sc_hd__mux2_1
X_8615_ _8909_/Q _8360_/C _8411_/X _8924_/Q _8614_/X VGND VGND VPWR VPWR _8625_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_167_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5758_ _5758_/A VGND VGND VPWR VPWR _8961_/D sky130_fd_sc_hd__clkbuf_1
X_8546_ _9382_/Q _8337_/X _8384_/X _9198_/Q _8545_/X VGND VGND VPWR VPWR _8549_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_154_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4709_ _8941_/Q _5704_/A _5918_/A _9038_/Q VGND VGND VPWR VPWR _4709_/X sky130_fd_sc_hd__a22o_1
X_8477_ _8477_/A0 _8476_/X _8653_/S VGND VGND VPWR VPWR _8478_/A sky130_fd_sc_hd__mux2_1
X_5689_ _5689_/A VGND VGND VPWR VPWR _8931_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7428_ _7359_/X hold133/X _7444_/S VGND VGND VPWR VPWR _7429_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold650 _7813_/X VGND VGND VPWR VPWR _7814_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7359_ hold37/X VGND VGND VPWR VPWR _7359_/X sky130_fd_sc_hd__buf_2
Xhold661 _5913_/X VGND VGND VPWR VPWR _9022_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap380 _4445_/Y VGND VGND VPWR VPWR _7623_/A sky130_fd_sc_hd__buf_8
Xhold672 _8911_/Q VGND VGND VPWR VPWR hold672/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap391 _4437_/Y VGND VGND VPWR VPWR _7712_/A sky130_fd_sc_hd__buf_8
Xhold683 _9206_/Q VGND VGND VPWR VPWR hold683/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 _9287_/Q VGND VGND VPWR VPWR hold694/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9029_ _9551_/CLK _9029_/D fanout499/X VGND VGND VPWR VPWR _9029_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4991_ _4991_/A _4991_/B VGND VGND VPWR VPWR _4991_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_91_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6730_ _6744_/A _6742_/B VGND VGND VPWR VPWR _6730_/X sky130_fd_sc_hd__or2_1
XFILLER_189_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6661_ _6661_/A _6661_/B _6661_/C _6660_/Y VGND VGND VPWR VPWR _6661_/X sky130_fd_sc_hd__or4b_1
X_5612_ _5306_/X hold535/X _5616_/S VGND VGND VPWR VPWR _5612_/X sky130_fd_sc_hd__mux2_1
X_8400_ _9184_/Q _8400_/B VGND VGND VPWR VPWR _8400_/X sky130_fd_sc_hd__or2_1
XFILLER_149_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9380_ _9420_/CLK _9380_/D fanout464/X VGND VGND VPWR VPWR _9380_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_176_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6592_ _6873_/B _6799_/A VGND VGND VPWR VPWR _6726_/A sky130_fd_sc_hd__nor2_1
X_8331_ _8331_/A VGND VGND VPWR VPWR _8331_/X sky130_fd_sc_hd__buf_6
XFILLER_164_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5543_ _5301_/X hold532/X _5549_/S VGND VGND VPWR VPWR _5544_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8262_ _5139_/A _9517_/Q _8013_/X VGND VGND VPWR VPWR _8262_/X sky130_fd_sc_hd__a21o_1
XFILLER_144_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5474_ _7158_/A _5474_/B _7158_/C _7158_/D VGND VGND VPWR VPWR _5475_/A sky130_fd_sc_hd__or4_4
X_7213_ _7213_/A VGND VGND VPWR VPWR _9200_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4425_ hold42/X _4425_/B VGND VGND VPWR VPWR _4878_/A sky130_fd_sc_hd__nand2_8
X_8193_ _8193_/A _8193_/B _8193_/C _8193_/D VGND VGND VPWR VPWR _8193_/X sky130_fd_sc_hd__or4_2
XFILLER_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout404 fanout406/X VGND VGND VPWR VPWR fanout404/X sky130_fd_sc_hd__clkbuf_4
X_7144_ _7144_/A _7284_/B VGND VGND VPWR VPWR _7156_/S sky130_fd_sc_hd__nand2_8
X_4356_ hold74/A hold30/X hold57/X VGND VGND VPWR VPWR hold58/A sky130_fd_sc_hd__o21bai_1
XFILLER_59_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout415 fanout416/X VGND VGND VPWR VPWR fanout415/X sky130_fd_sc_hd__buf_2
XFILLER_99_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout426 fanout457/X VGND VGND VPWR VPWR fanout426/X sky130_fd_sc_hd__clkbuf_4
Xfanout437 fanout439/X VGND VGND VPWR VPWR fanout437/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout448 fanout449/X VGND VGND VPWR VPWR fanout448/X sky130_fd_sc_hd__buf_2
X_7075_ _5947_/X _9140_/Q _7075_/S VGND VGND VPWR VPWR _7075_/X sky130_fd_sc_hd__mux2_1
Xfanout459 fanout462/X VGND VGND VPWR VPWR fanout459/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6026_ hold651/X _5683_/X _6030_/S VGND VGND VPWR VPWR _6026_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7977_ _7977_/A VGND VGND VPWR VPWR _7977_/X sky130_fd_sc_hd__buf_6
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6928_ _6937_/A _6928_/B _6928_/C VGND VGND VPWR VPWR _6929_/C sky130_fd_sc_hd__and3b_1
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6859_ _6859_/A _6859_/B _6859_/C _6628_/X VGND VGND VPWR VPWR _6964_/C sky130_fd_sc_hd__or4b_2
XFILLER_168_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9578_ _9578_/A _5090_/Y VGND VGND VPWR VPWR mgmt_gpio_out[24] sky130_fd_sc_hd__ebufn_8
XFILLER_183_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8529_ _9470_/Q _8354_/A _8376_/A _9430_/Q VGND VGND VPWR VPWR _8529_/X sky130_fd_sc_hd__a22o_1
XFILLER_13_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold480 _5509_/X VGND VGND VPWR VPWR _5510_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 _8870_/Q VGND VGND VPWR VPWR hold491/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1180 _9094_/Q VGND VGND VPWR VPWR hold862/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1191 _9434_/Q VGND VGND VPWR VPWR hold737/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_320 _9157_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_331 _5218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_342 _5947_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_353 _7319_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_364 _8379_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_375 input69/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_386 fanout457/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_397 _6015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_3_0_mgmt_gpio_in[4] clkbuf_2_3_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _5207_/A1
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_146_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5190_ _9483_/Q VGND VGND VPWR VPWR _5190_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_95_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7900_ _7902_/B _8352_/A _8392_/A VGND VGND VPWR VPWR _7900_/X sky130_fd_sc_hd__and3_1
XFILLER_83_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8880_ _9051_/CLK _8880_/D fanout447/X VGND VGND VPWR VPWR _8880_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_64_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7831_ _7831_/A VGND VGND VPWR VPWR _9479_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4974_ _8808_/Q _8807_/Q _8806_/Q VGND VGND VPWR VPWR _4975_/A sky130_fd_sc_hd__and3_1
X_7762_ hold209/X _7514_/A _7762_/S VGND VGND VPWR VPWR _7762_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9501_ _9501_/CLK _9501_/D fanout470/X VGND VGND VPWR VPWR _9501_/Q sky130_fd_sc_hd__dfstp_2
X_6713_ hold98/A _6908_/A _6584_/X _6712_/X VGND VGND VPWR VPWR _9105_/D sky130_fd_sc_hd__o22a_1
X_7693_ _7514_/X hold586/X _7693_/S VGND VGND VPWR VPWR _7693_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9432_ _9434_/CLK _9432_/D fanout450/X VGND VGND VPWR VPWR _9432_/Q sky130_fd_sc_hd__dfstp_1
X_6644_ _6973_/B _6462_/B _6726_/B VGND VGND VPWR VPWR _6644_/X sky130_fd_sc_hd__a21o_1
XFILLER_192_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9363_ _9427_/CLK _9363_/D fanout481/X VGND VGND VPWR VPWR _9363_/Q sky130_fd_sc_hd__dfrtp_4
X_6575_ _6331_/Y _6551_/Y _7002_/C _6574_/Y VGND VGND VPWR VPWR _6576_/D sky130_fd_sc_hd__a211o_1
XFILLER_118_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5526_ _5526_/A VGND VGND VPWR VPWR _8861_/D sky130_fd_sc_hd__clkbuf_1
X_8314_ _8354_/B VGND VGND VPWR VPWR _8314_/X sky130_fd_sc_hd__buf_6
X_9294_ _9461_/CLK _9294_/D fanout422/X VGND VGND VPWR VPWR _9294_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_118_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8245_ _9072_/Q _7979_/X _8077_/X _8936_/Q _8244_/X VGND VGND VPWR VPWR _8250_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_105_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5457_ _5301_/X hold471/X _5472_/S VGND VGND VPWR VPWR _5457_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4408_ _4555_/A _4425_/B VGND VGND VPWR VPWR _4861_/A sky130_fd_sc_hd__nand2_8
X_8176_ _8963_/Q _7960_/A _8001_/A _8863_/Q _8175_/X VGND VGND VPWR VPWR _8184_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_182_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5388_ _5388_/A hold20/A VGND VGND VPWR VPWR _5389_/A sky130_fd_sc_hd__and2_1
XFILLER_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7127_ hold689/X _7113_/A _7139_/B _7126_/X VGND VGND VPWR VPWR _7127_/X sky130_fd_sc_hd__o211a_1
XFILLER_87_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7058_ _9132_/Q _5761_/X _7072_/S VGND VGND VPWR VPWR _7058_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6009_ _6009_/A VGND VGND VPWR VPWR _9074_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_150 _7927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_161 _7949_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_172 _7962_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_183 _7981_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_194 _8001_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4690_ _4690_/A _4690_/B _4690_/C _4690_/D VGND VGND VPWR VPWR _4690_/X sky130_fd_sc_hd__or4_2
XFILLER_186_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6360_ _6315_/Y _6839_/A _6553_/B _6959_/B _6359_/X VGND VGND VPWR VPWR _6360_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_127_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5311_ _7648_/A VGND VGND VPWR VPWR _5311_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_142_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6291_ _6402_/A _6498_/B _6589_/D _6778_/A _6290_/X VGND VGND VPWR VPWR _6291_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_142_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8030_ _9313_/Q _8008_/B _8077_/A _9345_/Q _7984_/X VGND VGND VPWR VPWR _8030_/X
+ sky130_fd_sc_hd__a221o_1
X_5242_ _9235_/Q VGND VGND VPWR VPWR _5242_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_30_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _9427_/CLK sky130_fd_sc_hd__clkbuf_16
X_5173_ _5173_/A VGND VGND VPWR VPWR _5173_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput1 debug_mode VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__dlymetal6s2s_1
X_8932_ _9484_/CLK _8932_/D fanout432/X VGND VGND VPWR VPWR _8932_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_45_csclk _8954_/CLK VGND VGND VPWR VPWR _9291_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8863_ _9466_/CLK _8863_/D fanout471/X VGND VGND VPWR VPWR _8863_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7814_ _7814_/A VGND VGND VPWR VPWR _9471_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8794_ _5168_/A1 _8794_/D _5354_/X VGND VGND VPWR VPWR _8794_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7745_ _7745_/A VGND VGND VPWR VPWR _9439_/D sky130_fd_sc_hd__clkbuf_1
X_4957_ _8908_/Q _5630_/A _7074_/A _9140_/Q VGND VGND VPWR VPWR _4957_/X sky130_fd_sc_hd__a22o_1
XFILLER_101_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4888_ _4888_/A VGND VGND VPWR VPWR _9112_/D sky130_fd_sc_hd__clkbuf_1
X_7676_ _7514_/X hold603/X _7676_/S VGND VGND VPWR VPWR _7676_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9415_ _9461_/CLK _9415_/D fanout424/X VGND VGND VPWR VPWR _9415_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6627_ _6627_/A _6924_/C _6627_/C _6627_/D VGND VGND VPWR VPWR _6629_/C sky130_fd_sc_hd__or4_1
XFILLER_192_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9346_ _9370_/CLK _9346_/D fanout477/X VGND VGND VPWR VPWR _9346_/Q sky130_fd_sc_hd__dfrtp_4
X_6558_ _6790_/A _6558_/B _6558_/C VGND VGND VPWR VPWR _6559_/A sky130_fd_sc_hd__or3_1
XFILLER_180_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5509_ hold479/X _5392_/X _5515_/S VGND VGND VPWR VPWR _5509_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9277_ _9413_/CLK _9277_/D fanout458/X VGND VGND VPWR VPWR _9277_/Q sky130_fd_sc_hd__dfrtp_1
X_6489_ _6489_/A VGND VGND VPWR VPWR _6862_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_145_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8228_ _8228_/A _8228_/B _8228_/C _8228_/D VGND VGND VPWR VPWR _8228_/X sky130_fd_sc_hd__or4_1
XFILLER_106_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8159_ _9319_/Q _8275_/B VGND VGND VPWR VPWR _8159_/X sky130_fd_sc_hd__or2_1
XFILLER_87_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5860_ _5860_/A VGND VGND VPWR VPWR _9004_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4811_ _4811_/A VGND VGND VPWR VPWR _5897_/S sky130_fd_sc_hd__buf_8
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5791_ hold712/X _5687_/X _5793_/S VGND VGND VPWR VPWR _5792_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4742_ _8946_/Q _5715_/A _5642_/A _8916_/Q VGND VGND VPWR VPWR _4742_/X sky130_fd_sc_hd__a22o_1
X_7530_ _7439_/X hold238/X _7534_/S VGND VGND VPWR VPWR _7530_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7461_ _7299_/X hold520/X _7461_/S VGND VGND VPWR VPWR _7461_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4673_ _4673_/A _4673_/B _4673_/C _4673_/D VGND VGND VPWR VPWR _4689_/C sky130_fd_sc_hd__or4_2
X_9200_ _9461_/CLK _9200_/D fanout422/X VGND VGND VPWR VPWR _9200_/Q sky130_fd_sc_hd__dfstp_1
X_6412_ _6850_/B _6416_/A VGND VGND VPWR VPWR _6413_/B sky130_fd_sc_hd__nor2_2
X_7392_ _7302_/X hold938/X _7406_/S VGND VGND VPWR VPWR _7393_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9131_ _9487_/CLK _9131_/D fanout411/X VGND VGND VPWR VPWR _9131_/Q sky130_fd_sc_hd__dfrtp_1
X_6343_ _6507_/A _6510_/A _6343_/C VGND VGND VPWR VPWR _6560_/A sky130_fd_sc_hd__and3_1
XFILLER_127_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9062_ _9110_/CLK _9062_/D VGND VGND VPWR VPWR _9062_/Q sky130_fd_sc_hd__dfxtp_1
X_6274_ _6736_/A _6799_/A VGND VGND VPWR VPWR _6274_/X sky130_fd_sc_hd__or2_1
XFILLER_143_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8013_ _8013_/A VGND VGND VPWR VPWR _8013_/X sky130_fd_sc_hd__buf_2
X_5225_ _5225_/A VGND VGND VPWR VPWR _9569_/A sky130_fd_sc_hd__buf_1
XFILLER_130_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5156_ _9163_/Q _7902_/A _5155_/X VGND VGND VPWR VPWR _8996_/D sky130_fd_sc_hd__o21ai_1
XFILLER_69_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5087_ _9403_/Q VGND VGND VPWR VPWR _5087_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8915_ _9172_/CLK _8915_/D fanout492/X VGND VGND VPWR VPWR _8915_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_71_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8846_ _9172_/CLK _8846_/D fanout493/X VGND VGND VPWR VPWR _8846_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8777_ _5235__1/A _8777_/D _5319_/X VGND VGND VPWR VPWR hold17/A sky130_fd_sc_hd__dfrtn_1
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5989_ _5989_/A VGND VGND VPWR VPWR _9065_/D sky130_fd_sc_hd__buf_1
XFILLER_169_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7728_ _7728_/A VGND VGND VPWR VPWR _9431_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_50 _4852_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_61 _5067_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7659_ _7514_/X hold657/X hold84/X VGND VGND VPWR VPWR _7660_/A sky130_fd_sc_hd__mux2_1
XANTENNA_72 hold19/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_83 _5392_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_94 _5629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9329_ _9459_/CLK _9329_/D fanout479/X VGND VGND VPWR VPWR _9329_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold309 hold309/A VGND VGND VPWR VPWR hold309/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A VGND VGND VPWR VPWR _9110_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_97_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _5010_/A _5014_/S VGND VGND VPWR VPWR _5011_/B sky130_fd_sc_hd__nor2_1
XFILLER_39_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1009 _5128_/X VGND VGND VPWR VPWR _8827_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6961_ _6563_/A _6873_/Y _6874_/Y _6563_/B _6960_/X VGND VGND VPWR VPWR _7003_/C
+ sky130_fd_sc_hd__a221o_1
X_8700_ _8700_/A _8700_/B _8700_/C _8700_/D VGND VGND VPWR VPWR _8701_/D sky130_fd_sc_hd__or4_1
X_5912_ _5465_/X _9583_/A _5916_/S VGND VGND VPWR VPWR _5912_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6892_ _6891_/X _6781_/B _6967_/C _6967_/B VGND VGND VPWR VPWR _6892_/X sky130_fd_sc_hd__a31o_1
XFILLER_22_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8631_ _8960_/Q _8402_/X _8378_/X _8945_/Q _8630_/X VGND VGND VPWR VPWR _8631_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5843_ _9577_/A hold6/X hold43/X VGND VGND VPWR VPWR _5843_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8562_ _9319_/Q _8372_/X _8369_/X _9327_/Q _8561_/X VGND VGND VPWR VPWR _8563_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5774_ _5629_/X hold880/X _5782_/S VGND VGND VPWR VPWR _5775_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7513_ _7513_/A VGND VGND VPWR VPWR _9334_/D sky130_fd_sc_hd__clkbuf_1
X_4725_ _9403_/Q _7661_/A _5773_/A _8971_/Q VGND VGND VPWR VPWR _4725_/X sky130_fd_sc_hd__a22o_2
X_8493_ _9388_/Q _8292_/X _8294_/X _9292_/Q VGND VGND VPWR VPWR _8493_/X sky130_fd_sc_hd__a22o_1
XFILLER_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4656_ _4656_/A _5453_/B VGND VGND VPWR VPWR _5584_/A sky130_fd_sc_hd__nor2_4
XFILLER_107_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7444_ _7299_/X hold848/X _7444_/S VGND VGND VPWR VPWR _7445_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput70 mgmt_gpio_in[7] VGND VGND VPWR VPWR _5283_/B sky130_fd_sc_hd__buf_2
XFILLER_162_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold810 _7030_/X VGND VGND VPWR VPWR _7031_/A sky130_fd_sc_hd__dlygate4sd3_1
Xinput81 spi_sdo VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold821 _8838_/Q VGND VGND VPWR VPWR hold821/X sky130_fd_sc_hd__dlygate4sd3_1
X_7375_ _7302_/X hold853/X _7389_/S VGND VGND VPWR VPWR _7376_/A sky130_fd_sc_hd__mux2_1
X_4587_ _9469_/Q _7798_/A _7519_/A _9341_/Q _4586_/X VGND VGND VPWR VPWR _4590_/C
+ sky130_fd_sc_hd__a221o_1
Xinput92 spimemio_flash_io3_oeb VGND VGND VPWR VPWR input92/X sky130_fd_sc_hd__clkbuf_2
Xhold832 _9262_/Q VGND VGND VPWR VPWR hold832/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold843 _9074_/Q VGND VGND VPWR VPWR hold843/X sky130_fd_sc_hd__dlygate4sd3_1
X_9114_ _5235__1/A _9114_/D _7018_/X VGND VGND VPWR VPWR _9114_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_89_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold854 _7028_/X VGND VGND VPWR VPWR _7029_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6326_ _6666_/B VGND VGND VPWR VPWR _6874_/A sky130_fd_sc_hd__buf_4
Xhold865 hold865/A VGND VGND VPWR VPWR hold865/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold876 _9304_/Q VGND VGND VPWR VPWR hold876/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 _9384_/Q VGND VGND VPWR VPWR hold887/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold898 hold898/A VGND VGND VPWR VPWR hold898/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6257_ _6257_/A _6257_/B _6257_/C _6256_/X VGND VGND VPWR VPWR _6268_/A sky130_fd_sc_hd__or4b_1
X_9045_ _9541_/CLK _9045_/D VGND VGND VPWR VPWR _9045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5208_ _5208_/A VGND VGND VPWR VPWR _9563_/A sky130_fd_sc_hd__buf_1
XFILLER_190_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6188_ _6344_/B _6344_/A VGND VGND VPWR VPWR _6558_/C sky130_fd_sc_hd__nand2b_2
XFILLER_69_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5139_ _5139_/A _5160_/B VGND VGND VPWR VPWR _5139_/Y sky130_fd_sc_hd__nand2_1
XFILLER_123_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8829_ _8831_/CLK _8829_/D _5447_/X VGND VGND VPWR VPWR _8829_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_12_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4510_ _8791_/Q _8829_/Q VGND VGND VPWR VPWR _4964_/B sky130_fd_sc_hd__nand2_4
XFILLER_117_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5490_ _5471_/X hold469/X _5490_/S VGND VGND VPWR VPWR _5490_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4441_ input42/X _5867_/S _7712_/A _9431_/Q _4440_/X VGND VGND VPWR VPWR _4506_/A
+ sky130_fd_sc_hd__a221o_1
Xhold106 _7168_/X VGND VGND VPWR VPWR _7169_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 _9444_/Q VGND VGND VPWR VPWR hold117/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold128 _7502_/X VGND VGND VPWR VPWR _7503_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 _9078_/Q VGND VGND VPWR VPWR hold139/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7160_ _7128_/X hold814/X _7174_/S VGND VGND VPWR VPWR _7160_/X sky130_fd_sc_hd__mux2_1
X_4372_ hold77/X _5012_/A hold22/X VGND VGND VPWR VPWR _4372_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6111_ _6437_/A _6716_/A _6416_/A VGND VGND VPWR VPWR _6906_/B sky130_fd_sc_hd__or3_4
XFILLER_98_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7091_ _7091_/A _7284_/B VGND VGND VPWR VPWR _7106_/S sky130_fd_sc_hd__nand2_4
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6042_ _6042_/A VGND VGND VPWR VPWR _9088_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7993_ _7993_/A VGND VGND VPWR VPWR _7993_/X sky130_fd_sc_hd__buf_8
XFILLER_54_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6944_ _6944_/A _6944_/B _6944_/C _6943_/X VGND VGND VPWR VPWR _6994_/B sky130_fd_sc_hd__or4b_2
XFILLER_50_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6875_ _6345_/X _6873_/Y _6874_/Y _6563_/A VGND VGND VPWR VPWR _6937_/C sky130_fd_sc_hd__a22o_1
XFILLER_34_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8614_ _8929_/Q _8301_/A _8356_/C _8894_/Q _8613_/X VGND VGND VPWR VPWR _8614_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5826_ _5826_/A VGND VGND VPWR VPWR _5826_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8545_ _9438_/Q _7908_/X _8335_/X _9278_/Q VGND VGND VPWR VPWR _8545_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5757_ hold413/X _5687_/X _5759_/S VGND VGND VPWR VPWR _5758_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4708_ _8936_/Q _5693_/A _5596_/A _8896_/Q _4707_/X VGND VGND VPWR VPWR _4711_/C
+ sky130_fd_sc_hd__a221o_1
X_8476_ _9522_/Q _8475_/X _8627_/S VGND VGND VPWR VPWR _8476_/X sky130_fd_sc_hd__mux2_1
X_5688_ hold405/X _5687_/X _5691_/S VGND VGND VPWR VPWR _5689_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7427_ _7427_/A VGND VGND VPWR VPWR _9296_/D sky130_fd_sc_hd__clkbuf_1
X_4639_ _9244_/Q _4449_/Y _7781_/A _9460_/Q _4638_/X VGND VGND VPWR VPWR _4649_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_150_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold640 _7170_/X VGND VGND VPWR VPWR _7171_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold651 _9081_/Q VGND VGND VPWR VPWR hold651/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7358_ _7358_/A VGND VGND VPWR VPWR _9264_/D sky130_fd_sc_hd__clkbuf_1
Xhold662 hold662/A VGND VGND VPWR VPWR hold662/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap370 _4585_/Y VGND VGND VPWR VPWR _7144_/A sky130_fd_sc_hd__buf_8
XFILLER_116_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap381 _4438_/Y VGND VGND VPWR VPWR _7678_/A sky130_fd_sc_hd__buf_8
XFILLER_150_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold673 _5638_/X VGND VGND VPWR VPWR _5639_/A sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap392 _4389_/Y VGND VGND VPWR VPWR _7640_/A sky130_fd_sc_hd__buf_8
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold684 _7224_/X VGND VGND VPWR VPWR _7225_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6309_ _6309_/A _6558_/C VGND VGND VPWR VPWR _6314_/C sky130_fd_sc_hd__nor2_1
XFILLER_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold695 _7406_/X VGND VGND VPWR VPWR _7407_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7289_ _7233_/X hold769/X _7300_/S VGND VGND VPWR VPWR _7289_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9028_ _9551_/CLK _9028_/D fanout499/X VGND VGND VPWR VPWR _9028_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_89_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xnet499_2 _5207_/A1 VGND VGND VPWR VPWR _5236_/B sky130_fd_sc_hd__inv_2
X_4990_ _5040_/B _4997_/B hold80/A VGND VGND VPWR VPWR _4991_/B sky130_fd_sc_hd__o21a_1
XFILLER_51_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6660_ _6660_/A _6660_/B VGND VGND VPWR VPWR _6660_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5611_ _5611_/A VGND VGND VPWR VPWR _8899_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6591_ _6591_/A _6591_/B VGND VGND VPWR VPWR _6966_/C sky130_fd_sc_hd__nand2_1
X_8330_ _8392_/A _8398_/A _8357_/B VGND VGND VPWR VPWR _8331_/A sky130_fd_sc_hd__and3_2
X_5542_ _5542_/A VGND VGND VPWR VPWR _8868_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8261_ _8851_/Q _8010_/B _8250_/X _8260_/X _8105_/X VGND VGND VPWR VPWR _8261_/X
+ sky130_fd_sc_hd__o221a_1
X_5473_ _5473_/A VGND VGND VPWR VPWR _8839_/D sky130_fd_sc_hd__clkbuf_1
X_4424_ _4861_/A _4492_/B VGND VGND VPWR VPWR _4424_/Y sky130_fd_sc_hd__nor2_2
X_7212_ _7128_/X hold911/X _7226_/S VGND VGND VPWR VPWR _7213_/A sky130_fd_sc_hd__mux2_1
XFILLER_132_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8192_ _8943_/Q _8020_/X _7990_/X _8868_/Q _8191_/X VGND VGND VPWR VPWR _8193_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_99_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7143_ _7143_/A VGND VGND VPWR VPWR _9169_/D sky130_fd_sc_hd__clkbuf_1
X_4355_ hold29/X hold73/A hold56/X _4354_/X VGND VGND VPWR VPWR hold57/A sky130_fd_sc_hd__o31a_1
Xfanout405 fanout406/X VGND VGND VPWR VPWR fanout405/X sky130_fd_sc_hd__clkbuf_2
XFILLER_113_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout416 fanout457/X VGND VGND VPWR VPWR fanout416/X sky130_fd_sc_hd__clkbuf_4
Xfanout427 fanout429/X VGND VGND VPWR VPWR fanout427/X sky130_fd_sc_hd__clkbuf_4
XFILLER_59_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout438 fanout439/X VGND VGND VPWR VPWR fanout438/X sky130_fd_sc_hd__clkbuf_4
X_7074_ _7074_/A _7139_/B VGND VGND VPWR VPWR _7075_/S sky130_fd_sc_hd__nand2_1
Xfanout449 fanout457/X VGND VGND VPWR VPWR fanout449/X sky130_fd_sc_hd__buf_2
XFILLER_58_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6025_ _6025_/A VGND VGND VPWR VPWR _9080_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7976_ _9496_/Q _8000_/B _8002_/B VGND VGND VPWR VPWR _7977_/A sky130_fd_sc_hd__and3_2
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6927_ _6881_/A _6764_/A _6435_/A _6449_/B VGND VGND VPWR VPWR _6928_/C sky130_fd_sc_hd__o22a_1
XFILLER_23_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6858_ _6895_/A _6858_/B VGND VGND VPWR VPWR _6859_/A sky130_fd_sc_hd__nor2_1
X_5809_ _5951_/A VGND VGND VPWR VPWR _5809_/X sky130_fd_sc_hd__buf_6
X_9577_ _9577_/A _5091_/Y VGND VGND VPWR VPWR mgmt_gpio_out[23] sky130_fd_sc_hd__ebufn_8
X_6789_ _6939_/C _6939_/D VGND VGND VPWR VPWR _6807_/A sky130_fd_sc_hd__nand2_1
XFILLER_182_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8528_ hold983/X _8196_/S _8526_/X _8527_/X VGND VGND VPWR VPWR _9525_/D sky130_fd_sc_hd__o22a_1
XFILLER_182_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8459_ _9299_/Q _8314_/X _8331_/X _9403_/Q VGND VGND VPWR VPWR _8459_/X sky130_fd_sc_hd__a22o_1
XFILLER_123_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold470 _5490_/X VGND VGND VPWR VPWR _5491_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold481 _5916_/X VGND VGND VPWR VPWR _5917_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold492 _5545_/X VGND VGND VPWR VPWR _5546_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1170 _7118_/X VGND VGND VPWR VPWR hold591/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1181 _9188_/Q VGND VGND VPWR VPWR hold345/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1192 _8899_/Q VGND VGND VPWR VPWR hold494/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_310 _9503_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_321 _9162_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_332 _5291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_343 _5979_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_354 _7479_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_365 _8384_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_376 _5071_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_387 hold27/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_398 _6018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7830_ _5415_/X hold703/X _7830_/S VGND VGND VPWR VPWR _7830_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7761_ _7761_/A VGND VGND VPWR VPWR _9446_/D sky130_fd_sc_hd__clkbuf_1
X_4973_ _8827_/Q VGND VGND VPWR VPWR _5021_/A sky130_fd_sc_hd__clkinv_2
X_9500_ _9501_/CLK _9500_/D fanout470/X VGND VGND VPWR VPWR _9500_/Q sky130_fd_sc_hd__dfrtp_2
X_6712_ _6292_/X _6629_/X _6663_/X _8735_/A _6711_/X VGND VGND VPWR VPWR _6712_/X
+ sky130_fd_sc_hd__a2111o_1
X_7692_ _7692_/A VGND VGND VPWR VPWR _9414_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9431_ _9471_/CLK _9431_/D fanout421/X VGND VGND VPWR VPWR _9431_/Q sky130_fd_sc_hd__dfrtp_1
X_6643_ _6643_/A _6643_/B VGND VGND VPWR VPWR _6997_/A sky130_fd_sc_hd__or2_1
X_9362_ _9370_/CLK _9362_/D fanout477/X VGND VGND VPWR VPWR _9362_/Q sky130_fd_sc_hd__dfrtp_4
X_6574_ _7001_/A _6574_/B VGND VGND VPWR VPWR _6574_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8313_ _8375_/A _8389_/A _8357_/A VGND VGND VPWR VPWR _8354_/B sky130_fd_sc_hd__and3_4
X_5525_ _5311_/X hold400/X _5527_/S VGND VGND VPWR VPWR _5525_/X sky130_fd_sc_hd__mux2_1
X_9293_ _9413_/CLK _9293_/D fanout458/X VGND VGND VPWR VPWR _9293_/Q sky130_fd_sc_hd__dfrtp_1
X_8244_ _9082_/Q _7949_/X _8001_/X _8866_/Q VGND VGND VPWR VPWR _8244_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5456_ _5456_/A VGND VGND VPWR VPWR _8832_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4407_ hold60/X _4492_/A VGND VGND VPWR VPWR _4407_/Y sky130_fd_sc_hd__nor2_1
X_8175_ _8973_/Q _7947_/A _7981_/A _8913_/Q VGND VGND VPWR VPWR _8175_/X sky130_fd_sc_hd__a22o_1
X_5387_ _7517_/A VGND VGND VPWR VPWR _5387_/X sky130_fd_sc_hd__buf_6
XFILLER_99_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7126_ _7126_/A _7126_/B _7126_/C VGND VGND VPWR VPWR _7126_/X sky130_fd_sc_hd__or3_1
XFILLER_59_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7057_ _7057_/A VGND VGND VPWR VPWR _7072_/S sky130_fd_sc_hd__clkbuf_4
X_6008_ _5947_/X hold843/X _6019_/S VGND VGND VPWR VPWR _6008_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7959_ _7998_/A _7989_/B _7996_/B VGND VGND VPWR VPWR _7960_/A sky130_fd_sc_hd__and3_4
XFILLER_187_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_140 _7908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_151 _8000_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_162 _7949_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_173 _7962_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_184 _7990_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9503__504 VGND VGND VPWR VPWR _9503_/D _9503__504/LO sky130_fd_sc_hd__conb_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_195 _8001_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5310_ hold45/X VGND VGND VPWR VPWR _7648_/A sky130_fd_sc_hd__buf_4
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6290_ _6546_/A _6290_/B _6290_/C _6289_/Y VGND VGND VPWR VPWR _6290_/X sky130_fd_sc_hd__or4b_1
XFILLER_170_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5241_ _9227_/Q VGND VGND VPWR VPWR _5241_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5172_ _5172_/A VGND VGND VPWR VPWR _5173_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8931_ _9184_/CLK _8931_/D fanout438/X VGND VGND VPWR VPWR _8931_/Q sky130_fd_sc_hd__dfrtp_1
Xinput2 debug_oeb VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_opt_1_0_csclk _9210_/CLK VGND VGND VPWR VPWR clkbuf_opt_1_0_csclk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8862_ _9069_/CLK _8862_/D fanout433/X VGND VGND VPWR VPWR _8862_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_52_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7813_ _5415_/X hold649/X _7813_/S VGND VGND VPWR VPWR _7813_/X sky130_fd_sc_hd__mux2_1
X_8793_ _8831_/CLK _8793_/D _5352_/X VGND VGND VPWR VPWR _8793_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_52_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7744_ _5415_/X hold790/X hold86/X VGND VGND VPWR VPWR _7744_/X sky130_fd_sc_hd__mux2_1
X_4956_ _4956_/A _7111_/B VGND VGND VPWR VPWR _7074_/A sky130_fd_sc_hd__nor2_1
XFILLER_51_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7675_ _7675_/A VGND VGND VPWR VPWR _9406_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4887_ _4886_/X hold980/X _4964_/B VGND VGND VPWR VPWR _4888_/A sky130_fd_sc_hd__mux2_1
X_9414_ _9471_/CLK _9414_/D fanout421/X VGND VGND VPWR VPWR _9414_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_137_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6626_ _6950_/A _6626_/B _6626_/C _6626_/D VGND VGND VPWR VPWR _6627_/D sky130_fd_sc_hd__or4_1
XFILLER_165_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9345_ _9449_/CLK _9345_/D fanout479/X VGND VGND VPWR VPWR _9345_/Q sky130_fd_sc_hd__dfstp_2
X_6557_ _6227_/Y _6510_/Y _6232_/B VGND VGND VPWR VPWR _6822_/A sky130_fd_sc_hd__a21oi_1
X_5508_ _5508_/A VGND VGND VPWR VPWR _8853_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9276_ _9276_/CLK _9276_/D fanout462/X VGND VGND VPWR VPWR _9276_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6488_ _6748_/B _6887_/B VGND VGND VPWR VPWR _6489_/A sky130_fd_sc_hd__or2_1
X_8227_ _9037_/Q _7938_/X _7997_/X _8955_/Q _8226_/X VGND VGND VPWR VPWR _8228_/D
+ sky130_fd_sc_hd__a221o_1
X_5439_ _5439_/A VGND VGND VPWR VPWR _8825_/D sky130_fd_sc_hd__clkbuf_1
Xoutput350 _9540_/Q VGND VGND VPWR VPWR wb_dat_o[30] sky130_fd_sc_hd__buf_12
XFILLER_121_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8158_ _9215_/Q _7923_/X _7997_/X _9367_/Q _8157_/X VGND VGND VPWR VPWR _8162_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7109_ _5947_/X _9155_/Q _7109_/S VGND VGND VPWR VPWR _7109_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8089_ _9372_/Q _7960_/X _8001_/X _9268_/Q _8088_/X VGND VGND VPWR VPWR _8097_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4810_ _8811_/Q _5388_/A _7194_/A _9194_/Q _4809_/X VGND VGND VPWR VPWR _4816_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5790_ _5790_/A VGND VGND VPWR VPWR _8975_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4741_ _4741_/A _4741_/B _4741_/C _4741_/D VGND VGND VPWR VPWR _4752_/C sky130_fd_sc_hd__or4_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7460_ _7460_/A VGND VGND VPWR VPWR _9310_/D sky130_fd_sc_hd__clkbuf_1
X_4672_ input96/X _4488_/Y _4414_/Y _9340_/Q _4671_/X VGND VGND VPWR VPWR _4673_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_147_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6411_ _6597_/B VGND VGND VPWR VPWR _6503_/A sky130_fd_sc_hd__clkbuf_4
X_7391_ _7391_/A _7499_/B VGND VGND VPWR VPWR _7406_/S sky130_fd_sc_hd__nand2_4
XFILLER_162_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9130_ _9487_/CLK _9130_/D fanout411/X VGND VGND VPWR VPWR _9130_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_162_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6342_ _6603_/A _6764_/A VGND VGND VPWR VPWR _6352_/A sky130_fd_sc_hd__nor2_1
XFILLER_127_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9061_ _9110_/CLK _9061_/D VGND VGND VPWR VPWR _9061_/Q sky130_fd_sc_hd__dfxtp_1
X_6273_ _6279_/A VGND VGND VPWR VPWR _6736_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8012_ _8012_/A VGND VGND VPWR VPWR _8013_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_88_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5224_ _9007_/Q user_clock _9166_/Q VGND VGND VPWR VPWR _5225_/A sky130_fd_sc_hd__mux2_2
XFILLER_142_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5155_ _7916_/C _5155_/B VGND VGND VPWR VPWR _5155_/X sky130_fd_sc_hd__or2_1
XFILLER_96_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5086_ _9411_/Q VGND VGND VPWR VPWR _5086_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8914_ _9172_/CLK _8914_/D fanout492/X VGND VGND VPWR VPWR _8914_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_37_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8845_ _9172_/CLK _8845_/D fanout489/X VGND VGND VPWR VPWR _8845_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8776_ _9484_/CLK _8776_/D fanout430/X VGND VGND VPWR VPWR _8776_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5988_ _9065_/Q _5988_/A1 _5994_/S VGND VGND VPWR VPWR _5989_/A sky130_fd_sc_hd__mux2_2
X_7727_ _5415_/X hold655/X hold95/X VGND VGND VPWR VPWR _7727_/X sky130_fd_sc_hd__mux2_1
X_4939_ _4939_/A _4939_/B _4939_/C _4939_/D VGND VGND VPWR VPWR _4961_/B sky130_fd_sc_hd__or4_1
XANTENNA_40 _5630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7658_ _7658_/A VGND VGND VPWR VPWR _9398_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_51 _4884_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_62 _5067_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 hold19/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_84 _5395_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6609_ _6609_/A _6609_/B VGND VGND VPWR VPWR _6609_/Y sky130_fd_sc_hd__nand2_1
XFILLER_192_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_95 _5629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7589_ _7517_/X hold931/X hold75/X VGND VGND VPWR VPWR _7590_/A sky130_fd_sc_hd__mux2_1
X_9328_ _9328_/CLK _9328_/D fanout463/X VGND VGND VPWR VPWR _9328_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_4_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9259_ _9483_/CLK _9259_/D fanout473/X VGND VGND VPWR VPWR _9259_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_161_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_59_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _9087_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6960_ _6960_/A _6960_/B _6879_/X VGND VGND VPWR VPWR _6960_/X sky130_fd_sc_hd__or3b_1
XFILLER_81_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5911_ _5911_/A VGND VGND VPWR VPWR _5911_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_46_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6891_ _6891_/A _6891_/B VGND VGND VPWR VPWR _6891_/X sky130_fd_sc_hd__or2_1
XFILLER_179_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8630_ _8900_/Q _8312_/X _8376_/X _8950_/Q VGND VGND VPWR VPWR _8630_/X sky130_fd_sc_hd__a22o_1
X_5842_ _8839_/Q hold5/X _5842_/S VGND VGND VPWR VPWR hold6/A sky130_fd_sc_hd__mux2_1
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8561_ _9303_/Q _8314_/X _8331_/X _9407_/Q VGND VGND VPWR VPWR _8561_/X sky130_fd_sc_hd__a22o_1
X_5773_ _5773_/A _7043_/B VGND VGND VPWR VPWR _5782_/S sky130_fd_sc_hd__nand2_4
X_7512_ _7494_/X hold772/X _7515_/S VGND VGND VPWR VPWR _7512_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4724_ _4724_/A _4724_/B _4724_/C _4724_/D VGND VGND VPWR VPWR _4752_/A sky130_fd_sc_hd__or4_1
XFILLER_187_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8492_ _9236_/Q _8322_/X _8333_/X _9268_/Q _8491_/X VGND VGND VPWR VPWR _8499_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_147_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7443_ _7443_/A VGND VGND VPWR VPWR _9302_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4655_ _9196_/Q _7194_/A _4531_/Y _4650_/Y _4654_/X VGND VGND VPWR VPWR _4689_/B
+ sky130_fd_sc_hd__a2111o_1
Xinput60 mgmt_gpio_in[31] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__buf_4
Xhold800 _9194_/Q VGND VGND VPWR VPWR hold800/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput71 mgmt_gpio_in[8] VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold811 _8955_/Q VGND VGND VPWR VPWR hold811/X sky130_fd_sc_hd__dlygate4sd3_1
X_7374_ _7374_/A _7499_/B VGND VGND VPWR VPWR _7389_/S sky130_fd_sc_hd__nand2_8
Xinput82 spi_sdoenb VGND VGND VPWR VPWR input82/X sky130_fd_sc_hd__clkbuf_1
X_4586_ _9349_/Q _7536_/A _7144_/A _9555_/A VGND VGND VPWR VPWR _4586_/X sky130_fd_sc_hd__a22o_1
Xhold822 _5469_/X VGND VGND VPWR VPWR _5470_/A sky130_fd_sc_hd__dlygate4sd3_1
Xinput93 sram_ro_data[0] VGND VGND VPWR VPWR input93/X sky130_fd_sc_hd__clkbuf_2
X_9113_ _5235__1/A _9113_/D _7016_/X VGND VGND VPWR VPWR _9113_/Q sky130_fd_sc_hd__dfrtn_1
Xhold833 _7352_/X VGND VGND VPWR VPWR _7353_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 _6008_/X VGND VGND VPWR VPWR _6009_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6325_ _6325_/A VGND VGND VPWR VPWR _6666_/B sky130_fd_sc_hd__buf_2
Xhold855 _9048_/Q VGND VGND VPWR VPWR hold855/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold866 hold866/A VGND VGND VPWR VPWR hold866/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold877 hold877/A VGND VGND VPWR VPWR _5848_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 _9424_/Q VGND VGND VPWR VPWR hold888/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9044_ _9541_/CLK _9044_/D VGND VGND VPWR VPWR _9044_/Q sky130_fd_sc_hd__dfxtp_1
X_6256_ _6603_/A _6266_/A _6279_/A _6881_/A _6255_/X VGND VGND VPWR VPWR _6256_/X
+ sky130_fd_sc_hd__o221a_1
Xhold899 hold899/A VGND VGND VPWR VPWR hold899/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5207_ _9001_/Q _5207_/A1 _8796_/Q VGND VGND VPWR VPWR _5208_/A sky130_fd_sc_hd__mux2_2
X_6187_ _6317_/B _6187_/B VGND VGND VPWR VPWR _6344_/A sky130_fd_sc_hd__or2_2
XFILLER_191_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5138_ _5139_/A _5135_/X _5160_/B _9163_/Q _8996_/Q VGND VGND VPWR VPWR _8998_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_96_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5069_ _5035_/B _5068_/B _5067_/X _5068_/Y hold999/X VGND VGND VPWR VPWR _8780_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8828_ _8831_/CLK _8828_/D _5445_/X VGND VGND VPWR VPWR _8828_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8759_ _9032_/Q _8759_/A2 _8759_/B1 _5275_/A VGND VGND VPWR VPWR _8759_/X sky130_fd_sc_hd__a22o_1
XFILLER_40_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4440_ _9415_/Q _7678_/A _7695_/A _9423_/Q VGND VGND VPWR VPWR _4440_/X sky130_fd_sc_hd__a22o_1
Xhold107 _7169_/X VGND VGND VPWR VPWR _9180_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold118 _7756_/X VGND VGND VPWR VPWR _7757_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 _8972_/Q VGND VGND VPWR VPWR hold129/X sky130_fd_sc_hd__dlygate4sd3_1
X_4371_ hold9/X hold98/X hold74/A VGND VGND VPWR VPWR hold10/A sky130_fd_sc_hd__mux2_4
XFILLER_125_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6110_ _6181_/A _6721_/A VGND VGND VPWR VPWR _6416_/A sky130_fd_sc_hd__or2_4
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7090_ _7090_/A VGND VGND VPWR VPWR _9146_/D sky130_fd_sc_hd__clkbuf_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6041_ hold498/X _5690_/X _6041_/S VGND VGND VPWR VPWR _6042_/A sky130_fd_sc_hd__mux2_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7992_ _7998_/A _8000_/B _7992_/C VGND VGND VPWR VPWR _7993_/A sky130_fd_sc_hd__and3_4
X_6943_ _6850_/B _6416_/A _6862_/B _6274_/X VGND VGND VPWR VPWR _6943_/X sky130_fd_sc_hd__o31a_1
XFILLER_35_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6874_ _6874_/A _7001_/B VGND VGND VPWR VPWR _6874_/Y sky130_fd_sc_hd__nand2_1
XFILLER_179_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8613_ _8859_/Q _8391_/A _8367_/A _9095_/Q VGND VGND VPWR VPWR _8613_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5825_ _9571_/A _5824_/X hold43/X VGND VGND VPWR VPWR _5825_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8544_ _9230_/Q _8388_/X _8379_/X _9206_/Q _8543_/X VGND VGND VPWR VPWR _8549_/B
+ sky130_fd_sc_hd__a221o_1
X_5756_ _5756_/A VGND VGND VPWR VPWR _8960_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4707_ _9395_/Q _7640_/A _7194_/A _9195_/Q VGND VGND VPWR VPWR _4707_/X sky130_fd_sc_hd__a22o_1
X_8475_ _8455_/X _8461_/X _8474_/X _8399_/A _9187_/Q VGND VGND VPWR VPWR _8475_/X
+ sky130_fd_sc_hd__o32a_2
X_5687_ hold46/X VGND VGND VPWR VPWR _5687_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_135_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7426_ _7302_/X hold914/X _7444_/S VGND VGND VPWR VPWR _7427_/A sky130_fd_sc_hd__mux2_1
X_4638_ _9420_/Q _7695_/A _7605_/A _9380_/Q VGND VGND VPWR VPWR _4638_/X sky130_fd_sc_hd__a22o_1
Xhold630 hold630/A VGND VGND VPWR VPWR hold630/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7357_ _7302_/X hold922/X _7372_/S VGND VGND VPWR VPWR _7358_/A sky130_fd_sc_hd__mux2_1
Xhold641 hold641/A VGND VGND VPWR VPWR hold641/X sky130_fd_sc_hd__dlygate4sd3_1
X_4569_ _4569_/A _4569_/B _4569_/C _4569_/D VGND VGND VPWR VPWR _4573_/C sky130_fd_sc_hd__or4_1
Xmax_cap360 _4478_/Y VGND VGND VPWR VPWR _7536_/A sky130_fd_sc_hd__buf_8
Xhold652 _6026_/X VGND VGND VPWR VPWR _6027_/A sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap371 _4501_/Y VGND VGND VPWR VPWR _7408_/A sky130_fd_sc_hd__buf_8
Xhold663 _8940_/Q VGND VGND VPWR VPWR hold663/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold674 _9051_/Q VGND VGND VPWR VPWR hold674/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6308_ _6790_/B _6894_/B VGND VGND VPWR VPWR _6708_/B sky130_fd_sc_hd__nor2_1
Xhold685 _9463_/Q VGND VGND VPWR VPWR hold685/X sky130_fd_sc_hd__dlygate4sd3_1
X_7288_ _7288_/A VGND VGND VPWR VPWR _9233_/D sky130_fd_sc_hd__clkbuf_1
Xhold696 _7039_/X VGND VGND VPWR VPWR _7040_/A sky130_fd_sc_hd__dlygate4sd3_1
X_9027_ _9551_/CLK _9027_/D fanout499/X VGND VGND VPWR VPWR _9027_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_77_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6239_ _6562_/A _6556_/B VGND VGND VPWR VPWR _6241_/B sky130_fd_sc_hd__or2_2
XFILLER_94_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__1160_ clkbuf_0__1160_/X VGND VGND VPWR VPWR _5988_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_154_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5610_ _5301_/X hold494/X _5616_/S VGND VGND VPWR VPWR _5611_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6590_ _6897_/A _6609_/A _6195_/B VGND VGND VPWR VPWR _6626_/B sky130_fd_sc_hd__o21a_1
X_5541_ _5291_/X hold906/X _5549_/S VGND VGND VPWR VPWR _5542_/A sky130_fd_sc_hd__mux2_1
X_8260_ _8260_/A _8260_/B _8260_/C _8260_/D VGND VGND VPWR VPWR _8260_/X sky130_fd_sc_hd__or4_1
X_5472_ _5471_/X hold450/X _5472_/S VGND VGND VPWR VPWR _5472_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7211_ _7211_/A _7284_/B VGND VGND VPWR VPWR _7226_/S sky130_fd_sc_hd__nand2_8
X_4423_ _4635_/A _4748_/B VGND VGND VPWR VPWR _7746_/A sky130_fd_sc_hd__nor2_8
X_8191_ _8978_/Q _7931_/A _7933_/X _8923_/Q VGND VGND VPWR VPWR _8191_/X sky130_fd_sc_hd__a22o_1
XFILLER_144_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7142_ _5951_/X _9169_/Q _7142_/S VGND VGND VPWR VPWR _7142_/X sky130_fd_sc_hd__mux2_1
X_4354_ _9110_/Q hold73/A VGND VGND VPWR VPWR _4354_/X sky130_fd_sc_hd__or2b_1
XFILLER_99_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout406 fanout407/X VGND VGND VPWR VPWR fanout406/X sky130_fd_sc_hd__buf_2
Xfanout417 _5332_/A VGND VGND VPWR VPWR _5070_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout428 fanout429/X VGND VGND VPWR VPWR fanout428/X sky130_fd_sc_hd__clkbuf_2
XFILLER_140_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7073_ _7073_/A VGND VGND VPWR VPWR _9139_/D sky130_fd_sc_hd__clkbuf_1
Xfanout439 fanout449/X VGND VGND VPWR VPWR fanout439/X sky130_fd_sc_hd__buf_2
XFILLER_59_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6024_ hold483/X _5809_/X _6030_/S VGND VGND VPWR VPWR _6024_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7975_ _9408_/Q _7967_/X _7969_/X _9288_/Q _7974_/X VGND VGND VPWR VPWR _8006_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6926_ _6926_/A _6926_/B VGND VGND VPWR VPWR _6928_/B sky130_fd_sc_hd__or2_1
X_6857_ _6857_/A _6857_/B _6857_/C _6857_/D VGND VGND VPWR VPWR _6946_/C sky130_fd_sc_hd__or4_1
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5808_ _5808_/A VGND VGND VPWR VPWR _8983_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9576_ _9576_/A _5092_/Y VGND VGND VPWR VPWR mgmt_gpio_out[22] sky130_fd_sc_hd__ebufn_8
X_6788_ _6788_/A _6788_/B _6788_/C VGND VGND VPWR VPWR _6939_/D sky130_fd_sc_hd__or3_2
XFILLER_22_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8527_ _5139_/A hold954/X _8013_/X VGND VGND VPWR VPWR _8527_/X sky130_fd_sc_hd__a21o_1
X_5739_ _5629_/X hold869/X _5747_/S VGND VGND VPWR VPWR _5740_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8458_ _9451_/Q _8310_/X _8381_/X _9363_/Q _8457_/X VGND VGND VPWR VPWR _8458_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_163_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7409_ _7302_/X hold905/X _7423_/S VGND VGND VPWR VPWR _7410_/A sky130_fd_sc_hd__mux2_1
X_8389_ _8389_/A _8398_/A _8389_/C VGND VGND VPWR VPWR _8657_/B sky130_fd_sc_hd__and3_4
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold460 _7152_/X VGND VGND VPWR VPWR _7153_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold471 _8833_/Q VGND VGND VPWR VPWR hold471/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 _5917_/X VGND VGND VPWR VPWR _9024_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 _7060_/X VGND VGND VPWR VPWR _7061_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1160 _5747_/X VGND VGND VPWR VPWR _5748_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1171 _8921_/Q VGND VGND VPWR VPWR hold421/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1182 _8864_/Q VGND VGND VPWR VPWR hold495/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1193 _8895_/Q VGND VGND VPWR VPWR hold638/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_300 _5901_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_311 _9503_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_322 _9355_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_333 _5291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_344 _6015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_355 _7779_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_366 _9340_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_377 input42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_388 hold46/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_399 _7156_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7760_ hold379/X _7494_/A _7762_/S VGND VGND VPWR VPWR _7760_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4972_ _5068_/B _4972_/B VGND VGND VPWR VPWR _8806_/D sky130_fd_sc_hd__xor2_1
XFILLER_51_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6711_ _6754_/A _6754_/C _6964_/A _6710_/X _6382_/X VGND VGND VPWR VPWR _6711_/X
+ sky130_fd_sc_hd__o41a_1
X_7691_ _5410_/X hold201/X _7693_/S VGND VGND VPWR VPWR _7691_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9430_ _9471_/CLK _9430_/D fanout421/X VGND VGND VPWR VPWR _9430_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_149_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6642_ _6843_/C _6642_/B VGND VGND VPWR VPWR _6642_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9361_ _9475_/CLK _9361_/D fanout479/X VGND VGND VPWR VPWR _9361_/Q sky130_fd_sc_hd__dfstp_2
X_6573_ _6993_/A _6573_/B VGND VGND VPWR VPWR _7002_/C sky130_fd_sc_hd__or2_1
X_8312_ _8354_/A VGND VGND VPWR VPWR _8312_/X sky130_fd_sc_hd__buf_6
X_5524_ _5524_/A VGND VGND VPWR VPWR _8860_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9292_ _9436_/CLK _9292_/D fanout462/X VGND VGND VPWR VPWR _9292_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_173_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR clkbuf_2_3_0_mgmt_gpio_in[4]/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_8_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8243_ _8986_/Q _7993_/X _7999_/X _8951_/Q _8242_/X VGND VGND VPWR VPWR _8250_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_172_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5455_ _5291_/X hold828/X _5472_/S VGND VGND VPWR VPWR _5455_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4406_ _4492_/A _4499_/A VGND VGND VPWR VPWR _4406_/Y sky130_fd_sc_hd__nor2_4
XFILLER_132_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8174_ hold982/X _8017_/X _8173_/X VGND VGND VPWR VPWR _9514_/D sky130_fd_sc_hd__o21a_1
X_5386_ _5386_/A VGND VGND VPWR VPWR _5386_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7125_ _7125_/A VGND VGND VPWR VPWR _9162_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7056_ _7056_/A hold19/X VGND VGND VPWR VPWR _7057_/A sky130_fd_sc_hd__and2_1
XFILLER_74_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6007_ _6007_/A _7043_/B VGND VGND VPWR VPWR _6019_/S sky130_fd_sc_hd__nand2_2
XFILLER_74_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7958_ _7958_/A VGND VGND VPWR VPWR _7958_/X sky130_fd_sc_hd__buf_6
XFILLER_54_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6909_ _6824_/B _6889_/X _6905_/X _6908_/X VGND VGND VPWR VPWR _6909_/X sky130_fd_sc_hd__o31a_1
X_7889_ _7889_/A VGND VGND VPWR VPWR _9496_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9559_ _9559_/A _5109_/Y VGND VGND VPWR VPWR mgmt_gpio_out[5] sky130_fd_sc_hd__ebufn_8
XFILLER_183_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold290 _7293_/X VGND VGND VPWR VPWR _7294_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_130 _7517_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_141 _7908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_152 _7938_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_163 _7949_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 _7967_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_185 _7990_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_196 _8001_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5240_ _9219_/Q VGND VGND VPWR VPWR _5240_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5171_ _8795_/Q input86/X VGND VGND VPWR VPWR _5172_/A sky130_fd_sc_hd__or2b_1
XFILLER_123_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8930_ _9184_/CLK _8930_/D fanout439/X VGND VGND VPWR VPWR _8930_/Q sky130_fd_sc_hd__dfstp_1
Xinput3 debug_out VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8861_ _9184_/CLK _8861_/D fanout443/X VGND VGND VPWR VPWR _8861_/Q sky130_fd_sc_hd__dfrtp_4
X_7812_ _7812_/A VGND VGND VPWR VPWR _9470_/D sky130_fd_sc_hd__clkbuf_1
X_8792_ _8831_/CLK _8792_/D _5350_/X VGND VGND VPWR VPWR _8792_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7743_ _7743_/A VGND VGND VPWR VPWR _9438_/D sky130_fd_sc_hd__clkbuf_1
X_4955_ _9216_/Q _7249_/A _7176_/A _9184_/Q _4954_/X VGND VGND VPWR VPWR _4959_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_189_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7674_ _7494_/X hold740/X _7676_/S VGND VGND VPWR VPWR _7674_/X sky130_fd_sc_hd__mux2_1
X_4886_ _9111_/Q _4885_/X _4886_/S VGND VGND VPWR VPWR _4886_/X sky130_fd_sc_hd__mux2_1
X_9413_ _9413_/CLK _9413_/D fanout458/X VGND VGND VPWR VPWR _9413_/Q sky130_fd_sc_hd__dfrtp_1
X_6625_ _6716_/B _6243_/A _6623_/Y _6609_/A _6959_/A VGND VGND VPWR VPWR _6626_/D
+ sky130_fd_sc_hd__a41o_1
XFILLER_192_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9344_ _9416_/CLK _9344_/D fanout425/X VGND VGND VPWR VPWR _9344_/Q sky130_fd_sc_hd__dfstp_1
X_6556_ _6562_/A _6556_/B VGND VGND VPWR VPWR _6563_/A sky130_fd_sc_hd__nor2_2
X_5507_ hold917/X _5505_/X _5515_/S VGND VGND VPWR VPWR _5508_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9275_ _9291_/CLK _9275_/D fanout468/X VGND VGND VPWR VPWR _9275_/Q sky130_fd_sc_hd__dfrtp_4
X_6487_ _6858_/B _6435_/A _6524_/C _6894_/B VGND VGND VPWR VPWR _6978_/A sky130_fd_sc_hd__o22a_1
XFILLER_10_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8226_ _8880_/Q _7969_/X _7977_/X _8774_/Q VGND VGND VPWR VPWR _8226_/X sky130_fd_sc_hd__a22o_1
X_5438_ _5291_/X _8825_/Q _5440_/S VGND VGND VPWR VPWR _5438_/X sky130_fd_sc_hd__mux2_1
Xoutput340 _9045_/Q VGND VGND VPWR VPWR wb_dat_o[21] sky130_fd_sc_hd__buf_12
XFILLER_121_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput351 _9541_/Q VGND VGND VPWR VPWR wb_dat_o[31] sky130_fd_sc_hd__buf_12
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8157_ _9327_/Q _7962_/X _7988_/X _9439_/Q VGND VGND VPWR VPWR _8157_/X sky130_fd_sc_hd__a22o_1
X_5369_ _5375_/A _5378_/B VGND VGND VPWR VPWR _5370_/A sky130_fd_sc_hd__and2_1
XFILLER_114_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7108_ _7108_/A _7139_/B VGND VGND VPWR VPWR _7109_/S sky130_fd_sc_hd__nand2_1
X_8088_ _9380_/Q _7947_/X _7981_/X _9332_/Q VGND VGND VPWR VPWR _8088_/X sky130_fd_sc_hd__a22o_1
XFILLER_47_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7039_ _6015_/X _9124_/Q _7041_/S VGND VGND VPWR VPWR _7039_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ input38/X _4436_/A _5784_/A _8976_/Q _4739_/X VGND VGND VPWR VPWR _4741_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4671_ _9476_/Q _7815_/A _7032_/A _9125_/Q VGND VGND VPWR VPWR _4671_/X sky130_fd_sc_hd__a22o_1
X_6410_ _6504_/A _6739_/A VGND VGND VPWR VPWR _6597_/B sky130_fd_sc_hd__nor2_8
XFILLER_147_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7390_ _7390_/A VGND VGND VPWR VPWR _9279_/D sky130_fd_sc_hd__clkbuf_1
X_6341_ _6341_/A _6881_/A VGND VGND VPWR VPWR _6937_/A sky130_fd_sc_hd__nor2_1
XFILLER_115_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9060_ _9541_/CLK _9060_/D VGND VGND VPWR VPWR _9060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6272_ _6268_/X _6853_/A _6272_/C _6272_/D VGND VGND VPWR VPWR _6272_/X sky130_fd_sc_hd__and4bb_1
XFILLER_170_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8011_ _8015_/A _8015_/B VGND VGND VPWR VPWR _8012_/A sky130_fd_sc_hd__or2_1
XFILLER_88_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5223_ _5223_/A VGND VGND VPWR VPWR _5223_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_130_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5154_ _8999_/Q VGND VGND VPWR VPWR _7916_/C sky130_fd_sc_hd__inv_2
XFILLER_96_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5085_ _9419_/Q VGND VGND VPWR VPWR _5085_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8913_ _9427_/CLK _8913_/D fanout478/X VGND VGND VPWR VPWR _8913_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_37_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8844_ _9006_/CLK _8844_/D fanout493/X VGND VGND VPWR VPWR _8844_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_52_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8775_ _9184_/CLK _8775_/D fanout438/X VGND VGND VPWR VPWR _8775_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5987_ _5987_/A VGND VGND VPWR VPWR _9064_/D sky130_fd_sc_hd__clkbuf_1
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4938_ _9272_/Q _4938_/A2 _7781_/A _9456_/Q _4937_/X VGND VGND VPWR VPWR _4939_/D
+ sky130_fd_sc_hd__a221o_1
X_7726_ _7726_/A VGND VGND VPWR VPWR _9430_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_30 _4577_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7657_ _7494_/X hold732/X hold84/X VGND VGND VPWR VPWR _7658_/A sky130_fd_sc_hd__mux2_1
X_4869_ _8944_/Q _5715_/A _5795_/A _8979_/Q VGND VGND VPWR VPWR _4869_/X sky130_fd_sc_hd__a22o_1
XANTENNA_41 _5630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_52 _4883_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_63 _5067_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_74 hold19/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6608_ _6158_/B _6125_/A _6194_/B _6227_/Y VGND VGND VPWR VPWR _6608_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_21_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_85 _5690_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7588_ _7588_/A _7695_/B VGND VGND VPWR VPWR hold75/A sky130_fd_sc_hd__nand2_8
XANTENNA_96 _5629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9327_ _9367_/CLK _9327_/D fanout423/X VGND VGND VPWR VPWR _9327_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6539_ _6539_/A _6539_/B _6539_/C _6539_/D VGND VGND VPWR VPWR _6540_/D sky130_fd_sc_hd__and4_1
XFILLER_118_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9258_ _9466_/CLK _9258_/D fanout471/X VGND VGND VPWR VPWR _9258_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_97_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8209_ _8209_/A _8209_/B _8209_/C _8209_/D VGND VGND VPWR VPWR _8216_/B sky130_fd_sc_hd__or4_1
XFILLER_106_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9189_ _9486_/CLK _9189_/D fanout416/X VGND VGND VPWR VPWR _9189_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_102_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5910_ _5653_/X _9582_/A _5916_/S VGND VGND VPWR VPWR _5910_/X sky130_fd_sc_hd__mux2_1
X_6890_ _6894_/A _6895_/B _6926_/B VGND VGND VPWR VPWR _6890_/X sky130_fd_sc_hd__a21o_1
XFILLER_34_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5841_ _5841_/A VGND VGND VPWR VPWR _5841_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_61_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5772_ _5772_/A VGND VGND VPWR VPWR _8967_/D sky130_fd_sc_hd__clkbuf_1
X_8560_ _9335_/Q _8298_/X _8370_/X _9255_/Q _8559_/X VGND VGND VPWR VPWR _8563_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_15_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4723_ _4723_/A _4723_/B _4723_/C _4723_/D VGND VGND VPWR VPWR _4724_/D sky130_fd_sc_hd__or4_1
X_7511_ _7511_/A VGND VGND VPWR VPWR _9333_/D sky130_fd_sc_hd__clkbuf_1
X_8491_ _9284_/Q _8316_/X _8327_/X _9260_/Q VGND VGND VPWR VPWR _8491_/X sky130_fd_sc_hd__a22o_1
XFILLER_187_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7442_ _7279_/X hold836/X _7444_/S VGND VGND VPWR VPWR _7442_/X sky130_fd_sc_hd__mux2_1
X_4654_ _9428_/Q _7712_/A _5529_/A _8867_/Q _4653_/X VGND VGND VPWR VPWR _4654_/X
+ sky130_fd_sc_hd__a221o_1
Xinput50 mgmt_gpio_in[22] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__clkbuf_4
Xinput61 mgmt_gpio_in[32] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__clkbuf_2
X_7373_ _7373_/A VGND VGND VPWR VPWR _9271_/D sky130_fd_sc_hd__clkbuf_1
X_4585_ hold33/X _4956_/A VGND VGND VPWR VPWR _4585_/Y sky130_fd_sc_hd__nor2_2
Xhold801 _7199_/X VGND VGND VPWR VPWR _7200_/A sky130_fd_sc_hd__dlygate4sd3_1
Xinput72 mgmt_gpio_in[9] VGND VGND VPWR VPWR input72/X sky130_fd_sc_hd__clkbuf_1
Xhold812 _9037_/Q VGND VGND VPWR VPWR hold812/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_174_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold823 _8852_/Q VGND VGND VPWR VPWR hold823/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput83 spimemio_flash_clk VGND VGND VPWR VPWR input83/X sky130_fd_sc_hd__buf_2
Xinput94 sram_ro_data[10] VGND VGND VPWR VPWR input94/X sky130_fd_sc_hd__clkbuf_2
X_9112_ _5235__1/A _9112_/D _7014_/X VGND VGND VPWR VPWR _9112_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_116_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold834 _9286_/Q VGND VGND VPWR VPWR hold834/X sky130_fd_sc_hd__dlygate4sd3_1
X_6324_ _6324_/A _6828_/A VGND VGND VPWR VPWR _6325_/A sky130_fd_sc_hd__or2_1
XFILLER_143_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold845 hold845/A VGND VGND VPWR VPWR hold845/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 _5949_/X VGND VGND VPWR VPWR _5950_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 hold867/A VGND VGND VPWR VPWR _7141_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold878 _9376_/Q VGND VGND VPWR VPWR hold878/X sky130_fd_sc_hd__dlygate4sd3_1
X_9043_ _9541_/CLK _9043_/D VGND VGND VPWR VPWR _9043_/Q sky130_fd_sc_hd__dfxtp_1
Xhold889 _9352_/Q VGND VGND VPWR VPWR hold889/X sky130_fd_sc_hd__dlygate4sd3_1
X_6255_ _6881_/A _6610_/A VGND VGND VPWR VPWR _6255_/X sky130_fd_sc_hd__or2_1
XFILLER_115_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5206_ _5206_/A VGND VGND VPWR VPWR _9564_/A sky130_fd_sc_hd__clkbuf_1
X_6186_ _6175_/A _6633_/A _6437_/A VGND VGND VPWR VPWR _6187_/B sky130_fd_sc_hd__a21oi_1
XFILLER_57_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5137_ _7911_/B _7860_/A _9490_/Q _9491_/Q VGND VGND VPWR VPWR _5160_/B sky130_fd_sc_hd__and4b_1
X_5068_ _8808_/Q _5068_/B _5068_/C VGND VGND VPWR VPWR _5068_/Y sky130_fd_sc_hd__nand3_1
XFILLER_84_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8827_ _5168_/A1 _8827_/D _5443_/X VGND VGND VPWR VPWR _8827_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8758_ _8758_/A VGND VGND VPWR VPWR _9547_/D sky130_fd_sc_hd__clkbuf_1
X_7709_ _7709_/A VGND VGND VPWR VPWR _9422_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8689_ _8862_/Q _8391_/X _8367_/X _9098_/Q VGND VGND VPWR VPWR _8689_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold108 _9249_/Q VGND VGND VPWR VPWR hold108/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold119 _9257_/Q VGND VGND VPWR VPWR hold119/X sky130_fd_sc_hd__dlygate4sd3_1
X_4370_ hold8/X hold7/X hold94/X VGND VGND VPWR VPWR hold9/A sky130_fd_sc_hd__mux2_1
XFILLER_171_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6040_/A VGND VGND VPWR VPWR _9087_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7991_ _7998_/A _7991_/B _7996_/B VGND VGND VPWR VPWR _8077_/A sky130_fd_sc_hd__and3_2
X_6942_ _6942_/A _6942_/B VGND VGND VPWR VPWR _6953_/C sky130_fd_sc_hd__and2_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6873_ _6906_/A _6873_/B VGND VGND VPWR VPWR _6873_/Y sky130_fd_sc_hd__nand2_1
X_8612_ _8969_/Q _8506_/B _8607_/X _8609_/X _8611_/X VGND VGND VPWR VPWR _8612_/X
+ sky130_fd_sc_hd__a2111o_1
X_5824_ hold471/X hold37/X _5842_/S VGND VGND VPWR VPWR _5824_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8543_ _9390_/Q _8292_/X _8294_/X _9294_/Q VGND VGND VPWR VPWR _8543_/X sky130_fd_sc_hd__a22o_1
X_5755_ hold569/X _5683_/X _5759_/S VGND VGND VPWR VPWR _5756_/A sky130_fd_sc_hd__mux2_1
X_4706_ _9259_/Q _7339_/A _4477_/Y input29/X _4705_/X VGND VGND VPWR VPWR _4711_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8474_ _8474_/A _8474_/B _8474_/C _8474_/D VGND VGND VPWR VPWR _8474_/X sky130_fd_sc_hd__or4_1
XFILLER_147_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5686_ hold45/X VGND VGND VPWR VPWR hold46/A sky130_fd_sc_hd__buf_6
X_4637_ _9484_/Q _4898_/A2 _5573_/A _8887_/Q _4636_/X VGND VGND VPWR VPWR _4649_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7425_ _7425_/A _7499_/B VGND VGND VPWR VPWR _7444_/S sky130_fd_sc_hd__nand2_8
XFILLER_163_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold620 _8897_/Q VGND VGND VPWR VPWR hold620/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 _9199_/Q VGND VGND VPWR VPWR hold631/X sky130_fd_sc_hd__dlygate4sd3_1
X_4568_ _9293_/Q _7408_/A _4836_/A2 _9453_/Q _4567_/X VGND VGND VPWR VPWR _4569_/D
+ sky130_fd_sc_hd__a221o_2
X_7356_ _7356_/A _7499_/B VGND VGND VPWR VPWR _7372_/S sky130_fd_sc_hd__nand2_8
Xhold642 hold642/A VGND VGND VPWR VPWR hold642/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap361 _4459_/Y VGND VGND VPWR VPWR _7499_/A sky130_fd_sc_hd__buf_8
Xhold653 _9455_/Q VGND VGND VPWR VPWR hold653/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap372 _4491_/Y VGND VGND VPWR VPWR _5901_/A sky130_fd_sc_hd__buf_8
Xhold664 hold664/A VGND VGND VPWR VPWR hold664/X sky130_fd_sc_hd__dlygate4sd3_1
X_6307_ _6894_/B _6435_/A VGND VGND VPWR VPWR _6588_/B sky130_fd_sc_hd__nor2_1
Xmax_cap383 _4424_/Y VGND VGND VPWR VPWR _7194_/A sky130_fd_sc_hd__buf_8
Xhold675 _5956_/X VGND VGND VPWR VPWR _5957_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7287_ _7147_/X hold115/X _7300_/S VGND VGND VPWR VPWR _7287_/X sky130_fd_sc_hd__mux2_1
Xmax_cap394 _6376_/A VGND VGND VPWR VPWR _6547_/B sky130_fd_sc_hd__clkbuf_2
X_4499_ _4499_/A VGND VGND VPWR VPWR _7111_/B sky130_fd_sc_hd__buf_6
Xhold686 _7796_/X VGND VGND VPWR VPWR _7797_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold697 hold697/A VGND VGND VPWR VPWR _7382_/A sky130_fd_sc_hd__dlygate4sd3_1
X_9026_ _9551_/CLK _9026_/D fanout499/X VGND VGND VPWR VPWR _9026_/Q sky130_fd_sc_hd__dfrtp_1
X_6238_ _6603_/A _6279_/A VGND VGND VPWR VPWR _6857_/A sky130_fd_sc_hd__nor2_1
XFILLER_103_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6169_ _6169_/A _6175_/A _6633_/A VGND VGND VPWR VPWR _6317_/B sky130_fd_sc_hd__and3_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_43_csclk _8954_/CLK VGND VGND VPWR VPWR _9243_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_150_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_58_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _9084_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_40_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5540_ _5540_/A _5693_/B VGND VGND VPWR VPWR _5549_/S sky130_fd_sc_hd__nand2_2
XFILLER_192_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5471_ _7514_/A VGND VGND VPWR VPWR _5471_/X sky130_fd_sc_hd__buf_6
XFILLER_172_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4422_ _4675_/B VGND VGND VPWR VPWR _4635_/A sky130_fd_sc_hd__buf_12
X_7210_ _7210_/A VGND VGND VPWR VPWR _9199_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8190_ _9035_/Q _7938_/X _8077_/X _8933_/Q _8189_/X VGND VGND VPWR VPWR _8193_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_172_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7141_ _7141_/A VGND VGND VPWR VPWR _9168_/D sky130_fd_sc_hd__clkbuf_1
X_4353_ hold55/X hold22/X VGND VGND VPWR VPWR hold56/A sky130_fd_sc_hd__and2_1
Xfanout407 fanout410/X VGND VGND VPWR VPWR fanout407/X sky130_fd_sc_hd__clkbuf_2
XFILLER_99_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout418 fanout426/X VGND VGND VPWR VPWR _5332_/A sky130_fd_sc_hd__clkbuf_4
X_7072_ _9139_/Q _7514_/A _7072_/S VGND VGND VPWR VPWR _7072_/X sky130_fd_sc_hd__mux2_1
Xfanout429 fanout435/X VGND VGND VPWR VPWR fanout429/X sky130_fd_sc_hd__clkbuf_4
XFILLER_140_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6023_ _6023_/A VGND VGND VPWR VPWR _9079_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7974_ _9416_/Q _8224_/B _7973_/X _9192_/Q VGND VGND VPWR VPWR _7974_/X sky130_fd_sc_hd__a22o_1
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6925_ _6925_/A _6925_/B _6925_/C _6988_/B VGND VGND VPWR VPWR _6925_/X sky130_fd_sc_hd__or4_1
XFILLER_35_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6856_ _6856_/A _6856_/B _6855_/X VGND VGND VPWR VPWR _6969_/C sky130_fd_sc_hd__or3b_1
XFILLER_22_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5807_ hold895/X _5761_/X _5816_/S VGND VGND VPWR VPWR _5808_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9575_ _9575_/A _5093_/Y VGND VGND VPWR VPWR mgmt_gpio_out[21] sky130_fd_sc_hd__ebufn_8
X_6787_ _6790_/A _6764_/A _6624_/B VGND VGND VPWR VPWR _6939_/C sky130_fd_sc_hd__a21o_1
X_8526_ _9189_/Q _8400_/B _8512_/X _8525_/X _8105_/X VGND VGND VPWR VPWR _8526_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5738_ _5738_/A _7043_/B VGND VGND VPWR VPWR _5747_/S sky130_fd_sc_hd__nand2_4
XFILLER_6_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8457_ _9331_/Q _8298_/A _8370_/A _9251_/Q VGND VGND VPWR VPWR _8457_/X sky130_fd_sc_hd__a22o_1
XFILLER_175_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5669_ _5669_/A VGND VGND VPWR VPWR _8923_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7408_ _7408_/A _7499_/B VGND VGND VPWR VPWR _7423_/S sky130_fd_sc_hd__nand2_8
XFILLER_151_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8388_ _8388_/A VGND VGND VPWR VPWR _8388_/X sky130_fd_sc_hd__buf_8
XFILLER_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold450 _8839_/Q VGND VGND VPWR VPWR hold450/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold461 _7153_/X VGND VGND VPWR VPWR _9173_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7339_ _7339_/A _7499_/B VGND VGND VPWR VPWR _7354_/S sky130_fd_sc_hd__nand2_4
Xhold472 _5457_/X VGND VGND VPWR VPWR _5458_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 _9080_/Q VGND VGND VPWR VPWR hold483/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 hold494/A VGND VGND VPWR VPWR hold494/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9009_ _9464_/CLK _9009_/D fanout420/X VGND VGND VPWR VPWR _9009_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1150 _8888_/Q VGND VGND VPWR VPWR hold939/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1161 _5889_/X VGND VGND VPWR VPWR hold1161/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1172 _8919_/Q VGND VGND VPWR VPWR hold742/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1183 _8941_/Q VGND VGND VPWR VPWR hold505/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1194 _9088_/Q VGND VGND VPWR VPWR hold498/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_301 _4898_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_312 _9532_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_323 _9371_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_334 _5301_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_345 _6015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_356 _7933_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_367 _8962_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_378 input40/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_389 _8995_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_110_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4971_ _4971_/A _4971_/B VGND VGND VPWR VPWR _8807_/D sky130_fd_sc_hd__nor2_1
XFILLER_91_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6710_ _6710_/A _6948_/B _6710_/C _6710_/D VGND VGND VPWR VPWR _6710_/X sky130_fd_sc_hd__or4_1
XFILLER_51_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7690_ _7690_/A VGND VGND VPWR VPWR _9413_/D sky130_fd_sc_hd__clkbuf_1
X_6641_ _6850_/A _6640_/Y _6462_/B VGND VGND VPWR VPWR _6641_/X sky130_fd_sc_hd__a21o_1
XFILLER_177_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9360_ _9416_/CLK _9360_/D fanout425/X VGND VGND VPWR VPWR _9360_/Q sky130_fd_sc_hd__dfstp_1
X_6572_ _6340_/Y _6551_/Y _6882_/C _6937_/B VGND VGND VPWR VPWR _6576_/C sky130_fd_sc_hd__a211o_1
XFILLER_164_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8311_ _8355_/A _8392_/A _8392_/C VGND VGND VPWR VPWR _8354_/A sky130_fd_sc_hd__and3b_4
XFILLER_192_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5523_ _5306_/X hold508/X _5527_/S VGND VGND VPWR VPWR _5523_/X sky130_fd_sc_hd__mux2_1
X_9291_ _9291_/CLK _9291_/D fanout468/X VGND VGND VPWR VPWR _9291_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8242_ _9051_/Q _7923_/X _7938_/X _9038_/Q VGND VGND VPWR VPWR _8242_/X sky130_fd_sc_hd__a22o_1
X_5454_ _5454_/A VGND VGND VPWR VPWR _5472_/S sky130_fd_sc_hd__buf_4
X_4405_ _4405_/A VGND VGND VPWR VPWR _4499_/A sky130_fd_sc_hd__clkbuf_16
X_5385_ _7011_/A _7013_/B VGND VGND VPWR VPWR _5386_/A sky130_fd_sc_hd__and2_1
X_8173_ _5130_/A hold976/X _8013_/A _8172_/X VGND VGND VPWR VPWR _8173_/X sky130_fd_sc_hd__a211o_1
X_7124_ _5951_/X _9162_/Q _7124_/S VGND VGND VPWR VPWR _7124_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7055_ _7055_/A VGND VGND VPWR VPWR _9131_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6006_ _6006_/A VGND VGND VPWR VPWR _9073_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7957_ _8181_/B _8000_/B _7992_/C VGND VGND VPWR VPWR _7958_/A sky130_fd_sc_hd__and3_4
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6908_ _6908_/A _6978_/B VGND VGND VPWR VPWR _6908_/X sky130_fd_sc_hd__and2_1
X_7888_ _7887_/Y _8275_/B _7888_/S VGND VGND VPWR VPWR _7889_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6839_ _6839_/A _6839_/B VGND VGND VPWR VPWR _6839_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9558_ _9558_/A _5110_/Y VGND VGND VPWR VPWR mgmt_gpio_out[4] sky130_fd_sc_hd__ebufn_8
XFILLER_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8509_ _9453_/Q _8310_/X _8381_/X _9365_/Q _8508_/X VGND VGND VPWR VPWR _8512_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9489_ _9532_/CLK _9489_/D fanout442/X VGND VGND VPWR VPWR _9489_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_136_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold280 _7402_/X VGND VGND VPWR VPWR _7403_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 _9445_/Q VGND VGND VPWR VPWR hold291/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_120 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_131 _7517_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_142 _7908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_153 _7940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_164 _7949_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_175 _7969_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_186 _7993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_197 _8001_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5170_ _8794_/Q _5330_/A VGND VGND VPWR VPWR _5170_/Y sky130_fd_sc_hd__nor2_2
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput4 mask_rev_in[0] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8860_ _9184_/CLK _8860_/D fanout443/X VGND VGND VPWR VPWR _8860_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_92_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7811_ _5410_/X hold194/X _7813_/S VGND VGND VPWR VPWR _7811_/X sky130_fd_sc_hd__mux2_1
X_8791_ _5168_/A1 _8791_/D _5348_/X VGND VGND VPWR VPWR _8791_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_51_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7742_ _5410_/X hold335/X hold86/X VGND VGND VPWR VPWR _7743_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4954_ _9416_/Q _4439_/Y _5678_/A _8928_/Q VGND VGND VPWR VPWR _4954_/X sky130_fd_sc_hd__a22o_1
XFILLER_51_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7673_ _7673_/A VGND VGND VPWR VPWR _9405_/D sky130_fd_sc_hd__clkbuf_1
X_4885_ _4885_/A _4885_/B _4885_/C VGND VGND VPWR VPWR _4885_/X sky130_fd_sc_hd__or3_4
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9412_ _9468_/CLK _9412_/D fanout465/X VGND VGND VPWR VPWR _9412_/Q sky130_fd_sc_hd__dfrtp_4
X_6624_ _6873_/B _6624_/B VGND VGND VPWR VPWR _6959_/A sky130_fd_sc_hd__nor2_2
XFILLER_165_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9343_ _9471_/CLK _9343_/D _5332_/A VGND VGND VPWR VPWR _9343_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_118_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6555_ _6853_/A _6758_/A VGND VGND VPWR VPWR _6872_/C sky130_fd_sc_hd__or2_1
XFILLER_192_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5506_ _5506_/A _5715_/B VGND VGND VPWR VPWR _5515_/S sky130_fd_sc_hd__and2_2
XFILLER_146_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9274_ _9290_/CLK _9274_/D fanout468/X VGND VGND VPWR VPWR _9274_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6486_ _6486_/A VGND VGND VPWR VPWR _6809_/D sky130_fd_sc_hd__inv_2
XFILLER_133_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8225_ _8980_/Q _7931_/X _7979_/X _9071_/Q _8224_/X VGND VGND VPWR VPWR _8228_/C
+ sky130_fd_sc_hd__a221o_1
X_5437_ _5437_/A _7139_/B VGND VGND VPWR VPWR _5440_/S sky130_fd_sc_hd__nand2_1
XFILLER_105_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput330 _9057_/Q VGND VGND VPWR VPWR wb_dat_o[12] sky130_fd_sc_hd__buf_12
Xoutput341 _9046_/Q VGND VGND VPWR VPWR wb_dat_o[22] sky130_fd_sc_hd__buf_12
Xoutput352 _9064_/Q VGND VGND VPWR VPWR wb_dat_o[3] sky130_fd_sc_hd__buf_12
X_5368_ _5368_/A VGND VGND VPWR VPWR _5368_/X sky130_fd_sc_hd__clkbuf_1
X_8156_ _9255_/Q _7940_/X _7969_/X _9295_/Q _8155_/X VGND VGND VPWR VPWR _8162_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_126_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7107_ _7107_/A VGND VGND VPWR VPWR _9154_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8087_ _9356_/Q _8020_/X _7990_/X _9276_/Q _8086_/X VGND VGND VPWR VPWR _8104_/A
+ sky130_fd_sc_hd__a221o_1
X_5299_ hold36/X hold68/X _5413_/S VGND VGND VPWR VPWR hold69/A sky130_fd_sc_hd__mux2_8
X_7038_ _7038_/A VGND VGND VPWR VPWR _9123_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8989_ _9006_/CLK _8989_/D fanout493/X VGND VGND VPWR VPWR _9571_/A sky130_fd_sc_hd__dfrtp_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4670_ _4758_/A _4670_/B VGND VGND VPWR VPWR _7032_/A sky130_fd_sc_hd__nor2_4
XFILLER_174_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6340_ _6562_/A _6558_/B VGND VGND VPWR VPWR _6340_/Y sky130_fd_sc_hd__nor2_2
X_6271_ _6802_/A _6790_/B VGND VGND VPWR VPWR _6272_/D sky130_fd_sc_hd__or2_1
XFILLER_182_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8010_ _9184_/Q _8010_/B VGND VGND VPWR VPWR _8010_/X sky130_fd_sc_hd__or2_1
X_5222_ _5219_/Y input2/X input1/X VGND VGND VPWR VPWR _5223_/A sky130_fd_sc_hd__mux2_4
X_5153_ _8996_/Q VGND VGND VPWR VPWR _7902_/A sky130_fd_sc_hd__clkinv_2
XFILLER_130_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5084_ _9427_/Q VGND VGND VPWR VPWR _5084_/Y sky130_fd_sc_hd__inv_2
X_8912_ _9227_/CLK _8912_/D fanout450/X VGND VGND VPWR VPWR _8912_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8843_ _9172_/CLK _8843_/D fanout493/X VGND VGND VPWR VPWR _8843_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_37_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8774_ _9162_/CLK _8774_/D fanout438/X VGND VGND VPWR VPWR _8774_/Q sky130_fd_sc_hd__dfstp_2
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5986_ _9064_/Q _4752_/X _5994_/S VGND VGND VPWR VPWR _5987_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7725_ _5410_/X hold196/X hold95/X VGND VGND VPWR VPWR _7726_/A sky130_fd_sc_hd__mux2_1
X_4937_ _9440_/Q _7746_/A _4414_/Y _9336_/Q VGND VGND VPWR VPWR _4937_/X sky130_fd_sc_hd__a22o_1
XFILLER_177_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_20 _4506_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7656_ _7656_/A VGND VGND VPWR VPWR _9397_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_31 _5842_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4868_ _9257_/Q _7339_/A _5918_/A _9036_/Q _4867_/X VGND VGND VPWR VPWR _4873_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_138_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_42 _4702_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_53 _4885_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_64 _5067_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6607_ _6967_/A _6607_/B VGND VGND VPWR VPWR _6607_/Y sky130_fd_sc_hd__nor2_1
XFILLER_177_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_75 hold19/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7587_ _7587_/A VGND VGND VPWR VPWR _9367_/D sky130_fd_sc_hd__clkbuf_1
X_4799_ _9330_/Q _4459_/Y _5518_/A _8860_/Q _4798_/X VGND VGND VPWR VPWR _4806_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA_86 _5465_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_97 _5690_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9326_ _9367_/CLK _9326_/D fanout423/X VGND VGND VPWR VPWR _9326_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6538_ _6906_/C _6524_/C _6862_/A _6591_/B _6537_/X VGND VGND VPWR VPWR _6539_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_192_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9257_ _9483_/CLK _9257_/D fanout473/X VGND VGND VPWR VPWR _9257_/Q sky130_fd_sc_hd__dfstp_2
X_6469_ _6948_/A _6469_/B _6469_/C _6469_/D VGND VGND VPWR VPWR _6469_/X sky130_fd_sc_hd__or4_1
XFILLER_106_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8208_ _8859_/Q _7927_/X _8023_/B _8889_/Q _8207_/X VGND VGND VPWR VPWR _8209_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9188_ _9203_/CLK _9188_/D fanout450/X VGND VGND VPWR VPWR _9188_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_121_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8139_ _9222_/Q _7927_/A _7956_/A _9310_/Q _8138_/X VGND VGND VPWR VPWR _8140_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_87_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5840_ _9576_/A _5839_/X hold43/X VGND VGND VPWR VPWR _5840_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5771_ hold635/X _5690_/X _5771_/S VGND VGND VPWR VPWR _5772_/A sky130_fd_sc_hd__mux2_1
X_7510_ _7439_/X hold262/X _7515_/S VGND VGND VPWR VPWR _7510_/X sky130_fd_sc_hd__mux2_1
X_4722_ _9387_/Q _4445_/Y _5738_/A _8956_/Q _4721_/X VGND VGND VPWR VPWR _4723_/D
+ sky130_fd_sc_hd__a221o_1
X_8490_ _9460_/Q _8348_/X _8411_/X _9340_/Q _8489_/X VGND VGND VPWR VPWR _8500_/B
+ sky130_fd_sc_hd__a221o_1
X_7441_ _7441_/A VGND VGND VPWR VPWR _9301_/D sky130_fd_sc_hd__clkbuf_1
X_4653_ _9332_/Q _7499_/A _5715_/A _8947_/Q VGND VGND VPWR VPWR _4653_/X sky130_fd_sc_hd__a22o_1
Xinput40 mgmt_gpio_in[13] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__buf_2
Xinput51 mgmt_gpio_in[23] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__clkbuf_4
X_7372_ _7299_/X hold668/X _7372_/S VGND VGND VPWR VPWR _7372_/X sky130_fd_sc_hd__mux2_1
Xinput62 mgmt_gpio_in[33] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__clkbuf_2
Xhold802 hold802/A VGND VGND VPWR VPWR _7088_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4584_ _9301_/Q _7425_/A _5842_/S input49/X _4583_/X VGND VGND VPWR VPWR _4590_/B
+ sky130_fd_sc_hd__a221o_1
Xinput73 pad_flash_io0_di VGND VGND VPWR VPWR _5179_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_9111_ _5235__1/A _9111_/D _7012_/X VGND VGND VPWR VPWR _9111_/Q sky130_fd_sc_hd__dfrtn_1
Xhold813 _5923_/X VGND VGND VPWR VPWR _5924_/A sky130_fd_sc_hd__dlygate4sd3_1
Xinput84 spimemio_flash_csb VGND VGND VPWR VPWR input84/X sky130_fd_sc_hd__buf_2
Xinput95 sram_ro_data[11] VGND VGND VPWR VPWR input95/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6323_ _6334_/B _6800_/A VGND VGND VPWR VPWR _6869_/C sky130_fd_sc_hd__nor2_1
Xhold824 _9270_/Q VGND VGND VPWR VPWR hold824/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold835 _7404_/X VGND VGND VPWR VPWR _7405_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 hold846/A VGND VGND VPWR VPWR hold846/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 _9108_/Q VGND VGND VPWR VPWR hold857/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9042_ _9541_/CLK _9042_/D VGND VGND VPWR VPWR _9042_/Q sky130_fd_sc_hd__dfxtp_1
Xhold868 hold868/A VGND VGND VPWR VPWR _7138_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold879 _7607_/X VGND VGND VPWR VPWR _7608_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6254_ _6254_/A VGND VGND VPWR VPWR _6610_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_131_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5205_ _9002_/Q _5067_/B _8797_/Q VGND VGND VPWR VPWR _5206_/A sky130_fd_sc_hd__mux2_1
X_6185_ _6398_/B _6317_/B _6419_/A _6633_/A VGND VGND VPWR VPWR _6344_/B sky130_fd_sc_hd__a2bb2o_1
X_5136_ _9488_/Q _9489_/Q VGND VGND VPWR VPWR _7860_/A sky130_fd_sc_hd__nor2_1
X_5067_ _8808_/Q _5067_/B _5068_/C VGND VGND VPWR VPWR _5067_/X sky130_fd_sc_hd__and3_1
XFILLER_38_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8826_ _9474_/CLK _8826_/D fanout427/X VGND VGND VPWR VPWR _8826_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8757_ _8756_/X _8757_/A1 _8765_/S VGND VGND VPWR VPWR _8758_/A sky130_fd_sc_hd__mux2_1
X_5969_ _5969_/A VGND VGND VPWR VPWR _9056_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7708_ _5410_/X hold188/X _7710_/S VGND VGND VPWR VPWR _7708_/X sky130_fd_sc_hd__mux2_1
X_8688_ _8688_/A _8688_/B _8688_/C _8688_/D VGND VGND VPWR VPWR _8701_/B sky130_fd_sc_hd__or4_1
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7639_ _7639_/A VGND VGND VPWR VPWR _9391_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9309_ _9469_/CLK _9309_/D fanout458/X VGND VGND VPWR VPWR _9309_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_181_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold109 _9313_/Q VGND VGND VPWR VPWR hold109/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7990_ _7990_/A VGND VGND VPWR VPWR _7990_/X sky130_fd_sc_hd__buf_8
XFILLER_94_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6941_ _7000_/B _6941_/B _6958_/B VGND VGND VPWR VPWR _6942_/B sky130_fd_sc_hd__or3_1
XFILLER_35_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6872_ _6872_/A _6872_/B _6872_/C _6872_/D VGND VGND VPWR VPWR _6935_/C sky130_fd_sc_hd__or4_1
XFILLER_179_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8611_ _9100_/Q _8372_/A _8369_/A _8904_/Q _8610_/X VGND VGND VPWR VPWR _8611_/X
+ sky130_fd_sc_hd__a221o_1
X_5823_ _5823_/A VGND VGND VPWR VPWR _5823_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8542_ _9238_/Q _8322_/X _8333_/X _9270_/Q _8541_/X VGND VGND VPWR VPWR _8549_/A
+ sky130_fd_sc_hd__a221o_1
X_5754_ _5754_/A VGND VGND VPWR VPWR _8959_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4705_ _9467_/Q _7798_/A _7571_/A _9363_/Q VGND VGND VPWR VPWR _4705_/X sky130_fd_sc_hd__a22o_1
X_8473_ _8473_/A _8473_/B _8473_/C _8473_/D VGND VGND VPWR VPWR _8474_/D sky130_fd_sc_hd__or4_1
X_5685_ _5685_/A VGND VGND VPWR VPWR _8930_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7424_ _7424_/A VGND VGND VPWR VPWR _9295_/D sky130_fd_sc_hd__clkbuf_1
X_4636_ _9300_/Q _7425_/A _5773_/A _8972_/Q VGND VGND VPWR VPWR _4636_/X sky130_fd_sc_hd__a22o_1
XFILLER_135_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold610 _8905_/Q VGND VGND VPWR VPWR hold610/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_118_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold621 _9394_/Q VGND VGND VPWR VPWR hold621/X sky130_fd_sc_hd__dlygate4sd3_1
X_7355_ _7355_/A VGND VGND VPWR VPWR _9263_/D sky130_fd_sc_hd__clkbuf_1
X_4567_ _9285_/Q _7391_/A _7481_/A _9325_/Q VGND VGND VPWR VPWR _4567_/X sky130_fd_sc_hd__a22o_1
XFILLER_162_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold632 _7209_/X VGND VGND VPWR VPWR _7210_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold643 _9423_/Q VGND VGND VPWR VPWR hold643/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap362 _4458_/Y VGND VGND VPWR VPWR _7356_/A sky130_fd_sc_hd__buf_6
Xhold654 _7779_/X VGND VGND VPWR VPWR _7780_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6306_ _6858_/B _6435_/A VGND VGND VPWR VPWR _6948_/B sky130_fd_sc_hd__nor2_2
Xhold665 _9391_/Q VGND VGND VPWR VPWR hold665/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap384 _4419_/Y VGND VGND VPWR VPWR _7571_/A sky130_fd_sc_hd__buf_6
Xhold676 _9198_/Q VGND VGND VPWR VPWR hold676/X sky130_fd_sc_hd__dlygate4sd3_1
X_7286_ _7286_/A VGND VGND VPWR VPWR _9232_/D sky130_fd_sc_hd__clkbuf_1
X_4498_ _4748_/B _4667_/A VGND VGND VPWR VPWR _7321_/A sky130_fd_sc_hd__nor2_8
XFILLER_104_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold687 hold687/A VGND VGND VPWR VPWR _7274_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap395 _6345_/A VGND VGND VPWR VPWR _6795_/A sky130_fd_sc_hd__clkbuf_2
Xhold698 _7106_/X VGND VGND VPWR VPWR _7107_/A sky130_fd_sc_hd__dlygate4sd3_1
X_9025_ _9551_/CLK _9025_/D fanout499/X VGND VGND VPWR VPWR _9025_/Q sky130_fd_sc_hd__dfstp_1
X_6237_ _6237_/A VGND VGND VPWR VPWR _6279_/A sky130_fd_sc_hd__clkbuf_4
X_6168_ _6168_/A VGND VGND VPWR VPWR _6633_/A sky130_fd_sc_hd__buf_2
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5119_ _6079_/C _6079_/D _6078_/A _6078_/B VGND VGND VPWR VPWR _5120_/D sky130_fd_sc_hd__or4_1
XFILLER_85_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6099_ _6732_/A _6724_/A _6724_/B VGND VGND VPWR VPWR _6228_/A sky130_fd_sc_hd__or3_2
XFILLER_45_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A VGND VGND VPWR VPWR _9529_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_53_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8809_ _9480_/CLK _8809_/D fanout414/X VGND VGND VPWR VPWR _8809_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_43_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5470_ _5470_/A VGND VGND VPWR VPWR _8838_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4421_ _9343_/Q _4414_/Y _7605_/A _9383_/Q _4420_/X VGND VGND VPWR VPWR _4431_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_172_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7140_ _7128_/X _9168_/Q _7142_/S VGND VGND VPWR VPWR _7140_/X sky130_fd_sc_hd__mux2_1
X_4352_ hold29/X hold22/X _4351_/X VGND VGND VPWR VPWR hold30/A sky130_fd_sc_hd__a21oi_1
XFILLER_172_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout408 fanout410/X VGND VGND VPWR VPWR fanout408/X sky130_fd_sc_hd__clkbuf_4
X_7071_ _7071_/A VGND VGND VPWR VPWR _9138_/D sky130_fd_sc_hd__clkbuf_1
Xfanout419 fanout426/X VGND VGND VPWR VPWR fanout419/X sky130_fd_sc_hd__clkbuf_4
X_6022_ hold884/X _5761_/X _6030_/S VGND VGND VPWR VPWR _6023_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7973_ _7973_/A VGND VGND VPWR VPWR _7973_/X sky130_fd_sc_hd__buf_6
XFILLER_81_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6924_ _6976_/C _6924_/B _6924_/C _6924_/D VGND VGND VPWR VPWR _6988_/B sky130_fd_sc_hd__or4_1
XFILLER_35_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6855_ _6850_/A _6818_/A _6862_/B _6158_/B _6435_/A VGND VGND VPWR VPWR _6855_/X
+ sky130_fd_sc_hd__o32a_1
X_5806_ _5806_/A _7132_/B VGND VGND VPWR VPWR _5816_/S sky130_fd_sc_hd__and2_2
XFILLER_168_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9574_ _9574_/A _5094_/Y VGND VGND VPWR VPWR mgmt_gpio_out[20] sky130_fd_sc_hd__ebufn_8
XFILLER_167_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6786_ _6931_/A _6786_/B VGND VGND VPWR VPWR _6786_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8525_ _8701_/A _8525_/B _8525_/C VGND VGND VPWR VPWR _8525_/X sky130_fd_sc_hd__or3_1
XFILLER_148_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5737_ _5737_/A VGND VGND VPWR VPWR _8952_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8456_ _9371_/Q _8346_/X _8386_/X _9347_/Q VGND VGND VPWR VPWR _8456_/X sky130_fd_sc_hd__a22o_1
XFILLER_108_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5668_ _5629_/X hold847/X _5676_/S VGND VGND VPWR VPWR _5669_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7407_ _7407_/A VGND VGND VPWR VPWR _9287_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4619_ input48/X _4582_/A _5693_/A _8937_/Q VGND VGND VPWR VPWR _4619_/X sky130_fd_sc_hd__a22o_1
XFILLER_136_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8387_ _9192_/Q _8384_/X _8386_/X _9344_/Q VGND VGND VPWR VPWR _8387_/X sky130_fd_sc_hd__a22o_1
X_5599_ hold522/X _5587_/X _5605_/S VGND VGND VPWR VPWR _5600_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold440 _7291_/X VGND VGND VPWR VPWR _7292_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7338_ _7338_/A VGND VGND VPWR VPWR _9255_/D sky130_fd_sc_hd__clkbuf_1
Xhold451 _5472_/X VGND VGND VPWR VPWR _5473_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 _8773_/Q VGND VGND VPWR VPWR hold462/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold473 _8865_/Q VGND VGND VPWR VPWR hold473/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 _6024_/X VGND VGND VPWR VPWR _6025_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold495 hold495/A VGND VGND VPWR VPWR hold495/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7269_ _7147_/X hold134/X _7282_/S VGND VGND VPWR VPWR _7270_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9008_ _9532_/CLK _9008_/D fanout503/X VGND VGND VPWR VPWR hold73/A sky130_fd_sc_hd__dfrtp_4
XFILLER_38_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1140 _9426_/Q VGND VGND VPWR VPWR hold418/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1151 _8954_/Q VGND VGND VPWR VPWR hold850/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1162 _8784_/Q VGND VGND VPWR VPWR hold23/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1173 _9308_/Q VGND VGND VPWR VPWR hold326/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1184 _9366_/Q VGND VGND VPWR VPWR hold777/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_302 _4898_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1195 _9300_/Q VGND VGND VPWR VPWR hold288/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_313 hold5/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_324 _9427_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_335 _5315_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_346 _7147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_357 _8002_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_368 _9071_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_379 input33/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4970_ _5068_/B _4972_/B _4970_/B1 VGND VGND VPWR VPWR _4971_/B sky130_fd_sc_hd__a21oi_1
XFILLER_51_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6640_ _6850_/B _6887_/B VGND VGND VPWR VPWR _6640_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6571_ _6340_/Y _6281_/A _6839_/B _6345_/X VGND VGND VPWR VPWR _6937_/B sky130_fd_sc_hd__a22o_1
XFILLER_118_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8310_ _8360_/A VGND VGND VPWR VPWR _8310_/X sky130_fd_sc_hd__buf_6
X_5522_ _5522_/A VGND VGND VPWR VPWR _8859_/D sky130_fd_sc_hd__clkbuf_1
X_9290_ _9290_/CLK _9290_/D fanout468/X VGND VGND VPWR VPWR _9290_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_145_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8241_ hold987/X _8196_/S _8239_/X _8240_/X VGND VGND VPWR VPWR _9517_/D sky130_fd_sc_hd__o22a_1
XFILLER_118_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5453_ _7158_/A _5453_/B _5453_/C _7158_/D VGND VGND VPWR VPWR _5454_/A sky130_fd_sc_hd__or4_2
XFILLER_173_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4404_ hold58/X hold52/X VGND VGND VPWR VPWR _4405_/A sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_42_csclk _8954_/CLK VGND VGND VPWR VPWR _9167_/CLK sky130_fd_sc_hd__clkbuf_16
X_8172_ _9191_/Q _8010_/B _8162_/X _8171_/X _8627_/S VGND VGND VPWR VPWR _8172_/X
+ sky130_fd_sc_hd__o221a_2
X_5384_ _5384_/A VGND VGND VPWR VPWR _5384_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_160_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7123_ _7123_/A VGND VGND VPWR VPWR _7123_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7054_ _5465_/X _9131_/Q _7054_/S VGND VGND VPWR VPWR _7054_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6005_ hold609/X _5690_/X _6005_/S VGND VGND VPWR VPWR _6006_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_57_csclk _9090_/CLK VGND VGND VPWR VPWR _9051_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7956_ _7956_/A VGND VGND VPWR VPWR _8023_/B sky130_fd_sc_hd__buf_8
XFILLER_42_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6907_ _6824_/A _6907_/B _6907_/C VGND VGND VPWR VPWR _6978_/B sky130_fd_sc_hd__and3b_1
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7887_ _8275_/B _7887_/B VGND VGND VPWR VPWR _7887_/Y sky130_fd_sc_hd__nand2_1
X_6838_ _6838_/A _6838_/B VGND VGND VPWR VPWR _6841_/C sky130_fd_sc_hd__nor2_1
XFILLER_24_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9557_ _9557_/A _5111_/Y VGND VGND VPWR VPWR mgmt_gpio_out[3] sky130_fd_sc_hd__ebufn_8
XFILLER_149_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6769_ _7001_/A _6768_/Y _6433_/C VGND VGND VPWR VPWR _7006_/B sky130_fd_sc_hd__o21ba_1
XFILLER_7_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8508_ _9333_/Q _8298_/X _8370_/X _9253_/Q VGND VGND VPWR VPWR _8508_/X sky130_fd_sc_hd__a22o_1
X_9488_ _9529_/CLK _9488_/D fanout440/X VGND VGND VPWR VPWR _9488_/Q sky130_fd_sc_hd__dfrtp_2
X_8439_ _9218_/Q _8391_/X _8367_/X _9474_/Q _8438_/X VGND VGND VPWR VPWR _8439_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_136_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold270 hold270/A VGND VGND VPWR VPWR hold270/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 _7154_/X VGND VGND VPWR VPWR _7155_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 _7758_/X VGND VGND VPWR VPWR _7759_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_110 _6015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_121 _6262_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_132 _7645_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_143 _7984_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_154 _7940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 _8023_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_176 _7969_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_187 _7993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_198 _8001_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput5 mask_rev_in[10] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_1
X_7810_ _7810_/A VGND VGND VPWR VPWR _9469_/D sky130_fd_sc_hd__clkbuf_1
X_8790_ _5168_/A1 _8790_/D _5346_/X VGND VGND VPWR VPWR _8790_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7741_ _7741_/A VGND VGND VPWR VPWR _9437_/D sky130_fd_sc_hd__clkbuf_1
X_4953_ _9392_/Q _4389_/Y _5607_/A _8898_/Q _4952_/X VGND VGND VPWR VPWR _4960_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7672_ _7654_/X hold225/X _7676_/S VGND VGND VPWR VPWR _7672_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4884_ _4884_/A _4884_/B _4884_/C _4884_/D VGND VGND VPWR VPWR _4885_/C sky130_fd_sc_hd__or4_1
XFILLER_177_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9411_ _9475_/CLK _9411_/D fanout480/X VGND VGND VPWR VPWR _9411_/Q sky130_fd_sc_hd__dfrtp_4
X_6623_ _6623_/A _6967_/A VGND VGND VPWR VPWR _6623_/Y sky130_fd_sc_hd__nor2_2
XFILLER_20_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9342_ _9398_/CLK _9342_/D _5070_/A VGND VGND VPWR VPWR _9342_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_165_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6554_ _6281_/A _6328_/Y _6330_/Y VGND VGND VPWR VPWR _6935_/B sky130_fd_sc_hd__a21o_1
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5505_ _5761_/A VGND VGND VPWR VPWR _5505_/X sky130_fd_sc_hd__clkbuf_4
X_9273_ _9305_/CLK _9273_/D fanout467/X VGND VGND VPWR VPWR _9273_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_173_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6485_ _6811_/B _6811_/C _6441_/B _6543_/B VGND VGND VPWR VPWR _6486_/A sky130_fd_sc_hd__a31o_1
XFILLER_118_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8224_ _8960_/Q _8224_/B VGND VGND VPWR VPWR _8224_/X sky130_fd_sc_hd__and2_1
X_5436_ _5436_/A VGND VGND VPWR VPWR _8824_/D sky130_fd_sc_hd__clkbuf_1
Xoutput320 _9151_/Q VGND VGND VPWR VPWR sram_ro_addr[4] sky130_fd_sc_hd__buf_12
Xoutput331 _9058_/Q VGND VGND VPWR VPWR wb_dat_o[13] sky130_fd_sc_hd__buf_12
XFILLER_160_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput342 _9047_/Q VGND VGND VPWR VPWR wb_dat_o[23] sky130_fd_sc_hd__buf_12
Xoutput353 _9065_/Q VGND VGND VPWR VPWR wb_dat_o[4] sky130_fd_sc_hd__buf_12
X_8155_ _9287_/Q _7953_/B _8003_/X _9303_/Q VGND VGND VPWR VPWR _8155_/X sky130_fd_sc_hd__a22o_2
X_5367_ _5375_/A _5378_/B VGND VGND VPWR VPWR _5368_/A sky130_fd_sc_hd__and2_1
XFILLER_99_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7106_ _5471_/X _9154_/Q _7106_/S VGND VGND VPWR VPWR _7106_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8086_ _9404_/Q _7931_/X _7933_/X _9340_/Q VGND VGND VPWR VPWR _8086_/X sky130_fd_sc_hd__a22o_1
X_5298_ _5298_/A VGND VGND VPWR VPWR _8772_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7037_ _6012_/X _9123_/Q _7041_/S VGND VGND VPWR VPWR _7037_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8988_ _9178_/CLK _8988_/D fanout486/X VGND VGND VPWR VPWR _9570_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_27_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7939_ _8206_/B _7991_/B _8000_/B VGND VGND VPWR VPWR _7940_/A sky130_fd_sc_hd__and3_2
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6270_ _6802_/A _6790_/A VGND VGND VPWR VPWR _6272_/C sky130_fd_sc_hd__or2_1
XFILLER_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5221_ _5221_/A VGND VGND VPWR VPWR _5221_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5152_ _8778_/Q _5151_/Y _5068_/C _5016_/B hold949/X VGND VGND VPWR VPWR _5152_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_110_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5083_ _9435_/Q VGND VGND VPWR VPWR _5083_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8911_ _9051_/CLK _8911_/D fanout453/X VGND VGND VPWR VPWR _8911_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_37_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8842_ _9178_/CLK _8842_/D fanout486/X VGND VGND VPWR VPWR _8842_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_52_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8773_ _9162_/CLK _8773_/D fanout438/X VGND VGND VPWR VPWR _8773_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_52_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5985_ _5985_/A VGND VGND VPWR VPWR _9063_/D sky130_fd_sc_hd__clkbuf_1
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7724_ _7724_/A VGND VGND VPWR VPWR _9429_/D sky130_fd_sc_hd__clkbuf_1
X_4936_ _9132_/Q _7056_/A _6021_/A _9079_/Q _4935_/X VGND VGND VPWR VPWR _4939_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_52_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_10 _7081_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7655_ _7654_/X hold241/X hold84/X VGND VGND VPWR VPWR _7656_/A sky130_fd_sc_hd__mux2_1
X_4867_ _9148_/Q _7091_/A _5704_/A _8939_/Q VGND VGND VPWR VPWR _4867_/X sky130_fd_sc_hd__a22o_2
XANTENNA_21 _4460_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_32 _5727_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_43 _4741_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_54 _4885_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6606_ _6244_/X _6610_/A _6125_/A _6401_/A VGND VGND VPWR VPWR _6607_/B sky130_fd_sc_hd__o22a_1
XFILLER_193_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7586_ _7514_/X hold646/X hold78/X VGND VGND VPWR VPWR _7586_/X sky130_fd_sc_hd__mux2_1
XANTENNA_65 _5067_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 hold20/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4798_ _8925_/Q _5667_/A _5918_/A _9037_/Q VGND VGND VPWR VPWR _4798_/X sky130_fd_sc_hd__a22o_1
XANTENNA_87 _5465_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_98 _5809_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9325_ _9325_/CLK _9325_/D fanout460/X VGND VGND VPWR VPWR _9325_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_153_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6537_ _6906_/B _6781_/B _6655_/C _6898_/A _6748_/B VGND VGND VPWR VPWR _6537_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_21_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9256_ _9328_/CLK _9256_/D fanout463/X VGND VGND VPWR VPWR _9256_/Q sky130_fd_sc_hd__dfstp_2
X_6468_ _6468_/A _6468_/B _6468_/C _6468_/D VGND VGND VPWR VPWR _6469_/D sky130_fd_sc_hd__or4_1
XFILLER_133_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8207_ _8773_/Q _7977_/X _8206_/X _7983_/A VGND VGND VPWR VPWR _8207_/X sky130_fd_sc_hd__a22o_1
XFILLER_106_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5419_ _5419_/A VGND VGND VPWR VPWR _5435_/S sky130_fd_sc_hd__clkbuf_4
X_9187_ _9187_/CLK _9187_/D fanout456/X VGND VGND VPWR VPWR _9187_/Q sky130_fd_sc_hd__dfrtp_4
X_6399_ _6399_/A _6818_/A VGND VGND VPWR VPWR _6887_/A sky130_fd_sc_hd__or2_2
XFILLER_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8138_ _9398_/Q _7977_/A _8137_/X _7983_/A VGND VGND VPWR VPWR _8138_/X sky130_fd_sc_hd__a22o_1
XFILLER_99_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8069_ _9403_/Q _7931_/X _7933_/X _9339_/Q _8068_/X VGND VGND VPWR VPWR _8072_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_75_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5770_ _5770_/A VGND VGND VPWR VPWR _8966_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4721_ _8986_/Q _5806_/A _5630_/A _8911_/Q VGND VGND VPWR VPWR _4721_/X sky130_fd_sc_hd__a22o_1
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7440_ _7439_/X hold311/X _7444_/S VGND VGND VPWR VPWR _7440_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4652_ _4665_/A _4667_/B VGND VGND VPWR VPWR _5715_/A sky130_fd_sc_hd__nor2_8
XFILLER_147_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput30 mask_rev_in[4] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7371_ _7371_/A VGND VGND VPWR VPWR _9270_/D sky130_fd_sc_hd__clkbuf_1
Xinput41 mgmt_gpio_in[14] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__clkbuf_4
XFILLER_162_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput52 mgmt_gpio_in[24] VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4583_ _9333_/Q _7499_/A _7605_/A _9381_/Q VGND VGND VPWR VPWR _4583_/X sky130_fd_sc_hd__a22o_1
Xinput63 mgmt_gpio_in[34] VGND VGND VPWR VPWR _5279_/A sky130_fd_sc_hd__buf_4
Xhold803 hold803/A VGND VGND VPWR VPWR _7143_/A sky130_fd_sc_hd__dlygate4sd3_1
X_9110_ _9110_/CLK _9110_/D fanout503/X VGND VGND VPWR VPWR _9110_/Q sky130_fd_sc_hd__dfrtp_4
Xinput74 pad_flash_io1_di VGND VGND VPWR VPWR _5181_/B sky130_fd_sc_hd__clkbuf_1
Xhold814 _9176_/Q VGND VGND VPWR VPWR hold814/X sky130_fd_sc_hd__dlygate4sd3_1
X_6322_ _6334_/B _6624_/B VGND VGND VPWR VPWR _6959_/B sky130_fd_sc_hd__nor2_1
Xhold825 _7370_/X VGND VGND VPWR VPWR _7371_/A sky130_fd_sc_hd__dlygate4sd3_1
Xinput85 spimemio_flash_io0_do VGND VGND VPWR VPWR input85/X sky130_fd_sc_hd__buf_2
Xinput96 sram_ro_data[12] VGND VGND VPWR VPWR input96/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold836 _9302_/Q VGND VGND VPWR VPWR hold836/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 hold847/A VGND VGND VPWR VPWR hold847/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 _7229_/X VGND VGND VPWR VPWR _7230_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9041_ _9541_/CLK _9041_/D VGND VGND VPWR VPWR _9041_/Q sky130_fd_sc_hd__dfxtp_1
Xhold869 hold869/A VGND VGND VPWR VPWR hold869/X sky130_fd_sc_hd__dlygate4sd3_1
X_6253_ _6589_/C _6311_/B VGND VGND VPWR VPWR _6254_/A sky130_fd_sc_hd__or2_1
XFILLER_131_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5204_ _5204_/A VGND VGND VPWR VPWR _5204_/X sky130_fd_sc_hd__clkbuf_1
X_6184_ _6850_/A _6850_/B VGND VGND VPWR VPWR _6419_/A sky130_fd_sc_hd__nor2_8
XFILLER_97_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5135_ _8355_/A _8380_/A VGND VGND VPWR VPWR _5135_/X sky130_fd_sc_hd__or2_2
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5066_ _5066_/A VGND VGND VPWR VPWR _8781_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8825_ _9474_/CLK _8825_/D fanout427/X VGND VGND VPWR VPWR _8825_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_25_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8756_ _5271_/A _8756_/A2 _8756_/B1 _8727_/Y _8755_/X VGND VGND VPWR VPWR _8756_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_52_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5968_ _9056_/Q _4752_/X _5976_/S VGND VGND VPWR VPWR _5969_/A sky130_fd_sc_hd__mux2_1
X_4919_ _9472_/Q _7815_/A _5418_/A _8817_/Q VGND VGND VPWR VPWR _4919_/X sky130_fd_sc_hd__a22o_1
X_7707_ _7707_/A VGND VGND VPWR VPWR _9421_/D sky130_fd_sc_hd__clkbuf_1
X_5899_ _5899_/A VGND VGND VPWR VPWR _9016_/D sky130_fd_sc_hd__clkbuf_1
X_8687_ _9103_/Q _8372_/X _8369_/X _8907_/Q _8686_/X VGND VGND VPWR VPWR _8688_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7638_ _7514_/X hold665/X _7638_/S VGND VGND VPWR VPWR _7638_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7569_ _7514_/X hold841/X hold99/A VGND VGND VPWR VPWR _7570_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9308_ _9420_/CLK _9308_/D fanout465/X VGND VGND VPWR VPWR _9308_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9239_ _9398_/CLK _9239_/D fanout419/X VGND VGND VPWR VPWR _9239_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6940_ _6795_/A _6507_/A _6314_/C _6798_/D _6939_/Y VGND VGND VPWR VPWR _6958_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_66_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6871_ _6873_/B _6871_/B VGND VGND VPWR VPWR _6872_/A sky130_fd_sc_hd__nor2_1
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8610_ _8884_/Q _8354_/B _8331_/A _8979_/Q VGND VGND VPWR VPWR _8610_/X sky130_fd_sc_hd__a22o_1
X_5822_ _9570_/A _5818_/X hold43/X VGND VGND VPWR VPWR _5822_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8541_ _9286_/Q _8316_/X _8327_/X _9262_/Q VGND VGND VPWR VPWR _8541_/X sky130_fd_sc_hd__a22o_1
X_5753_ hold467/X _5587_/X _5759_/S VGND VGND VPWR VPWR _5754_/A sky130_fd_sc_hd__mux2_1
X_4704_ _4704_/A1 _4502_/Y _5388_/A _8812_/Q _4703_/X VGND VGND VPWR VPWR _4711_/A
+ sky130_fd_sc_hd__a221o_1
X_8472_ _9379_/Q _8337_/A _8384_/A _9195_/Q _8471_/X VGND VGND VPWR VPWR _8473_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5684_ hold605/X _5683_/X _5691_/S VGND VGND VPWR VPWR _5685_/A sky130_fd_sc_hd__mux2_1
X_7423_ _7299_/X hold530/X _7423_/S VGND VGND VPWR VPWR _7423_/X sky130_fd_sc_hd__mux2_1
X_4635_ _4635_/A _4685_/B VGND VGND VPWR VPWR _5773_/A sky130_fd_sc_hd__nor2_8
XFILLER_147_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold600 hold600/A VGND VGND VPWR VPWR hold600/X sky130_fd_sc_hd__dlygate4sd3_1
X_7354_ _7299_/X hold691/X _7354_/S VGND VGND VPWR VPWR _7354_/X sky130_fd_sc_hd__mux2_1
Xhold611 _8846_/Q VGND VGND VPWR VPWR hold611/X sky130_fd_sc_hd__dlygate4sd3_1
X_4566_ _9189_/Q _7176_/A _4477_/Y input31/X _4565_/X VGND VGND VPWR VPWR _4569_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold622 hold622/A VGND VGND VPWR VPWR hold622/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_118_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold633 _9482_/Q VGND VGND VPWR VPWR hold633/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 _7710_/X VGND VGND VPWR VPWR _7711_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6305_ _6461_/A VGND VGND VPWR VPWR _6435_/A sky130_fd_sc_hd__buf_4
XFILLER_150_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap363 _4454_/Y VGND VGND VPWR VPWR _7266_/A sky130_fd_sc_hd__buf_8
X_7285_ _7128_/X hold893/X _7300_/S VGND VGND VPWR VPWR _7286_/A sky130_fd_sc_hd__mux2_1
Xhold655 _9431_/Q VGND VGND VPWR VPWR hold655/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap374 _7832_/A VGND VGND VPWR VPWR _4898_/A2 sky130_fd_sc_hd__buf_8
X_4497_ _4748_/B _4499_/A VGND VGND VPWR VPWR _5388_/A sky130_fd_sc_hd__nor2_8
Xhold666 _7638_/X VGND VGND VPWR VPWR _7639_/A sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap385 _4416_/Y VGND VGND VPWR VPWR _7211_/A sky130_fd_sc_hd__buf_8
Xhold677 _7207_/X VGND VGND VPWR VPWR _7208_/A sky130_fd_sc_hd__dlygate4sd3_1
X_9024_ _9172_/CLK _9024_/D fanout492/X VGND VGND VPWR VPWR _9585_/A sky130_fd_sc_hd__dfrtp_1
Xhold688 _7237_/X VGND VGND VPWR VPWR _7238_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold699 hold699/A VGND VGND VPWR VPWR _7416_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6236_ _6317_/A _6906_/A VGND VGND VPWR VPWR _6237_/A sky130_fd_sc_hd__or2_1
XFILLER_131_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6167_ _6167_/A _6167_/B _6167_/C VGND VGND VPWR VPWR _6168_/A sky130_fd_sc_hd__and3_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _6078_/C _6078_/D _5118_/C input148/X VGND VGND VPWR VPWR _5120_/C sky130_fd_sc_hd__or4b_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6098_ _6175_/A _6095_/B _6097_/Y VGND VGND VPWR VPWR _6724_/B sky130_fd_sc_hd__a21oi_1
XFILLER_85_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5049_ _5047_/Y _5045_/Y _5048_/X VGND VGND VPWR VPWR _8789_/D sky130_fd_sc_hd__a21oi_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8808_ _5168_/A1 _8808_/D _5386_/X VGND VGND VPWR VPWR _8808_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_13_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8739_ _5287_/A _8739_/A2 _8739_/B1 _5275_/A VGND VGND VPWR VPWR _8739_/X sky130_fd_sc_hd__a22o_1
XFILLER_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4420_ _9207_/Q _7211_/A _7571_/A _9367_/Q VGND VGND VPWR VPWR _4420_/X sky130_fd_sc_hd__a22o_1
XFILLER_144_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4351_ _8805_/Q _5021_/B VGND VGND VPWR VPWR _4351_/X sky130_fd_sc_hd__and2_1
XFILLER_160_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout409 fanout410/X VGND VGND VPWR VPWR fanout409/X sky130_fd_sc_hd__clkbuf_4
X_7070_ _9138_/Q _7494_/A _7072_/S VGND VGND VPWR VPWR _7070_/X sky130_fd_sc_hd__mux2_1
X_6021_ _6021_/A _7132_/B VGND VGND VPWR VPWR _6030_/S sky130_fd_sc_hd__and2_2
XFILLER_86_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_1_csclk clkbuf_1_1_1_csclk/A VGND VGND VPWR VPWR clkbuf_2_3_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_140_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7972_ _8206_/B _7984_/C _7992_/C VGND VGND VPWR VPWR _7973_/A sky130_fd_sc_hd__and3_4
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6923_ _6923_/A _6982_/C VGND VGND VPWR VPWR _6923_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6854_ _6950_/B _6950_/C _6993_/C _6944_/C VGND VGND VPWR VPWR _6854_/X sky130_fd_sc_hd__or4_1
XFILLER_50_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5805_ _5805_/A VGND VGND VPWR VPWR _8982_/D sky130_fd_sc_hd__clkbuf_1
X_9573_ _9573_/A _5095_/Y VGND VGND VPWR VPWR mgmt_gpio_out[19] sky130_fd_sc_hd__ebufn_8
X_6785_ _6785_/A _6785_/B VGND VGND VPWR VPWR _6786_/B sky130_fd_sc_hd__nor2_1
XFILLER_10_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8524_ _8524_/A _8524_/B _8524_/C _8524_/D VGND VGND VPWR VPWR _8525_/C sky130_fd_sc_hd__or4_1
X_5736_ _5653_/X hold123/X _5736_/S VGND VGND VPWR VPWR _5736_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5667_ _5667_/A _5693_/B VGND VGND VPWR VPWR _5676_/S sky130_fd_sc_hd__nand2_2
X_8455_ _9419_/Q _8402_/X _8378_/X _9355_/Q _8454_/X VGND VGND VPWR VPWR _8455_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4618_ _4665_/A _4685_/B VGND VGND VPWR VPWR _5693_/A sky130_fd_sc_hd__nor2_8
X_7406_ _7299_/X hold694/X _7406_/S VGND VGND VPWR VPWR _7406_/X sky130_fd_sc_hd__mux2_1
X_8386_ _8386_/A VGND VGND VPWR VPWR _8386_/X sky130_fd_sc_hd__buf_6
X_5598_ _5598_/A VGND VGND VPWR VPWR _8893_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7337_ hold207/X _7514_/A _7337_/S VGND VGND VPWR VPWR _7337_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold430 hold430/A VGND VGND VPWR VPWR _7399_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold441 _5904_/X VGND VGND VPWR VPWR _5905_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4549_ _4549_/A _4549_/B _4549_/C _4549_/D VGND VGND VPWR VPWR _4549_/X sky130_fd_sc_hd__or4_4
Xhold452 _5393_/X VGND VGND VPWR VPWR _5394_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 _8859_/Q VGND VGND VPWR VPWR hold463/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold474 _5534_/X VGND VGND VPWR VPWR _5535_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7268_ _7268_/A VGND VGND VPWR VPWR _9224_/D sky130_fd_sc_hd__clkbuf_1
Xhold485 hold485/A VGND VGND VPWR VPWR hold485/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold496 _9474_/Q VGND VGND VPWR VPWR hold496/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9007_ _9172_/CLK _9007_/D fanout490/X VGND VGND VPWR VPWR _9007_/Q sky130_fd_sc_hd__dfrtp_1
X_6219_ _6219_/A VGND VGND VPWR VPWR _6790_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_89_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7199_ _6012_/X hold800/X _7209_/S VGND VGND VPWR VPWR _7199_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1130 _8884_/Q VGND VGND VPWR VPWR hold529/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1141 _9284_/Q VGND VGND VPWR VPWR hold285/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1152 _8882_/Q VGND VGND VPWR VPWR hold664/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1163 _7563_/X VGND VGND VPWR VPWR _7564_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1174 _9210_/Q VGND VGND VPWR VPWR hold865/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1185 _9346_/Q VGND VGND VPWR VPWR hold718/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1196 _8938_/Q VGND VGND VPWR VPWR hold903/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_303 _4898_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_314 hold15/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_325 _4531_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_336 _5387_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_347 _7147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_358 _7953_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_369 _9245_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6570_ _6851_/A _6759_/A VGND VGND VPWR VPWR _6882_/C sky130_fd_sc_hd__or2_1
X_5521_ _5301_/X hold463/X _5527_/S VGND VGND VPWR VPWR _5521_/X sky130_fd_sc_hd__mux2_1
X_8240_ _5139_/A hold978/X _8013_/X VGND VGND VPWR VPWR _8240_/X sky130_fd_sc_hd__a21o_1
XFILLER_117_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5452_ hold18/X _5413_/S hold104/X VGND VGND VPWR VPWR _5452_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_145_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4403_ hold82/X hold51/X VGND VGND VPWR VPWR hold52/A sky130_fd_sc_hd__or2_1
XFILLER_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8171_ _8171_/A _8171_/B _8171_/C _8171_/D VGND VGND VPWR VPWR _8171_/X sky130_fd_sc_hd__or4_1
X_5383_ _7011_/A _7013_/B VGND VGND VPWR VPWR _5384_/A sky130_fd_sc_hd__and2_1
XFILLER_99_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7122_ _5468_/X _9161_/Q _7124_/S VGND VGND VPWR VPWR _7122_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7053_ _7053_/A VGND VGND VPWR VPWR _9130_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6004_ _6004_/A VGND VGND VPWR VPWR _9072_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7955_ _8181_/B _7989_/B _8002_/C VGND VGND VPWR VPWR _7956_/A sky130_fd_sc_hd__and3_4
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6906_ _6906_/A _6906_/B _6906_/C VGND VGND VPWR VPWR _6907_/C sky130_fd_sc_hd__or3_1
X_7886_ _8181_/B VGND VGND VPWR VPWR _8275_/B sky130_fd_sc_hd__buf_6
X_6837_ _6566_/B _6481_/A _6693_/Y _6694_/Y _6446_/X VGND VGND VPWR VPWR _6838_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_50_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9556_ _9556_/A _5112_/Y VGND VGND VPWR VPWR mgmt_gpio_out[2] sky130_fd_sc_hd__ebufn_8
XFILLER_10_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6768_ _6768_/A VGND VGND VPWR VPWR _6768_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8507_ _9373_/Q _8346_/X _8386_/X _9349_/Q _8506_/X VGND VGND VPWR VPWR _8512_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5719_ _5719_/A VGND VGND VPWR VPWR _8944_/D sky130_fd_sc_hd__clkbuf_1
X_9487_ _9487_/CLK _9487_/D fanout411/X VGND VGND VPWR VPWR _9487_/Q sky130_fd_sc_hd__dfrtp_1
X_6699_ _6230_/X _6563_/A _6689_/X _6763_/A _6698_/X VGND VGND VPWR VPWR _6700_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_40_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8438_ _9442_/Q _8398_/B _8344_/X _9482_/Q VGND VGND VPWR VPWR _8438_/X sky130_fd_sc_hd__a22o_1
XFILLER_156_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8369_ _8369_/A VGND VGND VPWR VPWR _8369_/X sky130_fd_sc_hd__buf_6
XFILLER_123_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold260 _9221_/Q VGND VGND VPWR VPWR hold260/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 _9293_/Q VGND VGND VPWR VPWR hold271/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 _7155_/X VGND VGND VPWR VPWR _9174_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold293 _9253_/Q VGND VGND VPWR VPWR hold293/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_100 _5809_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 _6015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 _6964_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_133 _7645_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_144 _7923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_155 _7940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_166 _8023_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_177 _8224_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_188 _7997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_199 _8001_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput6 mask_rev_in[11] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4952_ _8825_/Q _5437_/A _7027_/A _9119_/Q VGND VGND VPWR VPWR _4952_/X sky130_fd_sc_hd__a22o_1
X_7740_ _7654_/X hold178/X hold86/X VGND VGND VPWR VPWR _7740_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4883_ _4883_/A _4883_/B _4883_/C _4883_/D VGND VGND VPWR VPWR _4884_/D sky130_fd_sc_hd__or4_1
X_7671_ _7671_/A VGND VGND VPWR VPWR _9404_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9410_ _9467_/CLK _9410_/D fanout475/X VGND VGND VPWR VPWR _9410_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_177_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6622_ _6609_/A _6462_/B _6966_/C _6620_/X _6869_/B VGND VGND VPWR VPWR _6626_/C
+ sky130_fd_sc_hd__a2111o_1
X_9341_ _9469_/CLK _9341_/D fanout458/X VGND VGND VPWR VPWR _9341_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_118_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6553_ _6966_/A _6553_/B VGND VGND VPWR VPWR _6959_/C sky130_fd_sc_hd__or2_1
XFILLER_146_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5504_ _5504_/A VGND VGND VPWR VPWR _5761_/A sky130_fd_sc_hd__buf_8
X_9272_ _9272_/CLK _9272_/D fanout421/X VGND VGND VPWR VPWR _9272_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_118_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6484_ _6484_/A _6484_/B VGND VGND VPWR VPWR _6484_/X sky130_fd_sc_hd__or2_1
XFILLER_173_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5435_ _8824_/Q _5415_/X _5435_/S VGND VGND VPWR VPWR _5435_/X sky130_fd_sc_hd__mux2_1
X_8223_ _8890_/Q _8023_/B _7958_/X _9091_/Q _8222_/X VGND VGND VPWR VPWR _8228_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput310 _5231_/X VGND VGND VPWR VPWR serial_resetn sky130_fd_sc_hd__buf_12
Xoutput321 _9152_/Q VGND VGND VPWR VPWR sram_ro_addr[5] sky130_fd_sc_hd__buf_12
Xoutput332 _9059_/Q VGND VGND VPWR VPWR wb_dat_o[14] sky130_fd_sc_hd__buf_12
Xoutput343 _9534_/Q VGND VGND VPWR VPWR wb_dat_o[24] sky130_fd_sc_hd__buf_12
XFILLER_160_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5366_ _5366_/A VGND VGND VPWR VPWR _5366_/X sky130_fd_sc_hd__clkbuf_1
X_8154_ _9375_/Q _7960_/X _8001_/X _9271_/Q _8153_/X VGND VGND VPWR VPWR _8162_/A
+ sky130_fd_sc_hd__a221o_1
Xoutput354 _9066_/Q VGND VGND VPWR VPWR wb_dat_o[5] sky130_fd_sc_hd__buf_12
X_7105_ _7105_/A VGND VGND VPWR VPWR _9153_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8085_ hold974/X _8017_/X _8084_/X VGND VGND VPWR VPWR _8085_/X sky130_fd_sc_hd__o21a_1
XFILLER_113_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5297_ _5291_/X hold820/X _5316_/S VGND VGND VPWR VPWR _5297_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7036_ _7036_/A VGND VGND VPWR VPWR _9122_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_752 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8987_ _9089_/CLK _8987_/D fanout433/X VGND VGND VPWR VPWR _8987_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_15_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7938_ _7938_/A VGND VGND VPWR VPWR _7938_/X sky130_fd_sc_hd__buf_6
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7869_ _8996_/Q _7902_/B VGND VGND VPWR VPWR _7869_/Y sky130_fd_sc_hd__nor2_2
XFILLER_50_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9539_ _9541_/CLK _9539_/D VGND VGND VPWR VPWR _9539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _9251_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_61_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_56_csclk _9090_/CLK VGND VGND VPWR VPWR _9092_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_174_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5220_ _5219_/Y _8779_/Q _7025_/B VGND VGND VPWR VPWR _5221_/A sky130_fd_sc_hd__mux2_4
XFILLER_170_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5151_ _8780_/Q VGND VGND VPWR VPWR _5151_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5082_ _9443_/Q VGND VGND VPWR VPWR _5082_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8910_ _9184_/CLK _8910_/D fanout438/X VGND VGND VPWR VPWR _8910_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8841_ _9172_/CLK _8841_/D fanout493/X VGND VGND VPWR VPWR _8841_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8772_ _9484_/CLK _8772_/D fanout427/X VGND VGND VPWR VPWR _8772_/Q sky130_fd_sc_hd__dfrtp_4
X_5984_ _9063_/Q _4817_/X _5994_/S VGND VGND VPWR VPWR _5985_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7723_ _7654_/X hold252/X hold95/A VGND VGND VPWR VPWR _7723_/X sky130_fd_sc_hd__mux2_1
X_4935_ _8923_/Q _5667_/A _5693_/A _8933_/Q VGND VGND VPWR VPWR _4935_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_3_7_0_csclk clkbuf_3_7_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_7_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_11 _9144_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7654_ hold15/X VGND VGND VPWR VPWR _7654_/X sky130_fd_sc_hd__buf_4
XANTENNA_22 _4460_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4866_ _9313_/Q _7463_/A _6066_/A _9100_/Q _4865_/X VGND VGND VPWR VPWR _4873_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA_33 _5693_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_44 _7132_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6605_ _6341_/A _6158_/B _6967_/B _6597_/Y _6250_/D VGND VGND VPWR VPWR _6605_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_193_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_55 _4939_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4797_ _4797_/A _4797_/B _4797_/C VGND VGND VPWR VPWR _4817_/B sky130_fd_sc_hd__or3_1
X_7585_ _7585_/A VGND VGND VPWR VPWR _9366_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_66 _5065_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_77 _5301_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_88 _5465_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9324_ _9420_/CLK _9324_/D fanout465/X VGND VGND VPWR VPWR _9324_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_99 _5809_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6536_ _6597_/A _6660_/A VGND VGND VPWR VPWR _6591_/B sky130_fd_sc_hd__nand2_1
XFILLER_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9255_ _9486_/CLK _9255_/D fanout416/X VGND VGND VPWR VPWR _9255_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_118_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6467_ _6467_/A _6467_/B _6976_/C _6467_/D VGND VGND VPWR VPWR _6468_/D sky130_fd_sc_hd__or4_1
XFILLER_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8206_ _9100_/Q _8206_/B VGND VGND VPWR VPWR _8206_/X sky130_fd_sc_hd__or2_1
X_5418_ _5418_/A hold19/X VGND VGND VPWR VPWR _5419_/A sky130_fd_sc_hd__and2_1
X_6398_ _6437_/A _6398_/B VGND VGND VPWR VPWR _6818_/A sky130_fd_sc_hd__or2_4
X_9186_ _9194_/CLK _9186_/D fanout456/X VGND VGND VPWR VPWR _9186_/Q sky130_fd_sc_hd__dfrtp_1
X_5349_ _5353_/A _5356_/B VGND VGND VPWR VPWR _5350_/A sky130_fd_sc_hd__and2_1
X_8137_ _9318_/Q _8181_/B VGND VGND VPWR VPWR _8137_/X sky130_fd_sc_hd__or2_1
XFILLER_99_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8068_ _9427_/Q _8068_/B VGND VGND VPWR VPWR _8068_/X sky130_fd_sc_hd__and2_1
XFILLER_153_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7019_ _7025_/A _7025_/B VGND VGND VPWR VPWR _7020_/A sky130_fd_sc_hd__and2_1
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4720_ _9219_/Q _7249_/A _5795_/A _8981_/Q _4719_/X VGND VGND VPWR VPWR _4723_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4651_ _4656_/A _4794_/B VGND VGND VPWR VPWR _5529_/A sky130_fd_sc_hd__nor2_8
XFILLER_187_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput20 mask_rev_in[24] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__clkbuf_2
Xinput31 mask_rev_in[5] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4582_ _4582_/A VGND VGND VPWR VPWR _5842_/S sky130_fd_sc_hd__buf_6
X_7370_ _7279_/X hold824/X _7372_/S VGND VGND VPWR VPWR _7370_/X sky130_fd_sc_hd__mux2_1
Xinput42 mgmt_gpio_in[15] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__clkbuf_4
Xinput53 mgmt_gpio_in[25] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__clkbuf_4
XFILLER_116_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput64 mgmt_gpio_in[35] VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__clkbuf_4
Xhold804 hold804/A VGND VGND VPWR VPWR hold804/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput75 porb VGND VGND VPWR VPWR input75/X sky130_fd_sc_hd__buf_2
X_6321_ _6535_/A _6839_/B _6481_/A VGND VGND VPWR VPWR _6553_/B sky130_fd_sc_hd__and3b_1
Xhold815 _7160_/X VGND VGND VPWR VPWR _7161_/A sky130_fd_sc_hd__dlygate4sd3_1
Xinput86 spimemio_flash_io0_oeb VGND VGND VPWR VPWR input86/X sky130_fd_sc_hd__buf_2
Xhold826 _9448_/Q VGND VGND VPWR VPWR hold826/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput97 sram_ro_data[13] VGND VGND VPWR VPWR input97/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold837 _7442_/X VGND VGND VPWR VPWR _7443_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold848 hold848/A VGND VGND VPWR VPWR hold848/X sky130_fd_sc_hd__dlygate4sd3_1
X_6252_ _6311_/B _6603_/A VGND VGND VPWR VPWR _6257_/C sky130_fd_sc_hd__nor2_1
X_9040_ _9541_/CLK _9040_/D VGND VGND VPWR VPWR _9040_/Q sky130_fd_sc_hd__dfxtp_1
Xhold859 _9480_/Q VGND VGND VPWR VPWR hold859/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5203_ _9173_/Q input81/X _5279_/B VGND VGND VPWR VPWR _5204_/A sky130_fd_sc_hd__mux2_8
X_6183_ _6183_/A VGND VGND VPWR VPWR _6850_/B sky130_fd_sc_hd__buf_6
XFILLER_130_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5134_ _8375_/A _8352_/A VGND VGND VPWR VPWR _8380_/A sky130_fd_sc_hd__nand2_2
XFILLER_57_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5065_ _5067_/B _5065_/A1 _5065_/S VGND VGND VPWR VPWR _5066_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8824_ _9487_/CLK _8824_/D fanout412/X VGND VGND VPWR VPWR _8824_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_25_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8755_ _5287_/A _8755_/A2 _8755_/B1 _5275_/A VGND VGND VPWR VPWR _8755_/X sky130_fd_sc_hd__a22o_1
XFILLER_40_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5967_ _5967_/A VGND VGND VPWR VPWR _9055_/D sky130_fd_sc_hd__clkbuf_1
X_7706_ _7654_/X hold212/X _7710_/S VGND VGND VPWR VPWR _7706_/X sky130_fd_sc_hd__mux2_1
X_4918_ _4918_/A1 _4502_/Y _7086_/A _9146_/Q _4917_/X VGND VGND VPWR VPWR _4921_/C
+ sky130_fd_sc_hd__a221o_1
X_8686_ _8887_/Q _8314_/X _8331_/X _8982_/Q VGND VGND VPWR VPWR _8686_/X sky130_fd_sc_hd__a22o_1
X_5898_ _9561_/A _5897_/X _5898_/S VGND VGND VPWR VPWR _5898_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7637_ _7637_/A VGND VGND VPWR VPWR _9390_/D sky130_fd_sc_hd__clkbuf_1
X_4849_ _9080_/Q _6021_/A _6032_/A _9085_/Q VGND VGND VPWR VPWR _4852_/C sky130_fd_sc_hd__a22o_1
XFILLER_166_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7568_ _7568_/A VGND VGND VPWR VPWR _9358_/D sky130_fd_sc_hd__clkbuf_1
X_9307_ _9459_/CLK _9307_/D fanout489/X VGND VGND VPWR VPWR _9307_/Q sky130_fd_sc_hd__dfrtp_4
X_6519_ _6887_/B _6926_/B VGND VGND VPWR VPWR _6520_/A sky130_fd_sc_hd__or2_1
XFILLER_4_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7499_ _7499_/A _7499_/B VGND VGND VPWR VPWR _7515_/S sky130_fd_sc_hd__nand2_8
X_9238_ _9272_/CLK _9238_/D fanout419/X VGND VGND VPWR VPWR _9238_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9169_ _9462_/CLK _9169_/D fanout408/X VGND VGND VPWR VPWR _9169_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_57_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6870_ _6870_/A _6870_/B VGND VGND VPWR VPWR _7000_/A sky130_fd_sc_hd__or2_1
X_5821_ _5453_/B _5453_/C _5819_/X _5842_/S hold21/A VGND VGND VPWR VPWR hold43/A
+ sky130_fd_sc_hd__o221a_4
X_8540_ _9462_/Q _8348_/X _8411_/X _9342_/Q _8539_/X VGND VGND VPWR VPWR _8550_/C
+ sky130_fd_sc_hd__a221o_1
X_5752_ _5752_/A VGND VGND VPWR VPWR _8958_/D sky130_fd_sc_hd__clkbuf_1
X_4703_ _9283_/Q _7391_/A _5540_/A _8871_/Q VGND VGND VPWR VPWR _4703_/X sky130_fd_sc_hd__a22o_2
XFILLER_187_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8471_ _9435_/Q _7908_/A _8358_/C _9275_/Q VGND VGND VPWR VPWR _8471_/X sky130_fd_sc_hd__a22o_1
X_5683_ _7645_/A VGND VGND VPWR VPWR _5683_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_147_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7422_ _7422_/A VGND VGND VPWR VPWR _9294_/D sky130_fd_sc_hd__clkbuf_1
X_4634_ _4656_/A _4956_/A VGND VGND VPWR VPWR _5573_/A sky130_fd_sc_hd__nor2_8
XFILLER_190_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold601 _8855_/Q VGND VGND VPWR VPWR hold601/X sky130_fd_sc_hd__dlygate4sd3_1
X_4565_ _9421_/Q _7695_/A _7446_/A _9309_/Q VGND VGND VPWR VPWR _4565_/X sky130_fd_sc_hd__a22o_2
X_7353_ _7353_/A VGND VGND VPWR VPWR _9262_/D sky130_fd_sc_hd__clkbuf_1
Xhold612 _5488_/X VGND VGND VPWR VPWR _5489_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold623 _5396_/X VGND VGND VPWR VPWR _5397_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold634 _7837_/X VGND VGND VPWR VPWR _7838_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6304_ _6635_/A _6440_/A VGND VGND VPWR VPWR _6461_/A sky130_fd_sc_hd__or2_1
Xhold645 _9071_/Q VGND VGND VPWR VPWR hold645/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap364 _4450_/Y VGND VGND VPWR VPWR _7781_/A sky130_fd_sc_hd__buf_8
X_4496_ _7126_/A _4748_/B VGND VGND VPWR VPWR _7176_/A sky130_fd_sc_hd__nor2_8
Xhold656 _7727_/X VGND VGND VPWR VPWR _7728_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7284_ _7284_/A _7284_/B VGND VGND VPWR VPWR _7300_/S sky130_fd_sc_hd__nand2_8
Xhold667 hold667/A VGND VGND VPWR VPWR hold667/X sky130_fd_sc_hd__dlygate4sd3_1
X_9023_ _9419_/CLK _9023_/D fanout492/X VGND VGND VPWR VPWR _9584_/A sky130_fd_sc_hd__dfrtp_1
Xmax_cap386 _4414_/Y VGND VGND VPWR VPWR _7519_/A sky130_fd_sc_hd__buf_8
Xhold678 hold678/A VGND VGND VPWR VPWR hold678/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap397 hold42/X VGND VGND VPWR VPWR _4489_/A sky130_fd_sc_hd__buf_4
Xhold689 _9163_/Q VGND VGND VPWR VPWR hold689/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6235_ _6235_/A VGND VGND VPWR VPWR _6906_/A sky130_fd_sc_hd__buf_2
XFILLER_103_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ _6166_/A VGND VGND VPWR VPWR _6311_/B sky130_fd_sc_hd__buf_4
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5117_ _6080_/C _6080_/D _6079_/A _6079_/B VGND VGND VPWR VPWR _5120_/B sky130_fd_sc_hd__or4_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6097_ _6181_/A _6095_/B _6721_/A VGND VGND VPWR VPWR _6097_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5048_ _5047_/A _5045_/A _5045_/B VGND VGND VPWR VPWR _5048_/X sky130_fd_sc_hd__o21a_1
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8807_ _8831_/CLK _8807_/D _5384_/X VGND VGND VPWR VPWR _8807_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_53_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6999_ _9110_/Q _8735_/A _6978_/X _6998_/X VGND VGND VPWR VPWR _7009_/B sky130_fd_sc_hd__a22o_1
XFILLER_41_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8738_ _8738_/A VGND VGND VPWR VPWR _9542_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8669_ _8986_/Q _8292_/X _8294_/X _8881_/Q VGND VGND VPWR VPWR _8669_/X sky130_fd_sc_hd__a22o_1
XFILLER_138_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4350_ hold22/X VGND VGND VPWR VPWR _5021_/B sky130_fd_sc_hd__clkinv_2
XFILLER_153_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6020_ _6020_/A VGND VGND VPWR VPWR _9078_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7971_ _7971_/A VGND VGND VPWR VPWR _8224_/B sky130_fd_sc_hd__buf_6
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6922_ _6922_/A _6922_/B _6922_/C VGND VGND VPWR VPWR _6982_/C sky130_fd_sc_hd__nor3_1
XFILLER_23_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6853_ _6853_/A _6853_/B _6853_/C _6853_/D VGND VGND VPWR VPWR _6944_/C sky130_fd_sc_hd__or4_1
XFILLER_120_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5804_ _5653_/X hold173/X _5804_/S VGND VGND VPWR VPWR _5804_/X sky130_fd_sc_hd__mux2_1
X_9572_ _9572_/A _5096_/Y VGND VGND VPWR VPWR mgmt_gpio_out[18] sky130_fd_sc_hd__ebufn_8
XFILLER_50_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6784_ _6784_/A _6922_/B _6784_/C _6784_/D VGND VGND VPWR VPWR _6785_/B sky130_fd_sc_hd__or4_1
X_8523_ _9229_/Q _8388_/X _8379_/X _9205_/Q _8522_/X VGND VGND VPWR VPWR _8524_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5735_ _5735_/A VGND VGND VPWR VPWR _8951_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8454_ _9467_/Q _8312_/X _8376_/X _9427_/Q VGND VGND VPWR VPWR _8454_/X sky130_fd_sc_hd__a22o_1
X_5666_ _5666_/A VGND VGND VPWR VPWR _8922_/D sky130_fd_sc_hd__clkbuf_1
X_7405_ _7405_/A VGND VGND VPWR VPWR _9286_/D sky130_fd_sc_hd__clkbuf_1
X_4617_ _4617_/A _4617_/B _4617_/C _4617_/D VGND VGND VPWR VPWR _4690_/B sky130_fd_sc_hd__or4_2
XFILLER_190_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8385_ _8385_/A _8385_/B VGND VGND VPWR VPWR _8386_/A sky130_fd_sc_hd__nor2_4
X_5597_ hold913/X _5505_/X _5605_/S VGND VGND VPWR VPWR _5598_/A sky130_fd_sc_hd__mux2_1
Xhold420 _5500_/X VGND VGND VPWR VPWR _5501_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7336_ _7336_/A VGND VGND VPWR VPWR _9254_/D sky130_fd_sc_hd__clkbuf_1
Xhold431 _9542_/Q VGND VGND VPWR VPWR hold431/X sky130_fd_sc_hd__dlygate4sd3_1
X_4548_ _4548_/A _4548_/B _4548_/C _4548_/D VGND VGND VPWR VPWR _4549_/D sky130_fd_sc_hd__or4_1
XFILLER_144_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold442 _5905_/X VGND VGND VPWR VPWR _9018_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold453 hold453/A VGND VGND VPWR VPWR hold453/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 _5521_/X VGND VGND VPWR VPWR _5522_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 _9473_/Q VGND VGND VPWR VPWR hold475/X sky130_fd_sc_hd__dlygate4sd3_1
X_7267_ _7128_/X hold912/X _7282_/S VGND VGND VPWR VPWR _7268_/A sky130_fd_sc_hd__mux2_1
Xhold486 _9178_/Q VGND VGND VPWR VPWR hold486/X sky130_fd_sc_hd__dlygate4sd3_1
X_4479_ hold33/X _7158_/B VGND VGND VPWR VPWR _4811_/A sky130_fd_sc_hd__nor2_8
XFILLER_104_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold497 _7820_/X VGND VGND VPWR VPWR _7821_/A sky130_fd_sc_hd__dlygate4sd3_1
X_9006_ _9006_/CLK _9006_/D fanout494/X VGND VGND VPWR VPWR _9006_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6218_ _6402_/A _6311_/B VGND VGND VPWR VPWR _6219_/A sky130_fd_sc_hd__or2_1
X_7198_ _7198_/A VGND VGND VPWR VPWR _9193_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1120 _9035_/Q VGND VGND VPWR VPWR hold890/A sky130_fd_sc_hd__dlygate4sd3_1
X_6149_ _6635_/A _6628_/B VGND VGND VPWR VPWR _6150_/A sky130_fd_sc_hd__or2_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1131 _8974_/Q VGND VGND VPWR VPWR hold768/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1142 _7400_/X VGND VGND VPWR VPWR _7401_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1153 _9072_/Q VGND VGND VPWR VPWR hold448/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1164 _9087_/Q VGND VGND VPWR VPWR hold500/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1175 _9370_/Q VGND VGND VPWR VPWR hold711/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1186 _5892_/X VGND VGND VPWR VPWR hold1186/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_304 _7304_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1197 _8943_/Q VGND VGND VPWR VPWR hold941/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_315 hold46/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_326 _4549_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_337 _5387_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_348 _7233_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_359 _8023_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5520_ _5520_/A VGND VGND VPWR VPWR _8858_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5451_ _5451_/A VGND VGND VPWR VPWR _5451_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_117_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4402_ _4418_/A _4402_/B VGND VGND VPWR VPWR _4492_/A sky130_fd_sc_hd__nand2_8
X_8170_ _9207_/Q _7938_/X _8077_/X _9351_/Q _8169_/X VGND VGND VPWR VPWR _8171_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_99_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5382_ _5382_/A VGND VGND VPWR VPWR _5382_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_160_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7121_ _7121_/A VGND VGND VPWR VPWR _7121_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7052_ _6018_/X _9130_/Q _7054_/S VGND VGND VPWR VPWR _7052_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6003_ hold448/X _5687_/X _6005_/S VGND VGND VPWR VPWR _6004_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7954_ _9376_/Q _7947_/X _7949_/X _9240_/Q _7953_/X VGND VGND VPWR VPWR _7965_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_54_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6905_ _6905_/A _6905_/B _6978_/C VGND VGND VPWR VPWR _6905_/X sky130_fd_sc_hd__or3b_1
XFILLER_35_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7885_ _9496_/Q VGND VGND VPWR VPWR _8181_/B sky130_fd_sc_hd__clkinv_4
XFILLER_35_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6836_ _6836_/A _6988_/A _6987_/D VGND VGND VPWR VPWR _6925_/C sky130_fd_sc_hd__or3_1
XFILLER_145_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9555_ _9555_/A VGND VGND VPWR VPWR _9555_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6767_ _6772_/A _6520_/A _6345_/X _6768_/A VGND VGND VPWR VPWR _6770_/C sky130_fd_sc_hd__a2bb2o_1
XFILLER_183_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8506_ _9413_/Q _8506_/B VGND VGND VPWR VPWR _8506_/X sky130_fd_sc_hd__and2_1
X_5718_ hold796/X _5587_/X _5724_/S VGND VGND VPWR VPWR _5719_/A sky130_fd_sc_hd__mux2_1
X_9486_ _9486_/CLK _9486_/D fanout416/X VGND VGND VPWR VPWR _9486_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6698_ _6673_/B _6481_/A _6693_/Y _6694_/Y _6697_/Y VGND VGND VPWR VPWR _6698_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_163_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8437_ _8437_/A _8437_/B _8437_/C _8437_/D VGND VGND VPWR VPWR _8437_/X sky130_fd_sc_hd__or4_4
X_5649_ _5649_/A VGND VGND VPWR VPWR _8915_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8368_ _8385_/A _8368_/B VGND VGND VPWR VPWR _8369_/A sky130_fd_sc_hd__nor2_4
XFILLER_151_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold250 _9413_/Q VGND VGND VPWR VPWR hold250/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 _7260_/X VGND VGND VPWR VPWR _7261_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7319_ _7299_/X hold527/X _7319_/S VGND VGND VPWR VPWR _7319_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold272 _7419_/X VGND VGND VPWR VPWR _7420_/A sky130_fd_sc_hd__dlygate4sd3_1
X_8299_ _9498_/Q _9497_/Q VGND VGND VPWR VPWR _8389_/C sky130_fd_sc_hd__nor2_2
Xhold283 _9332_/Q VGND VGND VPWR VPWR hold283/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 _7333_/X VGND VGND VPWR VPWR _7334_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 _5809_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_112 _6015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_123 _7147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 _7762_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 _7923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 _7947_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_167 _8023_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_178 _7973_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_189 _7997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_1_1_1_csclk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_167_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput7 mask_rev_in[12] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4951_ _9344_/Q _7536_/A _4483_/Y _4951_/B2 _4950_/X VGND VGND VPWR VPWR _4960_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_17_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7670_ _7651_/X hold373/X _7676_/S VGND VGND VPWR VPWR _7671_/A sky130_fd_sc_hd__mux2_1
X_4882_ _9369_/Q _7588_/A _5584_/A _8889_/Q _4881_/X VGND VGND VPWR VPWR _4883_/D
+ sky130_fd_sc_hd__a221o_1
X_6621_ _6873_/B _6800_/A VGND VGND VPWR VPWR _6869_/B sky130_fd_sc_hd__nor2_1
XFILLER_60_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9340_ _9468_/CLK _9340_/D fanout466/X VGND VGND VPWR VPWR _9340_/Q sky130_fd_sc_hd__dfrtp_4
X_6552_ _6736_/A _6624_/B VGND VGND VPWR VPWR _6966_/A sky130_fd_sc_hd__nor2_1
XFILLER_118_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5503_ _5503_/A VGND VGND VPWR VPWR _8852_/D sky130_fd_sc_hd__clkbuf_1
X_9271_ _9421_/CLK _9271_/D fanout460/X VGND VGND VPWR VPWR _9271_/Q sky130_fd_sc_hd__dfrtp_2
X_6483_ _6483_/A _6483_/B _6859_/B _6483_/D VGND VGND VPWR VPWR _6484_/B sky130_fd_sc_hd__or4_1
XFILLER_145_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8222_ _8965_/Q _7960_/X _7981_/X _8915_/Q VGND VGND VPWR VPWR _8222_/X sky130_fd_sc_hd__a22o_1
Xoutput300 _9141_/Q VGND VGND VPWR VPWR pwr_ctrl_out[0] sky130_fd_sc_hd__buf_12
X_5434_ _5434_/A VGND VGND VPWR VPWR _8823_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput311 _5280_/X VGND VGND VPWR VPWR spi_sdi sky130_fd_sc_hd__buf_12
XFILLER_160_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput322 _9153_/Q VGND VGND VPWR VPWR sram_ro_addr[6] sky130_fd_sc_hd__buf_12
XFILLER_105_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput333 _9060_/Q VGND VGND VPWR VPWR wb_dat_o[15] sky130_fd_sc_hd__buf_12
X_8153_ _9383_/Q _7947_/X _7981_/X _9335_/Q VGND VGND VPWR VPWR _8153_/X sky130_fd_sc_hd__a22o_1
Xoutput344 _9535_/Q VGND VGND VPWR VPWR wb_dat_o[25] sky130_fd_sc_hd__buf_12
X_5365_ _5375_/A _5378_/B VGND VGND VPWR VPWR _5366_/A sky130_fd_sc_hd__and2_1
Xoutput355 _9067_/Q VGND VGND VPWR VPWR wb_dat_o[6] sky130_fd_sc_hd__buf_12
X_7104_ _5468_/X _9153_/Q _7106_/S VGND VGND VPWR VPWR _7104_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_3_0_csclk clkbuf_3_3_0_csclk/A VGND VGND VPWR VPWR _9090_/CLK sky130_fd_sc_hd__clkbuf_8
X_8084_ _5130_/A _9509_/Q _8013_/A _8083_/X VGND VGND VPWR VPWR _8084_/X sky130_fd_sc_hd__a211o_1
X_5296_ _5296_/A _7139_/B VGND VGND VPWR VPWR _5316_/S sky130_fd_sc_hd__nand2_4
XFILLER_99_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7035_ _5951_/X _9122_/Q _7041_/S VGND VGND VPWR VPWR _7035_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8986_ _9084_/CLK _8986_/D fanout446/X VGND VGND VPWR VPWR _8986_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_55_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7937_ _8206_/B _7984_/C _8002_/B VGND VGND VPWR VPWR _7938_/A sky130_fd_sc_hd__and3_2
XFILLER_35_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
X_7868_ _7868_/A1 _7864_/A _7867_/Y VGND VGND VPWR VPWR _9491_/D sky130_fd_sc_hd__o21a_1
XFILLER_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6819_ _6898_/A _6818_/X _6812_/Y VGND VGND VPWR VPWR _6819_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_168_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7799_ _5387_/X hold921/X _7813_/S VGND VGND VPWR VPWR _7800_/A sky130_fd_sc_hd__mux2_1
X_9538_ _9541_/CLK _9538_/D VGND VGND VPWR VPWR _9538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9469_ _9469_/CLK _9469_/D fanout459/X VGND VGND VPWR VPWR _9469_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_10 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5150_ _8706_/A _8705_/B _5149_/Y VGND VGND VPWR VPWR _9025_/D sky130_fd_sc_hd__o21ai_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5081_ _9451_/Q VGND VGND VPWR VPWR _5081_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8840_ _9178_/CLK _8840_/D fanout486/X VGND VGND VPWR VPWR _8840_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_80_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8771_ _5292_/A _5149_/A _6908_/A _8770_/X VGND VGND VPWR VPWR _9551_/D sky130_fd_sc_hd__o31a_1
X_5983_ _5983_/A VGND VGND VPWR VPWR _9062_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7722_ _7722_/A VGND VGND VPWR VPWR _9428_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4934_ _9280_/Q _7391_/A _4650_/Y _4933_/X VGND VGND VPWR VPWR _4939_/B sky130_fd_sc_hd__a211o_2
XFILLER_178_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7653_ _7653_/A VGND VGND VPWR VPWR _9396_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4865_ _9289_/Q _7408_/A _4477_/Y input15/X VGND VGND VPWR VPWR _4865_/X sky130_fd_sc_hd__a22o_1
XANTENNA_12 _9339_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_23 _4460_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_34 _5784_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6604_ _6609_/A _6445_/Y _6603_/Y VGND VGND VPWR VPWR _6614_/C sky130_fd_sc_hd__a21o_1
X_7584_ _7494_/X hold777/X hold78/X VGND VGND VPWR VPWR _7585_/A sky130_fd_sc_hd__mux2_1
XANTENNA_45 _7132_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4796_ _9218_/Q _7249_/A _7571_/A _9362_/Q _4795_/X VGND VGND VPWR VPWR _4797_/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA_56 _4939_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_67 _5198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_78 _5311_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9323_ _9459_/CLK _9323_/D fanout489/X VGND VGND VPWR VPWR _9323_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_89 _5468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6535_ _6535_/A _6887_/B VGND VGND VPWR VPWR _6660_/A sky130_fd_sc_hd__nor2_2
XFILLER_192_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9254_ _9487_/CLK _9254_/D fanout411/X VGND VGND VPWR VPWR _9254_/Q sky130_fd_sc_hd__dfrtp_4
X_6466_ _6466_/A _6830_/A VGND VGND VPWR VPWR _6467_/D sky130_fd_sc_hd__nor2_1
XFILLER_118_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8205_ _9049_/Q _7923_/X _7997_/X _8954_/Q _8204_/X VGND VGND VPWR VPWR _8209_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5417_ _5417_/A VGND VGND VPWR VPWR _8816_/D sky130_fd_sc_hd__clkbuf_1
X_9185_ _9482_/CLK _9185_/D fanout433/X VGND VGND VPWR VPWR _9185_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_133_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6397_ _6466_/A VGND VGND VPWR VPWR _6781_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8136_ _9214_/Q _7923_/A _7997_/A _9366_/Q _8135_/X VGND VGND VPWR VPWR _8140_/C
+ sky130_fd_sc_hd__a221o_1
X_5348_ _5348_/A VGND VGND VPWR VPWR _5348_/X sky130_fd_sc_hd__clkbuf_1
X_8067_ _9235_/Q _8034_/X _7988_/X _9435_/Q _8066_/X VGND VGND VPWR VPWR _8072_/B
+ sky130_fd_sc_hd__a221o_1
X_5279_ _5279_/A _5279_/B VGND VGND VPWR VPWR _5280_/A sky130_fd_sc_hd__and2_1
XFILLER_87_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7018_ _7018_/A VGND VGND VPWR VPWR _7018_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_75_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8969_ _9419_/CLK _8969_/D fanout491/X VGND VGND VPWR VPWR _8969_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_71_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4650_ _7111_/B _7126_/B VGND VGND VPWR VPWR _4650_/Y sky130_fd_sc_hd__nor2_4
XFILLER_159_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput10 mask_rev_in[15] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__clkbuf_2
Xinput21 mask_rev_in[25] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__clkbuf_4
Xinput32 mask_rev_in[6] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__clkbuf_1
X_4581_ _9405_/Q _7661_/A _7781_/A _9461_/Q _4580_/X VGND VGND VPWR VPWR _4590_/A
+ sky130_fd_sc_hd__a221o_1
Xinput43 mgmt_gpio_in[16] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__clkbuf_4
Xinput54 mgmt_gpio_in[26] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6320_ _6392_/A _6392_/B VGND VGND VPWR VPWR _6481_/A sky130_fd_sc_hd__nor2_4
XFILLER_143_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold805 _9197_/Q VGND VGND VPWR VPWR hold805/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput65 mgmt_gpio_in[36] VGND VGND VPWR VPWR _9554_/A sky130_fd_sc_hd__buf_4
Xhold816 _8837_/Q VGND VGND VPWR VPWR hold816/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput76 qspi_enabled VGND VGND VPWR VPWR _5194_/S sky130_fd_sc_hd__buf_4
Xinput87 spimemio_flash_io1_do VGND VGND VPWR VPWR _9553_/A sky130_fd_sc_hd__clkbuf_4
Xhold827 _9184_/Q VGND VGND VPWR VPWR hold827/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput98 sram_ro_data[14] VGND VGND VPWR VPWR input98/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold838 _8840_/Q VGND VGND VPWR VPWR hold838/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 hold849/A VGND VGND VPWR VPWR hold849/X sky130_fd_sc_hd__dlygate4sd3_1
X_6251_ _6856_/A _6857_/A _6857_/B _6250_/X VGND VGND VPWR VPWR _6257_/B sky130_fd_sc_hd__or4b_2
XFILLER_107_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5202_ _5202_/A VGND VGND VPWR VPWR _9587_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6182_ _6182_/A _6169_/A VGND VGND VPWR VPWR _6183_/A sky130_fd_sc_hd__or2b_1
XFILLER_97_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5133_ _9500_/Q _9499_/Q VGND VGND VPWR VPWR _8352_/A sky130_fd_sc_hd__nor2b_2
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5064_ _5064_/A VGND VGND VPWR VPWR _8782_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8823_ _9487_/CLK _8823_/D fanout412/X VGND VGND VPWR VPWR _8823_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8754_ _8754_/A VGND VGND VPWR VPWR _9546_/D sky130_fd_sc_hd__clkbuf_1
X_5966_ _9055_/Q _4817_/X _5976_/S VGND VGND VPWR VPWR _5967_/A sky130_fd_sc_hd__mux2_1
X_7705_ _7705_/A VGND VGND VPWR VPWR _9420_/D sky130_fd_sc_hd__clkbuf_1
X_4917_ _9240_/Q _7304_/A _4915_/X _7108_/A VGND VGND VPWR VPWR _4917_/X sky130_fd_sc_hd__a22o_1
X_8685_ _8917_/Q _8298_/X _8370_/X _9088_/Q _8684_/X VGND VGND VPWR VPWR _8688_/C
+ sky130_fd_sc_hd__a221o_1
X_5897_ hold567/X hold5/X _5897_/S VGND VGND VPWR VPWR _5897_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7636_ _7494_/X hold735/X _7638_/S VGND VGND VPWR VPWR _7636_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4848_ _9297_/Q _7425_/A _7194_/A _9193_/Q _4847_/X VGND VGND VPWR VPWR _4852_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7567_ _7494_/X hold756/X hold99/A VGND VGND VPWR VPWR _7567_/X sky130_fd_sc_hd__mux2_1
X_4779_ _8819_/Q _5418_/A _5607_/A _8900_/Q VGND VGND VPWR VPWR _4779_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9306_ _9370_/CLK _9306_/D fanout475/X VGND VGND VPWR VPWR _9306_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_181_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6518_ _6518_/A _6527_/A VGND VGND VPWR VPWR _6518_/Y sky130_fd_sc_hd__nor2_4
XFILLER_174_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7498_ _7498_/A VGND VGND VPWR VPWR _9327_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9237_ _9421_/CLK _9237_/D fanout460/X VGND VGND VPWR VPWR _9237_/Q sky130_fd_sc_hd__dfrtp_1
X_6449_ _6466_/A _6449_/B VGND VGND VPWR VPWR _6759_/B sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_40_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _9181_/CLK sky130_fd_sc_hd__clkbuf_16
X_9168_ _9462_/CLK _9168_/D fanout408/X VGND VGND VPWR VPWR _9168_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_164_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8119_ _9229_/Q _7979_/X _8001_/X _9269_/Q _8118_/X VGND VGND VPWR VPWR _8127_/A
+ sky130_fd_sc_hd__a221o_1
Xclkbuf_2_0_0_csclk clkbuf_2_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_1_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
X_9099_ _9473_/CLK _9099_/D fanout431/X VGND VGND VPWR VPWR _9099_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_48_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_55_csclk clkbuf_opt_2_0_csclk/X VGND VGND VPWR VPWR _9088_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5820_ hold20/A VGND VGND VPWR VPWR hold21/A sky130_fd_sc_hd__buf_12
XFILLER_34_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5751_ hold870/X _5505_/X _5759_/S VGND VGND VPWR VPWR _5752_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4702_ _4702_/A _4702_/B _4702_/C _4702_/D VGND VGND VPWR VPWR _4724_/A sky130_fd_sc_hd__or4_1
X_8470_ _9227_/Q _8388_/A _8379_/A _9203_/Q _8469_/X VGND VGND VPWR VPWR _8473_/C
+ sky130_fd_sc_hd__a221o_1
X_5682_ _5682_/A VGND VGND VPWR VPWR _8929_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7421_ _7279_/X hold733/X _7423_/S VGND VGND VPWR VPWR _7421_/X sky130_fd_sc_hd__mux2_1
X_4633_ _4633_/A _4633_/B _4633_/C _4633_/D VGND VGND VPWR VPWR _4690_/C sky130_fd_sc_hd__or4_1
XFILLER_148_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7352_ _7279_/X hold832/X _7354_/S VGND VGND VPWR VPWR _7352_/X sky130_fd_sc_hd__mux2_1
XFILLER_162_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4564_ _9261_/Q _4409_/Y _7113_/A _4562_/X _4563_/X VGND VGND VPWR VPWR _4569_/B
+ sky130_fd_sc_hd__a221o_1
Xhold602 _5511_/X VGND VGND VPWR VPWR _5512_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold613 _8845_/Q VGND VGND VPWR VPWR hold613/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold624 _9231_/Q VGND VGND VPWR VPWR hold624/X sky130_fd_sc_hd__dlygate4sd3_1
X_6303_ _6303_/A VGND VGND VPWR VPWR _6440_/A sky130_fd_sc_hd__buf_4
Xhold635 hold635/A VGND VGND VPWR VPWR hold635/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7283_ _7283_/A VGND VGND VPWR VPWR _9231_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4495_ _4495_/A _4495_/B _4495_/C _4495_/D VGND VGND VPWR VPWR _4506_/C sky130_fd_sc_hd__or4_1
Xhold646 _9367_/Q VGND VGND VPWR VPWR hold646/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap365 _4427_/Y VGND VGND VPWR VPWR _7553_/A sky130_fd_sc_hd__buf_8
Xhold657 hold657/A VGND VGND VPWR VPWR hold657/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9022_ _9419_/CLK _9022_/D fanout491/X VGND VGND VPWR VPWR _9583_/A sky130_fd_sc_hd__dfrtp_1
Xmax_cap376 _4455_/Y VGND VGND VPWR VPWR _7481_/A sky130_fd_sc_hd__buf_8
Xhold668 _9271_/Q VGND VGND VPWR VPWR hold668/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap387 _4407_/Y VGND VGND VPWR VPWR _7391_/A sky130_fd_sc_hd__buf_6
Xhold679 _9205_/Q VGND VGND VPWR VPWR hold679/X sky130_fd_sc_hd__dlygate4sd3_1
X_6234_ _6248_/A _6420_/B VGND VGND VPWR VPWR _6235_/A sky130_fd_sc_hd__or2_1
Xmax_cap398 _4418_/A VGND VGND VPWR VPWR _4396_/A sky130_fd_sc_hd__buf_4
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _6248_/A _6317_/A _6167_/B VGND VGND VPWR VPWR _6166_/A sky130_fd_sc_hd__or3_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5116_ _6080_/A _6080_/B VGND VGND VPWR VPWR _5120_/A sky130_fd_sc_hd__or2_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096_ _6181_/B VGND VGND VPWR VPWR _6721_/A sky130_fd_sc_hd__buf_2
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5047_ _5047_/A VGND VGND VPWR VPWR _5047_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8806_ _5168_/A1 _8806_/D _5382_/X VGND VGND VPWR VPWR _8806_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6998_ _6998_/A _6998_/B VGND VGND VPWR VPWR _6998_/X sky130_fd_sc_hd__or2_1
XFILLER_53_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5949_ _5947_/X hold855/X _5958_/S VGND VGND VPWR VPWR _5949_/X sky130_fd_sc_hd__mux2_1
X_8737_ _8729_/X _8737_/A1 _8765_/S VGND VGND VPWR VPWR _8738_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8668_ _9077_/Q _8322_/X _8333_/X _8866_/Q _8667_/X VGND VGND VPWR VPWR _8675_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7619_ hold386/X _7494_/A _7621_/S VGND VGND VPWR VPWR _7620_/A sky130_fd_sc_hd__mux2_1
X_8599_ _8973_/Q _8337_/X _8384_/X _8853_/Q _8598_/X VGND VGND VPWR VPWR _8600_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput200 wb_sel_i[3] VGND VGND VPWR VPWR _8731_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_76_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7970_ _9496_/Q _7992_/C _8002_/C VGND VGND VPWR VPWR _7971_/A sky130_fd_sc_hd__and3_4
XFILLER_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6921_ _6799_/A _6828_/X _6926_/A _6852_/A VGND VGND VPWR VPWR _6922_/C sky130_fd_sc_hd__o22ai_1
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6852_ _6852_/A _6862_/B VGND VGND VPWR VPWR _6853_/B sky130_fd_sc_hd__nor2_1
XFILLER_23_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5803_ _5803_/A VGND VGND VPWR VPWR _8981_/D sky130_fd_sc_hd__clkbuf_1
X_9571_ _9571_/A _5097_/Y VGND VGND VPWR VPWR mgmt_gpio_out[17] sky130_fd_sc_hd__ebufn_8
X_6783_ _6955_/C _6867_/B _6782_/X VGND VGND VPWR VPWR _6784_/D sky130_fd_sc_hd__or3b_1
X_8522_ _9389_/Q _8292_/X _8294_/X _9293_/Q VGND VGND VPWR VPWR _8522_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5734_ _5650_/X hold390/X _5736_/S VGND VGND VPWR VPWR _5735_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8453_ hold968/X _8196_/S _8451_/X _8452_/X VGND VGND VPWR VPWR _8453_/X sky130_fd_sc_hd__o22a_1
X_5665_ hold662/X _5402_/X _5665_/S VGND VGND VPWR VPWR _5666_/A sky130_fd_sc_hd__mux2_1
XFILLER_176_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7404_ _7279_/X hold834/X _7406_/S VGND VGND VPWR VPWR _7404_/X sky130_fd_sc_hd__mux2_1
X_4616_ _9276_/Q _4938_/A2 _4483_/Y _4616_/B2 _4615_/X VGND VGND VPWR VPWR _4617_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_190_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8384_ _8384_/A VGND VGND VPWR VPWR _8384_/X sky130_fd_sc_hd__buf_8
XFILLER_135_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5596_ _5596_/A _5715_/B VGND VGND VPWR VPWR _5605_/S sky130_fd_sc_hd__and2_2
Xhold410 hold410/A VGND VGND VPWR VPWR hold410/X sky130_fd_sc_hd__dlygate4sd3_1
X_7335_ hold358/X _7494_/A _7337_/S VGND VGND VPWR VPWR _7335_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold421 hold421/A VGND VGND VPWR VPWR hold421/X sky130_fd_sc_hd__dlygate4sd3_1
X_4547_ _9310_/Q _7446_/A _7623_/A _9390_/Q _4546_/X VGND VGND VPWR VPWR _4548_/D
+ sky130_fd_sc_hd__a221o_1
Xhold432 _5289_/X VGND VGND VPWR VPWR _5504_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 _5399_/X VGND VGND VPWR VPWR _5400_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold454 hold454/A VGND VGND VPWR VPWR hold454/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold465 hold465/A VGND VGND VPWR VPWR _7083_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7266_ _7266_/A _7284_/B VGND VGND VPWR VPWR _7282_/S sky130_fd_sc_hd__nand2_8
X_4478_ _4492_/A _4665_/A VGND VGND VPWR VPWR _4478_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold476 _9457_/Q VGND VGND VPWR VPWR hold476/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 _7164_/X VGND VGND VPWR VPWR _7165_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold498 hold498/A VGND VGND VPWR VPWR hold498/X sky130_fd_sc_hd__dlygate4sd3_1
X_9005_ _9005_/CLK _9005_/D fanout490/X VGND VGND VPWR VPWR _9005_/Q sky130_fd_sc_hd__dfrtp_1
X_6217_ _6507_/A _6217_/B VGND VGND VPWR VPWR _6217_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7197_ _7147_/X hold316/X _7209_/S VGND VGND VPWR VPWR _7197_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6148_ _6324_/A VGND VGND VPWR VPWR _6635_/A sky130_fd_sc_hd__clkbuf_8
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1110 _9073_/Q VGND VGND VPWR VPWR hold609/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1121 _9378_/Q VGND VGND VPWR VPWR hold715/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1132 _9436_/Q VGND VGND VPWR VPWR hold381/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1143 _9420_/Q VGND VGND VPWR VPWR hold370/A sky130_fd_sc_hd__dlygate4sd3_1
X_6079_ _6079_/A _6079_/B _6079_/C _6079_/D VGND VGND VPWR VPWR _6170_/C sky130_fd_sc_hd__and4_1
XFILLER_57_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1154 _9085_/Q VGND VGND VPWR VPWR hold468/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1165 _8922_/Q VGND VGND VPWR VPWR hold662/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 _8874_/Q VGND VGND VPWR VPWR hold594/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1187 _8772_/Q VGND VGND VPWR VPWR hold820/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1198 _8947_/Q VGND VGND VPWR VPWR hold485/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_305 _7211_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_316 _7126_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_327 _4883_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_338 _5465_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_349 _7233_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5450_ _7011_/A _7013_/B VGND VGND VPWR VPWR _5451_/A sky130_fd_sc_hd__and2_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4401_ _4656_/A _5474_/B VGND VGND VPWR VPWR _7446_/A sky130_fd_sc_hd__nor2_8
X_5381_ _7011_/A _7013_/B VGND VGND VPWR VPWR _5382_/A sky130_fd_sc_hd__and2_1
XFILLER_172_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7120_ _5465_/X _9160_/Q _7124_/S VGND VGND VPWR VPWR _7120_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A VGND VGND VPWR VPWR _9532_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_99_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7051_ _7051_/A VGND VGND VPWR VPWR _9129_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6002_ _6002_/A VGND VGND VPWR VPWR _9071_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7953_ _9280_/Q _7953_/B VGND VGND VPWR VPWR _7953_/X sky130_fd_sc_hd__and2_1
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6904_ _6903_/X _6918_/A _6904_/C _6918_/B VGND VGND VPWR VPWR _6978_/C sky130_fd_sc_hd__and4b_1
X_7884_ _9495_/Q _7887_/B _7883_/B _7888_/S VGND VGND VPWR VPWR _9495_/D sky130_fd_sc_hd__a31o_1
XFILLER_23_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6835_ _6835_/A _6835_/B VGND VGND VPWR VPWR _6988_/A sky130_fd_sc_hd__or2_1
XFILLER_11_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6766_ _6779_/A _6874_/A VGND VGND VPWR VPWR _6768_/A sky130_fd_sc_hd__nand2_1
X_9554_ _9554_/A VGND VGND VPWR VPWR _9554_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5717_ _5717_/A VGND VGND VPWR VPWR _8943_/D sky130_fd_sc_hd__clkbuf_1
X_8505_ _9421_/Q _8402_/X _8378_/X _9357_/Q _8504_/X VGND VGND VPWR VPWR _8512_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_149_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9485_ _9485_/CLK _9485_/D fanout413/X VGND VGND VPWR VPWR _9485_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6697_ _6781_/C _6697_/B VGND VGND VPWR VPWR _6697_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5648_ _5647_/X hold572/X _5654_/S VGND VGND VPWR VPWR _5649_/A sky130_fd_sc_hd__mux2_1
X_8436_ _9314_/Q _8372_/X _8369_/X _9322_/Q _8435_/X VGND VGND VPWR VPWR _8437_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_163_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8367_ _8367_/A VGND VGND VPWR VPWR _8367_/X sky130_fd_sc_hd__clkbuf_8
X_5579_ _5579_/A VGND VGND VPWR VPWR _8885_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold240 _9340_/Q VGND VGND VPWR VPWR hold240/X sky130_fd_sc_hd__dlygate4sd3_1
X_7318_ _7318_/A VGND VGND VPWR VPWR _9246_/D sky130_fd_sc_hd__clkbuf_1
Xhold251 _7689_/X VGND VGND VPWR VPWR _7690_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 _9333_/Q VGND VGND VPWR VPWR hold262/X sky130_fd_sc_hd__dlygate4sd3_1
X_8298_ _8298_/A VGND VGND VPWR VPWR _8298_/X sky130_fd_sc_hd__buf_8
XFILLER_49_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold273 _9277_/Q VGND VGND VPWR VPWR hold273/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold284 _7508_/X VGND VGND VPWR VPWR _7509_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7249_ _7249_/A _7284_/B VGND VGND VPWR VPWR _7264_/S sky130_fd_sc_hd__nand2_8
Xhold295 _9209_/Q VGND VGND VPWR VPWR hold295/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_102 hold43/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_113 _6018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_124 _7233_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_135 _7796_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_146 _7923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_157 _7947_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 _8023_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_179 _7973_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 mask_rev_in[13] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4950_ _8983_/Q _5806_/A _6032_/A _9084_/Q VGND VGND VPWR VPWR _4950_/X sky130_fd_sc_hd__a22o_1
XFILLER_17_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4881_ _8899_/Q _5607_/A _7077_/A _9142_/Q VGND VGND VPWR VPWR _4881_/X sky130_fd_sc_hd__a22o_2
XFILLER_189_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6620_ _6726_/A _6726_/B _6863_/C _6620_/D VGND VGND VPWR VPWR _6620_/X sky130_fd_sc_hd__or4_1
XFILLER_177_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6551_ _6790_/A _6764_/A VGND VGND VPWR VPWR _6551_/Y sky130_fd_sc_hd__nand2_2
XFILLER_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5502_ hold823/X _5402_/X _5502_/S VGND VGND VPWR VPWR _5503_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9270_ _9421_/CLK _9270_/D fanout460/X VGND VGND VPWR VPWR _9270_/Q sky130_fd_sc_hd__dfrtp_4
X_6482_ _6482_/A _6772_/B VGND VGND VPWR VPWR _6483_/D sky130_fd_sc_hd__nor2_1
XFILLER_146_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8221_ _8860_/Q _7927_/X _8001_/X _8865_/Q _8220_/X VGND VGND VPWR VPWR _8228_/A
+ sky130_fd_sc_hd__a221o_1
X_5433_ _8823_/Q _7494_/A _5435_/S VGND VGND VPWR VPWR _5433_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput301 _9142_/Q VGND VGND VPWR VPWR pwr_ctrl_out[1] sky130_fd_sc_hd__buf_12
XFILLER_105_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput312 _5180_/X VGND VGND VPWR VPWR spimemio_flash_io0_di sky130_fd_sc_hd__buf_12
Xoutput323 _9154_/Q VGND VGND VPWR VPWR sram_ro_addr[7] sky130_fd_sc_hd__buf_12
X_8152_ hold976/X _8017_/X _8151_/X VGND VGND VPWR VPWR _8152_/X sky130_fd_sc_hd__o21a_1
X_5364_ _5364_/A VGND VGND VPWR VPWR _5364_/X sky130_fd_sc_hd__clkbuf_1
Xoutput334 _9040_/Q VGND VGND VPWR VPWR wb_dat_o[16] sky130_fd_sc_hd__buf_12
XFILLER_126_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput345 _9536_/Q VGND VGND VPWR VPWR wb_dat_o[26] sky130_fd_sc_hd__buf_12
Xoutput356 _9068_/Q VGND VGND VPWR VPWR wb_dat_o[7] sky130_fd_sc_hd__buf_12
X_7103_ _7103_/A VGND VGND VPWR VPWR _9152_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8083_ _9187_/Q _8010_/B _8072_/X _8082_/X _8627_/S VGND VGND VPWR VPWR _8083_/X
+ sky130_fd_sc_hd__o221a_1
X_5295_ hold20/X VGND VGND VPWR VPWR _7139_/B sky130_fd_sc_hd__buf_4
X_7034_ _7034_/A VGND VGND VPWR VPWR _9121_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8985_ _9084_/CLK _8985_/D fanout445/X VGND VGND VPWR VPWR _8985_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_82_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7936_ _9492_/Q _9493_/Q VGND VGND VPWR VPWR _8002_/B sky130_fd_sc_hd__and2b_4
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7867_ _7868_/A1 _7864_/A _7865_/A VGND VGND VPWR VPWR _7867_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6818_ _6818_/A _6887_/B _6416_/A VGND VGND VPWR VPWR _6818_/X sky130_fd_sc_hd__or3b_1
X_7798_ _7798_/A hold21/X VGND VGND VPWR VPWR _7813_/S sky130_fd_sc_hd__nand2_8
XFILLER_51_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9537_ _9541_/CLK _9537_/D VGND VGND VPWR VPWR _9537_/Q sky130_fd_sc_hd__dfxtp_1
X_6749_ _6906_/A _6736_/B _6858_/B VGND VGND VPWR VPWR _6861_/A sky130_fd_sc_hd__a21oi_1
XFILLER_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9468_ _9468_/CLK _9468_/D fanout465/X VGND VGND VPWR VPWR _9468_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_176_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8419_ _9433_/Q _7908_/A _8335_/X _9273_/Q VGND VGND VPWR VPWR _8419_/X sky130_fd_sc_hd__a22o_1
X_9399_ _9463_/CLK _9399_/D _5070_/A VGND VGND VPWR VPWR _9399_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5080_ _9459_/Q VGND VGND VPWR VPWR _5080_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8770_ _5149_/Y _8727_/Y _8734_/X _8769_/X _8732_/A VGND VGND VPWR VPWR _8770_/X
+ sky130_fd_sc_hd__a32o_1
X_5982_ _9062_/Q _4885_/X _5994_/S VGND VGND VPWR VPWR _5983_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4933_ _8863_/Q _5529_/A _7132_/A _9167_/Q _4932_/X VGND VGND VPWR VPWR _4933_/X
+ sky130_fd_sc_hd__a221o_1
X_7721_ _7651_/X hold354/X hold95/A VGND VGND VPWR VPWR _7722_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4864_ _4864_/A _4864_/B _4864_/C VGND VGND VPWR VPWR _4884_/B sky130_fd_sc_hd__or3_2
X_7652_ _7651_/X hold366/X hold84/X VGND VGND VPWR VPWR _7653_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_13 _9504_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_24 _4531_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6603_ _6603_/A _6610_/A VGND VGND VPWR VPWR _6603_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_35 _5529_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7583_ _7583_/A VGND VGND VPWR VPWR _9365_/D sky130_fd_sc_hd__clkbuf_1
X_4795_ _9149_/Q _7091_/A _4531_/Y _4794_/Y VGND VGND VPWR VPWR _4795_/X sky130_fd_sc_hd__a211o_1
XANTENNA_46 _4772_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_57 _4939_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_68 _5200_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6534_ _6850_/B _6887_/B _6533_/Y _6967_/C _6449_/B VGND VGND VPWR VPWR _6539_/C
+ sky130_fd_sc_hd__o32a_1
X_9322_ _9370_/CLK _9322_/D fanout475/X VGND VGND VPWR VPWR _9322_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_79 _5311_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9253_ _9487_/CLK _9253_/D fanout411/X VGND VGND VPWR VPWR _9253_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_137_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6465_ _6651_/A _6874_/A VGND VGND VPWR VPWR _6976_/C sky130_fd_sc_hd__nor2_2
X_5416_ _8816_/Q _5415_/X _5416_/S VGND VGND VPWR VPWR _5416_/X sky130_fd_sc_hd__mux2_1
X_8204_ _8904_/Q _7962_/X _7988_/X _8939_/Q VGND VGND VPWR VPWR _8204_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9184_ _9184_/CLK _9184_/D fanout443/X VGND VGND VPWR VPWR _9184_/Q sky130_fd_sc_hd__dfstp_2
X_6396_ _6402_/A _6396_/B VGND VGND VPWR VPWR _6466_/A sky130_fd_sc_hd__nand2_1
XFILLER_161_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8135_ _9326_/Q _7962_/A _7988_/A _9438_/Q VGND VGND VPWR VPWR _8135_/X sky130_fd_sc_hd__a22o_1
X_5347_ _5353_/A _5356_/B VGND VGND VPWR VPWR _5348_/A sky130_fd_sc_hd__and2_1
XFILLER_102_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8066_ _9203_/Q _7938_/A _7969_/X _9291_/Q VGND VGND VPWR VPWR _8066_/X sky130_fd_sc_hd__a22o_1
X_5278_ _5278_/A VGND VGND VPWR VPWR _5278_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7017_ _7025_/A _7025_/B VGND VGND VPWR VPWR _7018_/A sky130_fd_sc_hd__and2_1
XFILLER_87_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8968_ _9467_/CLK _8968_/D fanout476/X VGND VGND VPWR VPWR _8968_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7919_ _9163_/Q _7902_/A _7919_/A3 _5155_/X _7918_/X VGND VGND VPWR VPWR _9506_/D
+ sky130_fd_sc_hd__o311a_1
X_8899_ _9442_/CLK _8899_/D fanout436/X VGND VGND VPWR VPWR _8899_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_102_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput11 mask_rev_in[16] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__clkbuf_1
Xinput22 mask_rev_in[26] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4580_ _5277_/A _4811_/A _7211_/A _9205_/Q VGND VGND VPWR VPWR _4580_/X sky130_fd_sc_hd__a22o_1
XFILLER_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput33 mask_rev_in[7] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput44 mgmt_gpio_in[17] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__clkbuf_2
Xinput55 mgmt_gpio_in[27] VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput66 mgmt_gpio_in[37] VGND VGND VPWR VPWR _9555_/A sky130_fd_sc_hd__buf_4
Xinput77 ser_tx VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__clkbuf_1
Xhold806 _7205_/X VGND VGND VPWR VPWR _7206_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold817 _5466_/X VGND VGND VPWR VPWR _5467_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold828 _8832_/Q VGND VGND VPWR VPWR hold828/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput88 spimemio_flash_io1_oeb VGND VGND VPWR VPWR _5174_/B sky130_fd_sc_hd__buf_2
Xinput99 sram_ro_data[15] VGND VGND VPWR VPWR input99/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold839 _5476_/X VGND VGND VPWR VPWR _5477_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6250_ _6568_/A _6250_/B _6250_/C _6250_/D VGND VGND VPWR VPWR _6250_/X sky130_fd_sc_hd__and4b_1
X_5201_ _9171_/Q input78/X _5279_/B VGND VGND VPWR VPWR _5202_/A sky130_fd_sc_hd__mux2_4
XFILLER_131_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6181_ _6181_/A _6181_/B VGND VGND VPWR VPWR _6850_/A sky130_fd_sc_hd__nand2_8
XFILLER_170_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5132_ _9497_/Q _9498_/Q VGND VGND VPWR VPWR _8375_/A sky130_fd_sc_hd__nor2b_2
XFILLER_69_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5063_ _5065_/A1 hold11/X _5065_/S VGND VGND VPWR VPWR _5064_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8822_ _9487_/CLK _8822_/D fanout412/X VGND VGND VPWR VPWR _8822_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_65_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8753_ _8752_/X hold112/X _8765_/S VGND VGND VPWR VPWR _8754_/A sky130_fd_sc_hd__mux2_1
X_5965_ _5965_/A VGND VGND VPWR VPWR _9054_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7704_ _7651_/X hold370/X _7710_/S VGND VGND VPWR VPWR _7705_/A sky130_fd_sc_hd__mux2_1
X_4916_ _5453_/B _7111_/B VGND VGND VPWR VPWR _7108_/A sky130_fd_sc_hd__nor2_1
XFILLER_80_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8684_ _8922_/Q _8360_/A _8381_/A _8957_/Q VGND VGND VPWR VPWR _8684_/X sky130_fd_sc_hd__a22o_1
X_5896_ _5896_/A VGND VGND VPWR VPWR _5896_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7635_ _7635_/A VGND VGND VPWR VPWR _9389_/D sky130_fd_sc_hd__clkbuf_1
X_4847_ _9233_/Q _7284_/A _7605_/A _9377_/Q VGND VGND VPWR VPWR _4847_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4778_ _9298_/Q _7425_/A _7481_/A _9322_/Q _4777_/X VGND VGND VPWR VPWR _4781_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7566_ _7566_/A VGND VGND VPWR VPWR _9357_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9305_ _9305_/CLK _9305_/D fanout468/X VGND VGND VPWR VPWR _9305_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_165_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6517_ _6517_/A _6517_/B _6517_/C _6517_/D VGND VGND VPWR VPWR _6517_/X sky130_fd_sc_hd__or4_1
XFILLER_134_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7497_ _7299_/X hold564/X _7497_/S VGND VGND VPWR VPWR _7497_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9236_ _9328_/CLK _9236_/D fanout463/X VGND VGND VPWR VPWR _9236_/Q sky130_fd_sc_hd__dfrtp_4
X_6448_ _6436_/Y _6462_/B _6842_/B _6447_/X VGND VGND VPWR VPWR _6455_/C sky130_fd_sc_hd__a211o_1
XFILLER_134_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6379_ _6716_/A _6672_/B VGND VGND VPWR VPWR _6393_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9167_ _9167_/CLK _9167_/D fanout484/X VGND VGND VPWR VPWR _9167_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8118_ _9341_/Q _7933_/X _7988_/X _9437_/Q VGND VGND VPWR VPWR _8118_/X sky130_fd_sc_hd__a22o_1
XFILLER_102_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9098_ _9484_/CLK _9098_/D fanout428/X VGND VGND VPWR VPWR _9098_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_130_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8049_ _9218_/Q _7927_/A _7956_/A _9306_/Q _8048_/X VGND VGND VPWR VPWR _8050_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_180_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5750_ _5750_/A _7132_/B VGND VGND VPWR VPWR _5759_/S sky130_fd_sc_hd__and2_4
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4701_ _9483_/Q _4898_/A2 _7678_/A _9411_/Q _4700_/X VGND VGND VPWR VPWR _4702_/D
+ sky130_fd_sc_hd__a221o_2
X_5681_ hold588/X _5587_/X _5691_/S VGND VGND VPWR VPWR _5682_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4632_ _9452_/Q _4836_/A2 _5750_/A _8962_/Q _4631_/X VGND VGND VPWR VPWR _4633_/D
+ sky130_fd_sc_hd__a221o_1
X_7420_ _7420_/A VGND VGND VPWR VPWR _9293_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4563_ _9245_/Q _4449_/Y _7056_/A _9137_/Q VGND VGND VPWR VPWR _4563_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7351_ _7351_/A VGND VGND VPWR VPWR _9261_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold603 _9407_/Q VGND VGND VPWR VPWR hold603/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6302_ _6891_/A _6317_/A VGND VGND VPWR VPWR _6303_/A sky130_fd_sc_hd__or2_1
Xhold614 _5486_/X VGND VGND VPWR VPWR _5487_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7282_ _5471_/X hold624/X _7282_/S VGND VGND VPWR VPWR _7282_/X sky130_fd_sc_hd__mux2_1
Xhold625 _7282_/X VGND VGND VPWR VPWR _7283_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4494_ input99/X _4488_/Y _4582_/A input51/X _4493_/X VGND VGND VPWR VPWR _4495_/D
+ sky130_fd_sc_hd__a221o_1
Xhold636 _9335_/Q VGND VGND VPWR VPWR hold636/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 _7586_/X VGND VGND VPWR VPWR _7587_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap366 _4409_/Y VGND VGND VPWR VPWR _7339_/A sky130_fd_sc_hd__buf_8
Xhold658 _5914_/X VGND VGND VPWR VPWR _5915_/A sky130_fd_sc_hd__dlygate4sd3_1
X_9021_ _9419_/CLK _9021_/D fanout491/X VGND VGND VPWR VPWR _9582_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_89_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6233_ _6233_/A VGND VGND VPWR VPWR _6603_/A sky130_fd_sc_hd__buf_4
Xmax_cap377 _4449_/Y VGND VGND VPWR VPWR _7304_/A sky130_fd_sc_hd__buf_6
XFILLER_116_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold669 _7372_/X VGND VGND VPWR VPWR _7373_/A sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap388 _4484_/Y VGND VGND VPWR VPWR _7661_/A sky130_fd_sc_hd__buf_6
XFILLER_171_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap399 _4465_/B VGND VGND VPWR VPWR _4555_/B sky130_fd_sc_hd__buf_4
XFILLER_170_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6164_ _6895_/A _6894_/B VGND VGND VPWR VPWR _6708_/A sky130_fd_sc_hd__nor2_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5115_ _8793_/Q hold17/A _7025_/B VGND VGND VPWR VPWR _5115_/X sky130_fd_sc_hd__o21a_4
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6095_ _6181_/A _6095_/B VGND VGND VPWR VPWR _6724_/A sky130_fd_sc_hd__xor2_2
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5046_ _8790_/Q _5045_/A _5045_/Y _5047_/A VGND VGND VPWR VPWR _5046_/X sky130_fd_sc_hd__o22a_1
XFILLER_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8805_ _5168_/A1 _8805_/D _5379_/X VGND VGND VPWR VPWR _8805_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6997_ _6997_/A _6997_/B _6997_/C _6997_/D VGND VGND VPWR VPWR _6998_/B sky130_fd_sc_hd__or4_1
XFILLER_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8736_ _8736_/A VGND VGND VPWR VPWR _8765_/S sky130_fd_sc_hd__buf_2
XFILLER_41_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5948_ _5948_/A _7043_/B VGND VGND VPWR VPWR _5958_/S sky130_fd_sc_hd__nand2_4
XFILLER_179_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8667_ _8876_/Q _8316_/X _8327_/X _9092_/Q VGND VGND VPWR VPWR _8667_/X sky130_fd_sc_hd__a22o_1
X_5879_ _9177_/Q hold37/X _5897_/S VGND VGND VPWR VPWR hold70/A sky130_fd_sc_hd__mux2_1
XFILLER_178_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7618_ _7618_/A VGND VGND VPWR VPWR _9381_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8598_ _8938_/Q _7908_/X _8335_/X _8868_/Q VGND VGND VPWR VPWR _8598_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7549_ _7494_/X hold746/X _7551_/S VGND VGND VPWR VPWR _7549_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9219_ _9219_/CLK _9219_/D fanout469/X VGND VGND VPWR VPWR _9219_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_161_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput201 wb_stb_i VGND VGND VPWR VPWR _5123_/D sky130_fd_sc_hd__buf_2
XFILLER_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6920_ _9108_/Q _8735_/A _6908_/X _6919_/X VGND VGND VPWR VPWR _6953_/A sky130_fd_sc_hd__a22o_1
XFILLER_35_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6851_ _6851_/A _6851_/B _6851_/C _6851_/D VGND VGND VPWR VPWR _6993_/C sky130_fd_sc_hd__or4_1
XFILLER_35_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5802_ _5650_/X hold406/X _5804_/S VGND VGND VPWR VPWR _5803_/A sky130_fd_sc_hd__mux2_1
X_9570_ _9570_/A _5098_/Y VGND VGND VPWR VPWR mgmt_gpio_out[16] sky130_fd_sc_hd__ebufn_8
X_6782_ _6241_/B _6874_/A _6780_/X _6781_/X VGND VGND VPWR VPWR _6782_/X sky130_fd_sc_hd__o211a_1
X_8521_ _9237_/Q _8322_/X _8333_/X _9269_/Q _8520_/X VGND VGND VPWR VPWR _8524_/C
+ sky130_fd_sc_hd__a221o_1
X_5733_ _5733_/A VGND VGND VPWR VPWR _8950_/D sky130_fd_sc_hd__clkbuf_1
X_8452_ _5139_/A _9521_/Q _8013_/X VGND VGND VPWR VPWR _8452_/X sky130_fd_sc_hd__a21o_1
XFILLER_148_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5664_ _5664_/A VGND VGND VPWR VPWR _8921_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7403_ _7403_/A VGND VGND VPWR VPWR _9285_/D sky130_fd_sc_hd__clkbuf_1
X_4615_ _9444_/Q _7746_/A _5551_/A _8877_/Q VGND VGND VPWR VPWR _4615_/X sky130_fd_sc_hd__a22o_1
XFILLER_129_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5595_ _5595_/A VGND VGND VPWR VPWR _8892_/D sky130_fd_sc_hd__clkbuf_1
X_8383_ _9424_/Q _8376_/X _8378_/X _9352_/Q _8382_/X VGND VGND VPWR VPWR _8396_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold400 _8861_/Q VGND VGND VPWR VPWR hold400/X sky130_fd_sc_hd__dlygate4sd3_1
X_4546_ _9430_/Q _7712_/A _4406_/Y input9/X VGND VGND VPWR VPWR _4546_/X sky130_fd_sc_hd__a22o_1
X_7334_ _7334_/A VGND VGND VPWR VPWR _9253_/D sky130_fd_sc_hd__clkbuf_1
Xhold411 _9082_/Q VGND VGND VPWR VPWR hold411/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold422 hold422/A VGND VGND VPWR VPWR hold422/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold433 _5761_/A VGND VGND VPWR VPWR _7126_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 hold444/A VGND VGND VPWR VPWR hold444/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 hold455/A VGND VGND VPWR VPWR hold455/X sky130_fd_sc_hd__dlygate4sd3_1
X_4477_ _4499_/A _4667_/B VGND VGND VPWR VPWR _4477_/Y sky130_fd_sc_hd__nor2_8
X_7265_ _7265_/A VGND VGND VPWR VPWR _9223_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold466 hold466/A VGND VGND VPWR VPWR hold466/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 _8849_/Q VGND VGND VPWR VPWR hold477/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold488 _9450_/Q VGND VGND VPWR VPWR hold488/X sky130_fd_sc_hd__dlygate4sd3_1
X_9004_ _9006_/CLK _9004_/D fanout493/X VGND VGND VPWR VPWR _9566_/A sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_69_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _9069_/CLK sky130_fd_sc_hd__clkbuf_16
X_6216_ _6216_/A _6262_/A VGND VGND VPWR VPWR _6217_/B sky130_fd_sc_hd__nor2_2
Xhold499 _9449_/Q VGND VGND VPWR VPWR hold499/X sky130_fd_sc_hd__dlygate4sd3_1
X_7196_ _7196_/A VGND VGND VPWR VPWR _9192_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6147_ _6167_/B _6167_/C VGND VGND VPWR VPWR _6324_/A sky130_fd_sc_hd__nand2_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1100 _8893_/Q VGND VGND VPWR VPWR hold913/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1111 _8891_/Q VGND VGND VPWR VPWR hold667/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1122 _8944_/Q VGND VGND VPWR VPWR hold796/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1133 _9466_/Q VGND VGND VPWR VPWR hold725/A sky130_fd_sc_hd__dlygate4sd3_1
X_6078_ _6078_/A _6078_/B _6078_/C _6078_/D VGND VGND VPWR VPWR _6170_/B sky130_fd_sc_hd__and4_1
Xhold1144 _7137_/X VGND VGND VPWR VPWR hold868/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 _9398_/Q VGND VGND VPWR VPWR hold732/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1166 _9372_/Q VGND VGND VPWR VPWR hold270/A sky130_fd_sc_hd__dlygate4sd3_1
X_5029_ _8791_/Q _4972_/B _5029_/B1 VGND VGND VPWR VPWR _5031_/A sky130_fd_sc_hd__a21oi_1
Xhold1177 _8878_/Q VGND VGND VPWR VPWR hold932/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1188 _5297_/X VGND VGND VPWR VPWR _5298_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_306 _7391_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1199 _5898_/X VGND VGND VPWR VPWR hold1199/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_317 _5851_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_328 _5067_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_339 _5468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8719_ _9538_/Q _8719_/A1 _8725_/S VGND VGND VPWR VPWR _8720_/A sky130_fd_sc_hd__mux2_2
XFILLER_179_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4400_ _4425_/B _4465_/A VGND VGND VPWR VPWR _5474_/B sky130_fd_sc_hd__nand2_8
X_5380_ _5453_/C VGND VGND VPWR VPWR _7013_/B sky130_fd_sc_hd__buf_2
XFILLER_160_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7050_ _6015_/X _9129_/Q _7054_/S VGND VGND VPWR VPWR _7050_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6001_ hold645/X _5683_/X _6005_/S VGND VGND VPWR VPWR _6002_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7952_ _7952_/A VGND VGND VPWR VPWR _7953_/B sky130_fd_sc_hd__buf_6
XFILLER_82_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6903_ _6811_/B _6811_/C _6973_/B _6653_/A _6820_/Y VGND VGND VPWR VPWR _6903_/X
+ sky130_fd_sc_hd__a311o_1
X_7883_ _9495_/Q _7883_/B VGND VGND VPWR VPWR _7888_/S sky130_fd_sc_hd__nor2_1
XFILLER_23_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6834_ _6834_/A _6834_/B _6923_/A VGND VGND VPWR VPWR _6982_/B sky130_fd_sc_hd__and3_1
XFILLER_62_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9553_ _9553_/A VGND VGND VPWR VPWR _9553_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6765_ _6948_/A _6987_/B _6931_/B VGND VGND VPWR VPWR _6770_/B sky130_fd_sc_hd__or3_1
X_8504_ _9469_/Q _8312_/X _8376_/X _9429_/Q VGND VGND VPWR VPWR _8504_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5716_ hold941/X _5505_/X _5724_/S VGND VGND VPWR VPWR _5717_/A sky130_fd_sc_hd__mux2_1
X_9484_ _9484_/CLK _9484_/D fanout429/X VGND VGND VPWR VPWR _9484_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_148_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6696_ _6495_/B _6967_/B _6779_/C _6779_/A VGND VGND VPWR VPWR _6697_/B sky130_fd_sc_hd__o22a_1
XFILLER_109_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8435_ _9298_/Q _8314_/X _8331_/X _9402_/Q VGND VGND VPWR VPWR _8435_/X sky130_fd_sc_hd__a22o_1
X_5647_ _7645_/A VGND VGND VPWR VPWR _5647_/X sky130_fd_sc_hd__buf_4
XFILLER_191_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8366_ _8650_/A VGND VGND VPWR VPWR _8701_/A sky130_fd_sc_hd__clkbuf_8
X_5578_ _5306_/X hold542/X _5582_/S VGND VGND VPWR VPWR _5578_/X sky130_fd_sc_hd__mux2_1
Xhold230 _7634_/X VGND VGND VPWR VPWR _7635_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7317_ _7279_/X hold762/X _7319_/S VGND VGND VPWR VPWR _7317_/X sky130_fd_sc_hd__mux2_1
Xhold241 hold241/A VGND VGND VPWR VPWR hold241/X sky130_fd_sc_hd__dlygate4sd3_1
X_4529_ _4529_/A1 _4502_/Y _7781_/A _9462_/Q _4528_/X VGND VGND VPWR VPWR _4530_/D
+ sky130_fd_sc_hd__a221o_1
Xhold252 _9429_/Q VGND VGND VPWR VPWR hold252/X sky130_fd_sc_hd__dlygate4sd3_1
X_8297_ _8385_/A _8359_/B VGND VGND VPWR VPWR _8298_/A sky130_fd_sc_hd__nor2_2
Xhold263 _7510_/X VGND VGND VPWR VPWR _7511_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 _7385_/X VGND VGND VPWR VPWR _7386_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold285 hold285/A VGND VGND VPWR VPWR hold285/X sky130_fd_sc_hd__dlygate4sd3_1
X_7248_ _7248_/A VGND VGND VPWR VPWR _9215_/D sky130_fd_sc_hd__clkbuf_1
Xhold296 _7231_/X VGND VGND VPWR VPWR _7232_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7179_ _7179_/A VGND VGND VPWR VPWR _9184_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 _5951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_114 _6018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_125 _7233_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_136 _7830_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 _7923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_158 _7947_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_169 _7960_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 mask_rev_in[14] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4880_ input47/X _4811_/A _4502_/Y _4880_/B2 _4879_/X VGND VGND VPWR VPWR _4883_/C
+ sky130_fd_sc_hd__a221o_4
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6550_ _6894_/A _6894_/B VGND VGND VPWR VPWR _6582_/C sky130_fd_sc_hd__nor2_1
XFILLER_192_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5501_ _5501_/A VGND VGND VPWR VPWR _8851_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6481_ _6481_/A _6609_/B VGND VGND VPWR VPWR _6772_/B sky130_fd_sc_hd__nand2_1
XFILLER_146_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8220_ _9081_/Q _7949_/X _7988_/X _8940_/Q VGND VGND VPWR VPWR _8220_/X sky130_fd_sc_hd__a22o_1
X_5432_ hold27/X VGND VGND VPWR VPWR _7494_/A sky130_fd_sc_hd__buf_4
Xoutput302 _9143_/Q VGND VGND VPWR VPWR pwr_ctrl_out[2] sky130_fd_sc_hd__buf_12
XFILLER_133_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput313 _5182_/X VGND VGND VPWR VPWR spimemio_flash_io1_di sky130_fd_sc_hd__buf_12
Xoutput324 _9145_/Q VGND VGND VPWR VPWR sram_ro_clk sky130_fd_sc_hd__buf_12
X_5363_ _5375_/A _5378_/B VGND VGND VPWR VPWR _5364_/A sky130_fd_sc_hd__and2_1
X_8151_ _5130_/A _9512_/Q _8013_/A _8150_/X VGND VGND VPWR VPWR _8151_/X sky130_fd_sc_hd__a211o_1
XFILLER_126_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput335 _9041_/Q VGND VGND VPWR VPWR wb_dat_o[17] sky130_fd_sc_hd__buf_12
Xoutput346 _9537_/Q VGND VGND VPWR VPWR wb_dat_o[27] sky130_fd_sc_hd__buf_12
XFILLER_114_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7102_ _5465_/X _9152_/Q _7106_/S VGND VGND VPWR VPWR _7102_/X sky130_fd_sc_hd__mux2_1
Xoutput357 _9053_/Q VGND VGND VPWR VPWR wb_dat_o[8] sky130_fd_sc_hd__buf_12
X_5294_ hold19/X VGND VGND VPWR VPWR hold20/A sky130_fd_sc_hd__buf_8
XFILLER_87_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8082_ _8082_/A _8082_/B _8082_/C _8082_/D VGND VGND VPWR VPWR _8082_/X sky130_fd_sc_hd__or4_2
XFILLER_114_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7033_ _5947_/X _9121_/Q _7041_/S VGND VGND VPWR VPWR _7033_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8984_ _9084_/CLK _8984_/D fanout445/X VGND VGND VPWR VPWR _8984_/Q sky130_fd_sc_hd__dfrtp_4
X_7935_ _9208_/Q _7923_/X _7927_/X _9216_/Q _7934_/X VGND VGND VPWR VPWR _7965_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7866_ _7866_/A VGND VGND VPWR VPWR _9490_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6817_ _6918_/B _6917_/C VGND VGND VPWR VPWR _6817_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7797_ _7797_/A VGND VGND VPWR VPWR _9463_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9536_ _9541_/CLK _9536_/D VGND VGND VPWR VPWR _9536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6748_ _6876_/B _6748_/B VGND VGND VPWR VPWR _6859_/C sky130_fd_sc_hd__nor2_1
XFILLER_51_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9467_ _9467_/CLK _9467_/D fanout476/X VGND VGND VPWR VPWR _9467_/Q sky130_fd_sc_hd__dfrtp_4
X_6679_ _6503_/A _6441_/B _6460_/B _6935_/A VGND VGND VPWR VPWR _6704_/B sky130_fd_sc_hd__a31o_1
XFILLER_164_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8418_ _9225_/Q _8388_/X _8379_/X _9201_/Q _8417_/X VGND VGND VPWR VPWR _8423_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_164_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9398_ _9398_/CLK _9398_/D _5332_/A VGND VGND VPWR VPWR _9398_/Q sky130_fd_sc_hd__dfrtp_2
X_8349_ _9368_/Q _8346_/X _8348_/X _9456_/Q VGND VGND VPWR VPWR _8349_/X sky130_fd_sc_hd__a22o_1
XFILLER_105_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5981_ _5981_/A VGND VGND VPWR VPWR _9061_/D sky130_fd_sc_hd__clkbuf_1
X_7720_ _7720_/A VGND VGND VPWR VPWR _9427_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4932_ _8873_/Q _5551_/A _5727_/A _8948_/Q VGND VGND VPWR VPWR _4932_/X sky130_fd_sc_hd__a22o_1
XFILLER_33_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7651_ hold24/X VGND VGND VPWR VPWR _7651_/X sky130_fd_sc_hd__buf_4
XFILLER_32_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4863_ _9133_/Q _7056_/A _5437_/A _8826_/Q _4862_/X VGND VGND VPWR VPWR _4864_/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA_14 _7605_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6602_ _6345_/X _6507_/A _6597_/A _6518_/Y VGND VGND VPWR VPWR _6946_/A sky130_fd_sc_hd__a22o_1
XANTENNA_25 _4542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7582_ _7439_/X hold248/X hold78/X VGND VGND VPWR VPWR _7582_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4794_ _7111_/B _4794_/B VGND VGND VPWR VPWR _4794_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_36 _5529_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_47 _4791_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 _4939_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9321_ _9459_/CLK _9321_/D fanout479/X VGND VGND VPWR VPWR _9321_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA_69 _5204_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6533_ _6402_/A _6973_/A _6498_/B _6628_/A VGND VGND VPWR VPWR _6533_/Y sky130_fd_sc_hd__o211ai_2
X_9252_ _9420_/CLK _9252_/D fanout463/X VGND VGND VPWR VPWR _9252_/Q sky130_fd_sc_hd__dfrtp_1
X_6464_ _6495_/B _6815_/B _6898_/A VGND VGND VPWR VPWR _6467_/B sky130_fd_sc_hd__a21oi_1
X_8203_ _9085_/Q _7940_/X _7969_/X _8879_/Q _8202_/X VGND VGND VPWR VPWR _8209_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5415_ _7514_/A VGND VGND VPWR VPWR _5415_/X sky130_fd_sc_hd__clkbuf_4
X_9183_ _9251_/CLK _9183_/D fanout486/X VGND VGND VPWR VPWR _9183_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6395_ _6628_/A _6440_/A VGND VGND VPWR VPWR _6396_/B sky130_fd_sc_hd__nor2_1
X_8134_ _9254_/Q _7940_/A _7969_/A _9294_/Q _8133_/X VGND VGND VPWR VPWR _8140_/B
+ sky130_fd_sc_hd__a221o_1
X_5346_ _5346_/A VGND VGND VPWR VPWR _5346_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8065_ _9219_/Q _7927_/X _7977_/X _9395_/Q _8064_/X VGND VGND VPWR VPWR _8072_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_141_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5277_ _5277_/A _5277_/B VGND VGND VPWR VPWR _5278_/A sky130_fd_sc_hd__and2_1
XFILLER_102_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7016_ _7016_/A VGND VGND VPWR VPWR _7016_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8967_ _9482_/CLK _8967_/D fanout432/X VGND VGND VPWR VPWR _8967_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_71_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7918_ _8996_/Q _7916_/C _9506_/Q VGND VGND VPWR VPWR _7918_/X sky130_fd_sc_hd__a21o_1
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8898_ _9473_/CLK _8898_/D fanout436/X VGND VGND VPWR VPWR _8898_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_169_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7849_ _8997_/Q _8998_/Q VGND VGND VPWR VPWR _8015_/B sky130_fd_sc_hd__nor2_1
XFILLER_169_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9519_ _9529_/CLK _9519_/D fanout446/X VGND VGND VPWR VPWR _9519_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_7_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_0_mgmt_gpio_in[4] clkbuf_2_1_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _5168_/A1
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_59_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput12 mask_rev_in[17] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__clkbuf_1
Xinput23 mask_rev_in[27] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__clkbuf_1
Xinput34 mask_rev_in[8] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput45 mgmt_gpio_in[18] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__buf_2
Xinput56 mgmt_gpio_in[28] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold807 _7094_/X VGND VGND VPWR VPWR _7095_/A sky130_fd_sc_hd__dlygate4sd3_1
Xinput67 mgmt_gpio_in[3] VGND VGND VPWR VPWR _5071_/C sky130_fd_sc_hd__buf_6
Xinput78 spi_csb VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__clkbuf_1
Xhold818 _7156_/X VGND VGND VPWR VPWR _7157_/A sky130_fd_sc_hd__dlygate4sd3_1
Xinput89 spimemio_flash_io2_do VGND VGND VPWR VPWR input89/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold829 _5455_/X VGND VGND VPWR VPWR _5456_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5200_ _5200_/A VGND VGND VPWR VPWR _9586_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6180_ _6182_/A VGND VGND VPWR VPWR _6398_/B sky130_fd_sc_hd__inv_2
XFILLER_184_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5131_ _9501_/Q _9502_/Q VGND VGND VPWR VPWR _8355_/A sky130_fd_sc_hd__nand2b_4
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5062_ _5062_/A VGND VGND VPWR VPWR _8783_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8821_ _9484_/CLK _8821_/D fanout430/X VGND VGND VPWR VPWR _8821_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_65_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8752_ _5271_/A _8752_/A2 _8752_/B1 _8727_/Y _8751_/X VGND VGND VPWR VPWR _8752_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5964_ _9054_/Q _4885_/X _5976_/S VGND VGND VPWR VPWR _5965_/A sky130_fd_sc_hd__mux2_1
X_7703_ _7703_/A VGND VGND VPWR VPWR _9419_/D sky130_fd_sc_hd__clkbuf_1
X_4915_ _4915_/A VGND VGND VPWR VPWR _4915_/X sky130_fd_sc_hd__clkbuf_2
X_8683_ _8937_/Q _8386_/X _8506_/B _8972_/Q _8682_/X VGND VGND VPWR VPWR _8688_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5895_ _9015_/Q _5894_/X _5898_/S VGND VGND VPWR VPWR _5895_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7634_ _7439_/X hold229/X _7638_/S VGND VGND VPWR VPWR _7634_/X sky130_fd_sc_hd__mux2_1
X_4846_ _8934_/Q _5693_/A _5493_/A _8849_/Q VGND VGND VPWR VPWR _4852_/A sky130_fd_sc_hd__a22o_1
XFILLER_138_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7565_ _7439_/X hold233/X hold99/A VGND VGND VPWR VPWR _7565_/X sky130_fd_sc_hd__mux2_1
X_4777_ _8890_/Q _5584_/A _5750_/A _8960_/Q VGND VGND VPWR VPWR _4777_/X sky130_fd_sc_hd__a22o_1
X_9304_ _9464_/CLK _9304_/D fanout420/X VGND VGND VPWR VPWR _9304_/Q sky130_fd_sc_hd__dfstp_2
X_6516_ _6597_/A _6514_/Y _6643_/B VGND VGND VPWR VPWR _6517_/D sky130_fd_sc_hd__a21o_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7496_ _7496_/A VGND VGND VPWR VPWR _9326_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9235_ _9283_/CLK _9235_/D fanout484/X VGND VGND VPWR VPWR _9235_/Q sky130_fd_sc_hd__dfrtp_4
X_6447_ _6436_/Y _6445_/Y _6446_/X VGND VGND VPWR VPWR _6447_/X sky130_fd_sc_hd__a21o_1
XFILLER_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9166_ _9167_/CLK _9166_/D fanout484/X VGND VGND VPWR VPWR _9166_/Q sky130_fd_sc_hd__dfrtp_2
X_6378_ _6867_/A _6585_/B _6369_/X _6754_/C _6377_/X VGND VGND VPWR VPWR _6378_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_121_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8117_ _8117_/A _8117_/B _8117_/C _8117_/D VGND VGND VPWR VPWR _8117_/X sky130_fd_sc_hd__or4_1
XFILLER_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5329_ _5329_/A VGND VGND VPWR VPWR _5329_/X sky130_fd_sc_hd__clkbuf_1
X_9097_ _9473_/CLK _9097_/D fanout431/X VGND VGND VPWR VPWR _9097_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8048_ _9314_/Q _7983_/A _7977_/A _9394_/Q _7984_/X VGND VGND VPWR VPWR _8048_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_75_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4700_ _9339_/Q _7519_/A _7712_/A _9427_/Q VGND VGND VPWR VPWR _4700_/X sky130_fd_sc_hd__a22o_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ _5680_/A VGND VGND VPWR VPWR _8928_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4631_ _9188_/Q _7176_/A _5562_/A _8882_/Q VGND VGND VPWR VPWR _4631_/X sky130_fd_sc_hd__a22o_1
XFILLER_8_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7350_ _7242_/X hold297/X _7354_/S VGND VGND VPWR VPWR _7350_/X sky130_fd_sc_hd__mux2_1
X_4562_ _4562_/A VGND VGND VPWR VPWR _4562_/X sky130_fd_sc_hd__buf_2
XFILLER_116_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold604 _7676_/X VGND VGND VPWR VPWR _7677_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6301_ _6876_/B _6736_/A VGND VGND VPWR VPWR _6364_/A sky130_fd_sc_hd__nor2_1
XFILLER_190_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold615 _8970_/Q VGND VGND VPWR VPWR hold615/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold626 _9207_/Q VGND VGND VPWR VPWR hold626/X sky130_fd_sc_hd__dlygate4sd3_1
X_7281_ _7281_/A VGND VGND VPWR VPWR _9230_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4493_ input60/X _5901_/A _7249_/A _9223_/Q VGND VGND VPWR VPWR _4493_/X sky130_fd_sc_hd__a22o_1
Xhold637 _7515_/X VGND VGND VPWR VPWR _7516_/A sky130_fd_sc_hd__dlygate4sd3_1
X_9020_ _9419_/CLK _9020_/D fanout491/X VGND VGND VPWR VPWR _9581_/A sky130_fd_sc_hd__dfrtp_1
Xhold648 hold648/A VGND VGND VPWR VPWR hold648/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold659 _5915_/X VGND VGND VPWR VPWR _9023_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6232_ _6721_/A _6232_/B _6232_/C _6562_/A VGND VGND VPWR VPWR _6233_/A sky130_fd_sc_hd__or4_1
Xmax_cap378 _7374_/A VGND VGND VPWR VPWR _4938_/A2 sky130_fd_sc_hd__buf_6
Xmax_cap389 _7729_/A VGND VGND VPWR VPWR _4906_/A2 sky130_fd_sc_hd__buf_6
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6163_ _6635_/B VGND VGND VPWR VPWR _6894_/B sky130_fd_sc_hd__buf_2
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _5114_/A VGND VGND VPWR VPWR _7911_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_57_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6094_ _6716_/B _6243_/A VGND VGND VPWR VPWR _6732_/A sky130_fd_sc_hd__nand2_2
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _5045_/A _5045_/B VGND VGND VPWR VPWR _5045_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8804_ _5168_/A1 _8804_/D _5376_/X VGND VGND VPWR VPWR hold29/A sky130_fd_sc_hd__dfrtp_1
XFILLER_80_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6996_ _6419_/A _6521_/B _6812_/Y _6973_/C _6830_/Y VGND VGND VPWR VPWR _6997_/D
+ sky130_fd_sc_hd__a32o_1
X_8735_ _8735_/A _8735_/B _8735_/C _8734_/X VGND VGND VPWR VPWR _8736_/A sky130_fd_sc_hd__or4b_1
X_5947_ _7517_/A VGND VGND VPWR VPWR _5947_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_80_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8666_ _8911_/Q _8348_/X _8411_/X _8926_/Q _8665_/X VGND VGND VPWR VPWR _8676_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5878_ _5878_/A VGND VGND VPWR VPWR _5878_/X sky130_fd_sc_hd__clkbuf_1
X_7617_ hold305/X _5465_/A _7621_/S VGND VGND VPWR VPWR _7617_/X sky130_fd_sc_hd__mux2_1
X_4829_ _4829_/A _4829_/B _4829_/C _4829_/D VGND VGND VPWR VPWR _4885_/A sky130_fd_sc_hd__or4_2
XFILLER_21_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8597_ _9069_/Q _8388_/X _8379_/X _9035_/Q _8596_/X VGND VGND VPWR VPWR _8600_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_138_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7548_ _7548_/A VGND VGND VPWR VPWR _9349_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7479_ hold235/X _7514_/A _7479_/S VGND VGND VPWR VPWR _7480_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9218_ _9474_/CLK _9218_/D fanout429/X VGND VGND VPWR VPWR _9218_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_134_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9149_ _9485_/CLK _9149_/D fanout404/X VGND VGND VPWR VPWR _9149_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput202 wb_we_i VGND VGND VPWR VPWR _8732_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6850_ _6850_/A _6850_/B _6862_/B VGND VGND VPWR VPWR _6851_/B sky130_fd_sc_hd__nor3_1
X_5801_ _5801_/A VGND VGND VPWR VPWR _8980_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6781_ _6973_/A _6781_/B _6781_/C _6887_/A VGND VGND VPWR VPWR _6781_/X sky130_fd_sc_hd__or4_1
X_8520_ _9285_/Q _8316_/X _8327_/X _9261_/Q VGND VGND VPWR VPWR _8520_/X sky130_fd_sc_hd__a22o_1
X_5732_ _5647_/X hold597/X _5736_/S VGND VGND VPWR VPWR _5733_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8451_ _9186_/Q _8400_/B _8437_/X _8450_/X _8105_/X VGND VGND VPWR VPWR _8451_/X
+ sky130_fd_sc_hd__o221a_1
X_5663_ hold421/X _5398_/X _5665_/S VGND VGND VPWR VPWR _5664_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7402_ _7242_/X hold279/X _7406_/S VGND VGND VPWR VPWR _7402_/X sky130_fd_sc_hd__mux2_1
X_4614_ _4656_/A _4685_/B VGND VGND VPWR VPWR _5551_/A sky130_fd_sc_hd__nor2_8
X_8382_ _9200_/Q _8379_/X _8381_/X _9360_/Q VGND VGND VPWR VPWR _8382_/X sky130_fd_sc_hd__a22o_1
X_5594_ hold804/X _5402_/X _5594_/S VGND VGND VPWR VPWR _5595_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold401 _5525_/X VGND VGND VPWR VPWR _5526_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7333_ hold293/X _5465_/A _7337_/S VGND VGND VPWR VPWR _7333_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4545_ _9318_/Q _7463_/A _7321_/A _9254_/Q _4544_/X VGND VGND VPWR VPWR _4548_/C
+ sky130_fd_sc_hd__a221o_1
Xhold412 _6028_/X VGND VGND VPWR VPWR _6029_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 hold423/A VGND VGND VPWR VPWR hold423/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 hold434/A VGND VGND VPWR VPWR _9156_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 _9077_/Q VGND VGND VPWR VPWR hold445/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7264_ _5471_/X hold670/X _7264_/S VGND VGND VPWR VPWR _7264_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold456 _8834_/Q VGND VGND VPWR VPWR hold456/X sky130_fd_sc_hd__dlygate4sd3_1
X_4476_ _4476_/A _4536_/B VGND VGND VPWR VPWR _4667_/B sky130_fd_sc_hd__nand2_8
XFILLER_131_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold467 hold467/A VGND VGND VPWR VPWR hold467/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 _5496_/X VGND VGND VPWR VPWR _5497_/A sky130_fd_sc_hd__dlygate4sd3_1
X_9003_ _9006_/CLK _9003_/D fanout493/X VGND VGND VPWR VPWR _9565_/A sky130_fd_sc_hd__dfrtp_2
Xhold489 _7769_/X VGND VGND VPWR VPWR _7770_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6215_ _6215_/A VGND VGND VPWR VPWR _6507_/A sky130_fd_sc_hd__clkbuf_4
X_7195_ _7128_/X hold908/X _7209_/S VGND VGND VPWR VPWR _7196_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6146_ _6334_/B _6876_/B VGND VGND VPWR VPWR _6588_/A sky130_fd_sc_hd__nor2_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1101 _8918_/Q VGND VGND VPWR VPWR hold930/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1112 _8909_/Q VGND VGND VPWR VPWR hold728/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1123 _9418_/Q VGND VGND VPWR VPWR hold724/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6077_ _6192_/A _6312_/A VGND VGND VPWR VPWR _6739_/A sky130_fd_sc_hd__or2_4
XFILLER_58_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1134 _8959_/Q VGND VGND VPWR VPWR hold467/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1145 _8976_/Q VGND VGND VPWR VPWR hold712/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_180_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1156 _8946_/Q VGND VGND VPWR VPWR hold678/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1167 _8967_/Q VGND VGND VPWR VPWR hold635/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1178 _8858_/Q VGND VGND VPWR VPWR hold891/A sky130_fd_sc_hd__dlygate4sd3_1
X_5028_ _5019_/A _5021_/X _8794_/Q VGND VGND VPWR VPWR _5028_/X sky130_fd_sc_hd__a21o_1
XFILLER_38_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1189 _7112_/X VGND VGND VPWR VPWR hold434/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_307 _7661_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_318 _8992_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_329 _5067_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6979_ _6972_/X _6998_/A _6978_/X VGND VGND VPWR VPWR _6979_/X sky130_fd_sc_hd__o21a_1
XFILLER_41_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8718_ _8718_/A VGND VGND VPWR VPWR _9537_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8649_ _8649_/A _8649_/B _8649_/C _8649_/D VGND VGND VPWR VPWR _8650_/C sky130_fd_sc_hd__or4_1
XFILLER_182_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold990 _9527_/Q VGND VGND VPWR VPWR hold990/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6000_ _6000_/A VGND VGND VPWR VPWR _9070_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7951_ _8181_/B _7991_/B _8002_/C VGND VGND VPWR VPWR _7952_/A sky130_fd_sc_hd__and3_1
XFILLER_48_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6902_ _6902_/A _6972_/A _6915_/B _6997_/B VGND VGND VPWR VPWR _6905_/B sky130_fd_sc_hd__or4_1
XFILLER_47_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7882_ _7929_/B _7880_/Y _7883_/B VGND VGND VPWR VPWR _9494_/D sky130_fd_sc_hd__o21ai_1
XFILLER_50_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6833_ _6871_/B _6764_/A _6831_/Y _6832_/X VGND VGND VPWR VPWR _6923_/A sky130_fd_sc_hd__o211a_1
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6764_ _6764_/A _6764_/B VGND VGND VPWR VPWR _6931_/B sky130_fd_sc_hd__nor2_1
X_8503_ hold954/X _8017_/X _8502_/X VGND VGND VPWR VPWR _8503_/X sky130_fd_sc_hd__o21a_1
X_5715_ _5715_/A _5715_/B VGND VGND VPWR VPWR _5724_/S sky130_fd_sc_hd__and2_2
XFILLER_176_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9483_ _9483_/CLK _9483_/D fanout474/X VGND VGND VPWR VPWR _9483_/Q sky130_fd_sc_hd__dfrtp_4
X_6695_ _6695_/A _6695_/B VGND VGND VPWR VPWR _6779_/C sky130_fd_sc_hd__or2_1
X_8434_ _9450_/Q _8310_/X _8381_/X _9362_/Q _8433_/X VGND VGND VPWR VPWR _8437_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5646_ _5646_/A VGND VGND VPWR VPWR _8914_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8365_ _8398_/A _8398_/B _8398_/C _8398_/D VGND VGND VPWR VPWR _8474_/A sky130_fd_sc_hd__nor4_1
XFILLER_163_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5577_ _5577_/A VGND VGND VPWR VPWR _8884_/D sky130_fd_sc_hd__clkbuf_1
Xhold220 _9469_/Q VGND VGND VPWR VPWR hold220/X sky130_fd_sc_hd__dlygate4sd3_1
X_7316_ _7316_/A VGND VGND VPWR VPWR _9245_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4528_ _9470_/Q _4447_/Y _7764_/A _9454_/Q VGND VGND VPWR VPWR _4528_/X sky130_fd_sc_hd__a22o_1
Xhold231 _9309_/Q VGND VGND VPWR VPWR hold231/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold242 _9217_/Q VGND VGND VPWR VPWR hold242/X sky130_fd_sc_hd__dlygate4sd3_1
X_8296_ _8375_/A _8392_/C VGND VGND VPWR VPWR _8359_/B sky130_fd_sc_hd__nand2_2
XFILLER_104_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold253 _7723_/X VGND VGND VPWR VPWR _7724_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 _9364_/Q VGND VGND VPWR VPWR hold264/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7247_ _5471_/X hold716/X _7247_/S VGND VGND VPWR VPWR _7247_/X sky130_fd_sc_hd__mux2_1
Xhold275 _9485_/Q VGND VGND VPWR VPWR hold275/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 _9212_/Q VGND VGND VPWR VPWR hold286/X sky130_fd_sc_hd__dlygate4sd3_1
X_4459_ _4665_/A _4670_/B VGND VGND VPWR VPWR _4459_/Y sky130_fd_sc_hd__nor2_4
XFILLER_49_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold297 _9261_/Q VGND VGND VPWR VPWR hold297/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7178_ hold827/X _7126_/C _7192_/S VGND VGND VPWR VPWR _7179_/A sky130_fd_sc_hd__mux2_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6129_ _6141_/A _6732_/A _6128_/X VGND VGND VPWR VPWR _6130_/A sky130_fd_sc_hd__or3b_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_104 _5951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_115 _6018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 _7282_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_137 _7866_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_148 _7923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_159 _7947_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_53_csclk _8954_/CLK VGND VGND VPWR VPWR _8955_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_68_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _9474_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_189_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5500_ hold419/X _5398_/X _5502_/S VGND VGND VPWR VPWR _5500_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6480_ _6850_/A _6818_/A VGND VGND VPWR VPWR _6609_/B sky130_fd_sc_hd__nor2_1
XFILLER_146_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5431_ _5431_/A VGND VGND VPWR VPWR _8822_/D sky130_fd_sc_hd__clkbuf_1
Xoutput303 _9144_/Q VGND VGND VPWR VPWR pwr_ctrl_out[3] sky130_fd_sc_hd__buf_12
X_8150_ _9190_/Q _8010_/B _8149_/X _8105_/X VGND VGND VPWR VPWR _8150_/X sky130_fd_sc_hd__o211a_1
Xoutput314 _9554_/X VGND VGND VPWR VPWR spimemio_flash_io2_di sky130_fd_sc_hd__buf_12
X_5362_ _5362_/A VGND VGND VPWR VPWR _5362_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput325 _9146_/Q VGND VGND VPWR VPWR sram_ro_csb sky130_fd_sc_hd__buf_12
Xoutput336 _9042_/Q VGND VGND VPWR VPWR wb_dat_o[18] sky130_fd_sc_hd__buf_12
X_7101_ _7101_/A VGND VGND VPWR VPWR _9151_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput347 _9538_/Q VGND VGND VPWR VPWR wb_dat_o[28] sky130_fd_sc_hd__buf_12
Xoutput358 _9054_/Q VGND VGND VPWR VPWR wb_dat_o[9] sky130_fd_sc_hd__buf_12
X_8081_ _9371_/Q _7960_/X _7967_/X _9411_/Q _8080_/X VGND VGND VPWR VPWR _8082_/D
+ sky130_fd_sc_hd__a221o_1
X_5293_ hold18/X hold74/A _5292_/X VGND VGND VPWR VPWR hold19/A sky130_fd_sc_hd__o21a_4
XFILLER_87_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7032_ _7032_/A _7043_/B VGND VGND VPWR VPWR _7041_/S sky130_fd_sc_hd__nand2_2
XFILLER_101_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8983_ _9089_/CLK _8983_/D fanout433/X VGND VGND VPWR VPWR _8983_/Q sky130_fd_sc_hd__dfrtp_2
X_7934_ _9400_/Q _7931_/X _7933_/X _9336_/Q VGND VGND VPWR VPWR _7934_/X sky130_fd_sc_hd__a22o_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7865_ _7865_/A _7865_/B _7865_/C VGND VGND VPWR VPWR _7866_/A sky130_fd_sc_hd__and3_1
XFILLER_35_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6816_ _6891_/A _6976_/B _6976_/D VGND VGND VPWR VPWR _6917_/C sky130_fd_sc_hd__a21oi_1
X_7796_ _5415_/X hold685/X _7796_/S VGND VGND VPWR VPWR _7796_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6747_ _6623_/Y _6742_/Y _6607_/Y VGND VGND VPWR VPWR _6857_/D sky130_fd_sc_hd__a21o_1
X_9535_ _9541_/CLK _9535_/D VGND VGND VPWR VPWR _9535_/Q sky130_fd_sc_hd__dfxtp_1
X_9466_ _9466_/CLK _9466_/D fanout475/X VGND VGND VPWR VPWR _9466_/Q sky130_fd_sc_hd__dfrtp_2
X_6678_ _6897_/B _6503_/A _6460_/B _6673_/B _6217_/B VGND VGND VPWR VPWR _6704_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_164_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8417_ hold90/A _8292_/X _8294_/X _9289_/Q VGND VGND VPWR VPWR _8417_/X sky130_fd_sc_hd__a22o_1
X_5629_ _7517_/A VGND VGND VPWR VPWR _5629_/X sky130_fd_sc_hd__buf_4
X_9397_ _9453_/CLK _9397_/D fanout461/X VGND VGND VPWR VPWR _9397_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8348_ _8360_/C VGND VGND VPWR VPWR _8348_/X sky130_fd_sc_hd__buf_6
XFILLER_183_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8279_ _8947_/Q _8020_/X _8003_/X _8887_/Q _8278_/X VGND VGND VPWR VPWR _8282_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_104_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5980_ _9061_/Q _4961_/X _5994_/S VGND VGND VPWR VPWR _5981_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4931_ _4931_/A _4931_/B _4931_/C _4931_/D VGND VGND VPWR VPWR _4939_/A sky130_fd_sc_hd__or4_1
XFILLER_45_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7650_ _7650_/A VGND VGND VPWR VPWR _9395_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4862_ input12/X _4500_/Y _6007_/A _9075_/Q VGND VGND VPWR VPWR _4862_/X sky130_fd_sc_hd__a22o_1
XFILLER_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6601_ _6419_/A _6609_/A _6597_/B _6882_/A VGND VGND VPWR VPWR _6616_/B sky130_fd_sc_hd__a31o_1
XFILLER_33_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_15 _7605_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7581_ _7581_/A VGND VGND VPWR VPWR _9364_/D sky130_fd_sc_hd__clkbuf_1
X_4793_ _4793_/A1 _4444_/Y _4450_/Y _9458_/Q _4792_/X VGND VGND VPWR VPWR _4797_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA_26 _4569_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_37 _5584_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 _4807_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9320_ _9328_/CLK _9320_/D fanout464/X VGND VGND VPWR VPWR _9320_/Q sky130_fd_sc_hd__dfstp_2
X_6532_ _6628_/B _6828_/B _6531_/X _6425_/X _6895_/A VGND VGND VPWR VPWR _6539_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_158_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_59 _4939_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9251_ _9251_/CLK _9251_/D fanout485/X VGND VGND VPWR VPWR _9251_/Q sky130_fd_sc_hd__dfrtp_4
X_6463_ _6463_/A _6463_/B VGND VGND VPWR VPWR _6467_/A sky130_fd_sc_hd__nand2_1
XFILLER_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8202_ _8874_/Q _7953_/B _8003_/X _8884_/Q VGND VGND VPWR VPWR _8202_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5414_ hold5/X VGND VGND VPWR VPWR _7514_/A sky130_fd_sc_hd__buf_6
X_9182_ _9464_/CLK _9182_/D fanout420/X VGND VGND VPWR VPWR _9182_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6394_ _6673_/B _6670_/B _6672_/C _6925_/B VGND VGND VPWR VPWR _6987_/A sky130_fd_sc_hd__a31o_1
X_8133_ _9286_/Q _7952_/A _8003_/A _9302_/Q VGND VGND VPWR VPWR _8133_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5345_ _5353_/A _5356_/B VGND VGND VPWR VPWR _5346_/A sky130_fd_sc_hd__and2_1
XFILLER_114_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8064_ _9323_/Q _7962_/X _8023_/B _9307_/Q VGND VGND VPWR VPWR _8064_/X sky130_fd_sc_hd__a22o_1
X_5276_ _5276_/A VGND VGND VPWR VPWR _9027_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7015_ _7025_/A _7025_/B VGND VGND VPWR VPWR _7016_/A sky130_fd_sc_hd__and2_1
XFILLER_102_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8966_ _9184_/CLK _8966_/D fanout439/X VGND VGND VPWR VPWR _8966_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_43_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7917_ _9489_/Q _7916_/X _7914_/S _9505_/Q VGND VGND VPWR VPWR _7917_/X sky130_fd_sc_hd__a2bb2o_1
X_8897_ _9484_/CLK _8897_/D fanout430/X VGND VGND VPWR VPWR _8897_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_169_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7848_ _7848_/A VGND VGND VPWR VPWR _9487_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7779_ _5415_/X hold653/X _7779_/S VGND VGND VPWR VPWR _7779_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9518_ _9531_/CLK _9518_/D fanout452/X VGND VGND VPWR VPWR _9518_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9449_ _9449_/CLK _9449_/D fanout474/X VGND VGND VPWR VPWR _9449_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_124_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput13 mask_rev_in[18] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput24 mask_rev_in[28] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput35 mask_rev_in[9] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__clkbuf_1
Xinput46 mgmt_gpio_in[19] VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__buf_2
Xinput57 mgmt_gpio_in[29] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__buf_2
XFILLER_6_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput68 mgmt_gpio_in[5] VGND VGND VPWR VPWR _5277_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_116_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold808 _7075_/X VGND VGND VPWR VPWR _7076_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold819 _7157_/X VGND VGND VPWR VPWR _9175_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput79 spi_enabled VGND VGND VPWR VPWR _5279_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_184_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5130_ _5130_/A VGND VGND VPWR VPWR _5139_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_69_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5061_ hold11/X hold44/X _5065_/S VGND VGND VPWR VPWR _5062_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8820_ _9484_/CLK _8820_/D fanout430/X VGND VGND VPWR VPWR _8820_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_92_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8751_ _5287_/A _8751_/A2 _8751_/B1 _5275_/A VGND VGND VPWR VPWR _8751_/X sky130_fd_sc_hd__a22o_1
XFILLER_92_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5963_ _5963_/A VGND VGND VPWR VPWR _9053_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4914_ _8795_/Q _8780_/Q _9155_/Q VGND VGND VPWR VPWR _4915_/A sky130_fd_sc_hd__or3_1
X_7702_ _7648_/X _9419_/Q _7710_/S VGND VGND VPWR VPWR _7702_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8682_ _8967_/Q _8682_/B VGND VGND VPWR VPWR _8682_/X sky130_fd_sc_hd__and2_1
X_5894_ _9182_/Q hold27/X _5897_/S VGND VGND VPWR VPWR _5894_/X sky130_fd_sc_hd__mux2_1
X_4845_ hold96/A _4438_/Y _4531_/Y _4842_/X _4844_/X VGND VGND VPWR VPWR _4853_/C
+ sky130_fd_sc_hd__a2111o_1
X_7633_ _7633_/A VGND VGND VPWR VPWR _9388_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7564_ _7564_/A VGND VGND VPWR VPWR _9356_/D sky130_fd_sc_hd__clkbuf_1
X_4776_ input54/X _5901_/A _6055_/A _9096_/Q _4775_/X VGND VGND VPWR VPWR _4781_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6515_ _6732_/B _6900_/A VGND VGND VPWR VPWR _6643_/B sky130_fd_sc_hd__nor2_2
X_9303_ _9303_/CLK _9303_/D fanout464/X VGND VGND VPWR VPWR _9303_/Q sky130_fd_sc_hd__dfrtp_4
X_7495_ _7494_/X hold754/X _7497_/S VGND VGND VPWR VPWR _7495_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9234_ _9466_/CLK _9234_/D fanout471/X VGND VGND VPWR VPWR _9234_/Q sky130_fd_sc_hd__dfrtp_4
X_6446_ _6510_/A _6839_/B _6597_/B VGND VGND VPWR VPWR _6446_/X sky130_fd_sc_hd__and3_2
X_9165_ _9167_/CLK _9165_/D fanout484/X VGND VGND VPWR VPWR _9165_/Q sky130_fd_sc_hd__dfrtp_4
X_6377_ _6850_/A _6790_/B _6376_/Y _9032_/Q VGND VGND VPWR VPWR _6377_/X sky130_fd_sc_hd__o31a_1
XFILLER_164_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8116_ _9221_/Q _7927_/X _7947_/X _9381_/Q _8115_/X VGND VGND VPWR VPWR _8117_/D
+ sky130_fd_sc_hd__a221o_1
X_5328_ _5330_/A _5334_/B VGND VGND VPWR VPWR _5329_/A sky130_fd_sc_hd__and2_1
X_9096_ _9473_/CLK _9096_/D fanout431/X VGND VGND VPWR VPWR _9096_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_88_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8047_ _9210_/Q _7923_/A _7997_/A _9362_/Q _8046_/X VGND VGND VPWR VPWR _8050_/C
+ sky130_fd_sc_hd__a221o_1
X_5259_ _9371_/Q VGND VGND VPWR VPWR _5259_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8949_ _9283_/CLK _8949_/D fanout485/X VGND VGND VPWR VPWR _8949_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_71_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4630_ _4656_/A _4667_/B VGND VGND VPWR VPWR _5562_/A sky130_fd_sc_hd__nor2_8
XFILLER_30_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4561_ _9519_/Q _9160_/Q _9162_/Q VGND VGND VPWR VPWR _4562_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6300_ _6311_/B _6365_/B VGND VGND VPWR VPWR _6955_/B sky130_fd_sc_hd__nor2_2
Xhold605 _8930_/Q VGND VGND VPWR VPWR hold605/X sky130_fd_sc_hd__dlygate4sd3_1
X_7280_ _7279_/X hold765/X _7282_/S VGND VGND VPWR VPWR _7280_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold616 hold616/A VGND VGND VPWR VPWR hold616/X sky130_fd_sc_hd__dlygate4sd3_1
X_4492_ _4492_/A _4492_/B VGND VGND VPWR VPWR _7249_/A sky130_fd_sc_hd__nor2_8
Xhold627 _7226_/X VGND VGND VPWR VPWR _7227_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 hold638/A VGND VGND VPWR VPWR hold638/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold649 _9471_/Q VGND VGND VPWR VPWR hold649/X sky130_fd_sc_hd__dlygate4sd3_1
X_6231_ _6967_/A _6227_/Y _6228_/Y _6230_/X VGND VGND VPWR VPWR _6856_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_89_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap379 _4447_/Y VGND VGND VPWR VPWR _7798_/A sky130_fd_sc_hd__buf_6
XFILLER_131_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6162_ _6906_/C _6535_/A VGND VGND VPWR VPWR _6635_/B sky130_fd_sc_hd__or2_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _9504_/Q _9157_/Q _9162_/Q VGND VGND VPWR VPWR _5114_/A sky130_fd_sc_hd__mux2_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _6182_/A _6093_/B VGND VGND VPWR VPWR _6243_/A sky130_fd_sc_hd__xnor2_2
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5044_ _8788_/Q _5050_/B VGND VGND VPWR VPWR _5045_/B sky130_fd_sc_hd__nor2_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8803_ _5168_/A1 _8803_/D _5374_/X VGND VGND VPWR VPWR hold55/A sky130_fd_sc_hd__dfrtp_1
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6995_ _6951_/B _6970_/D _6993_/X _6965_/Y _6994_/Y VGND VGND VPWR VPWR _7009_/A
+ sky130_fd_sc_hd__o311a_1
X_8734_ _8732_/A _8734_/A2 _9030_/Q VGND VGND VPWR VPWR _8734_/X sky130_fd_sc_hd__a21bo_1
XFILLER_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5946_ _5946_/A VGND VGND VPWR VPWR _9047_/D sky130_fd_sc_hd__clkbuf_1
X_8665_ _8861_/Q _8391_/X _8367_/X _9097_/Q _8664_/X VGND VGND VPWR VPWR _8665_/X
+ sky130_fd_sc_hd__a221o_1
X_5877_ _9009_/Q _5875_/X _5898_/S VGND VGND VPWR VPWR _5877_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4828_ _9265_/Q _4458_/Y _5518_/A _8859_/Q _4827_/X VGND VGND VPWR VPWR _4829_/D
+ sky130_fd_sc_hd__a221o_1
X_7616_ _7616_/A VGND VGND VPWR VPWR _9380_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8596_ _8983_/Q _8292_/X _8294_/X _8878_/Q VGND VGND VPWR VPWR _8596_/X sky130_fd_sc_hd__a22o_1
XFILLER_138_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4759_ _4759_/A1 _4502_/Y _7132_/A _9165_/Q VGND VGND VPWR VPWR _4763_/B sky130_fd_sc_hd__a22o_1
X_7547_ _7439_/X hold236/X _7551_/S VGND VGND VPWR VPWR _7547_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7478_ _7478_/A VGND VGND VPWR VPWR _9318_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9217_ _9241_/CLK _9217_/D fanout456/X VGND VGND VPWR VPWR _9217_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_134_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6429_ _6597_/B _6429_/B VGND VGND VPWR VPWR _6492_/B sky130_fd_sc_hd__nand2_1
XFILLER_134_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9148_ _9456_/CLK _9148_/D fanout407/X VGND VGND VPWR VPWR _9148_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_191_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9079_ _9162_/CLK _9079_/D fanout440/X VGND VGND VPWR VPWR _9079_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5800_ _5647_/X hold582/X _5804_/S VGND VGND VPWR VPWR _5801_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6780_ _6895_/B _6781_/C _6967_/B _6779_/X VGND VGND VPWR VPWR _6780_/X sky130_fd_sc_hd__o31a_1
XFILLER_22_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5731_ _5731_/A VGND VGND VPWR VPWR _8949_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5662_ _5662_/A VGND VGND VPWR VPWR _8920_/D sky130_fd_sc_hd__clkbuf_1
X_8450_ _8701_/A _8450_/B _8450_/C VGND VGND VPWR VPWR _8450_/X sky130_fd_sc_hd__or3_1
XFILLER_175_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4613_ _5168_/A1 _4811_/A _4477_/Y input30/X _4612_/X VGND VGND VPWR VPWR _4617_/C
+ sky130_fd_sc_hd__a221o_2
X_7401_ _7401_/A VGND VGND VPWR VPWR _9284_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8381_ _8381_/A VGND VGND VPWR VPWR _8381_/X sky130_fd_sc_hd__buf_8
X_5593_ _5593_/A VGND VGND VPWR VPWR _8891_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7332_ _7332_/A VGND VGND VPWR VPWR _9252_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4544_ _9334_/Q _7499_/A _7661_/A _9406_/Q VGND VGND VPWR VPWR _4544_/X sky130_fd_sc_hd__a22o_1
XFILLER_128_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold402 _9298_/Q VGND VGND VPWR VPWR hold402/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 hold413/A VGND VGND VPWR VPWR hold413/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold424 _7346_/X VGND VGND VPWR VPWR _7347_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7263_ _7263_/A VGND VGND VPWR VPWR _9222_/D sky130_fd_sc_hd__clkbuf_1
Xhold435 hold435/A VGND VGND VPWR VPWR hold435/X sky130_fd_sc_hd__dlygate4sd3_1
X_4475_ _4475_/A VGND VGND VPWR VPWR _4536_/B sky130_fd_sc_hd__inv_4
Xhold446 _6016_/X VGND VGND VPWR VPWR _6017_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 _5459_/X VGND VGND VPWR VPWR _5460_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold468 hold468/A VGND VGND VPWR VPWR hold468/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9002_ _9178_/CLK _9002_/D fanout487/X VGND VGND VPWR VPWR _9002_/Q sky130_fd_sc_hd__dfrtp_1
X_6214_ _6794_/A _6633_/A VGND VGND VPWR VPWR _6215_/A sky130_fd_sc_hd__and2b_1
Xhold479 _8854_/Q VGND VGND VPWR VPWR hold479/X sky130_fd_sc_hd__dlygate4sd3_1
X_7194_ _7194_/A _7284_/B VGND VGND VPWR VPWR _7209_/S sky130_fd_sc_hd__nand2_8
XFILLER_143_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6145_ _6876_/B _6736_/B VGND VGND VPWR VPWR _6290_/B sky130_fd_sc_hd__nor2_1
XFILLER_38_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1102 _9092_/Q VGND VGND VPWR VPWR hold204/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1113 _9093_/Q VGND VGND VPWR VPWR hold337/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1124 _8987_/Q VGND VGND VPWR VPWR hold648/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _6076_/A VGND VGND VPWR VPWR _9103_/D sky130_fd_sc_hd__clkbuf_1
Xhold1135 _9383_/Q VGND VGND VPWR VPWR hold224/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 _9069_/Q VGND VGND VPWR VPWR hold901/A sky130_fd_sc_hd__dlygate4sd3_1
X_5027_ _5027_/A VGND VGND VPWR VPWR _8795_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1157 _8979_/Q VGND VGND VPWR VPWR hold454/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1168 _9038_/Q VGND VGND VPWR VPWR hold851/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1179 _7116_/X VGND VGND VPWR VPWR hold425/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_308 _7695_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_319 _8807_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6978_ _6978_/A _6978_/B _6978_/C _6978_/D VGND VGND VPWR VPWR _6978_/X sky130_fd_sc_hd__and4_1
XFILLER_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8717_ _9537_/Q _4752_/X _8725_/S VGND VGND VPWR VPWR _8718_/A sky130_fd_sc_hd__mux2_1
X_5929_ _9029_/Q _5929_/B VGND VGND VPWR VPWR _5930_/A sky130_fd_sc_hd__and2_1
XFILLER_179_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8648_ _9050_/Q _8356_/A _8360_/B _8890_/Q _8647_/X VGND VGND VPWR VPWR _8649_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_186_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8579_ hold990/X _8196_/S _8577_/X _8578_/X VGND VGND VPWR VPWR _8579_/X sky130_fd_sc_hd__o22a_1
XFILLER_166_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold980 _9112_/Q VGND VGND VPWR VPWR hold980/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold991 _8579_/X VGND VGND VPWR VPWR _9527_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7950_ _9495_/Q _9494_/Q VGND VGND VPWR VPWR _8002_/C sky130_fd_sc_hd__and2_2
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6901_ _6518_/Y _6812_/Y _6900_/Y _6642_/Y VGND VGND VPWR VPWR _6997_/B sky130_fd_sc_hd__a211o_1
X_7881_ _9494_/Q _7881_/B VGND VGND VPWR VPWR _7883_/B sky130_fd_sc_hd__or2_1
XFILLER_63_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6832_ _6334_/B _6871_/B _6524_/C _6830_/A _6463_/A VGND VGND VPWR VPWR _6832_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_35_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9551_ _9551_/CLK _9551_/D _8709_/B VGND VGND VPWR VPWR _9551_/Q sky130_fd_sc_hd__dfrtp_1
X_6763_ _6763_/A _6763_/B VGND VGND VPWR VPWR _6838_/A sky130_fd_sc_hd__or2_1
X_8502_ _5130_/A _9523_/Q _8013_/A _8501_/X VGND VGND VPWR VPWR _8502_/X sky130_fd_sc_hd__a211o_1
X_5714_ _5714_/A VGND VGND VPWR VPWR _8942_/D sky130_fd_sc_hd__clkbuf_1
X_9482_ _9482_/CLK _9482_/D fanout435/X VGND VGND VPWR VPWR _9482_/Q sky130_fd_sc_hd__dfrtp_1
X_6694_ _6227_/Y _6508_/A _6781_/C VGND VGND VPWR VPWR _6694_/Y sky130_fd_sc_hd__a21oi_1
X_8433_ _9330_/Q _8298_/X _8370_/X _9250_/Q VGND VGND VPWR VPWR _8433_/X sky130_fd_sc_hd__a22o_1
X_5645_ _5633_/X hold439/X _5654_/S VGND VGND VPWR VPWR _5646_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8364_ _8364_/A _8364_/B _8388_/A _8384_/A VGND VGND VPWR VPWR _8398_/D sky130_fd_sc_hd__or4_1
X_5576_ _5301_/X hold529/X _5582_/S VGND VGND VPWR VPWR _5577_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold210 _7762_/X VGND VGND VPWR VPWR _7763_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7315_ _7242_/X hold265/X _7319_/S VGND VGND VPWR VPWR _7315_/X sky130_fd_sc_hd__mux2_1
X_4527_ input98/X _4488_/Y _4500_/Y input18/X _4526_/X VGND VGND VPWR VPWR _4530_/C
+ sky130_fd_sc_hd__a221o_1
Xhold221 _7809_/X VGND VGND VPWR VPWR _7810_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold232 _7457_/X VGND VGND VPWR VPWR _7458_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8295_ _9502_/Q _9501_/Q VGND VGND VPWR VPWR _8385_/A sky130_fd_sc_hd__nand2b_4
Xhold243 _7252_/X VGND VGND VPWR VPWR _7253_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold254 _9388_/Q VGND VGND VPWR VPWR hold254/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 _9245_/Q VGND VGND VPWR VPWR hold265/X sky130_fd_sc_hd__dlygate4sd3_1
X_4458_ _4656_/A _4670_/B VGND VGND VPWR VPWR _4458_/Y sky130_fd_sc_hd__nor2_4
X_7246_ _7246_/A VGND VGND VPWR VPWR _9214_/D sky130_fd_sc_hd__clkbuf_1
Xhold276 _7843_/X VGND VGND VPWR VPWR _7844_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold287 _7240_/X VGND VGND VPWR VPWR _7241_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold298 _7350_/X VGND VGND VPWR VPWR _7351_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7177_ _7177_/A VGND VGND VPWR VPWR _7192_/S sky130_fd_sc_hd__buf_4
X_4389_ _4670_/B _4675_/B VGND VGND VPWR VPWR _4389_/Y sky130_fd_sc_hd__nor2_2
XFILLER_131_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6128_ _6399_/A _6724_/A VGND VGND VPWR VPWR _6128_/X sky130_fd_sc_hd__and2_2
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6059_ _6059_/A VGND VGND VPWR VPWR _9095_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 _6012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_116 _6018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 _7299_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 _8275_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_149 _7927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5430_ _8822_/Q _5465_/A _5435_/S VGND VGND VPWR VPWR _5430_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5361_ _5375_/A _5378_/B VGND VGND VPWR VPWR _5362_/A sky130_fd_sc_hd__and2_1
Xoutput304 _4915_/X VGND VGND VPWR VPWR reset sky130_fd_sc_hd__buf_12
XFILLER_161_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput315 _9555_/X VGND VGND VPWR VPWR spimemio_flash_io3_di sky130_fd_sc_hd__buf_12
XFILLER_114_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput326 _9533_/Q VGND VGND VPWR VPWR wb_ack_o sky130_fd_sc_hd__buf_12
Xoutput337 _9043_/Q VGND VGND VPWR VPWR wb_dat_o[19] sky130_fd_sc_hd__buf_12
X_7100_ _6018_/X _9151_/Q _7106_/S VGND VGND VPWR VPWR _7100_/X sky130_fd_sc_hd__mux2_1
X_8080_ _9211_/Q _7923_/X _7997_/X _9363_/Q VGND VGND VPWR VPWR _8080_/X sky130_fd_sc_hd__a22o_1
Xoutput348 _9539_/Q VGND VGND VPWR VPWR wb_dat_o[29] sky130_fd_sc_hd__buf_12
XFILLER_114_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5292_ _5292_/A hold74/X VGND VGND VPWR VPWR _5292_/X sky130_fd_sc_hd__or2b_1
X_7031_ _7031_/A VGND VGND VPWR VPWR _9120_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8982_ _9465_/CLK _8982_/D fanout471/X VGND VGND VPWR VPWR _8982_/Q sky130_fd_sc_hd__dfrtp_4
X_7933_ _7933_/A VGND VGND VPWR VPWR _7933_/X sky130_fd_sc_hd__buf_6
XFILLER_36_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7864_ _7864_/A VGND VGND VPWR VPWR _7865_/C sky130_fd_sc_hd__clkinv_2
XFILLER_51_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6815_ _6906_/C _6815_/B _6862_/A VGND VGND VPWR VPWR _6976_/D sky130_fd_sc_hd__nor3_1
XFILLER_168_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7795_ _7795_/A VGND VGND VPWR VPWR _9462_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9534_ _9541_/CLK _9534_/D VGND VGND VPWR VPWR _9534_/Q sky130_fd_sc_hd__dfxtp_1
X_6746_ _6728_/B _6730_/X _6745_/X VGND VGND VPWR VPWR _6969_/A sky130_fd_sc_hd__o21ai_1
XFILLER_50_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9465_ _9465_/CLK _9465_/D fanout472/X VGND VGND VPWR VPWR _9465_/Q sky130_fd_sc_hd__dfstp_1
X_6677_ _6897_/B _6521_/B _6413_/B _6673_/B _6328_/Y VGND VGND VPWR VPWR _6706_/B
+ sky130_fd_sc_hd__a32o_1
X_8416_ _9233_/Q _8356_/B _8364_/B _9265_/Q _8415_/X VGND VGND VPWR VPWR _8423_/A
+ sky130_fd_sc_hd__a221o_1
X_5628_ _5628_/A VGND VGND VPWR VPWR _8907_/D sky130_fd_sc_hd__clkbuf_1
X_9396_ _9420_/CLK _9396_/D fanout465/X VGND VGND VPWR VPWR _9396_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_164_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8347_ _8355_/A _8359_/B VGND VGND VPWR VPWR _8360_/C sky130_fd_sc_hd__nor2_4
XFILLER_164_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5559_ _5559_/A VGND VGND VPWR VPWR _8876_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8278_ _9039_/Q _7938_/A _7977_/X _8776_/Q VGND VGND VPWR VPWR _8278_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7229_ _7128_/X _9208_/Q _7247_/S VGND VGND VPWR VPWR _7229_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A VGND VGND VPWR VPWR _9520_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4930_ input93/X _4444_/Y _4501_/Y _9288_/Q _4929_/X VGND VGND VPWR VPWR _4931_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_33_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4861_ _4861_/A _7126_/A VGND VGND VPWR VPWR _5437_/A sky130_fd_sc_hd__nor2_1
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6600_ _6610_/A _7001_/A VGND VGND VPWR VPWR _6882_/A sky130_fd_sc_hd__nor2_1
XFILLER_178_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4792_ _9450_/Q _4836_/A2 _5704_/A _8940_/Q VGND VGND VPWR VPWR _4792_/X sky130_fd_sc_hd__a22o_1
XANTENNA_16 _7605_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7580_ _7436_/X hold264/X hold78/X VGND VGND VPWR VPWR _7581_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_27 _4569_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 _4676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_49 _4816_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6531_ _6887_/B _6862_/A VGND VGND VPWR VPWR _6531_/X sky130_fd_sc_hd__or2_1
XFILLER_146_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9250_ _9290_/CLK _9250_/D fanout467/X VGND VGND VPWR VPWR _9250_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6462_ _6973_/B _6462_/B VGND VGND VPWR VPWR _6463_/B sky130_fd_sc_hd__nand2_1
XFILLER_146_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8201_ _8964_/Q _7960_/X _8001_/X _8864_/Q _8200_/X VGND VGND VPWR VPWR _8209_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5413_ hold4/X _5413_/A1 _5413_/S VGND VGND VPWR VPWR _5413_/X sky130_fd_sc_hd__mux2_4
X_6393_ _6393_/A _6781_/C VGND VGND VPWR VPWR _6925_/B sky130_fd_sc_hd__nor2_1
X_9181_ _9181_/CLK _9181_/D fanout487/X VGND VGND VPWR VPWR _9181_/Q sky130_fd_sc_hd__dfrtp_1
X_5344_ _5344_/A VGND VGND VPWR VPWR _5344_/X sky130_fd_sc_hd__clkbuf_1
X_8132_ _9374_/Q _7960_/A _8001_/A _9270_/Q _8131_/X VGND VGND VPWR VPWR _8140_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5275_ _5275_/A _5287_/B VGND VGND VPWR VPWR _5276_/A sky130_fd_sc_hd__and2_1
X_8063_ _8063_/A VGND VGND VPWR VPWR _9509_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7014_ _7014_/A VGND VGND VPWR VPWR _7014_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8965_ _9184_/CLK _8965_/D fanout439/X VGND VGND VPWR VPWR _8965_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_71_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7916_ _9490_/Q _9491_/Q _7916_/C _9488_/Q VGND VGND VPWR VPWR _7916_/X sky130_fd_sc_hd__or4b_1
XFILLER_102_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8896_ _9473_/CLK _8896_/D fanout432/X VGND VGND VPWR VPWR _8896_/Q sky130_fd_sc_hd__dfstp_1
X_7847_ _5415_/X hold738/X _7847_/S VGND VGND VPWR VPWR _7847_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7778_ _7778_/A VGND VGND VPWR VPWR _9454_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9517_ _9531_/CLK _9517_/D fanout452/X VGND VGND VPWR VPWR _9517_/Q sky130_fd_sc_hd__dfrtp_1
X_6729_ _6869_/B _6729_/B _6729_/C VGND VGND VPWR VPWR _6966_/D sky130_fd_sc_hd__nand3b_1
XFILLER_149_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9448_ _9476_/CLK _9448_/D fanout414/X VGND VGND VPWR VPWR _9448_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_164_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_52_csclk _9090_/CLK VGND VGND VPWR VPWR _9091_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_164_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9379_ _9459_/CLK _9379_/D fanout480/X VGND VGND VPWR VPWR _9379_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_105_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_67_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _9484_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_59_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput14 mask_rev_in[19] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__clkbuf_1
Xinput25 mask_rev_in[29] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__clkbuf_2
Xinput36 mgmt_gpio_in[0] VGND VGND VPWR VPWR _5281_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_168_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput47 mgmt_gpio_in[1] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__buf_2
Xinput58 mgmt_gpio_in[2] VGND VGND VPWR VPWR _5012_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_183_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput69 mgmt_gpio_in[6] VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__buf_2
XFILLER_182_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold809 _8975_/Q VGND VGND VPWR VPWR hold809/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5060_ _5060_/A VGND VGND VPWR VPWR _8784_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8750_ _8750_/A VGND VGND VPWR VPWR _9545_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5962_ _9053_/Q _4961_/X _5976_/S VGND VGND VPWR VPWR _5963_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7701_ _7701_/A VGND VGND VPWR VPWR _9418_/D sky130_fd_sc_hd__clkbuf_1
X_4913_ input71/X _4436_/A _5795_/A _8978_/Q _4912_/X VGND VGND VPWR VPWR _4921_/B
+ sky130_fd_sc_hd__a221o_1
X_8681_ _8962_/Q _8402_/A _8378_/A _8947_/Q _8680_/X VGND VGND VPWR VPWR _8688_/A
+ sky130_fd_sc_hd__a221o_1
X_5893_ _5893_/A VGND VGND VPWR VPWR _9014_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7632_ _7436_/X hold254/X _7638_/S VGND VGND VPWR VPWR _7632_/X sky130_fd_sc_hd__mux2_1
X_4844_ _9353_/Q _4427_/Y _4406_/Y input35/X _4843_/X VGND VGND VPWR VPWR _4844_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_32_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7563_ _7436_/X hold258/X hold99/A VGND VGND VPWR VPWR _7563_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4775_ _9210_/Q _7228_/A _5738_/A _8955_/Q VGND VGND VPWR VPWR _4775_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9302_ _9325_/CLK _9302_/D fanout464/X VGND VGND VPWR VPWR _9302_/Q sky130_fd_sc_hd__dfrtp_4
X_6514_ _6514_/A VGND VGND VPWR VPWR _6514_/Y sky130_fd_sc_hd__inv_2
X_7494_ _7494_/A VGND VGND VPWR VPWR _7494_/X sky130_fd_sc_hd__buf_2
XFILLER_107_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9233_ _9483_/CLK _9233_/D fanout473/X VGND VGND VPWR VPWR _9233_/Q sky130_fd_sc_hd__dfstp_2
X_6445_ _6518_/A _6926_/B VGND VGND VPWR VPWR _6445_/Y sky130_fd_sc_hd__nor2_2
XFILLER_106_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9164_ _9383_/CLK _9164_/D fanout408/X VGND VGND VPWR VPWR _9164_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_164_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6376_ _6376_/A VGND VGND VPWR VPWR _6376_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8115_ _9245_/Q _7949_/X _7999_/X _9429_/Q VGND VGND VPWR VPWR _8115_/X sky130_fd_sc_hd__a22o_1
X_5327_ _5327_/A VGND VGND VPWR VPWR _5327_/X sky130_fd_sc_hd__clkbuf_1
X_9095_ _9473_/CLK _9095_/D fanout430/X VGND VGND VPWR VPWR _9095_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8046_ _9322_/Q _7962_/A _7988_/A _9434_/Q VGND VGND VPWR VPWR _8046_/X sky130_fd_sc_hd__a22o_1
XFILLER_102_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5258_ _9363_/Q VGND VGND VPWR VPWR _5258_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5189_ _5189_/A VGND VGND VPWR VPWR _5189_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8948_ _9467_/CLK _8948_/D fanout476/X VGND VGND VPWR VPWR _8948_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_189_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8879_ _9084_/CLK _8879_/D fanout447/X VGND VGND VPWR VPWR _8879_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4560_ _9429_/Q _4437_/Y _7815_/A _9477_/Q _4559_/X VGND VGND VPWR VPWR _4569_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_8_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold606 _8985_/Q VGND VGND VPWR VPWR hold606/X sky130_fd_sc_hd__dlygate4sd3_1
X_4491_ _7111_/A hold33/X VGND VGND VPWR VPWR _4491_/Y sky130_fd_sc_hd__nor2_2
XFILLER_155_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold617 _8920_/Q VGND VGND VPWR VPWR hold617/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 _7122_/X VGND VGND VPWR VPWR _7123_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold639 _9181_/Q VGND VGND VPWR VPWR hold639/X sky130_fd_sc_hd__dlygate4sd3_1
X_6230_ _6628_/A _6589_/C _6230_/C VGND VGND VPWR VPWR _6230_/X sky130_fd_sc_hd__and3_2
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6161_ _6437_/A _6716_/A _6428_/B VGND VGND VPWR VPWR _6535_/A sky130_fd_sc_hd__or3_4
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _9203_/Q VGND VGND VPWR VPWR _5112_/Y sky130_fd_sc_hd__inv_2
X_6092_ _6093_/B _6092_/B VGND VGND VPWR VPWR _6716_/B sky130_fd_sc_hd__or2_2
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _5127_/A _4977_/B _5065_/S _5042_/Y VGND VGND VPWR VPWR _5050_/B sky130_fd_sc_hd__o31a_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_wbbd_sck _9550_/Q VGND VGND VPWR VPWR clkbuf_0_wbbd_sck/X sky130_fd_sc_hd__clkbuf_16
X_8802_ _5168_/A1 _8802_/D _5372_/X VGND VGND VPWR VPWR hold80/A sky130_fd_sc_hd__dfrtp_1
XFILLER_65_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6994_ _6994_/A _6994_/B _6994_/C VGND VGND VPWR VPWR _6994_/Y sky130_fd_sc_hd__nor3_1
X_8733_ _9034_/Q _8731_/Y _8732_/Y _9032_/Q VGND VGND VPWR VPWR _8735_/C sky130_fd_sc_hd__a22o_1
XFILLER_80_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5945_ _9047_/Q _4507_/X _5945_/S VGND VGND VPWR VPWR _5946_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8664_ _8931_/Q _8398_/B _8344_/X _8896_/Q VGND VGND VPWR VPWR _8664_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5876_ _7158_/B _5453_/C _5819_/X _5897_/S hold21/A VGND VGND VPWR VPWR _5898_/S
+ sky130_fd_sc_hd__o221a_4
XFILLER_178_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7615_ hold310/X _5690_/A _7621_/S VGND VGND VPWR VPWR _7615_/X sky130_fd_sc_hd__mux2_1
X_4827_ _8974_/Q _5784_/A _6043_/A _9090_/Q VGND VGND VPWR VPWR _4827_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8595_ _9079_/Q _8324_/X _8341_/X _8888_/Q VGND VGND VPWR VPWR _8600_/B sky130_fd_sc_hd__a22o_1
X_7546_ _7546_/A VGND VGND VPWR VPWR _9348_/D sky130_fd_sc_hd__clkbuf_1
X_4758_ _4758_/A _5453_/B VGND VGND VPWR VPWR _7132_/A sky130_fd_sc_hd__nor2_4
XFILLER_193_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7477_ hold398/X _7494_/A _7479_/S VGND VGND VPWR VPWR _7478_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4689_ _4689_/A _4689_/B _4689_/C _4689_/D VGND VGND VPWR VPWR _4690_/D sky130_fd_sc_hd__or4_1
XFILLER_146_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9216_ _9383_/CLK _9216_/D fanout409/X VGND VGND VPWR VPWR _9216_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_107_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6428_ _6850_/B _6428_/B VGND VGND VPWR VPWR _6429_/B sky130_fd_sc_hd__nor2_1
XFILLER_134_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9147_ _9456_/CLK _9147_/D fanout407/X VGND VGND VPWR VPWR _9147_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_68_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6359_ _6869_/C _6869_/D _6359_/C VGND VGND VPWR VPWR _6359_/X sky130_fd_sc_hd__or3_1
XFILLER_88_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9078_ _9484_/CLK _9078_/D fanout430/X VGND VGND VPWR VPWR _9078_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_102_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8029_ _9249_/Q _7940_/X _8001_/X _9265_/Q _8028_/X VGND VGND VPWR VPWR _8037_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_84_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5730_ _5633_/X hold455/X _5736_/S VGND VGND VPWR VPWR _5731_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5661_ hold617/X _5395_/X _5665_/S VGND VGND VPWR VPWR _5662_/A sky130_fd_sc_hd__mux2_1
XFILLER_176_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7400_ _7239_/X hold285/X _7406_/S VGND VGND VPWR VPWR _7400_/X sky130_fd_sc_hd__mux2_1
X_4612_ _9228_/Q _4454_/Y _5678_/A _8932_/Q VGND VGND VPWR VPWR _4612_/X sky130_fd_sc_hd__a22o_1
X_8380_ _8380_/A _8385_/A VGND VGND VPWR VPWR _8381_/A sky130_fd_sc_hd__nor2_8
XFILLER_191_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5592_ hold667/X _5398_/X _5594_/S VGND VGND VPWR VPWR _5593_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7331_ hold309/X _5690_/A _7337_/S VGND VGND VPWR VPWR _7331_/X sky130_fd_sc_hd__mux2_1
X_4543_ input69/X _4811_/A _7571_/A _9366_/Q _4542_/X VGND VGND VPWR VPWR _4548_/B
+ sky130_fd_sc_hd__a221o_1
Xhold403 _7431_/X VGND VGND VPWR VPWR _7432_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold414 _9402_/Q VGND VGND VPWR VPWR hold414/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 hold425/A VGND VGND VPWR VPWR _7117_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 hold436/A VGND VGND VPWR VPWR hold436/X sky130_fd_sc_hd__dlygate4sd3_1
X_7262_ _5468_/X hold794/X _7264_/S VGND VGND VPWR VPWR _7262_/X sky130_fd_sc_hd__mux2_1
X_4474_ _4675_/B _5474_/B VGND VGND VPWR VPWR _7729_/A sky130_fd_sc_hd__nor2_8
Xhold447 _5422_/X VGND VGND VPWR VPWR _5423_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 _8969_/Q VGND VGND VPWR VPWR hold458/X sky130_fd_sc_hd__dlygate4sd3_1
X_9001_ _9006_/CLK _9001_/D fanout493/X VGND VGND VPWR VPWR _9001_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_116_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6213_ _6213_/A VGND VGND VPWR VPWR _6871_/B sky130_fd_sc_hd__clkbuf_4
Xhold469 _8847_/Q VGND VGND VPWR VPWR hold469/X sky130_fd_sc_hd__dlygate4sd3_1
X_7193_ _7193_/A VGND VGND VPWR VPWR _9191_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6144_ _6144_/A VGND VGND VPWR VPWR _6736_/B sky130_fd_sc_hd__buf_4
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1103 _9274_/Q VGND VGND VPWR VPWR hold782/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1114 _6053_/X VGND VGND VPWR VPWR _6054_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ hold159/X _5690_/A _6075_/S VGND VGND VPWR VPWR _6075_/X sky130_fd_sc_hd__mux2_1
Xhold1125 _8986_/Q VGND VGND VPWR VPWR hold436/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1136 _8928_/Q VGND VGND VPWR VPWR hold918/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1147 _9095_/Q VGND VGND VPWR VPWR hold630/A sky130_fd_sc_hd__dlygate4sd3_1
X_5026_ _8795_/Q hold999/X _5026_/S VGND VGND VPWR VPWR _5027_/A sky130_fd_sc_hd__mux2_1
Xhold1158 _9266_/Q VGND VGND VPWR VPWR hold778/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 _8901_/Q VGND VGND VPWR VPWR hold399/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_309 fanout498/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6977_ _6987_/C _6977_/B _6977_/C VGND VGND VPWR VPWR _6978_/D sky130_fd_sc_hd__nor3_1
XFILLER_80_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8716_ _8716_/A VGND VGND VPWR VPWR _9536_/D sky130_fd_sc_hd__clkbuf_1
X_5928_ _5928_/A VGND VGND VPWR VPWR _9039_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8647_ _8774_/Q _8304_/A _8354_/C _9081_/Q VGND VGND VPWR VPWR _8647_/X sky130_fd_sc_hd__a22o_1
X_5859_ _9566_/A _5858_/X _5868_/S VGND VGND VPWR VPWR _5859_/X sky130_fd_sc_hd__mux2_1
X_8578_ _5139_/A _9526_/Q _8013_/X VGND VGND VPWR VPWR _8578_/X sky130_fd_sc_hd__a21o_1
XFILLER_119_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7529_ _7529_/A VGND VGND VPWR VPWR _9340_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold970 _9531_/Q VGND VGND VPWR VPWR hold970/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 _9027_/Q VGND VGND VPWR VPWR _5870_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold992 _9031_/Q VGND VGND VPWR VPWR _5149_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6900_ _6900_/A _6900_/B VGND VGND VPWR VPWR _6900_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7880_ _7881_/B _7887_/B VGND VGND VPWR VPWR _7880_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6831_ _6897_/B _6830_/Y _6467_/D _6758_/B _6758_/A VGND VGND VPWR VPWR _6831_/Y
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9550_ _9550_/CLK _9550_/D _8709_/B VGND VGND VPWR VPWR _9550_/Q sky130_fd_sc_hd__dfrtp_2
X_6762_ _6230_/X _6973_/B _6481_/A _6811_/B VGND VGND VPWR VPWR _6763_/B sky130_fd_sc_hd__o211a_1
X_8501_ _9188_/Q _8400_/B _8487_/X _8500_/X _8627_/S VGND VGND VPWR VPWR _8501_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_188_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5713_ hold616/X _5690_/X _5713_/S VGND VGND VPWR VPWR _5714_/A sky130_fd_sc_hd__mux2_1
X_9481_ _9482_/CLK _9481_/D fanout435/X VGND VGND VPWR VPWR _9481_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_50_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6693_ _6695_/B _6775_/C VGND VGND VPWR VPWR _6693_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8432_ _9370_/Q _8346_/X _8386_/X _9346_/Q _8431_/X VGND VGND VPWR VPWR _8437_/B
+ sky130_fd_sc_hd__a221o_1
X_5644_ _5644_/A VGND VGND VPWR VPWR _8913_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8363_ _8363_/A _8368_/B VGND VGND VPWR VPWR _8384_/A sky130_fd_sc_hd__nor2_2
X_5575_ _5575_/A VGND VGND VPWR VPWR _8883_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold200 hold200/A VGND VGND VPWR VPWR _5887_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 hold211/A VGND VGND VPWR VPWR _5857_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7314_ _7314_/A VGND VGND VPWR VPWR _9244_/D sky130_fd_sc_hd__clkbuf_1
X_4526_ _9286_/Q _4407_/Y _7678_/A _9414_/Q VGND VGND VPWR VPWR _4526_/X sky130_fd_sc_hd__a22o_1
XFILLER_117_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold222 _9229_/Q VGND VGND VPWR VPWR hold222/X sky130_fd_sc_hd__dlygate4sd3_1
X_8294_ _8358_/A VGND VGND VPWR VPWR _8294_/X sky130_fd_sc_hd__buf_6
Xhold233 _9357_/Q VGND VGND VPWR VPWR hold233/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 _9453_/Q VGND VGND VPWR VPWR hold244/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 _7632_/X VGND VGND VPWR VPWR _7633_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7245_ _5468_/X hold785/X _7247_/S VGND VGND VPWR VPWR _7245_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4457_ hold60/X _7111_/A VGND VGND VPWR VPWR _4457_/Y sky130_fd_sc_hd__nor2_2
Xhold266 _7315_/X VGND VGND VPWR VPWR _7316_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold277 _9268_/Q VGND VGND VPWR VPWR hold277/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold288 hold288/A VGND VGND VPWR VPWR hold288/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 _9454_/Q VGND VGND VPWR VPWR hold299/X sky130_fd_sc_hd__dlygate4sd3_1
X_7176_ _7176_/A hold19/X VGND VGND VPWR VPWR _7177_/A sky130_fd_sc_hd__and2_1
XFILLER_131_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4388_ hold83/X VGND VGND VPWR VPWR _4675_/B sky130_fd_sc_hd__buf_6
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6127_ _6721_/A VGND VGND VPWR VPWR _6399_/A sky130_fd_sc_hd__clkinv_2
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6058_ _5951_/X hold630/X _6064_/S VGND VGND VPWR VPWR _6059_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5009_ _5009_/A VGND VGND VPWR VPWR _5010_/A sky130_fd_sc_hd__inv_2
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 _6012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_117 _6048_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_128 _7299_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_139 _7908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5360_ _5360_/A VGND VGND VPWR VPWR _5360_/X sky130_fd_sc_hd__clkbuf_1
Xoutput305 _5278_/X VGND VGND VPWR VPWR ser_rx sky130_fd_sc_hd__buf_12
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput316 _9147_/Q VGND VGND VPWR VPWR sram_ro_addr[0] sky130_fd_sc_hd__buf_12
Xoutput327 _9061_/Q VGND VGND VPWR VPWR wb_dat_o[0] sky130_fd_sc_hd__buf_12
XFILLER_114_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput338 _9062_/Q VGND VGND VPWR VPWR wb_dat_o[1] sky130_fd_sc_hd__buf_12
Xoutput349 _9063_/Q VGND VGND VPWR VPWR wb_dat_o[2] sky130_fd_sc_hd__buf_12
XFILLER_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5291_ _7517_/A VGND VGND VPWR VPWR _5291_/X sky130_fd_sc_hd__buf_6
XFILLER_114_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7030_ _5951_/X _9120_/Q _7030_/S VGND VGND VPWR VPWR _7030_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8981_ _9283_/CLK _8981_/D fanout484/X VGND VGND VPWR VPWR _8981_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_95_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7932_ _7998_/A _7989_/B _7984_/C VGND VGND VPWR VPWR _7933_/A sky130_fd_sc_hd__and3_1
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7863_ _9488_/Q _9489_/Q _9490_/Q _7863_/D VGND VGND VPWR VPWR _7864_/A sky130_fd_sc_hd__and4_1
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6814_ _6535_/A _6862_/B _6655_/C _6510_/Y _6660_/Y VGND VGND VPWR VPWR _6918_/B
+ sky130_fd_sc_hd__o221a_1
X_7794_ _5410_/X hold324/X _7796_/S VGND VGND VPWR VPWR _7794_/X sky130_fd_sc_hd__mux2_1
X_9533_ _9551_/CLK _9533_/D _8709_/B VGND VGND VPWR VPWR _9533_/Q sky130_fd_sc_hd__dfrtp_4
X_6745_ _6609_/Y _6744_/X _6967_/A VGND VGND VPWR VPWR _6745_/X sky130_fd_sc_hd__a21o_1
XFILLER_50_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9464_ _9464_/CLK _9464_/D fanout421/X VGND VGND VPWR VPWR _9464_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_31_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6676_ _6315_/Y _6673_/B _6897_/B _6462_/B VGND VGND VPWR VPWR _6706_/A sky130_fd_sc_hd__a22o_1
XFILLER_149_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8415_ _9281_/Q _8358_/B _8364_/A _9257_/Q VGND VGND VPWR VPWR _8415_/X sky130_fd_sc_hd__a22o_1
X_5627_ hold622/X _5402_/X _5627_/S VGND VGND VPWR VPWR _5628_/A sky130_fd_sc_hd__mux2_1
X_9395_ _9475_/CLK _9395_/D fanout480/X VGND VGND VPWR VPWR _9395_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_191_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8346_ _8682_/B VGND VGND VPWR VPWR _8346_/X sky130_fd_sc_hd__buf_8
XFILLER_164_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5558_ _5311_/X hold453/X _5560_/S VGND VGND VPWR VPWR _5559_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4509_ hold963/X _4507_/X _4886_/S VGND VGND VPWR VPWR _4509_/X sky130_fd_sc_hd__mux2_1
X_8277_ _8977_/Q _7947_/X _7973_/X _8857_/Q _8276_/X VGND VGND VPWR VPWR _8282_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5489_ _5489_/A VGND VGND VPWR VPWR _8846_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7228_ _7228_/A _7284_/B VGND VGND VPWR VPWR _7247_/S sky130_fd_sc_hd__nand2_8
XFILLER_116_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7159_ _7159_/A VGND VGND VPWR VPWR _7174_/S sky130_fd_sc_hd__buf_6
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4860_ _9425_/Q _4437_/Y _7086_/A _9145_/Q _4859_/X VGND VGND VPWR VPWR _4864_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4791_ _4791_/A _4791_/B _4791_/C _4791_/D VGND VGND VPWR VPWR _4797_/A sky130_fd_sc_hd__or4_1
XANTENNA_17 _7746_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 _4570_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 _5540_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6530_ _6917_/B _6642_/B _6729_/B _6530_/D VGND VGND VPWR VPWR _6539_/A sky130_fd_sc_hd__and4_1
XFILLER_118_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6461_ _6461_/A _6898_/A VGND VGND VPWR VPWR _6463_/A sky130_fd_sc_hd__or2_1
XFILLER_185_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8200_ _8974_/Q _7947_/X _7981_/X _8914_/Q VGND VGND VPWR VPWR _8200_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5412_ _5412_/A VGND VGND VPWR VPWR _8815_/D sky130_fd_sc_hd__clkbuf_1
X_9180_ _9181_/CLK _9180_/D fanout486/X VGND VGND VPWR VPWR _9180_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6392_ _6392_/A _6392_/B VGND VGND VPWR VPWR _6781_/C sky130_fd_sc_hd__or2_2
XFILLER_133_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8131_ _9382_/Q _7947_/A _7981_/A _9334_/Q VGND VGND VPWR VPWR _8131_/X sky130_fd_sc_hd__a22o_1
X_5343_ _5353_/A _5356_/B VGND VGND VPWR VPWR _5344_/A sky130_fd_sc_hd__and2_1
XFILLER_114_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8062_ _8062_/A0 _8061_/X _8196_/S VGND VGND VPWR VPWR _8063_/A sky130_fd_sc_hd__mux2_1
X_5274_ _5274_/A VGND VGND VPWR VPWR _9028_/D sky130_fd_sc_hd__clkbuf_1
X_7013_ _7025_/A _7013_/B VGND VGND VPWR VPWR _7014_/A sky130_fd_sc_hd__and2_1
XFILLER_28_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8964_ _9184_/CLK _8964_/D fanout443/X VGND VGND VPWR VPWR _8964_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_71_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7915_ _7915_/A VGND VGND VPWR VPWR _9504_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8895_ _9473_/CLK _8895_/D fanout432/X VGND VGND VPWR VPWR _8895_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_102_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7846_ _7846_/A VGND VGND VPWR VPWR _9486_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7777_ _5410_/X hold299/X _7779_/S VGND VGND VPWR VPWR _7777_/X sky130_fd_sc_hd__mux2_1
X_4989_ _4989_/A VGND VGND VPWR VPWR _8804_/D sky130_fd_sc_hd__clkbuf_1
X_9516_ _9531_/CLK _9516_/D fanout452/X VGND VGND VPWR VPWR _9516_/Q sky130_fd_sc_hd__dfrtp_1
X_6728_ _6732_/A _6728_/B _6742_/B VGND VGND VPWR VPWR _6729_/C sky130_fd_sc_hd__or3_1
XFILLER_137_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9447_ _9486_/CLK _9447_/D fanout413/X VGND VGND VPWR VPWR _9447_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6659_ _6738_/A _6659_/B _6659_/C _6809_/C VGND VGND VPWR VPWR _6661_/C sky130_fd_sc_hd__or4b_1
XFILLER_164_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9378_ _9466_/CLK _9378_/D fanout471/X VGND VGND VPWR VPWR _9378_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8329_ _9232_/Q _8322_/X _8324_/X _9240_/Q _8328_/X VGND VGND VPWR VPWR _8351_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput15 mask_rev_in[1] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__clkbuf_2
Xinput26 mask_rev_in[2] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput37 mgmt_gpio_in[10] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput48 mgmt_gpio_in[20] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__clkbuf_2
Xinput59 mgmt_gpio_in[30] VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__buf_4
XFILLER_10_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5961_ _5961_/A VGND VGND VPWR VPWR _5976_/S sky130_fd_sc_hd__clkbuf_4
X_7700_ _7645_/X hold724/X _7710_/S VGND VGND VPWR VPWR _7701_/A sky130_fd_sc_hd__mux2_1
X_4912_ _9464_/Q _7798_/A _7678_/A _9408_/Q VGND VGND VPWR VPWR _4912_/X sky130_fd_sc_hd__a22o_1
X_8680_ _8902_/Q _8354_/A _8376_/A _8952_/Q VGND VGND VPWR VPWR _8680_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5892_ _9559_/A _5891_/X _5898_/S VGND VGND VPWR VPWR _5892_/X sky130_fd_sc_hd__mux2_1
X_7631_ _7631_/A VGND VGND VPWR VPWR _9387_/D sky130_fd_sc_hd__clkbuf_1
X_4843_ _9441_/Q _7746_/A _5762_/A _8964_/Q VGND VGND VPWR VPWR _4843_/X sky130_fd_sc_hd__a22o_1
XFILLER_33_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7562_ _7562_/A VGND VGND VPWR VPWR _9355_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4774_ _9346_/Q _7536_/A _7321_/A _9250_/Q _4773_/X VGND VGND VPWR VPWR _4781_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_165_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9301_ _9325_/CLK _9301_/D fanout460/X VGND VGND VPWR VPWR _9301_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_193_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6513_ _6748_/B _6900_/A VGND VGND VPWR VPWR _6517_/C sky130_fd_sc_hd__nor2_1
XFILLER_158_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7493_ _7493_/A VGND VGND VPWR VPWR _9325_/D sky130_fd_sc_hd__clkbuf_1
X_9232_ _9437_/CLK _9232_/D fanout419/X VGND VGND VPWR VPWR _9232_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_146_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6444_ _6444_/A VGND VGND VPWR VPWR _6926_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_134_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9163_ _9452_/CLK _9163_/D fanout415/X VGND VGND VPWR VPWR _9163_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_115_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6375_ _6811_/B _6811_/C _6422_/B VGND VGND VPWR VPWR _6754_/C sky130_fd_sc_hd__and3_1
X_8114_ _9253_/Q _7940_/X _8113_/X VGND VGND VPWR VPWR _8117_/C sky130_fd_sc_hd__a21o_1
XFILLER_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5326_ _5330_/A _5334_/B VGND VGND VPWR VPWR _5327_/A sky130_fd_sc_hd__and2_1
X_9094_ _9484_/CLK _9094_/D fanout428/X VGND VGND VPWR VPWR _9094_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_130_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8045_ _9250_/Q _7940_/A _7969_/A _9290_/Q _8044_/X VGND VGND VPWR VPWR _8050_/B
+ sky130_fd_sc_hd__a221o_1
X_5257_ _9355_/Q VGND VGND VPWR VPWR _5257_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5188_ _9174_/Q input89/X _5194_/S VGND VGND VPWR VPWR _5189_/A sky130_fd_sc_hd__mux2_2
XFILLER_28_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8947_ _9088_/CLK _8947_/D fanout454/X VGND VGND VPWR VPWR _8947_/Q sky130_fd_sc_hd__dfrtp_4
X_8878_ _9089_/CLK _8878_/D fanout433/X VGND VGND VPWR VPWR _8878_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_24_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7829_ _7829_/A VGND VGND VPWR VPWR _9478_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4490_ _7158_/A _5453_/B VGND VGND VPWR VPWR _4582_/A sky130_fd_sc_hd__nor2_8
Xhold607 _8857_/Q VGND VGND VPWR VPWR hold607/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold618 _5424_/X VGND VGND VPWR VPWR _5425_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold629 _7123_/X VGND VGND VPWR VPWR _9161_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap359 _7764_/A VGND VGND VPWR VPWR _4836_/A2 sky130_fd_sc_hd__buf_6
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6160_ _6973_/A _6399_/A VGND VGND VPWR VPWR _6428_/B sky130_fd_sc_hd__or2_4
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5111_ _9211_/Q VGND VGND VPWR VPWR _5111_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _6175_/A _6095_/B _6437_/A VGND VGND VPWR VPWR _6092_/B sky130_fd_sc_hd__a21oi_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5042_ _5051_/C VGND VGND VPWR VPWR _5042_/Y sky130_fd_sc_hd__inv_2
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8801_ _5168_/A1 _8801_/D _5370_/X VGND VGND VPWR VPWR _8801_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6993_ _6993_/A _6993_/B _6993_/C _6993_/D VGND VGND VPWR VPWR _6993_/X sky130_fd_sc_hd__or4_1
XFILLER_92_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8732_ _8732_/A _8732_/B VGND VGND VPWR VPWR _8732_/Y sky130_fd_sc_hd__nand2_1
X_5944_ _5944_/A VGND VGND VPWR VPWR _9046_/D sky130_fd_sc_hd__clkbuf_1
X_8663_ _8663_/A _8663_/B _8663_/C _8663_/D VGND VGND VPWR VPWR _8663_/X sky130_fd_sc_hd__or4_1
XFILLER_33_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5875_ hold814/X _7517_/A _5897_/S VGND VGND VPWR VPWR _5875_/X sky130_fd_sc_hd__mux2_1
X_4826_ _9122_/Q _7032_/A _5948_/A _9049_/Q _4825_/X VGND VGND VPWR VPWR _4829_/C
+ sky130_fd_sc_hd__a221o_1
X_7614_ _7614_/A VGND VGND VPWR VPWR _9379_/D sky130_fd_sc_hd__clkbuf_1
X_8594_ _9048_/Q _8289_/X _8304_/X _8772_/Q VGND VGND VPWR VPWR _8600_/A sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_66_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _9473_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_166_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7545_ _7436_/X hold267/X _7551_/S VGND VGND VPWR VPWR _7546_/A sky130_fd_sc_hd__mux2_1
X_4757_ _9274_/Q _4938_/A2 _7605_/A _9378_/Q _4756_/X VGND VGND VPWR VPWR _4763_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_147_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7476_ _7476_/A VGND VGND VPWR VPWR _9317_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4688_ _4688_/A _4688_/B _4688_/C _4688_/D VGND VGND VPWR VPWR _4689_/D sky130_fd_sc_hd__or4_1
X_9215_ _9383_/CLK _9215_/D fanout409/X VGND VGND VPWR VPWR _9215_/Q sky130_fd_sc_hd__dfrtp_2
X_6427_ _6440_/A _6891_/B VGND VGND VPWR VPWR _6524_/C sky130_fd_sc_hd__or2_4
XFILLER_162_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9146_ _9462_/CLK _9146_/D fanout408/X VGND VGND VPWR VPWR _9146_/Q sky130_fd_sc_hd__dfstp_2
X_6358_ _6328_/Y _6839_/A _6935_/A _6357_/X VGND VGND VPWR VPWR _6359_/C sky130_fd_sc_hd__a211o_1
XFILLER_103_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5309_ hold44/X hold197/X hold74/A VGND VGND VPWR VPWR _5309_/X sky130_fd_sc_hd__mux2_1
X_9077_ _9162_/CLK _9077_/D fanout437/X VGND VGND VPWR VPWR _9077_/Q sky130_fd_sc_hd__dfrtp_4
X_6289_ _6589_/D _6597_/A _6710_/A VGND VGND VPWR VPWR _6289_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_88_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8028_ hold88/A _8224_/B _7967_/X hold96/A VGND VGND VPWR VPWR _8028_/X sky130_fd_sc_hd__a22o_1
XFILLER_29_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_19_csclk _9303_/CLK VGND VGND VPWR VPWR _9325_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_140_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold4 hold4/A VGND VGND VPWR VPWR hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5660_ _5660_/A VGND VGND VPWR VPWR _8919_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4611_ _4635_/A _7158_/B VGND VGND VPWR VPWR _5678_/A sky130_fd_sc_hd__nor2_2
X_5591_ _5591_/A VGND VGND VPWR VPWR _8890_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7330_ hold67/X VGND VGND VPWR VPWR _9251_/D sky130_fd_sc_hd__clkbuf_1
X_4542_ input27/X _4460_/Y _4477_/Y input32/X VGND VGND VPWR VPWR _4542_/X sky130_fd_sc_hd__a22o_1
XFILLER_129_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold404 _8971_/Q VGND VGND VPWR VPWR hold404/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire390 _4439_/Y VGND VGND VPWR VPWR _7695_/A sky130_fd_sc_hd__buf_8
X_7261_ _7261_/A VGND VGND VPWR VPWR _9221_/D sky130_fd_sc_hd__clkbuf_1
Xhold415 _7666_/X VGND VGND VPWR VPWR _7667_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4473_ _9487_/Q _7832_/A _5418_/A _8824_/Q _4472_/X VGND VGND VPWR VPWR _4495_/A
+ sky130_fd_sc_hd__a221o_1
Xhold426 _9410_/Q VGND VGND VPWR VPWR hold426/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 _8856_/Q VGND VGND VPWR VPWR hold437/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 hold448/A VGND VGND VPWR VPWR hold448/X sky130_fd_sc_hd__dlygate4sd3_1
X_9000_ _9178_/CLK _9000_/D fanout486/X VGND VGND VPWR VPWR _9000_/Q sky130_fd_sc_hd__dfrtp_2
Xhold459 hold459/A VGND VGND VPWR VPWR hold459/X sky130_fd_sc_hd__dlygate4sd3_1
X_6212_ _6216_/A _6262_/A VGND VGND VPWR VPWR _6213_/A sky130_fd_sc_hd__or2_1
XFILLER_143_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7192_ hold205/X _7514_/A _7192_/S VGND VGND VPWR VPWR _7192_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6143_ _6628_/B _6420_/B VGND VGND VPWR VPWR _6144_/A sky130_fd_sc_hd__or2_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ hold72/X VGND VGND VPWR VPWR _9102_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1104 _9258_/Q VGND VGND VPWR VPWR hold781/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1115 _5859_/X VGND VGND VPWR VPWR hold1115/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1126 _8956_/Q VGND VGND VPWR VPWR hold710/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 _9319_/Q VGND VGND VPWR VPWR hold235/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5025_ _5068_/B _5025_/B VGND VGND VPWR VPWR _5026_/S sky130_fd_sc_hd__nor2_1
XFILLER_85_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1148 _9399_/Q VGND VGND VPWR VPWR hold657/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 _8957_/Q VGND VGND VPWR VPWR hold336/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6976_ _8735_/A _6976_/B _6976_/C _6976_/D VGND VGND VPWR VPWR _6977_/C sky130_fd_sc_hd__or4_1
X_8715_ _9536_/Q _4817_/X _8725_/S VGND VGND VPWR VPWR _8716_/A sky130_fd_sc_hd__mux2_1
X_5927_ _5653_/X hold360/X _5927_/S VGND VGND VPWR VPWR _5927_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8646_ _8975_/Q _8337_/A _8384_/A _8855_/Q _8645_/X VGND VGND VPWR VPWR _8649_/C
+ sky130_fd_sc_hd__a221o_1
X_5858_ hold137/X hold24/X _5867_/S VGND VGND VPWR VPWR _5858_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4809_ _9394_/Q _4389_/Y _5996_/A _9071_/Q VGND VGND VPWR VPWR _4809_/X sky130_fd_sc_hd__a22o_1
XFILLER_186_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8577_ _9191_/Q _8400_/B _8576_/X _8105_/X VGND VGND VPWR VPWR _8577_/X sky130_fd_sc_hd__o211a_2
X_5789_ hold809/X _5683_/X _5793_/S VGND VGND VPWR VPWR _5790_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7528_ _7436_/X hold240/X _7534_/S VGND VGND VPWR VPWR _7529_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7459_ _7279_/X hold759/X _7461_/S VGND VGND VPWR VPWR _7459_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold960 _8604_/X VGND VGND VPWR VPWR _9528_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 _8679_/X VGND VGND VPWR VPWR _9531_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold982 _9514_/Q VGND VGND VPWR VPWR hold982/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold993 _9499_/Q VGND VGND VPWR VPWR hold993/X sky130_fd_sc_hd__dlygate4sd3_1
X_9129_ _9487_/CLK _9129_/D fanout411/X VGND VGND VPWR VPWR _9129_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6830_ _6830_/A VGND VGND VPWR VPWR _6830_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6761_ _6761_/A _6761_/B _6761_/C VGND VGND VPWR VPWR _6785_/A sky130_fd_sc_hd__or3_1
X_5712_ _5712_/A VGND VGND VPWR VPWR _8941_/D sky130_fd_sc_hd__clkbuf_1
X_8500_ _8701_/A _8500_/B _8500_/C VGND VGND VPWR VPWR _8500_/X sky130_fd_sc_hd__or3_1
XFILLER_149_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6692_ _6721_/A _6692_/B VGND VGND VPWR VPWR _6775_/C sky130_fd_sc_hd__nand2_1
X_9480_ _9480_/CLK _9480_/D fanout415/X VGND VGND VPWR VPWR _9480_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8431_ _9410_/Q _8506_/B VGND VGND VPWR VPWR _8431_/X sky130_fd_sc_hd__and2_1
X_5643_ _5629_/X hold830/X _5654_/S VGND VGND VPWR VPWR _5644_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8362_ _8363_/A _8377_/B VGND VGND VPWR VPWR _8388_/A sky130_fd_sc_hd__nor2_2
X_5574_ _5291_/X hold846/X _5582_/S VGND VGND VPWR VPWR _5575_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7313_ _7239_/X hold307/X _7319_/S VGND VGND VPWR VPWR _7313_/X sky130_fd_sc_hd__mux2_1
X_4525_ input50/X _4582_/A _7553_/A _9358_/Q _4524_/X VGND VGND VPWR VPWR _4530_/B
+ sky130_fd_sc_hd__a221o_1
Xhold201 _9414_/Q VGND VGND VPWR VPWR hold201/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 _9421_/Q VGND VGND VPWR VPWR hold212/X sky130_fd_sc_hd__dlygate4sd3_1
X_8293_ _8342_/B _8389_/A _8357_/A VGND VGND VPWR VPWR _8358_/A sky130_fd_sc_hd__and3_2
XFILLER_172_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold223 _7277_/X VGND VGND VPWR VPWR _7278_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 _7565_/X VGND VGND VPWR VPWR _7566_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7244_ _7244_/A VGND VGND VPWR VPWR _9213_/D sky130_fd_sc_hd__clkbuf_1
Xhold245 _7775_/X VGND VGND VPWR VPWR _7776_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold256 _9477_/Q VGND VGND VPWR VPWR hold256/X sky130_fd_sc_hd__dlygate4sd3_1
X_4456_ _9231_/Q _7266_/A _4455_/Y _9327_/Q VGND VGND VPWR VPWR _4463_/C sky130_fd_sc_hd__a22o_1
XFILLER_117_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold267 _9348_/Q VGND VGND VPWR VPWR hold267/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold278 _7366_/X VGND VGND VPWR VPWR _7367_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold289 _9236_/Q VGND VGND VPWR VPWR hold289/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7175_ _7175_/A VGND VGND VPWR VPWR _9183_/D sky130_fd_sc_hd__clkbuf_1
X_4387_ hold31/X hold82/X hold51/X VGND VGND VPWR VPWR hold83/A sky130_fd_sc_hd__or3b_1
XFILLER_86_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6126_ _6479_/A _6732_/B VGND VGND VPWR VPWR _6585_/A sky130_fd_sc_hd__nor2_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6057_ _6057_/A VGND VGND VPWR VPWR _9094_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5008_ _5068_/C _5021_/B hold8/A VGND VGND VPWR VPWR _5011_/A sky130_fd_sc_hd__o21ai_1
XFILLER_73_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 _6012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 _6416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_129 _7302_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6959_ _6959_/A _6959_/B _6959_/C _6959_/D VGND VGND VPWR VPWR _7000_/C sky130_fd_sc_hd__or4_1
XFILLER_186_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8629_ _8629_/A VGND VGND VPWR VPWR _9529_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold790 _9439_/Q VGND VGND VPWR VPWR hold790/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput306 _7911_/B VGND VGND VPWR VPWR serial_clock sky130_fd_sc_hd__buf_12
Xoutput317 _9148_/Q VGND VGND VPWR VPWR sram_ro_addr[1] sky130_fd_sc_hd__buf_12
Xoutput328 _9055_/Q VGND VGND VPWR VPWR wb_dat_o[10] sky130_fd_sc_hd__buf_12
XFILLER_114_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput339 _9044_/Q VGND VGND VPWR VPWR wb_dat_o[20] sky130_fd_sc_hd__buf_12
X_5290_ _5504_/A VGND VGND VPWR VPWR _7517_/A sky130_fd_sc_hd__buf_6
XFILLER_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8980_ _9005_/CLK _8980_/D fanout485/X VGND VGND VPWR VPWR _8980_/Q sky130_fd_sc_hd__dfstp_4
X_7931_ _7931_/A VGND VGND VPWR VPWR _7931_/X sky130_fd_sc_hd__buf_8
XFILLER_36_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7862_ _9488_/Q _9489_/Q _7863_/D _9490_/Q VGND VGND VPWR VPWR _7865_/B sky130_fd_sc_hd__a31o_1
XFILLER_63_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6813_ _6596_/B _6640_/Y _6518_/Y VGND VGND VPWR VPWR _6813_/X sky130_fd_sc_hd__a21o_1
X_7793_ _7793_/A VGND VGND VPWR VPWR _9461_/D sky130_fd_sc_hd__clkbuf_1
X_9532_ _9532_/CLK _9532_/D fanout446/X VGND VGND VPWR VPWR _9532_/Q sky130_fd_sc_hd__dfrtp_1
X_6744_ _6744_/A _6744_/B _6873_/B VGND VGND VPWR VPWR _6744_/X sky130_fd_sc_hd__or3_1
X_9463_ _9463_/CLK _9463_/D fanout410/X VGND VGND VPWR VPWR _9463_/Q sky130_fd_sc_hd__dfrtp_1
X_6675_ _6862_/A _6926_/A _6959_/B VGND VGND VPWR VPWR _6707_/C sky130_fd_sc_hd__o21bai_1
X_8414_ _9457_/Q _8348_/X _8411_/X _9337_/Q _8413_/X VGND VGND VPWR VPWR _8424_/B
+ sky130_fd_sc_hd__a221o_1
X_5626_ _5626_/A VGND VGND VPWR VPWR _8906_/D sky130_fd_sc_hd__clkbuf_1
X_9394_ _9471_/CLK _9394_/D _5070_/A VGND VGND VPWR VPWR _9394_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_164_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8345_ _8352_/A _8392_/A _8398_/A VGND VGND VPWR VPWR _8682_/B sky130_fd_sc_hd__and3_4
X_5557_ _5557_/A VGND VGND VPWR VPWR _8875_/D sky130_fd_sc_hd__clkbuf_1
X_4508_ _8808_/Q _8807_/Q _8806_/Q VGND VGND VPWR VPWR _4550_/S sky130_fd_sc_hd__nor3_2
X_8276_ _9078_/Q _8034_/A _8008_/B _8275_/X VGND VGND VPWR VPWR _8276_/X sky130_fd_sc_hd__a22o_1
XFILLER_2_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5488_ _5468_/X hold611/X _5490_/S VGND VGND VPWR VPWR _5488_/X sky130_fd_sc_hd__mux2_1
X_4439_ _4878_/A _4675_/B VGND VGND VPWR VPWR _4439_/Y sky130_fd_sc_hd__nor2_2
X_7227_ _7227_/A VGND VGND VPWR VPWR _9207_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout500 _8709_/B VGND VGND VPWR VPWR fanout500/X sky130_fd_sc_hd__clkbuf_2
XFILLER_160_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7158_ _7158_/A _7158_/B _7158_/C _7158_/D VGND VGND VPWR VPWR _7159_/A sky130_fd_sc_hd__or4_1
XFILLER_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6109_ _6182_/A VGND VGND VPWR VPWR _6716_/A sky130_fd_sc_hd__buf_4
XFILLER_86_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7089_ _5947_/X _9146_/Q _7089_/S VGND VGND VPWR VPWR _7089_/X sky130_fd_sc_hd__mux2_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4790_ _9442_/Q _7746_/A _6007_/A _9076_/Q _4789_/X VGND VGND VPWR VPWR _4791_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_18 _7746_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_29 _4570_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6460_ _6597_/B _6460_/B VGND VGND VPWR VPWR _6898_/A sky130_fd_sc_hd__nand2_2
XFILLER_9_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5411_ _8815_/Q _5410_/X _5416_/S VGND VGND VPWR VPWR _5411_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6391_ _6788_/B _6391_/B VGND VGND VPWR VPWR _6672_/C sky130_fd_sc_hd__nor2_2
XFILLER_173_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8130_ hold997/X _8017_/X _8128_/X _8129_/X VGND VGND VPWR VPWR _9512_/D sky130_fd_sc_hd__o22a_1
XFILLER_161_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5342_ _5342_/A VGND VGND VPWR VPWR _5342_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8061_ _9508_/Q _7920_/Y _8060_/X _8997_/Q VGND VGND VPWR VPWR _8061_/X sky130_fd_sc_hd__o22a_1
X_5273_ _9030_/Q _5287_/B VGND VGND VPWR VPWR _5274_/A sky130_fd_sc_hd__and2_1
XFILLER_99_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7012_ _7012_/A VGND VGND VPWR VPWR _7012_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8963_ _9482_/CLK _8963_/D fanout432/X VGND VGND VPWR VPWR _8963_/Q sky130_fd_sc_hd__dfrtp_4
X_7914_ _8015_/A _7914_/A1 _7914_/S VGND VGND VPWR VPWR _7915_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8894_ _9184_/CLK _8894_/D fanout432/X VGND VGND VPWR VPWR _8894_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_24_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7845_ _5410_/X hold320/X _7847_/S VGND VGND VPWR VPWR _7845_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7776_ _7776_/A VGND VGND VPWR VPWR _9453_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4988_ _4987_/X hold29/A _5014_/S VGND VGND VPWR VPWR _4989_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9515_ _9531_/CLK _9515_/D fanout452/X VGND VGND VPWR VPWR _9515_/Q sky130_fd_sc_hd__dfrtp_1
X_6727_ _6967_/A _6744_/B VGND VGND VPWR VPWR _6728_/B sky130_fd_sc_hd__or2_1
XFILLER_177_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9446_ _9486_/CLK _9446_/D fanout413/X VGND VGND VPWR VPWR _9446_/Q sky130_fd_sc_hd__dfrtp_1
X_6658_ _6658_/A _6781_/B VGND VGND VPWR VPWR _6809_/C sky130_fd_sc_hd__or2_1
XFILLER_192_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5609_ _5609_/A VGND VGND VPWR VPWR _8898_/D sky130_fd_sc_hd__clkbuf_1
X_9377_ _9483_/CLK _9377_/D fanout473/X VGND VGND VPWR VPWR _9377_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6589_ _6891_/A _6628_/A _6589_/C _6589_/D VGND VGND VPWR VPWR _6627_/C sky130_fd_sc_hd__and4_1
X_8328_ _9416_/Q _8402_/A _8327_/X _9256_/Q VGND VGND VPWR VPWR _8328_/X sky130_fd_sc_hd__a22o_1
XFILLER_105_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8259_ _9087_/Q _7940_/X _8003_/X _8886_/Q _8258_/X VGND VGND VPWR VPWR _8260_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput16 mask_rev_in[20] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput27 mask_rev_in[30] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput38 mgmt_gpio_in[11] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__clkbuf_4
Xinput49 mgmt_gpio_in[21] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__buf_2
XFILLER_6_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5960_ _9027_/Q _8709_/B VGND VGND VPWR VPWR _5961_/A sky130_fd_sc_hd__and2_1
X_4911_ _9400_/Q _4484_/Y _7043_/A _9126_/Q _4910_/X VGND VGND VPWR VPWR _4921_/A
+ sky130_fd_sc_hd__a221o_1
X_5891_ hold639/X hold15/X _5897_/S VGND VGND VPWR VPWR _5891_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7630_ _7433_/X _9387_/Q _7638_/S VGND VGND VPWR VPWR _7630_/X sky130_fd_sc_hd__mux2_1
X_4842_ hold92/A _4484_/Y _7815_/A _9473_/Q VGND VGND VPWR VPWR _4842_/X sky130_fd_sc_hd__a22o_1
XANTENNA_290 _4786_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7561_ _7433_/X _9355_/Q hold99/X VGND VGND VPWR VPWR _7561_/X sky130_fd_sc_hd__mux2_1
X_4773_ input26/X _4477_/Y _5806_/A _8985_/Q VGND VGND VPWR VPWR _4773_/X sky130_fd_sc_hd__a22o_2
XFILLER_193_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9300_ _9420_/CLK _9300_/D fanout465/X VGND VGND VPWR VPWR _9300_/Q sky130_fd_sc_hd__dfrtp_2
X_6512_ _6521_/B _6506_/Y _6508_/Y _6511_/Y VGND VGND VPWR VPWR _6517_/B sky130_fd_sc_hd__o22a_1
X_7492_ _7439_/X hold301/X _7497_/S VGND VGND VPWR VPWR _7492_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9231_ _9437_/CLK _9231_/D fanout419/X VGND VGND VPWR VPWR _9231_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6443_ _6596_/B _6818_/A VGND VGND VPWR VPWR _6444_/A sky130_fd_sc_hd__or2_1
XFILLER_134_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9162_ _9162_/CLK _9162_/D fanout440/X VGND VGND VPWR VPWR _9162_/Q sky130_fd_sc_hd__dfrtp_4
X_6374_ _6589_/C _6815_/B VGND VGND VPWR VPWR _6422_/B sky130_fd_sc_hd__nor2_4
X_8113_ _9349_/Q _8077_/X _7997_/X _9365_/Q VGND VGND VPWR VPWR _8113_/X sky130_fd_sc_hd__a22o_1
X_5325_ _5325_/A VGND VGND VPWR VPWR _5325_/X sky130_fd_sc_hd__clkbuf_1
X_9093_ _9194_/CLK _9093_/D fanout450/X VGND VGND VPWR VPWR _9093_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_115_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5256_ _9347_/Q VGND VGND VPWR VPWR _5256_/Y sky130_fd_sc_hd__inv_2
X_8044_ _9282_/Q _7952_/A _8003_/A _9298_/Q VGND VGND VPWR VPWR _8044_/X sky130_fd_sc_hd__a22o_1
XFILLER_87_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5187_ _5187_/A VGND VGND VPWR VPWR _5187_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8946_ _9051_/CLK _8946_/D fanout453/X VGND VGND VPWR VPWR _8946_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8877_ _9465_/CLK _8877_/D fanout471/X VGND VGND VPWR VPWR _8877_/Q sky130_fd_sc_hd__dfrtp_4
X_7828_ _5410_/X hold246/X _7830_/S VGND VGND VPWR VPWR _7828_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7759_ _7759_/A VGND VGND VPWR VPWR _9445_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9429_ _9453_/CLK _9429_/D fanout461/X VGND VGND VPWR VPWR _9429_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_164_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold608 _5515_/X VGND VGND VPWR VPWR _5516_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold619 _8965_/Q VGND VGND VPWR VPWR hold619/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5110_ _9219_/Q VGND VGND VPWR VPWR _5110_/Y sky130_fd_sc_hd__inv_2
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6090_ _6739_/A _6739_/B VGND VGND VPWR VPWR _6141_/A sky130_fd_sc_hd__or2_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _5041_/A VGND VGND VPWR VPWR _5065_/S sky130_fd_sc_hd__buf_6
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8800_ _5168_/A1 _8800_/D _5368_/X VGND VGND VPWR VPWR hold39/A sky130_fd_sc_hd__dfrtp_1
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR rebuffer3/A sky130_fd_sc_hd__clkbuf_16
XFILLER_38_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6992_ _6830_/A _6967_/C _6266_/X VGND VGND VPWR VPWR _6993_/D sky130_fd_sc_hd__o21ai_1
X_8731_ _8731_/A _8732_/A VGND VGND VPWR VPWR _8731_/Y sky130_fd_sc_hd__nand2_1
XFILLER_92_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5943_ _9046_/Q _4549_/X _5945_/S VGND VGND VPWR VPWR _5944_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8662_ hold71/A _8372_/X _8369_/X _8906_/Q _8661_/X VGND VGND VPWR VPWR _8663_/D
+ sky130_fd_sc_hd__a221o_1
X_5874_ _5413_/S _8706_/A _5149_/A _5870_/X _6908_/A VGND VGND VPWR VPWR _9008_/D
+ sky130_fd_sc_hd__a2111o_4
XFILLER_139_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7613_ _9379_/Q hold46/X _7621_/S VGND VGND VPWR VPWR _7613_/X sky130_fd_sc_hd__mux2_1
X_4825_ input53/X _4491_/Y _4898_/A2 _9481_/Q VGND VGND VPWR VPWR _4825_/X sky130_fd_sc_hd__a22o_1
X_8593_ _9074_/Q _8322_/X _8333_/X _8863_/Q _8592_/X VGND VGND VPWR VPWR _8601_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_193_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7544_ _7544_/A VGND VGND VPWR VPWR _9347_/D sky130_fd_sc_hd__clkbuf_1
X_4756_ _9290_/Q _7408_/A _5762_/A _8965_/Q VGND VGND VPWR VPWR _4756_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7475_ hold332/X _5465_/A _7479_/S VGND VGND VPWR VPWR _7475_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4687_ _9372_/Q _7588_/A _5630_/A _8912_/Q _4686_/X VGND VGND VPWR VPWR _4688_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9214_ _9462_/CLK _9214_/D fanout408/X VGND VGND VPWR VPWR _9214_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_146_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6426_ _6435_/A _6900_/A VGND VGND VPWR VPWR _6843_/C sky130_fd_sc_hd__or2_1
XFILLER_162_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9145_ _9462_/CLK _9145_/D fanout408/X VGND VGND VPWR VPWR _9145_/Q sky130_fd_sc_hd__dfrtp_4
X_6357_ _6217_/B _6839_/A _6330_/Y _6356_/X VGND VGND VPWR VPWR _6357_/X sky130_fd_sc_hd__a211o_1
XFILLER_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5308_ _5308_/A VGND VGND VPWR VPWR _8774_/D sky130_fd_sc_hd__clkbuf_1
X_9076_ _9162_/CLK _9076_/D fanout437/X VGND VGND VPWR VPWR _9076_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_88_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6288_ _6895_/A _6906_/C _6524_/B VGND VGND VPWR VPWR _6710_/A sky130_fd_sc_hd__nor3_1
XFILLER_102_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8027_ _8027_/A _8027_/B _8027_/C _8027_/D VGND VGND VPWR VPWR _8027_/X sky130_fd_sc_hd__or4_2
X_5239_ _9203_/Q VGND VGND VPWR VPWR _5239_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8929_ _9473_/CLK _8929_/D fanout438/X VGND VGND VPWR VPWR _8929_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_140_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold5 hold5/A VGND VGND VPWR VPWR hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_181_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4610_ _8907_/Q _5618_/A _5795_/A _8982_/Q _4609_/X VGND VGND VPWR VPWR _4617_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_175_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5590_ hold784/X _5395_/X _5594_/S VGND VGND VPWR VPWR _5591_/A sky130_fd_sc_hd__mux2_1
X_4541_ _9342_/Q _4414_/Y _4938_/A2 _9278_/Q _4540_/X VGND VGND VPWR VPWR _4548_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold405 hold405/A VGND VGND VPWR VPWR hold405/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold416 _7150_/X VGND VGND VPWR VPWR _7151_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7260_ _7242_/X hold260/X _7264_/S VGND VGND VPWR VPWR _7260_/X sky130_fd_sc_hd__mux2_1
X_4472_ _9479_/Q _7815_/A _7056_/A _9139_/Q VGND VGND VPWR VPWR _4472_/X sky130_fd_sc_hd__a22o_1
XFILLER_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold427 _7683_/X VGND VGND VPWR VPWR _7684_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 _5513_/X VGND VGND VPWR VPWR _5514_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 _8896_/Q VGND VGND VPWR VPWR hold449/X sky130_fd_sc_hd__dlygate4sd3_1
X_6211_ _6345_/A _6345_/B VGND VGND VPWR VPWR _6216_/A sky130_fd_sc_hd__nand2_2
X_7191_ _7191_/A VGND VGND VPWR VPWR _9190_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6142_ _6142_/A VGND VGND VPWR VPWR _6876_/B sky130_fd_sc_hd__clkbuf_4
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ hold71/X hold46/X _6075_/S VGND VGND VPWR VPWR hold72/A sky130_fd_sc_hd__mux2_1
XFILLER_97_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1105 _7135_/X VGND VGND VPWR VPWR hold793/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1116 _9089_/Q VGND VGND VPWR VPWR hold883/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1127 _8929_/Q VGND VGND VPWR VPWR hold588/A sky130_fd_sc_hd__dlygate4sd3_1
X_5024_ _5068_/C _5039_/B VGND VGND VPWR VPWR _5025_/B sky130_fd_sc_hd__nand2_1
XFILLER_57_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1138 _8953_/Q VGND VGND VPWR VPWR hold869/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 _5853_/X VGND VGND VPWR VPWR hold1149/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6975_ _6887_/Y _6973_/X _6974_/Y _6889_/X VGND VGND VPWR VPWR _6998_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8714_ _8714_/A VGND VGND VPWR VPWR _9535_/D sky130_fd_sc_hd__clkbuf_1
X_5926_ _5926_/A VGND VGND VPWR VPWR _9038_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8645_ _8940_/Q _7908_/A _8358_/C _8870_/Q VGND VGND VPWR VPWR _8645_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5857_ _5857_/A VGND VGND VPWR VPWR _9003_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4808_ _9186_/Q _7176_/A _7446_/A _9306_/Q _4807_/X VGND VGND VPWR VPWR _4816_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_166_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8576_ _8701_/A _8576_/B _8576_/C _8576_/D VGND VGND VPWR VPWR _8576_/X sky130_fd_sc_hd__or4_1
X_5788_ _5788_/A VGND VGND VPWR VPWR _8974_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7527_ _7527_/A VGND VGND VPWR VPWR _9339_/D sky130_fd_sc_hd__clkbuf_1
X_4739_ _4739_/A1 _4444_/Y _4406_/Y input6/X VGND VGND VPWR VPWR _4739_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7458_ _7458_/A VGND VGND VPWR VPWR _9309_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6409_ _6628_/B _6409_/B VGND VGND VPWR VPWR _6469_/B sky130_fd_sc_hd__nor2_1
Xhold950 _5152_/X VGND VGND VPWR VPWR _8828_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold961 _9113_/Q VGND VGND VPWR VPWR hold961/X sky130_fd_sc_hd__dlygate4sd3_1
X_7389_ _7299_/X hold533/X _7389_/S VGND VGND VPWR VPWR _7389_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold972 _9116_/Q VGND VGND VPWR VPWR hold972/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9128_ _9485_/CLK _9128_/D fanout405/X VGND VGND VPWR VPWR _9128_/Q sky130_fd_sc_hd__dfrtp_4
Xhold983 _9525_/Q VGND VGND VPWR VPWR hold983/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 _8778_/Q VGND VGND VPWR VPWR hold994/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9059_ _9541_/CLK _9059_/D VGND VGND VPWR VPWR _9059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_50_csclk _9090_/CLK VGND VGND VPWR VPWR _9187_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_141_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_65_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _9482_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_48_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6760_ _6422_/B _6462_/B _6706_/A _6553_/B VGND VGND VPWR VPWR _6761_/C sky130_fd_sc_hd__a211o_1
XFILLER_62_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5711_ hold505/X _5687_/X _5713_/S VGND VGND VPWR VPWR _5712_/A sky130_fd_sc_hd__mux2_1
X_6691_ _6691_/A _6470_/A VGND VGND VPWR VPWR _6695_/B sky130_fd_sc_hd__or2b_1
X_8430_ _9418_/Q _8402_/X _8378_/X _9354_/Q _8429_/X VGND VGND VPWR VPWR _8437_/A
+ sky130_fd_sc_hd__a221o_1
X_5642_ _5642_/A _5693_/B VGND VGND VPWR VPWR _5654_/S sky130_fd_sc_hd__nand2_4
X_8361_ _8361_/A _8361_/B _8361_/C _8361_/D VGND VGND VPWR VPWR _8398_/C sky130_fd_sc_hd__or4_1
XFILLER_176_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5573_ _5573_/A _5693_/B VGND VGND VPWR VPWR _5582_/S sky130_fd_sc_hd__nand2_2
XFILLER_129_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7312_ _7312_/A VGND VGND VPWR VPWR _9243_/D sky130_fd_sc_hd__clkbuf_1
X_4524_ _9422_/Q _4439_/Y _7056_/A _9138_/Q VGND VGND VPWR VPWR _4524_/X sky130_fd_sc_hd__a22o_1
Xhold202 _7691_/X VGND VGND VPWR VPWR _7692_/A sky130_fd_sc_hd__dlygate4sd3_1
X_8292_ _8292_/A VGND VGND VPWR VPWR _8292_/X sky130_fd_sc_hd__buf_6
Xhold213 _7706_/X VGND VGND VPWR VPWR _7707_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 hold224/A VGND VGND VPWR VPWR hold224/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_18_csclk _9303_/CLK VGND VGND VPWR VPWR _9328_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold235 hold235/A VGND VGND VPWR VPWR hold235/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 _9478_/Q VGND VGND VPWR VPWR hold246/X sky130_fd_sc_hd__dlygate4sd3_1
X_7243_ _7242_/X hold180/X _7247_/S VGND VGND VPWR VPWR _7243_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4455_ _4861_/A _4674_/A VGND VGND VPWR VPWR _4455_/Y sky130_fd_sc_hd__nor2_2
Xhold257 _7826_/X VGND VGND VPWR VPWR _7827_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 _9241_/Q VGND VGND VPWR VPWR hold268/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 _9285_/Q VGND VGND VPWR VPWR hold279/X sky130_fd_sc_hd__dlygate4sd3_1
X_4386_ hold74/A hold30/X hold57/X VGND VGND VPWR VPWR hold31/A sky130_fd_sc_hd__o21ai_1
X_7174_ _5471_/X hold567/X _7174_/S VGND VGND VPWR VPWR _7174_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6125_ _6125_/A VGND VGND VPWR VPWR _6732_/B sky130_fd_sc_hd__buf_6
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _5947_/X hold862/X _6064_/S VGND VGND VPWR VPWR _6057_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5007_ _8827_/Q VGND VGND VPWR VPWR _5068_/C sky130_fd_sc_hd__buf_2
XFILLER_45_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_108 _6012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_119 _6850_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6958_ _6958_/A _6958_/B _6958_/C VGND VGND VPWR VPWR _7004_/A sky130_fd_sc_hd__nor3_1
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5909_ _5909_/A VGND VGND VPWR VPWR _5909_/X sky130_fd_sc_hd__clkbuf_1
X_6889_ _6521_/B _6508_/Y _6822_/X _6888_/X VGND VGND VPWR VPWR _6889_/X sky130_fd_sc_hd__a211o_1
XFILLER_22_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8628_ _8628_/A0 _8627_/X _8653_/S VGND VGND VPWR VPWR _8629_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8559_ _9455_/Q _8360_/A _8381_/A _9367_/Q VGND VGND VPWR VPWR _8559_/X sky130_fd_sc_hd__a22o_1
XFILLER_108_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold780 _7216_/X VGND VGND VPWR VPWR _7217_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold791 _7744_/X VGND VGND VPWR VPWR _7745_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput307 _4562_/X VGND VGND VPWR VPWR serial_data_1 sky130_fd_sc_hd__buf_12
Xoutput318 _9149_/Q VGND VGND VPWR VPWR sram_ro_addr[2] sky130_fd_sc_hd__buf_12
Xoutput329 _9056_/Q VGND VGND VPWR VPWR wb_dat_o[11] sky130_fd_sc_hd__buf_12
XFILLER_114_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7930_ _7998_/A _7989_/B _8000_/B VGND VGND VPWR VPWR _7931_/A sky130_fd_sc_hd__and3_1
X_7861_ _7861_/A1 _7857_/Y _7860_/Y _7851_/Y VGND VGND VPWR VPWR _9489_/D sky130_fd_sc_hd__a22o_1
XFILLER_63_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6812_ _6815_/B _6967_/C VGND VGND VPWR VPWR _6812_/Y sky130_fd_sc_hd__nand2_2
X_7792_ _7654_/X hold176/X _7796_/S VGND VGND VPWR VPWR _7792_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9531_ _9531_/CLK _9531_/D fanout446/X VGND VGND VPWR VPWR _9531_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_189_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6743_ _6719_/Y _6128_/X _6742_/Y _6657_/B _6603_/Y VGND VGND VPWR VPWR _6946_/B
+ sky130_fd_sc_hd__a311o_1
X_9462_ _9462_/CLK _9462_/D fanout408/X VGND VGND VPWR VPWR _9462_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6674_ _6895_/B _6425_/X _6939_/A VGND VGND VPWR VPWR _6835_/B sky130_fd_sc_hd__o21ai_1
X_8413_ _9441_/Q _8301_/A _8344_/X _9481_/Q _8412_/X VGND VGND VPWR VPWR _8413_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_191_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5625_ hold435/X _5398_/X _5627_/S VGND VGND VPWR VPWR _5626_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9393_ _9427_/CLK _9393_/D fanout476/X VGND VGND VPWR VPWR _9393_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_191_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8344_ _8356_/C VGND VGND VPWR VPWR _8344_/X sky130_fd_sc_hd__buf_4
XFILLER_117_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5556_ _5306_/X hold540/X _5560_/S VGND VGND VPWR VPWR _5556_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4507_ _4507_/A _4507_/B VGND VGND VPWR VPWR _4507_/X sky130_fd_sc_hd__or2_4
XFILLER_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8275_ _9103_/Q _8275_/B VGND VGND VPWR VPWR _8275_/X sky130_fd_sc_hd__or2_1
X_5487_ _5487_/A VGND VGND VPWR VPWR _8845_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7226_ _5471_/X hold626/X _7226_/S VGND VGND VPWR VPWR _7226_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4438_ _4492_/A _4635_/A VGND VGND VPWR VPWR _4438_/Y sky130_fd_sc_hd__nor2_2
XFILLER_116_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout501 _5929_/B VGND VGND VPWR VPWR _8709_/B sky130_fd_sc_hd__buf_2
XFILLER_132_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7157_ _7157_/A VGND VGND VPWR VPWR _7157_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4369_ hold63/X hold41/X VGND VGND VPWR VPWR _4402_/B sky130_fd_sc_hd__nor2b_4
XFILLER_116_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6108_ _6479_/A _6779_/A VGND VGND VPWR VPWR _6754_/A sky130_fd_sc_hd__nor2_1
X_7088_ _7088_/A VGND VGND VPWR VPWR _9145_/D sky130_fd_sc_hd__clkbuf_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6039_ hold500/X _5687_/X _6041_/S VGND VGND VPWR VPWR _6040_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_19 _7158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5410_ hold27/X VGND VGND VPWR VPWR _5410_/X sky130_fd_sc_hd__buf_4
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6390_ _6470_/A _6691_/A _6667_/A _6471_/C VGND VGND VPWR VPWR _6670_/B sky130_fd_sc_hd__and4_1
XFILLER_126_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5341_ _5353_/A _5356_/B VGND VGND VPWR VPWR _5342_/A sky130_fd_sc_hd__and2_1
XFILLER_142_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8060_ _9186_/Q _8009_/A _8050_/X _8059_/X VGND VGND VPWR VPWR _8060_/X sky130_fd_sc_hd__o22a_1
X_5272_ _5272_/A VGND VGND VPWR VPWR _9029_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7011_ _7011_/A _7013_/B VGND VGND VPWR VPWR _7012_/A sky130_fd_sc_hd__and2_1
XFILLER_114_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8962_ _9087_/CLK _8962_/D fanout446/X VGND VGND VPWR VPWR _8962_/Q sky130_fd_sc_hd__dfrtp_4
X_7913_ _7858_/Y _7869_/Y _7912_/X _8999_/Q VGND VGND VPWR VPWR _7914_/S sky130_fd_sc_hd__a22o_1
X_8893_ _9484_/CLK _8893_/D fanout430/X VGND VGND VPWR VPWR _8893_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_70_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7844_ _7844_/A VGND VGND VPWR VPWR _9485_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7775_ _7654_/X hold244/X _7779_/S VGND VGND VPWR VPWR _7775_/X sky130_fd_sc_hd__mux2_1
X_4987_ _5021_/B _4983_/S _4986_/X hold56/A VGND VGND VPWR VPWR _4987_/X sky130_fd_sc_hd__a31o_1
XFILLER_168_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9514_ _9531_/CLK _9514_/D fanout452/X VGND VGND VPWR VPWR _9514_/Q sky130_fd_sc_hd__dfrtp_1
X_6726_ _6726_/A _6726_/B _6726_/C VGND VGND VPWR VPWR _6863_/D sky130_fd_sc_hd__or3_1
XFILLER_149_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9445_ _9485_/CLK _9445_/D fanout411/X VGND VGND VPWR VPWR _9445_/Q sky130_fd_sc_hd__dfrtp_1
X_6657_ _6657_/A _6657_/B _6915_/A _6657_/D VGND VGND VPWR VPWR _6659_/C sky130_fd_sc_hd__or4_1
XFILLER_177_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5608_ _5291_/X hold845/X _5616_/S VGND VGND VPWR VPWR _5609_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9376_ _9376_/CLK _9376_/D fanout416/X VGND VGND VPWR VPWR _9376_/Q sky130_fd_sc_hd__dfstp_1
X_6588_ _6588_/A _6588_/B VGND VGND VPWR VPWR _6924_/C sky130_fd_sc_hd__or2_2
XFILLER_191_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8327_ _8364_/A VGND VGND VPWR VPWR _8327_/X sky130_fd_sc_hd__buf_8
XFILLER_152_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5539_ _5539_/A VGND VGND VPWR VPWR _8867_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8258_ _8906_/Q _7962_/X _7977_/X _8775_/Q VGND VGND VPWR VPWR _8258_/X sky130_fd_sc_hd__a22o_1
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7209_ _5471_/X hold631/X _7209_/S VGND VGND VPWR VPWR _7209_/X sky130_fd_sc_hd__mux2_1
X_8189_ _8968_/Q _7967_/A _8068_/B _8948_/Q VGND VGND VPWR VPWR _8189_/X sky130_fd_sc_hd__a22o_1
XFILLER_120_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput17 mask_rev_in[21] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__buf_2
Xinput28 mask_rev_in[31] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput39 mgmt_gpio_in[12] VGND VGND VPWR VPWR _5285_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_183_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4910_ _9200_/Q _7211_/A _5738_/A _8953_/Q VGND VGND VPWR VPWR _4910_/X sky130_fd_sc_hd__a22o_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5890_ _5890_/A VGND VGND VPWR VPWR _9013_/D sky130_fd_sc_hd__clkbuf_1
X_4841_ _4841_/A _4841_/B _4841_/C _4841_/D VGND VGND VPWR VPWR _4853_/B sky130_fd_sc_hd__or4_1
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_280 input38/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_291 _9123_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7560_ _7560_/A VGND VGND VPWR VPWR _9354_/D sky130_fd_sc_hd__clkbuf_1
X_4772_ _4772_/A _4772_/B _4772_/C _4772_/D VGND VGND VPWR VPWR _4782_/B sky130_fd_sc_hd__or4_2
XFILLER_159_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6511_ _6887_/A _6499_/B _6509_/X _6510_/Y VGND VGND VPWR VPWR _6511_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_186_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7491_ _7491_/A VGND VGND VPWR VPWR _9324_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9230_ _9437_/CLK _9230_/D fanout419/X VGND VGND VPWR VPWR _9230_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6442_ _6527_/A _6926_/A VGND VGND VPWR VPWR _6842_/B sky130_fd_sc_hd__nor2_1
XFILLER_146_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9161_ _9161_/CLK _9161_/D fanout442/X VGND VGND VPWR VPWR _9161_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6373_ _6373_/A VGND VGND VPWR VPWR _6815_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_173_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A VGND VGND VPWR VPWR _9531_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8112_ _9405_/Q _7931_/X _7990_/X _9277_/Q _8111_/X VGND VGND VPWR VPWR _8117_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_114_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5324_ _5330_/A _5334_/B VGND VGND VPWR VPWR _5325_/A sky130_fd_sc_hd__and2_1
X_9092_ _9092_/CLK _9092_/D fanout451/X VGND VGND VPWR VPWR _9092_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_115_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8043_ _9370_/Q _7960_/A _8001_/A _9266_/Q _8042_/X VGND VGND VPWR VPWR _8050_/A
+ sky130_fd_sc_hd__a221o_1
X_5255_ _9339_/Q VGND VGND VPWR VPWR _5255_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5186_ _9175_/Q input91/X _5194_/S VGND VGND VPWR VPWR _5187_/A sky130_fd_sc_hd__mux2_2
XFILLER_3_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8945_ _9088_/CLK _8945_/D fanout454/X VGND VGND VPWR VPWR _8945_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_113_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8876_ _9251_/CLK _8876_/D fanout486/X VGND VGND VPWR VPWR _8876_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_36_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7827_ _7827_/A VGND VGND VPWR VPWR _9477_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7758_ hold291/X _5465_/A _7762_/S VGND VGND VPWR VPWR _7758_/X sky130_fd_sc_hd__mux2_1
X_6709_ _6924_/B _6709_/B _6709_/C _6709_/D VGND VGND VPWR VPWR _6710_/D sky130_fd_sc_hd__or4_1
X_7689_ _7654_/X hold250/X _7693_/S VGND VGND VPWR VPWR _7689_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9428_ _9468_/CLK _9428_/D fanout465/X VGND VGND VPWR VPWR _9428_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_164_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9359_ _9359_/CLK _9359_/D fanout422/X VGND VGND VPWR VPWR _9359_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold609 hold609/A VGND VGND VPWR VPWR hold609/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _8827_/Q _5040_/B _5040_/C VGND VGND VPWR VPWR _5041_/A sky130_fd_sc_hd__or3_1
XFILLER_69_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6991_ _7004_/A _6962_/X _6980_/X _6990_/Y VGND VGND VPWR VPWR _9109_/D sky130_fd_sc_hd__a211o_1
XFILLER_93_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8730_ _8732_/A _8769_/A2 _9033_/Q VGND VGND VPWR VPWR _8735_/B sky130_fd_sc_hd__a21boi_1
XFILLER_92_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5942_ _5942_/A VGND VGND VPWR VPWR _9045_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8661_ _8886_/Q _8314_/X _8331_/X _8981_/Q VGND VGND VPWR VPWR _8661_/X sky130_fd_sc_hd__a22o_1
X_5873_ _5873_/A VGND VGND VPWR VPWR _6908_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_34_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7612_ _7612_/A VGND VGND VPWR VPWR _9378_/D sky130_fd_sc_hd__clkbuf_1
X_4824_ _8810_/Q _5388_/A _7113_/A _9162_/Q _4823_/X VGND VGND VPWR VPWR _4829_/B
+ sky130_fd_sc_hd__a221o_1
X_8592_ _8873_/Q _8316_/X _8327_/X _9089_/Q VGND VGND VPWR VPWR _8592_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7543_ _7433_/X _9347_/Q _7551_/S VGND VGND VPWR VPWR _7543_/X sky130_fd_sc_hd__mux2_1
X_4755_ _4755_/A VGND VGND VPWR VPWR _9114_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7474_ _7474_/A VGND VGND VPWR VPWR _9316_/D sky130_fd_sc_hd__clkbuf_1
X_4686_ _9324_/Q _7481_/A _6055_/A _9098_/Q VGND VGND VPWR VPWR _4686_/X sky130_fd_sc_hd__a22o_1
X_9213_ _9437_/CLK _9213_/D fanout419/X VGND VGND VPWR VPWR _9213_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6425_ _6535_/A _6887_/B VGND VGND VPWR VPWR _6425_/X sky130_fd_sc_hd__or2_1
XFILLER_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9144_ _9162_/CLK _9144_/D fanout440/X VGND VGND VPWR VPWR _9144_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6356_ _6331_/Y _6839_/A _6758_/A _6872_/B _6355_/X VGND VGND VPWR VPWR _6356_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_161_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5307_ _5306_/X hold514/X _5316_/S VGND VGND VPWR VPWR _5307_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9075_ _9162_/CLK _9075_/D fanout436/X VGND VGND VPWR VPWR _9075_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_170_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6287_ _6437_/A _6716_/A _6596_/B VGND VGND VPWR VPWR _6524_/B sky130_fd_sc_hd__or3_2
XFILLER_102_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8026_ _9217_/Q _7927_/X _7962_/X _9321_/Q _8025_/X VGND VGND VPWR VPWR _8027_/D
+ sky130_fd_sc_hd__a221o_1
X_5238_ _9211_/Q VGND VGND VPWR VPWR _5238_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5169_ _5169_/A VGND VGND VPWR VPWR _5169_/X sky130_fd_sc_hd__buf_1
XFILLER_56_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8928_ _9484_/CLK _8928_/D fanout432/X VGND VGND VPWR VPWR _8928_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8859_ _9184_/CLK _8859_/D fanout443/X VGND VGND VPWR VPWR _8859_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_40_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold6 hold6/A VGND VGND VPWR VPWR hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4540_ _9374_/Q _7588_/A _7113_/A _4539_/X VGND VGND VPWR VPWR _4540_/X sky130_fd_sc_hd__a22o_1
XFILLER_190_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4471_ _4499_/A _4891_/B VGND VGND VPWR VPWR _7056_/A sky130_fd_sc_hd__nor2_8
Xhold406 hold406/A VGND VGND VPWR VPWR hold406/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold417 _7151_/X VGND VGND VPWR VPWR _9172_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold428 _5426_/X VGND VGND VPWR VPWR _5427_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 _8914_/Q VGND VGND VPWR VPWR hold439/X sky130_fd_sc_hd__dlygate4sd3_1
X_6210_ _6721_/A _6232_/C VGND VGND VPWR VPWR _6345_/B sky130_fd_sc_hd__nor2_1
XFILLER_116_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7190_ hold322/X _7494_/A _7192_/S VGND VGND VPWR VPWR _7190_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6141_ _6141_/A _6732_/A _6623_/A VGND VGND VPWR VPWR _6142_/A sky130_fd_sc_hd__or3_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ _6072_/A VGND VGND VPWR VPWR _9101_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1106 _9316_/Q VGND VGND VPWR VPWR hold334/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1117 _9282_/Q VGND VGND VPWR VPWR hold771/A sky130_fd_sc_hd__dlygate4sd3_1
X_5023_ _8808_/Q _8807_/Q VGND VGND VPWR VPWR _5039_/B sky130_fd_sc_hd__and2_1
Xhold1128 _9290_/Q VGND VGND VPWR VPWR hold787/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1139 _5403_/X VGND VGND VPWR VPWR hold576/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6974_ _6891_/A _6628_/A _6973_/A _6736_/B VGND VGND VPWR VPWR _6974_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_41_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5925_ _5650_/X hold851/X _5927_/S VGND VGND VPWR VPWR _5926_/A sky130_fd_sc_hd__mux2_1
X_8713_ _9535_/Q _4885_/X _8725_/S VGND VGND VPWR VPWR _8714_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8644_ _9071_/Q _8388_/A _8379_/A _9037_/Q _8643_/X VGND VGND VPWR VPWR _8649_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_110_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5856_ _9565_/A _5855_/X _5868_/S VGND VGND VPWR VPWR _5856_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4807_ _9410_/Q _7678_/A _5773_/A _8970_/Q VGND VGND VPWR VPWR _4807_/X sky130_fd_sc_hd__a22o_1
X_8575_ _8575_/A _8575_/B _8575_/C _8575_/D VGND VGND VPWR VPWR _8576_/D sky130_fd_sc_hd__or4_1
X_5787_ hold768/X _5587_/X _5793_/S VGND VGND VPWR VPWR _5788_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7526_ _7433_/X _9339_/Q _7534_/S VGND VGND VPWR VPWR _7526_/X sky130_fd_sc_hd__mux2_1
X_4738_ _9331_/Q _7499_/A _7481_/A _9323_/Q _4737_/X VGND VGND VPWR VPWR _4741_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_147_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7457_ _7439_/X hold231/X _7461_/S VGND VGND VPWR VPWR _7457_/X sky130_fd_sc_hd__mux2_1
XFILLER_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4669_ _9039_/Q _5918_/A _5642_/A _8917_/Q _4668_/X VGND VGND VPWR VPWR _4673_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_107_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_646 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6408_ _6635_/A _6894_/B VGND VGND VPWR VPWR _6409_/B sky130_fd_sc_hd__or2_1
Xhold940 hold940/A VGND VGND VPWR VPWR hold940/X sky130_fd_sc_hd__dlygate4sd3_1
X_7388_ _7388_/A VGND VGND VPWR VPWR _9278_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold951 _8831_/Q VGND VGND VPWR VPWR _5019_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 _4819_/X VGND VGND VPWR VPWR _4820_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9127_ _9485_/CLK _9127_/D fanout405/X VGND VGND VPWR VPWR _9127_/Q sky130_fd_sc_hd__dfstp_2
Xhold973 _4593_/X VGND VGND VPWR VPWR _4594_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_134_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold984 _9118_/Q VGND VGND VPWR VPWR hold984/X sky130_fd_sc_hd__dlygate4sd3_1
X_6339_ _6881_/A _6666_/B VGND VGND VPWR VPWR _6759_/A sky130_fd_sc_hd__nor2_1
XFILLER_150_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold995 _5163_/Y VGND VGND VPWR VPWR _8830_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9058_ _9541_/CLK _9058_/D VGND VGND VPWR VPWR _9058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8009_ _8009_/A VGND VGND VPWR VPWR _8010_/B sky130_fd_sc_hd__buf_4
XFILLER_130_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5710_ _5710_/A VGND VGND VPWR VPWR _8940_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6690_ _6673_/B _6481_/A _6670_/B _6483_/B VGND VGND VPWR VPWR _6763_/A sky130_fd_sc_hd__a31o_1
XFILLER_188_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5641_ _5641_/A VGND VGND VPWR VPWR _8912_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8360_ _8360_/A _8360_/B _8360_/C _8379_/A VGND VGND VPWR VPWR _8361_/D sky130_fd_sc_hd__or4_1
X_5572_ _5572_/A VGND VGND VPWR VPWR _8882_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_1_csclk clkbuf_1_0_1_csclk/A VGND VGND VPWR VPWR clkbuf_2_1_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
X_7311_ _7236_/X _9243_/Q _7319_/S VGND VGND VPWR VPWR _7311_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4523_ _9198_/Q _4424_/Y _5418_/A _8823_/Q _4522_/X VGND VGND VPWR VPWR _4530_/A
+ sky130_fd_sc_hd__a221o_1
X_8291_ _8342_/B _8336_/A _8357_/B VGND VGND VPWR VPWR _8292_/A sky130_fd_sc_hd__and3_2
XFILLER_144_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold203 hold203/A VGND VGND VPWR VPWR _7185_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 _9204_/Q VGND VGND VPWR VPWR hold214/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 _9405_/Q VGND VGND VPWR VPWR hold225/X sky130_fd_sc_hd__dlygate4sd3_1
X_7242_ hold15/X VGND VGND VPWR VPWR _7242_/X sky130_fd_sc_hd__buf_4
X_4454_ _4878_/A _4667_/A VGND VGND VPWR VPWR _4454_/Y sky130_fd_sc_hd__nor2_4
Xhold236 _9349_/Q VGND VGND VPWR VPWR hold236/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold247 _7828_/X VGND VGND VPWR VPWR _7829_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 _9356_/Q VGND VGND VPWR VPWR hold258/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 _7307_/X VGND VGND VPWR VPWR _7308_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7173_ _7173_/A VGND VGND VPWR VPWR _9182_/D sky130_fd_sc_hd__clkbuf_1
X_4385_ _4396_/A _4555_/A VGND VGND VPWR VPWR _4670_/B sky130_fd_sc_hd__nand2_8
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6124_ _6498_/B _6828_/B VGND VGND VPWR VPWR _6125_/A sky130_fd_sc_hd__nand2_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _6055_/A _7043_/B VGND VGND VPWR VPWR _6064_/S sky130_fd_sc_hd__nand2_2
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _5006_/A VGND VGND VPWR VPWR _8800_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_109 _6015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6957_ _6957_/A _6957_/B _6957_/C VGND VGND VPWR VPWR _6958_/C sky130_fd_sc_hd__or3_1
XFILLER_54_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5908_ _5650_/X _9581_/A _5916_/S VGND VGND VPWR VPWR _5908_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6888_ _6973_/A _6897_/B _6887_/Y _6446_/X VGND VGND VPWR VPWR _6888_/X sky130_fd_sc_hd__a31o_1
X_5839_ hold821/X hold27/X _5842_/S VGND VGND VPWR VPWR _5839_/X sky130_fd_sc_hd__mux2_1
X_8627_ _9528_/Q _8626_/X _8627_/S VGND VGND VPWR VPWR _8627_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8558_ _9351_/Q _8386_/X _8506_/B _9415_/Q _8557_/X VGND VGND VPWR VPWR _8563_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_108_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7509_ _7509_/A VGND VGND VPWR VPWR _9332_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8489_ _9220_/Q _8391_/X _8367_/X _9476_/Q _8488_/X VGND VGND VPWR VPWR _8489_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_108_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold770 _7289_/X VGND VGND VPWR VPWR _7290_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 hold781/A VGND VGND VPWR VPWR hold781/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold792 _7035_/X VGND VGND VPWR VPWR _7036_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput308 _4539_/X VGND VGND VPWR VPWR serial_data_2 sky130_fd_sc_hd__buf_12
Xoutput319 _9150_/Q VGND VGND VPWR VPWR sram_ro_addr[3] sky130_fd_sc_hd__buf_12
XFILLER_5_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7860_ _7860_/A _7860_/B VGND VGND VPWR VPWR _7860_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6811_ _6811_/A _6811_/B _6811_/C VGND VGND VPWR VPWR _6824_/C sky130_fd_sc_hd__and3_1
X_7791_ _7791_/A VGND VGND VPWR VPWR _9460_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9530_ _9531_/CLK _9530_/D fanout448/X VGND VGND VPWR VPWR _9530_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_51_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6742_ _6744_/A _6742_/B VGND VGND VPWR VPWR _6742_/Y sky130_fd_sc_hd__nor2_1
XFILLER_189_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9461_ _9461_/CLK _9461_/D fanout423/X VGND VGND VPWR VPWR _9461_/Q sky130_fd_sc_hd__dfrtp_1
X_6673_ _6673_/A _6673_/B VGND VGND VPWR VPWR _6939_/A sky130_fd_sc_hd__nand2_1
XFILLER_176_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8412_ _9217_/Q _8391_/A _8367_/A _9473_/Q VGND VGND VPWR VPWR _8412_/X sky130_fd_sc_hd__a22o_1
XFILLER_31_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5624_ _5624_/A VGND VGND VPWR VPWR _8905_/D sky130_fd_sc_hd__clkbuf_1
X_9392_ _9392_/CLK _9392_/D fanout425/X VGND VGND VPWR VPWR _9392_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_176_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8343_ _8355_/A _8377_/B VGND VGND VPWR VPWR _8356_/C sky130_fd_sc_hd__nor2_4
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5555_ _5555_/A VGND VGND VPWR VPWR _8874_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4506_ _4506_/A _4506_/B _4506_/C _4506_/D VGND VGND VPWR VPWR _4507_/B sky130_fd_sc_hd__or4_1
X_8274_ _9088_/Q _7940_/X _7997_/X _8957_/Q _8273_/X VGND VGND VPWR VPWR _8282_/A
+ sky130_fd_sc_hd__a221o_1
X_5486_ _5465_/X hold613/X _5490_/S VGND VGND VPWR VPWR _5486_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7225_ _7225_/A VGND VGND VPWR VPWR _9206_/D sky130_fd_sc_hd__clkbuf_1
X_4437_ _7111_/A _4675_/B VGND VGND VPWR VPWR _4437_/Y sky130_fd_sc_hd__nor2_4
XFILLER_144_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout502 fanout503/X VGND VGND VPWR VPWR _5929_/B sky130_fd_sc_hd__clkbuf_4
X_7156_ _5465_/X _9175_/Q _7156_/S VGND VGND VPWR VPWR _7156_/X sky130_fd_sc_hd__mux2_1
X_4368_ hold40/X hold363/X hold73/X VGND VGND VPWR VPWR hold41/A sky130_fd_sc_hd__mux2_4
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6107_ _6107_/A VGND VGND VPWR VPWR _6779_/A sky130_fd_sc_hd__buf_4
XFILLER_59_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7087_ _5951_/X _9145_/Q _7089_/S VGND VGND VPWR VPWR _7087_/X sky130_fd_sc_hd__mux2_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6038_ _6038_/A VGND VGND VPWR VPWR _9086_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7989_ _8275_/B _7989_/B _8000_/B VGND VGND VPWR VPWR _7990_/A sky130_fd_sc_hd__and3_2
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_64_csclk _9090_/CLK VGND VGND VPWR VPWR _8852_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_157_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_79_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _9480_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_173_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_17_csclk _9303_/CLK VGND VGND VPWR VPWR _9420_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5340_ _5340_/A VGND VGND VPWR VPWR _5340_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5271_ _5271_/A _5287_/B VGND VGND VPWR VPWR _5272_/A sky130_fd_sc_hd__and2_1
XFILLER_99_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7010_ _7010_/A VGND VGND VPWR VPWR _9110_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8961_ _9162_/CLK _8961_/D fanout441/X VGND VGND VPWR VPWR _8961_/Q sky130_fd_sc_hd__dfrtp_4
X_7912_ _9488_/Q _9489_/Q _9490_/Q _9491_/Q VGND VGND VPWR VPWR _7912_/X sky130_fd_sc_hd__a211o_1
X_8892_ _9051_/CLK _8892_/D fanout444/X VGND VGND VPWR VPWR _8892_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_64_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7843_ _5465_/A hold275/X _7847_/S VGND VGND VPWR VPWR _7843_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7774_ _7774_/A VGND VGND VPWR VPWR _9452_/D sky130_fd_sc_hd__clkbuf_1
X_4986_ hold55/A hold80/A _4997_/B hold29/A VGND VGND VPWR VPWR _4986_/X sky130_fd_sc_hd__a31o_1
X_9513_ _9531_/CLK _9513_/D fanout452/X VGND VGND VPWR VPWR _9513_/Q sky130_fd_sc_hd__dfrtp_1
X_6725_ _6725_/A _6725_/B VGND VGND VPWR VPWR _6726_/C sky130_fd_sc_hd__nor2_1
XFILLER_149_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9444_ _9484_/CLK _9444_/D fanout429/X VGND VGND VPWR VPWR _9444_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_137_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6656_ _6887_/A _6528_/B _6918_/A VGND VGND VPWR VPWR _6657_/D sky130_fd_sc_hd__o21ai_1
XFILLER_192_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5607_ _5607_/A _5693_/B VGND VGND VPWR VPWR _5616_/S sky130_fd_sc_hd__nand2_2
XFILLER_176_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9375_ _9461_/CLK _9375_/D fanout423/X VGND VGND VPWR VPWR _9375_/Q sky130_fd_sc_hd__dfrtp_2
X_6587_ _6876_/B _6732_/B VGND VGND VPWR VPWR _6627_/A sky130_fd_sc_hd__nor2_1
XFILLER_191_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8326_ _8342_/B _8357_/A _8357_/B VGND VGND VPWR VPWR _8364_/A sky130_fd_sc_hd__and3_2
X_5538_ _5315_/X _5538_/A1 _5538_/S VGND VGND VPWR VPWR _5538_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8257_ _8861_/Q _7927_/X _7990_/X _8871_/Q _8256_/X VGND VGND VPWR VPWR _8260_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_117_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5469_ _5468_/X hold821/X _5472_/S VGND VGND VPWR VPWR _5469_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7208_ _7208_/A VGND VGND VPWR VPWR _9198_/D sky130_fd_sc_hd__clkbuf_1
X_8188_ _9074_/Q _8034_/X _8185_/X _8187_/X VGND VGND VPWR VPWR _8193_/B sky130_fd_sc_hd__a211o_1
X_7139_ _7139_/A _7139_/B VGND VGND VPWR VPWR _7142_/S sky130_fd_sc_hd__nand2_1
XFILLER_101_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput18 mask_rev_in[22] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__buf_2
Xinput29 mask_rev_in[3] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__clkbuf_2
XFILLER_168_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4840_ input72/X _4436_/A _5667_/A _8924_/Q _4839_/X VGND VGND VPWR VPWR _4841_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_270 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_281 _5281_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_292 _9124_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4771_ _9258_/Q _7339_/A _7144_/A _5279_/A _4770_/X VGND VGND VPWR VPWR _4772_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_60_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6510_ _6510_/A _6973_/B VGND VGND VPWR VPWR _6510_/Y sky130_fd_sc_hd__nand2_2
XFILLER_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7490_ _7436_/X hold303/X _7497_/S VGND VGND VPWR VPWR _7490_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6441_ _6597_/B _6441_/B VGND VGND VPWR VPWR _6926_/A sky130_fd_sc_hd__nand2_2
XFILLER_146_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9160_ _9161_/CLK _9160_/D fanout442/X VGND VGND VPWR VPWR _9160_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_174_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6372_ _6628_/A _6440_/A VGND VGND VPWR VPWR _6373_/A sky130_fd_sc_hd__or2_1
X_8111_ _9285_/Q _7953_/B _7981_/X _9333_/Q VGND VGND VPWR VPWR _8111_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5323_ _5323_/A VGND VGND VPWR VPWR _5323_/X sky130_fd_sc_hd__clkbuf_1
X_9091_ _9091_/CLK _9091_/D fanout455/X VGND VGND VPWR VPWR _9091_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_142_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8042_ _9378_/Q _7947_/A _7981_/A _9330_/Q VGND VGND VPWR VPWR _8042_/X sky130_fd_sc_hd__a22o_1
X_5254_ _9331_/Q VGND VGND VPWR VPWR _5254_/Y sky130_fd_sc_hd__inv_2
X_5185_ _9395_/Q VGND VGND VPWR VPWR _5185_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_3_6_0_csclk clkbuf_3_7_0_csclk/A VGND VGND VPWR VPWR _8954_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8944_ _9243_/CLK _8944_/D fanout469/X VGND VGND VPWR VPWR _8944_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_71_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8875_ _9251_/CLK _8875_/D fanout485/X VGND VGND VPWR VPWR _8875_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_36_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7826_ _7654_/X hold256/X _7830_/S VGND VGND VPWR VPWR _7826_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7757_ _7757_/A VGND VGND VPWR VPWR _9444_/D sky130_fd_sc_hd__clkbuf_1
X_4969_ _4969_/A _4971_/A VGND VGND VPWR VPWR _8808_/D sky130_fd_sc_hd__xor2_1
XFILLER_11_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6708_ _6708_/A _6708_/B VGND VGND VPWR VPWR _6709_/D sky130_fd_sc_hd__or2_1
XFILLER_165_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7688_ _7688_/A VGND VGND VPWR VPWR _9412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9427_ _9427_/CLK _9427_/D fanout478/X VGND VGND VPWR VPWR _9427_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6639_ _6894_/B _6781_/B _6917_/B VGND VGND VPWR VPWR _6977_/B sky130_fd_sc_hd__o21ai_1
XFILLER_192_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9358_ _9367_/CLK _9358_/D fanout422/X VGND VGND VPWR VPWR _9358_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8309_ _8355_/A _8368_/B VGND VGND VPWR VPWR _8360_/A sky130_fd_sc_hd__nor2_8
XFILLER_133_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9289_ _9305_/CLK _9289_/D fanout468/X VGND VGND VPWR VPWR _9289_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6990_ _6982_/X _7007_/B _7008_/A VGND VGND VPWR VPWR _6990_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_53_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5941_ _9045_/Q _4591_/X _5945_/S VGND VGND VPWR VPWR _5942_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5872_ _9030_/Q _6543_/B VGND VGND VPWR VPWR _5873_/A sky130_fd_sc_hd__or2_1
X_8660_ _8921_/Q _8310_/X _8381_/X _8956_/Q _8659_/X VGND VGND VPWR VPWR _8663_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4823_ _9127_/Q _7043_/A _5996_/A _9070_/Q VGND VGND VPWR VPWR _4823_/X sky130_fd_sc_hd__a22o_1
X_7611_ hold715/X _6048_/X _7621_/S VGND VGND VPWR VPWR _7612_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8591_ _8908_/Q _8348_/X _8411_/X _8923_/Q _8590_/X VGND VGND VPWR VPWR _8601_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_166_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7542_ _7542_/A VGND VGND VPWR VPWR _9346_/D sky130_fd_sc_hd__clkbuf_1
X_4754_ _4753_/X hold956/X _4964_/B VGND VGND VPWR VPWR _4754_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7473_ hold334/X _5690_/A _7479_/S VGND VGND VPWR VPWR _7473_/X sky130_fd_sc_hd__mux2_1
X_4685_ hold33/X _4685_/B VGND VGND VPWR VPWR _6055_/A sky130_fd_sc_hd__nor2_8
X_9212_ _9462_/CLK _9212_/D fanout408/X VGND VGND VPWR VPWR _9212_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_162_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6424_ _6518_/A VGND VGND VPWR VPWR _6887_/B sky130_fd_sc_hd__buf_2
XFILLER_146_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9143_ _9162_/CLK _9143_/D fanout437/X VGND VGND VPWR VPWR _9143_/Q sky130_fd_sc_hd__dfrtp_4
X_6355_ _7002_/B _6573_/B _6355_/C _6355_/D VGND VGND VPWR VPWR _6355_/X sky130_fd_sc_hd__or4_1
XFILLER_103_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5306_ _7645_/A VGND VGND VPWR VPWR _5306_/X sky130_fd_sc_hd__clkbuf_8
X_9074_ _9484_/CLK _9074_/D fanout428/X VGND VGND VPWR VPWR _9074_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_130_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6286_ _6973_/A _6399_/A VGND VGND VPWR VPWR _6596_/B sky130_fd_sc_hd__nand2_4
XFILLER_130_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8025_ _9377_/Q _7947_/X _7977_/X _9393_/Q VGND VGND VPWR VPWR _8025_/X sky130_fd_sc_hd__a22o_1
X_5237_ _5413_/S _5237_/A2 _5334_/B _5236_/Y VGND VGND VPWR VPWR _5237_/X sky130_fd_sc_hd__a22o_2
XFILLER_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5168_ input83/X _5168_/A1 _8794_/Q VGND VGND VPWR VPWR _5169_/A sky130_fd_sc_hd__mux2_2
XFILLER_29_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5099_ _9307_/Q VGND VGND VPWR VPWR _5099_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8927_ _9467_/CLK _8927_/D fanout475/X VGND VGND VPWR VPWR _8927_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_71_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8858_ _9069_/CLK _8858_/D fanout434/X VGND VGND VPWR VPWR _8858_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7809_ _7654_/X hold220/X _7813_/S VGND VGND VPWR VPWR _7809_/X sky130_fd_sc_hd__mux2_1
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8789_ _8831_/CLK _8789_/D _5344_/X VGND VGND VPWR VPWR _8789_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_12_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold7 hold7/A VGND VGND VPWR VPWR hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4470_ _4470_/A VGND VGND VPWR VPWR _4891_/B sky130_fd_sc_hd__buf_6
Xhold407 _8966_/Q VGND VGND VPWR VPWR hold407/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire382 _4428_/Y VGND VGND VPWR VPWR _7284_/A sky130_fd_sc_hd__buf_8
Xwire393 _8474_/A VGND VGND VPWR VPWR _8650_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold418 hold418/A VGND VGND VPWR VPWR hold418/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold429 _7364_/X VGND VGND VPWR VPWR _7365_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6140_ _6724_/A _6724_/B VGND VGND VPWR VPWR _6623_/A sky130_fd_sc_hd__or2b_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ hold512/X _6048_/X _6075_/S VGND VGND VPWR VPWR _6071_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5022_ hold949/X _5019_/Y _5021_/X _8796_/Q VGND VGND VPWR VPWR _8796_/D sky130_fd_sc_hd__a31o_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1107 _7473_/X VGND VGND VPWR VPWR _7474_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1118 _9252_/Q VGND VGND VPWR VPWR hold309/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1129 _5856_/X VGND VGND VPWR VPWR hold211/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6973_ _6973_/A _6973_/B _6973_/C VGND VGND VPWR VPWR _6973_/X sky130_fd_sc_hd__or3_1
XFILLER_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8712_ _8712_/A VGND VGND VPWR VPWR _9534_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5924_ _5924_/A VGND VGND VPWR VPWR _9037_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8643_ _8985_/Q _8292_/A _8358_/A _8880_/Q VGND VGND VPWR VPWR _8643_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5855_ _8843_/Q _7648_/A _5867_/S VGND VGND VPWR VPWR _5855_/X sky130_fd_sc_hd__mux2_1
X_4806_ _4806_/A _4806_/B _4806_/C _4806_/D VGND VGND VPWR VPWR _4817_/C sky130_fd_sc_hd__or4_1
XFILLER_166_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8574_ _9215_/Q _8289_/X _8341_/X _9311_/Q _8573_/X VGND VGND VPWR VPWR _8575_/D
+ sky130_fd_sc_hd__a221o_1
X_5786_ _5786_/A VGND VGND VPWR VPWR _8973_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7525_ _7525_/A VGND VGND VPWR VPWR _9338_/D sky130_fd_sc_hd__clkbuf_1
X_4737_ _9443_/Q _7746_/A _5551_/A _8876_/Q VGND VGND VPWR VPWR _4737_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4668_ _9083_/Q _6021_/A _5996_/A _9073_/Q VGND VGND VPWR VPWR _4668_/X sky130_fd_sc_hd__a22o_1
X_7456_ _7456_/A VGND VGND VPWR VPWR _9308_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6407_ _6895_/A _6651_/A VGND VGND VPWR VPWR _6948_/A sky130_fd_sc_hd__nor2_1
Xhold930 hold930/A VGND VGND VPWR VPWR hold930/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4599_ input24/X _4460_/Y _4458_/Y _9268_/Q VGND VGND VPWR VPWR _4599_/X sky130_fd_sc_hd__a22o_1
Xhold941 hold941/A VGND VGND VPWR VPWR hold941/X sky130_fd_sc_hd__dlygate4sd3_1
X_7387_ _7279_/X hold750/X _7389_/S VGND VGND VPWR VPWR _7387_/X sky130_fd_sc_hd__mux2_1
Xhold952 _5028_/X VGND VGND VPWR VPWR _8794_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold963 _9117_/Q VGND VGND VPWR VPWR hold963/X sky130_fd_sc_hd__dlygate4sd3_1
X_9126_ _9485_/CLK _9126_/D fanout405/X VGND VGND VPWR VPWR _9126_/Q sky130_fd_sc_hd__dfrtp_4
Xhold974 _9510_/Q VGND VGND VPWR VPWR hold974/X sky130_fd_sc_hd__dlygate4sd3_1
X_6338_ _6338_/A _6764_/A VGND VGND VPWR VPWR _6354_/B sky130_fd_sc_hd__nor2_1
Xhold985 _9518_/Q VGND VGND VPWR VPWR hold985/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 _9025_/Q VGND VGND VPWR VPWR _8705_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6269_ _6279_/A _6871_/B VGND VGND VPWR VPWR _6853_/A sky130_fd_sc_hd__nor2_1
X_9057_ _9110_/CLK _9057_/D VGND VGND VPWR VPWR _9057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8008_ _8275_/B _8008_/B VGND VGND VPWR VPWR _8009_/A sky130_fd_sc_hd__nand2_2
Xclkbuf_2_3_0_csclk clkbuf_2_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_7_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_151_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5640_ _5315_/X hold328/X _5640_/S VGND VGND VPWR VPWR _5640_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5571_ hold664/X _5402_/X _5571_/S VGND VGND VPWR VPWR _5572_/A sky130_fd_sc_hd__mux2_1
X_7310_ _7310_/A VGND VGND VPWR VPWR _9242_/D sky130_fd_sc_hd__clkbuf_1
X_4522_ _9246_/Q _4449_/Y _4436_/A input41/X VGND VGND VPWR VPWR _4522_/X sky130_fd_sc_hd__a22o_1
X_8290_ _9499_/Q _9500_/Q VGND VGND VPWR VPWR _8357_/B sky130_fd_sc_hd__and2b_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold204 hold204/A VGND VGND VPWR VPWR hold204/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold215 _7220_/X VGND VGND VPWR VPWR _7221_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7241_ _7241_/A VGND VGND VPWR VPWR _9212_/D sky130_fd_sc_hd__clkbuf_1
X_4453_ _4492_/B VGND VGND VPWR VPWR _4667_/A sky130_fd_sc_hd__buf_12
XFILLER_7_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold226 _7672_/X VGND VGND VPWR VPWR _7673_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold237 _7547_/X VGND VGND VPWR VPWR _7548_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold248 _9365_/Q VGND VGND VPWR VPWR hold248/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold259 hold259/A VGND VGND VPWR VPWR hold259/X sky130_fd_sc_hd__dlygate4sd3_1
X_7172_ _5468_/X hold681/X _7174_/S VGND VGND VPWR VPWR _7172_/X sky130_fd_sc_hd__mux2_1
X_4384_ hold63/X hold41/X VGND VGND VPWR VPWR _4555_/A sky130_fd_sc_hd__nor2_8
XFILLER_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6123_ _6891_/B VGND VGND VPWR VPWR _6828_/B sky130_fd_sc_hd__inv_2
XFILLER_98_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _6054_/A VGND VGND VPWR VPWR _9093_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _5004_/X hold39/A _5014_/S VGND VGND VPWR VPWR _5006_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6956_ _6956_/A _6987_/C _6956_/C VGND VGND VPWR VPWR _6957_/C sky130_fd_sc_hd__or3_1
X_5907_ _5907_/A VGND VGND VPWR VPWR _5907_/X sky130_fd_sc_hd__clkbuf_1
X_6887_ _6887_/A _6887_/B VGND VGND VPWR VPWR _6887_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8626_ _8606_/X _8612_/X _8625_/X _8399_/A _8849_/Q VGND VGND VPWR VPWR _8626_/X
+ sky130_fd_sc_hd__o32a_1
X_5838_ _5838_/A VGND VGND VPWR VPWR _5838_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8557_ _9375_/Q _8682_/B VGND VGND VPWR VPWR _8557_/X sky130_fd_sc_hd__and2_1
X_5769_ hold407/X _5687_/X _5771_/S VGND VGND VPWR VPWR _5770_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7508_ _7436_/X hold283/X _7515_/S VGND VGND VPWR VPWR _7508_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8488_ _9444_/Q _8398_/B _8344_/X _9484_/Q VGND VGND VPWR VPWR _8488_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7439_ hold15/X VGND VGND VPWR VPWR _7439_/X sky130_fd_sc_hd__buf_2
XFILLER_146_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold760 _7459_/X VGND VGND VPWR VPWR _7460_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_146_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold771 hold771/A VGND VGND VPWR VPWR hold771/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 hold782/A VGND VGND VPWR VPWR hold782/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9109_ _9110_/CLK _9109_/D fanout503/X VGND VGND VPWR VPWR _9109_/Q sky130_fd_sc_hd__dfrtp_4
Xhold793 hold793/A VGND VGND VPWR VPWR _7136_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput309 _5233_/X VGND VGND VPWR VPWR serial_load sky130_fd_sc_hd__buf_12
XFILLER_153_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6810_ _6948_/A _6925_/A _6948_/B VGND VGND VPWR VPWR _6824_/B sky130_fd_sc_hd__or3_1
XFILLER_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7790_ _7651_/X hold184/X _7796_/S VGND VGND VPWR VPWR _7790_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6741_ _6924_/C _6856_/B _6741_/C _6741_/D VGND VGND VPWR VPWR _6751_/B sky130_fd_sc_hd__or4_1
XFILLER_189_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9460_ _9476_/CLK _9460_/D fanout414/X VGND VGND VPWR VPWR _9460_/Q sky130_fd_sc_hd__dfrtp_4
X_6672_ _6716_/A _6672_/B _6672_/C VGND VGND VPWR VPWR _6835_/A sky130_fd_sc_hd__and3_1
XFILLER_149_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8411_ _8411_/A VGND VGND VPWR VPWR _8411_/X sky130_fd_sc_hd__buf_6
X_5623_ hold610/X _5395_/X _5627_/S VGND VGND VPWR VPWR _5624_/A sky130_fd_sc_hd__mux2_1
X_9391_ _9463_/CLK _9391_/D _5332_/A VGND VGND VPWR VPWR _9391_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8342_ _8352_/A _8342_/B VGND VGND VPWR VPWR _8377_/B sky130_fd_sc_hd__nand2_2
XFILLER_145_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5554_ _5301_/X hold594/X _5560_/S VGND VGND VPWR VPWR _5555_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4505_ _9191_/Q _7176_/A _5388_/A _8816_/Q _4504_/X VGND VGND VPWR VPWR _4506_/D
+ sky130_fd_sc_hd__a221o_1
X_8273_ _8962_/Q _8224_/B _7981_/X _8917_/Q VGND VGND VPWR VPWR _8273_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5485_ _5485_/A VGND VGND VPWR VPWR _8844_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7224_ _5468_/X hold683/X _7226_/S VGND VGND VPWR VPWR _7224_/X sky130_fd_sc_hd__mux2_1
X_4436_ _4436_/A VGND VGND VPWR VPWR _5867_/S sky130_fd_sc_hd__buf_8
XFILLER_104_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout503 input196/X VGND VGND VPWR VPWR fanout503/X sky130_fd_sc_hd__buf_4
X_7155_ _7155_/A VGND VGND VPWR VPWR _7155_/X sky130_fd_sc_hd__clkbuf_1
X_4367_ hold39/X hold8/X hold22/X VGND VGND VPWR VPWR hold40/A sky130_fd_sc_hd__mux2_1
XFILLER_86_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6106_ _6891_/B _6828_/A VGND VGND VPWR VPWR _6107_/A sky130_fd_sc_hd__or2_1
X_7086_ _7086_/A _7139_/B VGND VGND VPWR VPWR _7089_/S sky130_fd_sc_hd__nand2_1
XFILLER_86_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6037_ hold551/X _5683_/X _6041_/S VGND VGND VPWR VPWR _6037_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7988_ _7988_/A VGND VGND VPWR VPWR _7988_/X sky130_fd_sc_hd__buf_8
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6939_ _6939_/A _6939_/B _6939_/C _6939_/D VGND VGND VPWR VPWR _6939_/Y sky130_fd_sc_hd__nand4_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8609_ _8919_/Q _8310_/X _8381_/X _8954_/Q _8608_/X VGND VGND VPWR VPWR _8609_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_csclk _5237_/X VGND VGND VPWR VPWR clkbuf_0_csclk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_136_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold590 _7121_/X VGND VGND VPWR VPWR _9160_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_1_0_1_csclk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_18_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5270_ _8793_/Q hold18/A _7025_/B VGND VGND VPWR VPWR _5270_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_99_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8960_ _9088_/CLK _8960_/D fanout454/X VGND VGND VPWR VPWR _8960_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7911_ _8652_/S _7911_/B VGND VGND VPWR VPWR _8015_/A sky130_fd_sc_hd__nor2_1
X_8891_ _9051_/CLK _8891_/D fanout453/X VGND VGND VPWR VPWR _8891_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7842_ _7842_/A VGND VGND VPWR VPWR _9484_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7773_ _7651_/X hold192/X _7779_/S VGND VGND VPWR VPWR _7773_/X sky130_fd_sc_hd__mux2_1
X_4985_ hold944/X _5014_/S _4984_/Y VGND VGND VPWR VPWR _8805_/D sky130_fd_sc_hd__a21o_1
X_9512_ _9531_/CLK _9512_/D fanout451/X VGND VGND VPWR VPWR _9512_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6724_ _6724_/A _6724_/B _6967_/A VGND VGND VPWR VPWR _6725_/A sky130_fd_sc_hd__or3_2
Xclkbuf_3_2_0_csclk clkbuf_3_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_2_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
X_9443_ _9459_/CLK hold48/X fanout489/X VGND VGND VPWR VPWR _9443_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_176_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6655_ _6906_/B _6815_/B _6655_/C VGND VGND VPWR VPWR _6918_/A sky130_fd_sc_hd__or3_1
XFILLER_31_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5606_ _5606_/A VGND VGND VPWR VPWR _8897_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9374_ _9461_/CLK _9374_/D fanout423/X VGND VGND VPWR VPWR _9374_/Q sky130_fd_sc_hd__dfrtp_4
X_6586_ _6754_/B _6867_/A VGND VGND VPWR VPWR _6865_/A sky130_fd_sc_hd__or2_1
XFILLER_11_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8325_ _8342_/B _8389_/A _8398_/A VGND VGND VPWR VPWR _8402_/A sky130_fd_sc_hd__and3_4
XFILLER_191_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5537_ _5537_/A VGND VGND VPWR VPWR _8866_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8256_ _9092_/Q _7958_/X _8224_/B _8961_/Q VGND VGND VPWR VPWR _8256_/X sky130_fd_sc_hd__a22o_1
X_5468_ _7494_/A VGND VGND VPWR VPWR _5468_/X sky130_fd_sc_hd__buf_12
XFILLER_132_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7207_ _5468_/X hold676/X _7209_/S VGND VGND VPWR VPWR _7207_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4419_ _7111_/A _4674_/A VGND VGND VPWR VPWR _4419_/Y sky130_fd_sc_hd__nor2_1
X_8187_ _9079_/Q _7949_/A _7973_/A _8853_/Q _8186_/X VGND VGND VPWR VPWR _8187_/X
+ sky130_fd_sc_hd__a221o_1
X_5399_ _8812_/Q _5398_/X _5416_/S VGND VGND VPWR VPWR _5399_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7138_ _7138_/A VGND VGND VPWR VPWR _9167_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7069_ _7069_/A VGND VGND VPWR VPWR _9137_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput19 mask_rev_in[23] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_754 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_260 _5174_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_271 _9555_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_282 _5281_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_293 _9127_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4770_ _8895_/Q _5596_/A _6032_/A _9086_/Q VGND VGND VPWR VPWR _4770_/X sky130_fd_sc_hd__a22o_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6440_ _6440_/A _6891_/B VGND VGND VPWR VPWR _6441_/B sky130_fd_sc_hd__nor2_4
X_6371_ _6415_/A _6739_/A VGND VGND VPWR VPWR _6811_/C sky130_fd_sc_hd__nor2_2
XFILLER_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8110_ _9413_/Q _7967_/X _7993_/X _9389_/Q _8109_/X VGND VGND VPWR VPWR _8117_/A
+ sky130_fd_sc_hd__a221o_1
X_5322_ _5330_/A _5334_/B VGND VGND VPWR VPWR _5323_/A sky130_fd_sc_hd__and2_1
X_9090_ _9090_/CLK _9090_/D fanout454/X VGND VGND VPWR VPWR _9090_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8041_ hold947/X _8017_/X _8040_/X VGND VGND VPWR VPWR _8041_/X sky130_fd_sc_hd__o21a_1
X_5253_ _9323_/Q VGND VGND VPWR VPWR _5253_/Y sky130_fd_sc_hd__inv_2
X_5184_ _8829_/Q _5183_/Y _4964_/B VGND VGND VPWR VPWR _8779_/D sky130_fd_sc_hd__o21a_1
XFILLER_3_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_63_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _9184_/CLK sky130_fd_sc_hd__clkbuf_16
X_8943_ _9051_/CLK _8943_/D fanout444/X VGND VGND VPWR VPWR _8943_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_83_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8874_ _9251_/CLK _8874_/D fanout486/X VGND VGND VPWR VPWR _8874_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_24_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7825_ _7825_/A VGND VGND VPWR VPWR _9476_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_78_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _9476_/CLK sky130_fd_sc_hd__clkbuf_16
X_7756_ hold117/X _5690_/A _7762_/S VGND VGND VPWR VPWR _7756_/X sky130_fd_sc_hd__mux2_1
X_4968_ _8807_/Q _5068_/B _4972_/B VGND VGND VPWR VPWR _4971_/A sky130_fd_sc_hd__and3_1
XFILLER_11_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6707_ _6835_/A _6835_/B _6707_/C _6707_/D VGND VGND VPWR VPWR _6709_/C sky130_fd_sc_hd__or4_1
XFILLER_177_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7687_ _7651_/X hold372/X _7693_/S VGND VGND VPWR VPWR _7688_/A sky130_fd_sc_hd__mux2_1
X_4899_ _9424_/Q _4437_/Y _5715_/A _8943_/Q _4898_/X VGND VGND VPWR VPWR _4899_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_137_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9426_ _9467_/CLK _9426_/D fanout475/X VGND VGND VPWR VPWR _9426_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6638_ _6948_/A _6925_/A VGND VGND VPWR VPWR _6987_/C sky130_fd_sc_hd__or2_1
XFILLER_164_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9357_ _9421_/CLK _9357_/D fanout460/X VGND VGND VPWR VPWR _9357_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_180_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6569_ _6563_/A _6839_/B _6551_/Y _6345_/X _6568_/X VGND VGND VPWR VPWR _6576_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_164_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8308_ _8342_/B _8392_/C VGND VGND VPWR VPWR _8368_/B sky130_fd_sc_hd__nand2_4
XFILLER_180_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9288_ _9288_/CLK _9288_/D fanout425/X VGND VGND VPWR VPWR _9288_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_133_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_16_csclk _9303_/CLK VGND VGND VPWR VPWR _9468_/CLK sky130_fd_sc_hd__clkbuf_16
X_8239_ _8850_/Q _8010_/B _8228_/X _8238_/X _8105_/X VGND VGND VPWR VPWR _8239_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_160_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5940_ _5940_/A VGND VGND VPWR VPWR _9044_/D sky130_fd_sc_hd__buf_1
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5871_ _5871_/A _5871_/B _9034_/Q VGND VGND VPWR VPWR _6543_/B sky130_fd_sc_hd__or3_4
XFILLER_61_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7610_ _7610_/A VGND VGND VPWR VPWR _9377_/D sky130_fd_sc_hd__clkbuf_1
X_4822_ _9217_/Q _7249_/A _5618_/A _8904_/Q _4821_/X VGND VGND VPWR VPWR _4829_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8590_ _8858_/Q _8391_/X _8367_/X _9094_/Q _8589_/X VGND VGND VPWR VPWR _8590_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7541_ _7430_/X hold718/X _7551_/S VGND VGND VPWR VPWR _7542_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4753_ _9113_/Q _4752_/X _4886_/S VGND VGND VPWR VPWR _4753_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7472_ _7472_/A VGND VGND VPWR VPWR _9315_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4684_ hold33/X _4794_/B VGND VGND VPWR VPWR _5630_/A sky130_fd_sc_hd__nor2_8
X_9211_ _9227_/CLK _9211_/D fanout467/X VGND VGND VPWR VPWR _9211_/Q sky130_fd_sc_hd__dfrtp_4
X_6423_ _6900_/A _6772_/A VGND VGND VPWR VPWR _6433_/C sky130_fd_sc_hd__nor2_1
XFILLER_134_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9142_ _9161_/CLK _9142_/D fanout440/X VGND VGND VPWR VPWR _9142_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6354_ _6882_/B _6354_/B _6759_/A _6354_/D VGND VGND VPWR VPWR _6355_/D sky130_fd_sc_hd__or4_1
XFILLER_161_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5305_ hold12/X VGND VGND VPWR VPWR _7645_/A sky130_fd_sc_hd__buf_6
X_9073_ _9482_/CLK _9073_/D fanout433/X VGND VGND VPWR VPWR _9073_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_130_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6285_ _6628_/B _6420_/B VGND VGND VPWR VPWR _6597_/A sky130_fd_sc_hd__nor2_8
X_8024_ _9369_/Q _7960_/X _7973_/X _9193_/Q _8023_/X VGND VGND VPWR VPWR _8027_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5236_ _5413_/S _5236_/B VGND VGND VPWR VPWR _5236_/Y sky130_fd_sc_hd__nor2_2
XFILLER_124_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5167_ _8795_/Q _5330_/A VGND VGND VPWR VPWR _5167_/Y sky130_fd_sc_hd__nor2_2
XFILLER_84_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5098_ _9315_/Q VGND VGND VPWR VPWR _5098_/Y sky130_fd_sc_hd__inv_2
X_8926_ _9005_/CLK _8926_/D fanout489/X VGND VGND VPWR VPWR _8926_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_56_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8857_ _9184_/CLK _8857_/D fanout443/X VGND VGND VPWR VPWR _8857_/Q sky130_fd_sc_hd__dfstp_2
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7808_ _7808_/A VGND VGND VPWR VPWR _9468_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8788_ _5168_/A1 _8788_/D _5342_/X VGND VGND VPWR VPWR _8788_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_24_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7739_ _7739_/A VGND VGND VPWR VPWR _9436_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9409_ _9459_/CLK _9409_/D fanout480/X VGND VGND VPWR VPWR hold96/A sky130_fd_sc_hd__dfstp_4
XFILLER_138_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold8 hold8/A VGND VGND VPWR VPWR hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_47_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold408 _9386_/Q VGND VGND VPWR VPWR hold408/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold419 _8851_/Q VGND VGND VPWR VPWR hold419/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_109_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _6070_/A VGND VGND VPWR VPWR _9100_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _5021_/A _5021_/B _5040_/C VGND VGND VPWR VPWR _5021_/X sky130_fd_sc_hd__and3_1
Xhold1108 _8931_/Q VGND VGND VPWR VPWR hold405/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1119 _7331_/X VGND VGND VPWR VPWR _7332_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6972_ _6972_/A _6972_/B _6972_/C VGND VGND VPWR VPWR _6972_/X sky130_fd_sc_hd__or3_1
XFILLER_53_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8711_ _9534_/Q _4961_/X _8725_/S VGND VGND VPWR VPWR _8712_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5923_ _5647_/X hold812/X _5927_/S VGND VGND VPWR VPWR _5923_/X sky130_fd_sc_hd__mux2_1
X_8642_ _9076_/Q _8356_/B _8364_/B _8865_/Q _8641_/X VGND VGND VPWR VPWR _8649_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5854_ _5854_/A VGND VGND VPWR VPWR _9002_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4805_ _9159_/Q _7113_/A _5948_/A _9050_/Q _4804_/X VGND VGND VPWR VPWR _4806_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_167_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8573_ _9399_/Q _8304_/X _8324_/X _9247_/Q VGND VGND VPWR VPWR _8573_/X sky130_fd_sc_hd__a22o_1
X_5785_ hold915/X _5761_/X _5793_/S VGND VGND VPWR VPWR _5786_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7524_ _7430_/X hold713/X _7534_/S VGND VGND VPWR VPWR _7525_/A sky130_fd_sc_hd__mux2_1
X_4736_ _9299_/Q _7425_/A _4734_/Y _4736_/B2 _4735_/X VGND VGND VPWR VPWR _4741_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_159_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7455_ _7436_/X hold326/X _7461_/S VGND VGND VPWR VPWR _7456_/A sky130_fd_sc_hd__mux2_1
X_4667_ _4667_/A _4667_/B VGND VGND VPWR VPWR _5996_/A sky130_fd_sc_hd__nor2_4
X_6406_ _6406_/A VGND VGND VPWR VPWR _6651_/A sky130_fd_sc_hd__clkbuf_2
Xhold920 _9240_/Q VGND VGND VPWR VPWR hold920/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_134_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold931 _9368_/Q VGND VGND VPWR VPWR hold931/X sky130_fd_sc_hd__dlygate4sd3_1
X_7386_ _7386_/A VGND VGND VPWR VPWR _9277_/D sky130_fd_sc_hd__clkbuf_1
X_4598_ _9348_/Q _4478_/Y _7056_/A _9136_/Q _4597_/X VGND VGND VPWR VPWR _4598_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold942 _9026_/Q VGND VGND VPWR VPWR _9031_/D sky130_fd_sc_hd__dlygate4sd3_1
X_9125_ _9485_/CLK _9125_/D fanout405/X VGND VGND VPWR VPWR _9125_/Q sky130_fd_sc_hd__dfrtp_2
Xhold953 _9507_/Q VGND VGND VPWR VPWR hold953/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold964 _4551_/X VGND VGND VPWR VPWR _4552_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6337_ _6341_/A _6338_/A VGND VGND VPWR VPWR _6882_/B sky130_fd_sc_hd__nor2_1
Xhold975 _8085_/X VGND VGND VPWR VPWR _9510_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 _8263_/X VGND VGND VPWR VPWR _9518_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 _9512_/Q VGND VGND VPWR VPWR hold997/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9056_ _9110_/CLK _9056_/D VGND VGND VPWR VPWR _9056_/Q sky130_fd_sc_hd__dfxtp_1
X_6268_ _6268_/A _6851_/A _6268_/C _6268_/D VGND VGND VPWR VPWR _6268_/X sky130_fd_sc_hd__or4_1
X_8007_ _8007_/A _8007_/B VGND VGND VPWR VPWR _8007_/X sky130_fd_sc_hd__or2_1
X_5219_ _9187_/Q VGND VGND VPWR VPWR _5219_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6199_ _6199_/A VGND VGND VPWR VPWR _6800_/A sky130_fd_sc_hd__buf_2
XFILLER_28_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8909_ _8955_/CLK _8909_/D fanout469/X VGND VGND VPWR VPWR _8909_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_44_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5570_ _5570_/A VGND VGND VPWR VPWR _8881_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4521_ _4521_/A _4521_/B _4521_/C _4521_/D VGND VGND VPWR VPWR _4549_/A sky130_fd_sc_hd__or4_1
XFILLER_144_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold205 _9191_/Q VGND VGND VPWR VPWR hold205/X sky130_fd_sc_hd__dlygate4sd3_1
X_7240_ _7239_/X hold286/X _7247_/S VGND VGND VPWR VPWR _7240_/X sky130_fd_sc_hd__mux2_1
X_4452_ _9471_/Q _7798_/A _7374_/A _9279_/Q _4451_/X VGND VGND VPWR VPWR _4463_/B
+ sky130_fd_sc_hd__a221o_1
Xhold216 _9269_/Q VGND VGND VPWR VPWR hold216/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold227 hold227/A VGND VGND VPWR VPWR hold227/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold238 _9341_/Q VGND VGND VPWR VPWR hold238/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold249 _7582_/X VGND VGND VPWR VPWR _7583_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7171_ _7171_/A VGND VGND VPWR VPWR _9181_/D sky130_fd_sc_hd__clkbuf_1
X_4383_ _4468_/B hold10/X VGND VGND VPWR VPWR _4418_/A sky130_fd_sc_hd__nor2b_4
XFILLER_131_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6122_ _6248_/A _6794_/A VGND VGND VPWR VPWR _6498_/B sky130_fd_sc_hd__and2_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ hold337/X _5690_/A _6053_/S VGND VGND VPWR VPWR _6053_/X sky130_fd_sc_hd__mux2_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5004_ hold8/A _5040_/B _5002_/Y _5003_/X VGND VGND VPWR VPWR _5004_/X sky130_fd_sc_hd__a22o_1
XFILLER_38_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6955_ _6955_/A _6955_/B _6955_/C _6955_/D VGND VGND VPWR VPWR _6957_/B sky130_fd_sc_hd__or4_1
XFILLER_53_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5906_ _5647_/X _9580_/A _5916_/S VGND VGND VPWR VPWR _5906_/X sky130_fd_sc_hd__mux2_1
X_6886_ _7000_/A _6935_/C _6886_/C _6886_/D VGND VGND VPWR VPWR _6886_/X sky130_fd_sc_hd__or4_1
XFILLER_179_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8625_ _8650_/A _8625_/B _8625_/C VGND VGND VPWR VPWR _8625_/X sky130_fd_sc_hd__or3_1
X_5837_ _9575_/A _5836_/X hold43/X VGND VGND VPWR VPWR _5837_/X sky130_fd_sc_hd__mux2_1
XFILLER_167_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8556_ _9423_/Q _8402_/X _8378_/A _9359_/Q _8555_/X VGND VGND VPWR VPWR _8563_/A
+ sky130_fd_sc_hd__a221o_1
X_5768_ _5768_/A VGND VGND VPWR VPWR _8965_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7507_ _7507_/A VGND VGND VPWR VPWR _9331_/D sky130_fd_sc_hd__clkbuf_1
X_4719_ _9087_/Q _6032_/A _6007_/A _9077_/Q VGND VGND VPWR VPWR _4719_/X sky130_fd_sc_hd__a22o_1
X_8487_ _8487_/A _8487_/B _8487_/C _8487_/D VGND VGND VPWR VPWR _8487_/X sky130_fd_sc_hd__or4_4
X_5699_ _5699_/A VGND VGND VPWR VPWR _8935_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7438_ _7438_/A VGND VGND VPWR VPWR _9300_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold750 _9278_/Q VGND VGND VPWR VPWR hold750/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7369_ _7369_/A VGND VGND VPWR VPWR _9269_/D sky130_fd_sc_hd__clkbuf_1
Xhold761 _5435_/X VGND VGND VPWR VPWR _5436_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold772 _9334_/Q VGND VGND VPWR VPWR hold772/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 _7046_/X VGND VGND VPWR VPWR _7047_/A sky130_fd_sc_hd__dlygate4sd3_1
X_9108_ _9110_/CLK _9108_/D fanout503/X VGND VGND VPWR VPWR _9108_/Q sky130_fd_sc_hd__dfrtp_4
Xhold794 _9222_/Q VGND VGND VPWR VPWR hold794/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9039_ _9187_/CLK _9039_/D fanout450/X VGND VGND VPWR VPWR _9039_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_39_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6740_ _6739_/Y _6721_/X _6732_/Y _6469_/B VGND VGND VPWR VPWR _6741_/D sky130_fd_sc_hd__a31o_1
XFILLER_189_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6671_ _6925_/B _6836_/A VGND VGND VPWR VPWR _6709_/B sky130_fd_sc_hd__or2_1
XFILLER_31_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8410_ hold96/A _8506_/B _8405_/X _8407_/X _8409_/X VGND VGND VPWR VPWR _8410_/X
+ sky130_fd_sc_hd__a2111o_2
X_5622_ _5622_/A VGND VGND VPWR VPWR _8904_/D sky130_fd_sc_hd__clkbuf_1
X_9390_ _9398_/CLK _9390_/D _5332_/A VGND VGND VPWR VPWR _9390_/Q sky130_fd_sc_hd__dfrtp_2
X_8341_ _8360_/B VGND VGND VPWR VPWR _8341_/X sky130_fd_sc_hd__buf_6
XFILLER_129_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5553_ _5553_/A VGND VGND VPWR VPWR _8873_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4504_ _9255_/Q _7321_/A _4500_/Y input19/X _4503_/X VGND VGND VPWR VPWR _4504_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_144_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8272_ _8272_/A _8272_/B _8272_/C _8272_/D VGND VGND VPWR VPWR _8272_/X sky130_fd_sc_hd__or4_1
X_5484_ _5315_/X hold137/X _5490_/S VGND VGND VPWR VPWR _5484_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7223_ _7223_/A VGND VGND VPWR VPWR _9205_/D sky130_fd_sc_hd__clkbuf_1
X_4435_ _7158_/A _5474_/B VGND VGND VPWR VPWR _4436_/A sky130_fd_sc_hd__nor2_8
XFILLER_172_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7154_ _6018_/X _9174_/Q _7156_/S VGND VGND VPWR VPWR _7154_/X sky130_fd_sc_hd__mux2_1
X_4366_ _4365_/X hold62/X hold74/A VGND VGND VPWR VPWR hold63/A sky130_fd_sc_hd__mux2_4
XFILLER_86_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6105_ _6891_/A _6317_/A VGND VGND VPWR VPWR _6828_/A sky130_fd_sc_hd__nand2_8
X_7085_ hold66/X VGND VGND VPWR VPWR _9144_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _6036_/A VGND VGND VPWR VPWR _9085_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7987_ _9496_/Q _7989_/B _8002_/C VGND VGND VPWR VPWR _7988_/A sky130_fd_sc_hd__and3_2
XFILLER_42_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6938_ _6956_/A _6987_/C _6956_/C _7003_/B VGND VGND VPWR VPWR _6941_/B sky130_fd_sc_hd__or4_1
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6869_ _6869_/A _6869_/B _6869_/C _6869_/D VGND VGND VPWR VPWR _6870_/B sky130_fd_sc_hd__or4_1
XFILLER_22_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8608_ _8914_/Q _8298_/A _8370_/A _9085_/Q VGND VGND VPWR VPWR _8608_/X sky130_fd_sc_hd__a22o_1
X_9588_ _9588_/A _5080_/Y VGND VGND VPWR VPWR mgmt_gpio_out[34] sky130_fd_sc_hd__ebufn_8
XFILLER_22_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8539_ _9222_/Q _8391_/X _8367_/X _9478_/Q _8538_/X VGND VGND VPWR VPWR _8539_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_157_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold580 _5954_/X VGND VGND VPWR VPWR _5955_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 hold591/A VGND VGND VPWR VPWR _7119_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1280 _9314_/Q VGND VGND VPWR VPWR hold566/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7910_ _7902_/B _7908_/X _7909_/Y _7910_/B2 VGND VGND VPWR VPWR _9502_/D sky130_fd_sc_hd__a22o_1
X_8890_ _9051_/CLK _8890_/D fanout451/X VGND VGND VPWR VPWR _8890_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7841_ _5402_/X hold573/X _7847_/S VGND VGND VPWR VPWR _7842_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7772_ _7772_/A VGND VGND VPWR VPWR _9451_/D sky130_fd_sc_hd__clkbuf_1
X_4984_ _5014_/S _4984_/B VGND VGND VPWR VPWR _4984_/Y sky130_fd_sc_hd__nor2_1
XFILLER_168_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9511_ _9531_/CLK _9511_/D fanout451/X VGND VGND VPWR VPWR _9511_/Q sky130_fd_sc_hd__dfrtp_1
X_6723_ _6853_/D _6944_/B _6993_/B VGND VGND VPWR VPWR _6752_/A sky130_fd_sc_hd__or3_1
X_9442_ _9442_/CLK _9442_/D fanout438/X VGND VGND VPWR VPWR _9442_/Q sky130_fd_sc_hd__dfrtp_1
X_6654_ _6922_/A _6530_/D VGND VGND VPWR VPWR _6915_/A sky130_fd_sc_hd__or2b_1
XFILLER_176_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5605_ hold620/X _5402_/X _5605_/S VGND VGND VPWR VPWR _5606_/A sky130_fd_sc_hd__mux2_1
X_9373_ _9469_/CLK _9373_/D fanout458/X VGND VGND VPWR VPWR _9373_/Q sky130_fd_sc_hd__dfrtp_4
X_6585_ _6585_/A _6585_/B VGND VGND VPWR VPWR _6714_/B sky130_fd_sc_hd__or2_1
XFILLER_118_721 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8324_ _8354_/C VGND VGND VPWR VPWR _8324_/X sky130_fd_sc_hd__buf_6
XFILLER_118_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5536_ _5311_/X hold422/X _5538_/S VGND VGND VPWR VPWR _5537_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8255_ _8981_/Q _7931_/X _8034_/X _9077_/Q _8254_/X VGND VGND VPWR VPWR _8260_/B
+ sky130_fd_sc_hd__a221o_1
X_5467_ _5467_/A VGND VGND VPWR VPWR _8837_/D sky130_fd_sc_hd__clkbuf_1
X_7206_ _7206_/A VGND VGND VPWR VPWR _9197_/D sky130_fd_sc_hd__clkbuf_1
X_4418_ _4418_/A hold42/X VGND VGND VPWR VPWR _7111_/A sky130_fd_sc_hd__nand2_8
X_8186_ _9089_/Q _7958_/A _7971_/A _8958_/Q VGND VGND VPWR VPWR _8186_/X sky130_fd_sc_hd__a22o_1
X_5398_ _7648_/A VGND VGND VPWR VPWR _5398_/X sky130_fd_sc_hd__buf_6
X_7137_ _9167_/Q _7126_/C _7137_/S VGND VGND VPWR VPWR _7137_/X sky130_fd_sc_hd__mux2_1
X_4349_ hold73/X VGND VGND VPWR VPWR hold74/A sky130_fd_sc_hd__buf_6
X_7068_ _9137_/Q _5465_/A _7072_/S VGND VGND VPWR VPWR _7068_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6019_ _6018_/X hold139/X _6019_/S VGND VGND VPWR VPWR _6019_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_250 wb_sel_i[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_261 _5174_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_272 _5279_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_283 input25/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_294 _4539_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6370_ _6510_/A VGND VGND VPWR VPWR _6811_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_161_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5321_ _5321_/A VGND VGND VPWR VPWR _5321_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_142_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8040_ _5130_/A _9507_/Q _8013_/A _8039_/X VGND VGND VPWR VPWR _8040_/X sky130_fd_sc_hd__a211o_1
XFILLER_130_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5252_ _9315_/Q VGND VGND VPWR VPWR _5252_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5183_ _8828_/Q _8831_/Q VGND VGND VPWR VPWR _5183_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8942_ _9482_/CLK _8942_/D fanout433/X VGND VGND VPWR VPWR _8942_/Q sky130_fd_sc_hd__dfrtp_2
X_8873_ _9465_/CLK _8873_/D fanout471/X VGND VGND VPWR VPWR _8873_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_36_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7824_ _7651_/X hold190/X _7830_/S VGND VGND VPWR VPWR _7824_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4967_ _8827_/Q _5040_/B _8829_/Q VGND VGND VPWR VPWR _4972_/B sky130_fd_sc_hd__or3_2
X_7755_ hold47/X VGND VGND VPWR VPWR hold48/A sky130_fd_sc_hd__clkbuf_1
XFILLER_149_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6706_ _6706_/A _6706_/B _6706_/C _6706_/D VGND VGND VPWR VPWR _6707_/D sky130_fd_sc_hd__or4_1
X_7686_ _7686_/A VGND VGND VPWR VPWR _9411_/D sky130_fd_sc_hd__clkbuf_1
X_4898_ _9480_/Q _4898_/A2 _5784_/A _8973_/Q VGND VGND VPWR VPWR _4898_/X sky130_fd_sc_hd__a22o_1
X_6637_ _6891_/A _6976_/B _6636_/Y VGND VGND VPWR VPWR _6646_/A sky130_fd_sc_hd__a21o_1
X_9425_ _9427_/CLK _9425_/D fanout476/X VGND VGND VPWR VPWR _9425_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_192_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9356_ _9468_/CLK _9356_/D fanout466/X VGND VGND VPWR VPWR _9356_/Q sky130_fd_sc_hd__dfrtp_4
X_6568_ _6568_/A _6822_/A _6960_/A _6567_/X VGND VGND VPWR VPWR _6568_/X sky130_fd_sc_hd__or4b_1
XFILLER_152_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5519_ _5291_/X hold891/X _5527_/S VGND VGND VPWR VPWR _5520_/A sky130_fd_sc_hd__mux2_1
X_8307_ _9208_/Q _8289_/X _8292_/X _9384_/Q _8306_/X VGND VGND VPWR VPWR _8397_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_105_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9287_ _9325_/CLK _9287_/D fanout464/X VGND VGND VPWR VPWR _9287_/Q sky130_fd_sc_hd__dfrtp_1
X_6499_ _6828_/B _6499_/B VGND VGND VPWR VPWR _6500_/A sky130_fd_sc_hd__or2_1
XFILLER_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8238_ _8238_/A _8238_/B _8238_/C _8238_/D VGND VGND VPWR VPWR _8238_/X sky130_fd_sc_hd__or4_2
XFILLER_160_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8169_ _9415_/Q _7967_/A _7999_/X _9431_/Q VGND VGND VPWR VPWR _8169_/X sky130_fd_sc_hd__a22o_1
XFILLER_87_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_727 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5870_ _9031_/D _5870_/B _5870_/C _5870_/D VGND VGND VPWR VPWR _5870_/X sky130_fd_sc_hd__or4_1
XFILLER_178_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4821_ _4821_/A1 _4488_/Y _5806_/A _8984_/Q VGND VGND VPWR VPWR _4821_/X sky130_fd_sc_hd__a22o_1
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7540_ _7540_/A VGND VGND VPWR VPWR _9345_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4752_ _4752_/A _4752_/B _4752_/C _4752_/D VGND VGND VPWR VPWR _4752_/X sky130_fd_sc_hd__or4_4
X_7471_ _9315_/Q hold46/X _7479_/S VGND VGND VPWR VPWR _7471_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4683_ _9396_/Q _7640_/A _7321_/A _9252_/Q _4682_/X VGND VGND VPWR VPWR _4688_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9210_ _9210_/CLK _9210_/D fanout467/X VGND VGND VPWR VPWR _9210_/Q sky130_fd_sc_hd__dfrtp_1
X_6422_ _6897_/B _6422_/B VGND VGND VPWR VPWR _6772_/A sky130_fd_sc_hd__nor2_2
XFILLER_147_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9141_ _9161_/CLK _9141_/D fanout440/X VGND VGND VPWR VPWR _9141_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_127_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6353_ _6340_/Y _6839_/A _6937_/A _6352_/X VGND VGND VPWR VPWR _6354_/D sky130_fd_sc_hd__a211o_1
XFILLER_161_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5304_ hold11/X hold557/X hold74/A VGND VGND VPWR VPWR _5304_/X sky130_fd_sc_hd__mux2_2
X_9072_ _9084_/CLK _9072_/D fanout445/X VGND VGND VPWR VPWR _9072_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_142_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6284_ _6588_/A _6950_/A _6708_/A _6283_/X VGND VGND VPWR VPWR _6290_/C sky130_fd_sc_hd__or4b_1
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8023_ _9305_/Q _8023_/B VGND VGND VPWR VPWR _8023_/X sky130_fd_sc_hd__and2_1
XFILLER_130_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5166_ _5166_/A VGND VGND VPWR VPWR _5166_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5097_ _9323_/Q VGND VGND VPWR VPWR _5097_/Y sky130_fd_sc_hd__inv_2
X_8925_ _9283_/CLK _8925_/D fanout489/X VGND VGND VPWR VPWR _8925_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_71_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8856_ _9084_/CLK _8856_/D fanout445/X VGND VGND VPWR VPWR _8856_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_25_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7807_ _7651_/X hold350/X _7813_/S VGND VGND VPWR VPWR _7808_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5999_ hold546/X _5809_/X _6005_/S VGND VGND VPWR VPWR _6000_/A sky130_fd_sc_hd__mux2_1
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8787_ _5207_/A1 _8787_/D _5340_/X VGND VGND VPWR VPWR hold4/A sky130_fd_sc_hd__dfrtp_1
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7738_ _7651_/X hold381/X hold86/X VGND VGND VPWR VPWR _7739_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7669_ _7669_/A VGND VGND VPWR VPWR _9403_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9408_ _9464_/CLK _9408_/D fanout420/X VGND VGND VPWR VPWR _9408_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_125_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9339_ _9475_/CLK _9339_/D fanout481/X VGND VGND VPWR VPWR _9339_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput290 _8825_/Q VGND VGND VPWR VPWR pll_trim[24] sky130_fd_sc_hd__buf_12
XFILLER_58_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold9 hold9/A VGND VGND VPWR VPWR hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_101_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_62_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _9442_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire373 _4485_/Y VGND VGND VPWR VPWR _7588_/A sky130_fd_sc_hd__buf_6
Xhold409 _7628_/X VGND VGND VPWR VPWR _7629_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_77_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _9452_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _8829_/Q VGND VGND VPWR VPWR _5040_/C sky130_fd_sc_hd__inv_2
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1109 _8983_/Q VGND VGND VPWR VPWR hold895/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6971_ _6462_/B _6812_/Y _6973_/C _6660_/A _6661_/B VGND VGND VPWR VPWR _6972_/C
+ sky130_fd_sc_hd__a221o_1
X_8710_ _8710_/A VGND VGND VPWR VPWR _8725_/S sky130_fd_sc_hd__buf_2
XFILLER_34_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5922_ _5922_/A VGND VGND VPWR VPWR _9036_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8641_ _8875_/Q _8358_/B _8364_/A _9091_/Q VGND VGND VPWR VPWR _8641_/X sky130_fd_sc_hd__a22o_1
X_5853_ _9002_/Q _5852_/X _5868_/S VGND VGND VPWR VPWR _5853_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4804_ _9101_/Q _6066_/A _5618_/A _8905_/Q VGND VGND VPWR VPWR _4804_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5784_ _5784_/A _7132_/B VGND VGND VPWR VPWR _5793_/S sky130_fd_sc_hd__and2_2
X_8572_ _9383_/Q _8337_/X _8384_/X _9199_/Q _8571_/X VGND VGND VPWR VPWR _8575_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4735_ _9072_/Q _5996_/A _5678_/A _8931_/Q VGND VGND VPWR VPWR _4735_/X sky130_fd_sc_hd__a22o_2
X_7523_ _7523_/A VGND VGND VPWR VPWR _9337_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7454_ _7454_/A VGND VGND VPWR VPWR _9307_/D sky130_fd_sc_hd__clkbuf_1
X_4666_ _5453_/B _4667_/A VGND VGND VPWR VPWR _6021_/A sky130_fd_sc_hd__nor2_8
XFILLER_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6405_ _6906_/C _6524_/B VGND VGND VPWR VPWR _6406_/A sky130_fd_sc_hd__or2_1
Xhold910 _7110_/X VGND VGND VPWR VPWR _9155_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7385_ _7242_/X hold273/X _7389_/S VGND VGND VPWR VPWR _7385_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4597_ _9236_/Q _7284_/A _6043_/A _9093_/Q VGND VGND VPWR VPWR _4597_/X sky130_fd_sc_hd__a22o_1
Xhold921 _9464_/Q VGND VGND VPWR VPWR hold921/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold932 hold932/A VGND VGND VPWR VPWR hold932/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 _9111_/Q VGND VGND VPWR VPWR hold943/X sky130_fd_sc_hd__dlygate4sd3_1
X_9124_ _9485_/CLK _9124_/D fanout404/X VGND VGND VPWR VPWR _9124_/Q sky130_fd_sc_hd__dfrtp_4
Xhold954 _9524_/Q VGND VGND VPWR VPWR hold954/X sky130_fd_sc_hd__dlygate4sd3_1
X_6336_ _7001_/A _6779_/A VGND VGND VPWR VPWR _6355_/C sky130_fd_sc_hd__nor2_1
XFILLER_89_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold965 _8789_/Q VGND VGND VPWR VPWR _5047_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold976 _9513_/Q VGND VGND VPWR VPWR hold976/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 _9517_/Q VGND VGND VPWR VPWR hold987/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 _8704_/X VGND VGND VPWR VPWR _9532_/D sky130_fd_sc_hd__dlygate4sd3_1
X_9055_ _9110_/CLK _9055_/D VGND VGND VPWR VPWR _9055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6267_ _7002_/A _6993_/A _6266_/X VGND VGND VPWR VPWR _6268_/D sky130_fd_sc_hd__or3b_1
XFILLER_130_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5218_ _5218_/A VGND VGND VPWR VPWR _5218_/X sky130_fd_sc_hd__clkbuf_1
X_8006_ _8006_/A _8006_/B _8006_/C _8006_/D VGND VGND VPWR VPWR _8007_/B sky130_fd_sc_hd__or4_1
XFILLER_130_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6198_ _6562_/B _6558_/C VGND VGND VPWR VPWR _6199_/A sky130_fd_sc_hd__or2_1
XFILLER_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5149_ _5149_/A VGND VGND VPWR VPWR _5149_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8908_ _9069_/CLK _8908_/D fanout429/X VGND VGND VPWR VPWR _8908_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_72_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8839_ _9475_/CLK _8839_/D fanout481/X VGND VGND VPWR VPWR _8839_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_40_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4520_ _9230_/Q _7266_/A _7605_/A _9382_/Q _4519_/X VGND VGND VPWR VPWR _4521_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_144_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold206 _7192_/X VGND VGND VPWR VPWR _7193_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4451_ _9247_/Q _7304_/A _7781_/A _9463_/Q VGND VGND VPWR VPWR _4451_/X sky130_fd_sc_hd__a22o_1
XFILLER_156_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold217 _7368_/X VGND VGND VPWR VPWR _7369_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 _7072_/X VGND VGND VPWR VPWR _7073_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold239 _7530_/X VGND VGND VPWR VPWR _7531_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7170_ _5465_/X hold639/X _7174_/S VGND VGND VPWR VPWR _7170_/X sky130_fd_sc_hd__mux2_1
X_4382_ _4858_/B _4492_/B VGND VGND VPWR VPWR _7228_/A sky130_fd_sc_hd__nor2_8
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6121_ _6906_/B _6748_/B _6906_/C VGND VGND VPWR VPWR _6754_/B sky130_fd_sc_hd__nor3_2
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ _6052_/A VGND VGND VPWR VPWR _9092_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ hold8/A hold76/A hold39/A VGND VGND VPWR VPWR _5003_/X sky130_fd_sc_hd__a21o_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6954_ _6954_/A VGND VGND VPWR VPWR _9108_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5905_ _5905_/A VGND VGND VPWR VPWR _5905_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6885_ _7003_/A _6939_/B _6885_/C VGND VGND VPWR VPWR _6886_/D sky130_fd_sc_hd__nand3b_1
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8624_ _8624_/A _8624_/B _8624_/C _8624_/D VGND VGND VPWR VPWR _8625_/C sky130_fd_sc_hd__or4_1
XFILLER_167_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5836_ hold816/X hold15/X _5842_/S VGND VGND VPWR VPWR _5836_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5767_ hold619/X _5683_/X _5771_/S VGND VGND VPWR VPWR _5768_/A sky130_fd_sc_hd__mux2_1
X_8555_ _9471_/Q _8354_/A _8376_/A _9431_/Q VGND VGND VPWR VPWR _8555_/X sky130_fd_sc_hd__a22o_1
X_7506_ _7433_/X _9331_/Q _7515_/S VGND VGND VPWR VPWR _7506_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4718_ _9315_/Q _7463_/A _7091_/A _9150_/Q _4717_/X VGND VGND VPWR VPWR _4723_/B
+ sky130_fd_sc_hd__a221o_1
X_8486_ _9316_/Q _8372_/X _8369_/X _9324_/Q _8485_/X VGND VGND VPWR VPWR _8487_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_175_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5698_ _5647_/X hold578/X _5702_/S VGND VGND VPWR VPWR _5699_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4649_ _4649_/A _4649_/B _4649_/C _4649_/D VGND VGND VPWR VPWR _4689_/A sky130_fd_sc_hd__or4_1
X_7437_ _7436_/X hold288/X _7444_/S VGND VGND VPWR VPWR _7438_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold740 _9406_/Q VGND VGND VPWR VPWR hold740/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold751 _7387_/X VGND VGND VPWR VPWR _7388_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7368_ _7242_/X hold216/X _7372_/S VGND VGND VPWR VPWR _7368_/X sky130_fd_sc_hd__mux2_1
Xhold762 _9246_/Q VGND VGND VPWR VPWR hold762/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 _7512_/X VGND VGND VPWR VPWR _7513_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9107_ _9110_/CLK _9107_/D fanout503/X VGND VGND VPWR VPWR hold62/A sky130_fd_sc_hd__dfrtp_4
X_6319_ _6151_/Y _6152_/X _6380_/B VGND VGND VPWR VPWR _6392_/B sky130_fd_sc_hd__mux2_1
Xhold784 _8890_/Q VGND VGND VPWR VPWR hold784/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold795 _7262_/X VGND VGND VPWR VPWR _7263_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7299_ _7514_/A VGND VGND VPWR VPWR _7299_/X sky130_fd_sc_hd__buf_4
XFILLER_39_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9038_ _9090_/CLK _9038_/D fanout453/X VGND VGND VPWR VPWR _9038_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_89_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6670_ _6673_/B _6670_/B _6672_/C VGND VGND VPWR VPWR _6836_/A sky130_fd_sc_hd__and3_1
XFILLER_149_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5621_ hold525/X _5587_/X _5627_/S VGND VGND VPWR VPWR _5622_/A sky130_fd_sc_hd__mux2_1
X_8340_ _8392_/A _8389_/A _8357_/A VGND VGND VPWR VPWR _8360_/B sky130_fd_sc_hd__and3_2
X_5552_ _5291_/X hold899/X _5560_/S VGND VGND VPWR VPWR _5553_/A sky130_fd_sc_hd__mux2_1
X_4503_ _9295_/Q _7408_/A _4502_/Y _4503_/B2 VGND VGND VPWR VPWR _4503_/X sky130_fd_sc_hd__a22o_1
XFILLER_157_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8271_ _8967_/Q _7960_/X _7967_/X _8972_/Q _8270_/X VGND VGND VPWR VPWR _8272_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_172_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5483_ _5483_/A VGND VGND VPWR VPWR _8843_/D sky130_fd_sc_hd__clkbuf_1
X_4434_ hold33/X VGND VGND VPWR VPWR _7158_/A sky130_fd_sc_hd__clkbuf_16
X_7222_ _5465_/X hold679/X _7226_/S VGND VGND VPWR VPWR _7222_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7153_ _7153_/A VGND VGND VPWR VPWR _7153_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4365_ hold49/X hold39/X hold22/X VGND VGND VPWR VPWR _4365_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6104_ _6104_/A VGND VGND VPWR VPWR _6891_/B sky130_fd_sc_hd__buf_4
XFILLER_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7084_ _9144_/Q hold46/X hold65/X VGND VGND VPWR VPWR _7084_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6035_ hold468/X _5809_/X _6041_/S VGND VGND VPWR VPWR _6036_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7986_ _9392_/Q _7977_/X _7979_/X _9224_/Q _7985_/X VGND VGND VPWR VPWR _8006_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6937_ _6937_/A _6937_/B _6937_/C _6937_/D VGND VGND VPWR VPWR _7003_/B sky130_fd_sc_hd__or4_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6868_ _6958_/A VGND VGND VPWR VPWR _6942_/A sky130_fd_sc_hd__inv_2
XFILLER_10_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8607_ _8964_/Q _8346_/X _8386_/A _8934_/Q VGND VGND VPWR VPWR _8607_/X sky130_fd_sc_hd__a22o_1
X_5819_ _5453_/C _5901_/A VGND VGND VPWR VPWR _5819_/X sky130_fd_sc_hd__and2b_1
X_9587_ _9587_/A _5081_/Y VGND VGND VPWR VPWR mgmt_gpio_out[33] sky130_fd_sc_hd__ebufn_8
XFILLER_50_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6799_ _6799_/A _7001_/B VGND VGND VPWR VPWR _6870_/A sky130_fd_sc_hd__nor2_1
XFILLER_10_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8538_ _9446_/Q _8301_/A _8344_/X _9486_/Q VGND VGND VPWR VPWR _8538_/X sky130_fd_sc_hd__a22o_1
XFILLER_6_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8469_ _9387_/Q _8292_/A _8358_/A _9291_/Q VGND VGND VPWR VPWR _8469_/X sky130_fd_sc_hd__a22o_1
XFILLER_163_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold570 _9218_/Q VGND VGND VPWR VPWR hold570/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold581 _5428_/X VGND VGND VPWR VPWR _5429_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 _8850_/Q VGND VGND VPWR VPWR hold592/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1270 _8876_/Q VGND VGND VPWR VPWR hold453/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1281 _8934_/Q VGND VGND VPWR VPWR hold466/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput190 wb_dat_i[4] VGND VGND VPWR VPWR _8752_/B1 sky130_fd_sc_hd__clkbuf_1
X_7840_ _7840_/A VGND VGND VPWR VPWR _9483_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7771_ _7648_/X _9451_/Q _7779_/S VGND VGND VPWR VPWR _7771_/X sky130_fd_sc_hd__mux2_1
X_4983_ _4351_/X hold30/A _4983_/S VGND VGND VPWR VPWR _4984_/B sky130_fd_sc_hd__mux2_1
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9510_ _9531_/CLK _9510_/D fanout454/X VGND VGND VPWR VPWR _9510_/Q sky130_fd_sc_hd__dfrtp_1
X_6722_ _6719_/Y _6721_/X _6717_/Y _6643_/B _6882_/A VGND VGND VPWR VPWR _6993_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_177_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9441_ _9482_/CLK _9441_/D fanout432/X VGND VGND VPWR VPWR _9441_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_149_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6653_ _6653_/A _6822_/B VGND VGND VPWR VPWR _6659_/B sky130_fd_sc_hd__or2_1
X_5604_ _5604_/A VGND VGND VPWR VPWR _8896_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9372_ _9468_/CLK _9372_/D fanout465/X VGND VGND VPWR VPWR _9372_/Q sky130_fd_sc_hd__dfrtp_4
X_6584_ _6754_/A _6585_/B _6583_/X _6377_/X VGND VGND VPWR VPWR _6584_/X sky130_fd_sc_hd__o31a_1
XFILLER_191_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_733 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8323_ _8352_/A _8392_/A _8357_/A VGND VGND VPWR VPWR _8354_/C sky130_fd_sc_hd__and3_2
X_5535_ _5535_/A VGND VGND VPWR VPWR _8865_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5466_ _5465_/X hold816/X _5472_/S VGND VGND VPWR VPWR _5466_/X sky130_fd_sc_hd__mux2_1
X_8254_ _8971_/Q _7967_/X _8008_/B _8253_/X VGND VGND VPWR VPWR _8254_/X sky130_fd_sc_hd__a22o_1
XFILLER_132_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_747 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4417_ hold41/X hold63/X VGND VGND VPWR VPWR hold42/A sky130_fd_sc_hd__nor2b_4
XFILLER_105_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7205_ _5465_/X hold805/X _7209_/S VGND VGND VPWR VPWR _7205_/X sky130_fd_sc_hd__mux2_1
X_5397_ _5397_/A VGND VGND VPWR VPWR _8811_/D sky130_fd_sc_hd__clkbuf_1
X_8185_ _9069_/Q _7979_/A _7993_/A _8983_/Q VGND VGND VPWR VPWR _8185_/X sky130_fd_sc_hd__a22o_1
XFILLER_120_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7136_ _7136_/A VGND VGND VPWR VPWR _9166_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7067_ _7067_/A VGND VGND VPWR VPWR _9136_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6018_ hold24/X VGND VGND VPWR VPWR _6018_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_39_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7969_ _7969_/A VGND VGND VPWR VPWR _7969_/X sky130_fd_sc_hd__buf_6
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_240 _9164_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_251 wb_sel_i[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_262 _5174_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_273 _5012_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_284 input18/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_295 _4836_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer1 _5226_/A1 VGND VGND VPWR VPWR _9550_/CLK sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_174_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5320_ _5330_/A _5334_/B VGND VGND VPWR VPWR _5321_/A sky130_fd_sc_hd__and2_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5251_ _9307_/Q VGND VGND VPWR VPWR _5251_/Y sky130_fd_sc_hd__inv_2
X_5182_ _5182_/A VGND VGND VPWR VPWR _5182_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_68_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8941_ _9087_/CLK _8941_/D fanout445/X VGND VGND VPWR VPWR _8941_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_113_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8872_ _9483_/CLK _8872_/D fanout474/X VGND VGND VPWR VPWR _8872_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_37_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7823_ _7823_/A VGND VGND VPWR VPWR _9475_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7754_ _9443_/Q hold46/X _7762_/S VGND VGND VPWR VPWR hold47/A sky130_fd_sc_hd__mux2_1
X_4966_ hold94/A VGND VGND VPWR VPWR _5040_/B sky130_fd_sc_hd__buf_2
X_6705_ _6521_/B _6413_/B _6441_/B _6869_/C VGND VGND VPWR VPWR _6706_/D sky130_fd_sc_hd__a31o_1
XFILLER_20_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7685_ _7648_/X _9411_/Q _7693_/S VGND VGND VPWR VPWR _7685_/X sky130_fd_sc_hd__mux2_1
X_4897_ _9069_/Q _5996_/A _7139_/A _9168_/Q VGND VGND VPWR VPWR _4897_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9424_ _9471_/CLK _9424_/D _5070_/A VGND VGND VPWR VPWR _9424_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_165_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6636_ _6732_/B _6830_/A _6463_/A VGND VGND VPWR VPWR _6636_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_165_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9355_ _9475_/CLK _9355_/D fanout478/X VGND VGND VPWR VPWR _9355_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6567_ _6874_/A _6561_/X _6792_/A _6574_/B VGND VGND VPWR VPWR _6567_/X sky130_fd_sc_hd__o22a_1
XFILLER_192_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8306_ _9288_/Q _8294_/X _8298_/X _9328_/Q _8305_/X VGND VGND VPWR VPWR _8306_/X
+ sky130_fd_sc_hd__a221o_1
X_5518_ _5518_/A _5693_/B VGND VGND VPWR VPWR _5527_/S sky130_fd_sc_hd__nand2_2
XFILLER_106_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9286_ _9325_/CLK _9286_/D fanout464/X VGND VGND VPWR VPWR _9286_/Q sky130_fd_sc_hd__dfrtp_4
X_6498_ _6635_/A _6498_/B VGND VGND VPWR VPWR _6499_/B sky130_fd_sc_hd__nand2_1
XFILLER_145_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8237_ _9076_/Q _8034_/X _7999_/X _8950_/Q _8236_/X VGND VGND VPWR VPWR _8238_/D
+ sky130_fd_sc_hd__a221o_1
X_5449_ _5449_/A VGND VGND VPWR VPWR _5449_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_78_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8168_ _9239_/Q _8034_/X _8165_/X _8167_/X VGND VGND VPWR VPWR _8171_/C sky130_fd_sc_hd__a211o_1
X_7119_ _7119_/A VGND VGND VPWR VPWR _9159_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8099_ _9260_/Q _7958_/X _8224_/B _9420_/Q VGND VGND VPWR VPWR _8099_/X sky130_fd_sc_hd__a22o_1
XFILLER_19_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _8767_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_43_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4820_ _4820_/A VGND VGND VPWR VPWR _9113_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ _4751_/A _4751_/B _4751_/C _4751_/D VGND VGND VPWR VPWR _4752_/D sky130_fd_sc_hd__or4_2
XFILLER_193_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7470_ _7470_/A VGND VGND VPWR VPWR _9314_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4682_ input56/X _5901_/A _5540_/A _8872_/Q VGND VGND VPWR VPWR _4682_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6421_ _6421_/A VGND VGND VPWR VPWR _6897_/B sky130_fd_sc_hd__buf_4
XFILLER_162_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9140_ _9474_/CLK _9140_/D fanout427/X VGND VGND VPWR VPWR _9140_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_127_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6352_ _6352_/A _6560_/A _6352_/C _6352_/D VGND VGND VPWR VPWR _6352_/X sky130_fd_sc_hd__or4_1
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5303_ _5303_/A VGND VGND VPWR VPWR _8773_/D sky130_fd_sc_hd__clkbuf_1
X_9071_ _9161_/CLK _9071_/D fanout445/X VGND VGND VPWR VPWR _9071_/Q sky130_fd_sc_hd__dfstp_4
X_6283_ _6311_/B _6624_/B _6195_/Y _6282_/X VGND VGND VPWR VPWR _6283_/X sky130_fd_sc_hd__o211a_1
XFILLER_115_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8022_ _9353_/Q _8020_/X _7958_/X _9257_/Q _8021_/X VGND VGND VPWR VPWR _8027_/B
+ sky130_fd_sc_hd__a221o_1
X_5234_ hold74/X VGND VGND VPWR VPWR _5413_/S sky130_fd_sc_hd__buf_6
XFILLER_69_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5165_ input84/X _5071_/C _8795_/Q VGND VGND VPWR VPWR _5166_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5096_ _9331_/Q VGND VGND VPWR VPWR _5096_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8924_ _9005_/CLK _8924_/D fanout489/X VGND VGND VPWR VPWR _8924_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8855_ _9084_/CLK _8855_/D fanout445/X VGND VGND VPWR VPWR _8855_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_25_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7806_ _7806_/A VGND VGND VPWR VPWR _9467_/D sky130_fd_sc_hd__clkbuf_1
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8786_ _5207_/A1 _8786_/D _5338_/X VGND VGND VPWR VPWR _8786_/Q sky130_fd_sc_hd__dfrtp_1
X_5998_ _5998_/A VGND VGND VPWR VPWR _9069_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7737_ _7737_/A VGND VGND VPWR VPWR _9435_/D sky130_fd_sc_hd__clkbuf_1
X_4949_ _4949_/A _4949_/B _4949_/C _4949_/D VGND VGND VPWR VPWR _4960_/A sky130_fd_sc_hd__or4_1
XFILLER_184_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7668_ _7648_/X _9403_/Q _7676_/S VGND VGND VPWR VPWR _7668_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9407_ _9461_/CLK _9407_/D fanout423/X VGND VGND VPWR VPWR _9407_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6619_ _6619_/A _6944_/A _6853_/C _6619_/D VGND VGND VPWR VPWR _6620_/D sky130_fd_sc_hd__or4_1
XFILLER_137_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7599_ _7439_/X hold227/X hold75/X VGND VGND VPWR VPWR _7600_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9338_ _9370_/CLK _9338_/D fanout478/X VGND VGND VPWR VPWR _9338_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_146_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9269_ _9421_/CLK _9269_/D fanout460/X VGND VGND VPWR VPWR _9269_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput280 _8816_/Q VGND VGND VPWR VPWR pll_trim[15] sky130_fd_sc_hd__buf_12
XFILLER_58_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput291 _8826_/Q VGND VGND VPWR VPWR pll_trim[25] sky130_fd_sc_hd__buf_12
XFILLER_101_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire396 _5270_/Y VGND VGND VPWR VPWR _5287_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6970_ _6994_/A _6994_/B _6994_/C _6970_/D VGND VGND VPWR VPWR _6970_/X sky130_fd_sc_hd__or4_1
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5921_ _5633_/X hold707/X _5927_/S VGND VGND VPWR VPWR _5921_/X sky130_fd_sc_hd__mux2_1
X_8640_ _8910_/Q _8360_/C _8411_/A _8925_/Q _8639_/X VGND VGND VPWR VPWR _8650_/B
+ sky130_fd_sc_hd__a221o_1
X_5852_ hold506/X hold12/X _5867_/S VGND VGND VPWR VPWR _5852_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4803_ input45/X _4582_/A _5529_/A _8865_/Q _4802_/X VGND VGND VPWR VPWR _4806_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_167_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8571_ _9439_/Q _7908_/X _8335_/X _9279_/Q VGND VGND VPWR VPWR _8571_/X sky130_fd_sc_hd__a22o_1
X_5783_ _5783_/A VGND VGND VPWR VPWR _8972_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7522_ _7359_/X hold148/X _7534_/S VGND VGND VPWR VPWR _7523_/A sky130_fd_sc_hd__mux2_1
X_4734_ _7111_/A _4758_/A VGND VGND VPWR VPWR _4734_/Y sky130_fd_sc_hd__nor2_4
XFILLER_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7453_ _7433_/X _9307_/Q _7461_/S VGND VGND VPWR VPWR _7453_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4665_ _4665_/A _4794_/B VGND VGND VPWR VPWR _5642_/A sky130_fd_sc_hd__nor2_8
XFILLER_175_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6404_ _6334_/B _6906_/B _6403_/X VGND VGND VPWR VPWR _6404_/Y sky130_fd_sc_hd__o21ai_1
Xhold900 _9432_/Q VGND VGND VPWR VPWR hold900/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold911 _9200_/Q VGND VGND VPWR VPWR hold911/X sky130_fd_sc_hd__dlygate4sd3_1
X_7384_ _7384_/A VGND VGND VPWR VPWR _9276_/D sky130_fd_sc_hd__clkbuf_1
X_4596_ _4667_/A _4891_/B VGND VGND VPWR VPWR _6043_/A sky130_fd_sc_hd__nor2_4
Xhold922 _9264_/Q VGND VGND VPWR VPWR hold922/X sky130_fd_sc_hd__dlygate4sd3_1
X_9123_ _9485_/CLK _9123_/D fanout404/X VGND VGND VPWR VPWR _9123_/Q sky130_fd_sc_hd__dfstp_2
Xhold933 _7145_/X VGND VGND VPWR VPWR _7146_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_127_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold944 _8805_/Q VGND VGND VPWR VPWR hold944/X sky130_fd_sc_hd__dlygate4sd3_1
X_6335_ _7001_/A _6666_/B VGND VGND VPWR VPWR _6573_/B sky130_fd_sc_hd__nor2_1
XFILLER_162_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold955 _8503_/X VGND VGND VPWR VPWR _9524_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 _5046_/X VGND VGND VPWR VPWR _8790_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 _8152_/X VGND VGND VPWR VPWR _9513_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold988 _8285_/X VGND VGND VPWR VPWR _9519_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9054_ _9110_/CLK _9054_/D VGND VGND VPWR VPWR _9054_/Q sky130_fd_sc_hd__dfxtp_1
Xhold999 _8780_/Q VGND VGND VPWR VPWR hold999/X sky130_fd_sc_hd__dlygate4sd3_1
X_6266_ _6266_/A _7001_/A VGND VGND VPWR VPWR _6266_/X sky130_fd_sc_hd__or2_1
XFILLER_142_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8005_ _9360_/Q _7997_/X _7999_/X _9424_/Q _8004_/X VGND VGND VPWR VPWR _8006_/D
+ sky130_fd_sc_hd__a221o_1
X_5217_ _9009_/Q input3/X input1/X VGND VGND VPWR VPWR _5218_/A sky130_fd_sc_hd__mux2_4
XFILLER_57_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6197_ _6795_/A _6197_/B VGND VGND VPWR VPWR _6562_/B sky130_fd_sc_hd__nand2_1
XFILLER_28_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5148_ _8705_/A VGND VGND VPWR VPWR _8706_/A sky130_fd_sc_hd__inv_2
XFILLER_29_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5079_ _8792_/Q hold17/X _8829_/Q _5016_/B VGND VGND VPWR VPWR _8777_/D sky130_fd_sc_hd__o211a_1
XFILLER_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8907_ _9442_/CLK _8907_/D fanout436/X VGND VGND VPWR VPWR _8907_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_37_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8838_ _9370_/CLK _8838_/D fanout477/X VGND VGND VPWR VPWR _8838_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_71_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8769_ _5275_/A _8769_/A2 _8768_/X VGND VGND VPWR VPWR _8769_/X sky130_fd_sc_hd__a21o_1
XFILLER_40_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4450_ _7158_/A _4670_/B VGND VGND VPWR VPWR _4450_/Y sky130_fd_sc_hd__nor2_2
XFILLER_156_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold207 _9255_/Q VGND VGND VPWR VPWR hold207/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold218 _9237_/Q VGND VGND VPWR VPWR hold218/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 _9389_/Q VGND VGND VPWR VPWR hold229/X sky130_fd_sc_hd__dlygate4sd3_1
X_4381_ _4381_/A VGND VGND VPWR VPWR _4492_/B sky130_fd_sc_hd__buf_8
XFILLER_98_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6120_ _6504_/A _6415_/B VGND VGND VPWR VPWR _6906_/C sky130_fd_sc_hd__nand2_4
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ hold204/X hold46/X _6053_/S VGND VGND VPWR VPWR _6052_/A sky130_fd_sc_hd__mux2_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _5040_/B _5002_/B VGND VGND VPWR VPWR _5002_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6953_ _6953_/A _6953_/B _6953_/C _6952_/X VGND VGND VPWR VPWR _6954_/A sky130_fd_sc_hd__or4b_1
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5904_ _5633_/X _9579_/A _5916_/S VGND VGND VPWR VPWR _5904_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6884_ _6624_/B _6574_/B _6939_/D _6939_/A VGND VGND VPWR VPWR _6885_/C sky130_fd_sc_hd__o211a_1
X_8623_ _9049_/Q _8356_/A _8360_/B _8889_/Q _8622_/X VGND VGND VPWR VPWR _8624_/D
+ sky130_fd_sc_hd__a221o_1
X_5835_ _5835_/A VGND VGND VPWR VPWR _5835_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8554_ _8554_/A VGND VGND VPWR VPWR _9526_/D sky130_fd_sc_hd__clkbuf_1
X_5766_ _5766_/A VGND VGND VPWR VPWR _8964_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7505_ _7505_/A VGND VGND VPWR VPWR _9330_/D sky130_fd_sc_hd__clkbuf_1
X_4717_ _9129_/Q _7043_/A _5762_/A _8966_/Q VGND VGND VPWR VPWR _4717_/X sky130_fd_sc_hd__a22o_1
XFILLER_108_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8485_ _9300_/Q _8314_/X _8331_/X _9404_/Q VGND VGND VPWR VPWR _8485_/X sky130_fd_sc_hd__a22o_1
XFILLER_175_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5697_ _5697_/A VGND VGND VPWR VPWR _8934_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7436_ hold24/X VGND VGND VPWR VPWR _7436_/X sky130_fd_sc_hd__clkbuf_2
X_4648_ _8957_/Q _5738_/A _6032_/A _9088_/Q _4647_/X VGND VGND VPWR VPWR _4649_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold730 _9342_/Q VGND VGND VPWR VPWR hold730/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 _7674_/X VGND VGND VPWR VPWR _7675_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7367_ _7367_/A VGND VGND VPWR VPWR _9268_/D sky130_fd_sc_hd__clkbuf_1
X_4579_ _4579_/A1 _4502_/Y _7228_/A _9213_/Q _4578_/X VGND VGND VPWR VPWR _4591_/B
+ sky130_fd_sc_hd__a221o_1
Xhold752 _7104_/X VGND VGND VPWR VPWR _7105_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold763 _7317_/X VGND VGND VPWR VPWR _7318_/A sky130_fd_sc_hd__dlygate4sd3_1
X_9106_ _9110_/CLK _9106_/D _5929_/B VGND VGND VPWR VPWR _9106_/Q sky130_fd_sc_hd__dfrtp_4
X_6318_ _6318_/A _6672_/B VGND VGND VPWR VPWR _6380_/B sky130_fd_sc_hd__nand2_1
Xhold774 _9109_/Q VGND VGND VPWR VPWR hold774/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 _9214_/Q VGND VGND VPWR VPWR hold785/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7298_ _7298_/A VGND VGND VPWR VPWR _9238_/D sky130_fd_sc_hd__clkbuf_1
Xhold796 hold796/A VGND VGND VPWR VPWR hold796/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9037_ _9187_/CLK _9037_/D fanout455/X VGND VGND VPWR VPWR _9037_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_130_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6249_ _6249_/A _6266_/A _6610_/B VGND VGND VPWR VPWR _6250_/D sky130_fd_sc_hd__or3_1
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_61_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _9162_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_76_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _9376_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_40_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_14_csclk clkbuf_opt_1_0_csclk/X VGND VGND VPWR VPWR _9173_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_29_csclk _9303_/CLK VGND VGND VPWR VPWR _9370_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold90 hold90/A VGND VGND VPWR VPWR hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_90_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5620_ _5620_/A VGND VGND VPWR VPWR _8903_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5551_ _5551_/A _5693_/B VGND VGND VPWR VPWR _5560_/S sky130_fd_sc_hd__nand2_2
XFILLER_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4502_ _4758_/A _4667_/B VGND VGND VPWR VPWR _4502_/Y sky130_fd_sc_hd__nor2_8
X_8270_ _9083_/Q _7949_/X _7962_/X _8907_/Q VGND VGND VPWR VPWR _8270_/X sky130_fd_sc_hd__a22o_1
X_5482_ _5311_/X hold367/X _5490_/S VGND VGND VPWR VPWR _5482_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7221_ _7221_/A VGND VGND VPWR VPWR _9204_/D sky130_fd_sc_hd__clkbuf_1
X_4433_ hold32/X VGND VGND VPWR VPWR hold33/A sky130_fd_sc_hd__buf_12
X_7152_ _6015_/X _9173_/Q _7156_/S VGND VGND VPWR VPWR _7152_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4364_ _4364_/A VGND VGND VPWR VPWR _4758_/A sky130_fd_sc_hd__buf_8
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6103_ _6167_/B _6402_/A VGND VGND VPWR VPWR _6104_/A sky130_fd_sc_hd__or2_1
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7083_ _7083_/A VGND VGND VPWR VPWR _9143_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6034_ _6034_/A VGND VGND VPWR VPWR _9084_/D sky130_fd_sc_hd__clkbuf_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7985_ _9328_/Q _7981_/X _8008_/B _9312_/Q _7984_/X VGND VGND VPWR VPWR _7985_/X
+ sky130_fd_sc_hd__a221o_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6936_ _6603_/A _7001_/B _6255_/X VGND VGND VPWR VPWR _6937_/D sky130_fd_sc_hd__o21ai_1
XFILLER_35_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6867_ _6867_/A _6867_/B _6808_/X _6809_/C VGND VGND VPWR VPWR _6958_/A sky130_fd_sc_hd__or4bb_2
XFILLER_179_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8606_ _8959_/Q _8402_/X _8378_/X _8944_/Q _8605_/X VGND VGND VPWR VPWR _8606_/X
+ sky130_fd_sc_hd__a221o_1
X_5818_ hold828/X _7517_/A _5842_/S VGND VGND VPWR VPWR _5818_/X sky130_fd_sc_hd__mux2_1
X_9586_ _9586_/A _5082_/Y VGND VGND VPWR VPWR mgmt_gpio_out[32] sky130_fd_sc_hd__ebufn_8
XFILLER_10_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6798_ _6867_/A _6955_/D _6880_/A _6798_/D VGND VGND VPWR VPWR _6806_/C sky130_fd_sc_hd__or4_1
X_8537_ _8537_/A _8537_/B _8537_/C _8537_/D VGND VGND VPWR VPWR _8550_/B sky130_fd_sc_hd__or4_1
X_5749_ hold19/X VGND VGND VPWR VPWR _7132_/B sky130_fd_sc_hd__buf_4
XFILLER_6_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8468_ _9243_/Q _8324_/X _8360_/B _9307_/Q VGND VGND VPWR VPWR _8473_/B sky130_fd_sc_hd__a22o_1
XFILLER_108_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7419_ _7242_/X hold271/X _7423_/S VGND VGND VPWR VPWR _7419_/X sky130_fd_sc_hd__mux2_1
X_8399_ _8399_/A VGND VGND VPWR VPWR _8400_/B sky130_fd_sc_hd__buf_6
XFILLER_151_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold560 _9242_/Q VGND VGND VPWR VPWR hold560/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold571 _7254_/X VGND VGND VPWR VPWR _7255_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold582 _8980_/Q VGND VGND VPWR VPWR hold582/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 _5498_/X VGND VGND VPWR VPWR _5499_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1260 _8867_/Q VGND VGND VPWR VPWR _5538_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1271 _8881_/Q VGND VGND VPWR VPWR hold410/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1282 _7381_/X VGND VGND VPWR VPWR hold697/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_400 _7302_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput180 wb_dat_i[24] VGND VGND VPWR VPWR _8729_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput191 wb_dat_i[5] VGND VGND VPWR VPWR _8756_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7770_ _7770_/A VGND VGND VPWR VPWR _9450_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4982_ hold29/A hold55/A hold80/A _4997_/B VGND VGND VPWR VPWR _4983_/S sky130_fd_sc_hd__nand4_1
X_6721_ _6721_/A _6724_/A VGND VGND VPWR VPWR _6721_/X sky130_fd_sc_hd__and2_2
XFILLER_32_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9440_ _9480_/CLK _9440_/D fanout414/X VGND VGND VPWR VPWR _9440_/Q sky130_fd_sc_hd__dfstp_1
X_6652_ _6811_/B _6422_/B _6521_/B _6506_/Y VGND VGND VPWR VPWR _6822_/B sky130_fd_sc_hd__a31o_1
X_5603_ hold449/X _5398_/X _5605_/S VGND VGND VPWR VPWR _5604_/A sky130_fd_sc_hd__mux2_1
X_9371_ _9475_/CLK _9371_/D fanout481/X VGND VGND VPWR VPWR _9371_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_164_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6583_ _6778_/A _6867_/A _6955_/B _6583_/D VGND VGND VPWR VPWR _6583_/X sky130_fd_sc_hd__or4_1
XFILLER_176_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8322_ _8356_/B VGND VGND VPWR VPWR _8322_/X sky130_fd_sc_hd__buf_8
X_5534_ _5306_/X hold473/X _5538_/S VGND VGND VPWR VPWR _5534_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8253_ hold71/A _8275_/B VGND VGND VPWR VPWR _8253_/X sky130_fd_sc_hd__or2_1
XFILLER_127_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5465_ _5465_/A VGND VGND VPWR VPWR _5465_/X sky130_fd_sc_hd__clkbuf_16
X_7204_ _7204_/A VGND VGND VPWR VPWR _9196_/D sky130_fd_sc_hd__clkbuf_1
X_4416_ _4670_/B _4492_/B VGND VGND VPWR VPWR _4416_/Y sky130_fd_sc_hd__nor2_2
XFILLER_133_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8184_ _8184_/A _8184_/B _8184_/C _8184_/D VGND VGND VPWR VPWR _8193_/A sky130_fd_sc_hd__or4_1
X_5396_ _8811_/Q _5395_/X _5416_/S VGND VGND VPWR VPWR _5396_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7135_ _9166_/Q _5809_/X _7137_/S VGND VGND VPWR VPWR _7135_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7066_ _9136_/Q _5690_/A _7072_/S VGND VGND VPWR VPWR _7066_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6017_ _6017_/A VGND VGND VPWR VPWR _9077_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _5237_/A2 sky130_fd_sc_hd__clkbuf_16
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7968_ _8206_/B _7992_/C _8002_/C VGND VGND VPWR VPWR _7969_/A sky130_fd_sc_hd__and3_2
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6919_ _6997_/C _6972_/B _6918_/X VGND VGND VPWR VPWR _6919_/X sky130_fd_sc_hd__or3b_1
X_7899_ _9498_/Q _9497_/Q VGND VGND VPWR VPWR _8392_/A sky130_fd_sc_hd__and2_2
XFILLER_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9569_ _9569_/A _5099_/Y VGND VGND VPWR VPWR mgmt_gpio_out[15] sky130_fd_sc_hd__ebufn_2
XFILLER_109_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold390 _8951_/Q VGND VGND VPWR VPWR hold390/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1090 _7736_/X VGND VGND VPWR VPWR _7737_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_230 _9433_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_241 _9000_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_252 input93/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_263 _5174_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_274 _5285_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_285 _4759_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_296 _7499_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer2 _5226_/A1 VGND VGND VPWR VPWR _9501_/CLK sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_173_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_586 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5250_ _9299_/Q VGND VGND VPWR VPWR _5250_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5181_ _8794_/Q _5181_/B VGND VGND VPWR VPWR _5182_/A sky130_fd_sc_hd__and2b_1
XFILLER_68_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8940_ _9087_/CLK _8940_/D fanout445/X VGND VGND VPWR VPWR _8940_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_56_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8871_ _9181_/CLK _8871_/D fanout488/X VGND VGND VPWR VPWR _8871_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7822_ _7648_/X _9475_/Q _7830_/S VGND VGND VPWR VPWR _7822_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7753_ _7753_/A VGND VGND VPWR VPWR _9442_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4965_ hold943/X _4964_/B _4961_/X _4964_/Y VGND VGND VPWR VPWR _9111_/D sky130_fd_sc_hd__a22o_1
XFILLER_51_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6704_ _6704_/A _6704_/B _6704_/C _6704_/D VGND VGND VPWR VPWR _6706_/C sky130_fd_sc_hd__or4_1
XFILLER_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7684_ _7684_/A VGND VGND VPWR VPWR _9410_/D sky130_fd_sc_hd__clkbuf_1
X_4896_ _4896_/A _4896_/B _4896_/C _4896_/D VGND VGND VPWR VPWR _4922_/A sky130_fd_sc_hd__or4_1
X_9423_ _9461_/CLK _9423_/D fanout421/X VGND VGND VPWR VPWR _9423_/Q sky130_fd_sc_hd__dfrtp_1
X_6635_ _6635_/A _6635_/B VGND VGND VPWR VPWR _6976_/B sky130_fd_sc_hd__nor2_2
XFILLER_149_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9354_ _9370_/CLK _9354_/D fanout477/X VGND VGND VPWR VPWR _9354_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6566_ _6715_/B _6566_/B VGND VGND VPWR VPWR _6574_/B sky130_fd_sc_hd__nor2_2
XFILLER_138_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8305_ _9440_/Q _8398_/B _8304_/X _9392_/Q VGND VGND VPWR VPWR _8305_/X sky130_fd_sc_hd__a22o_1
XFILLER_152_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5517_ hold20/X VGND VGND VPWR VPWR _5693_/B sky130_fd_sc_hd__buf_8
X_9285_ _9325_/CLK _9285_/D fanout464/X VGND VGND VPWR VPWR _9285_/Q sky130_fd_sc_hd__dfrtp_1
X_6497_ _6732_/B _6514_/A VGND VGND VPWR VPWR _6726_/B sky130_fd_sc_hd__nor2_2
XFILLER_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8236_ _8925_/Q _7933_/X _7973_/X _8855_/Q VGND VGND VPWR VPWR _8236_/X sky130_fd_sc_hd__a22o_1
X_5448_ _7011_/A _7013_/B VGND VGND VPWR VPWR _5449_/A sky130_fd_sc_hd__and2_1
XFILLER_160_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8167_ _9247_/Q _7949_/A _7973_/A _9199_/Q _8166_/X VGND VGND VPWR VPWR _8167_/X
+ sky130_fd_sc_hd__a221o_1
X_5379_ _5379_/A VGND VGND VPWR VPWR _5379_/X sky130_fd_sc_hd__clkbuf_1
X_7118_ _6012_/X _9159_/Q _7124_/S VGND VGND VPWR VPWR _7118_/X sky130_fd_sc_hd__mux2_1
X_8098_ _9228_/Q _7979_/X _7993_/X _9388_/Q VGND VGND VPWR VPWR _8098_/X sky130_fd_sc_hd__a22o_1
XFILLER_87_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7049_ _7049_/A VGND VGND VPWR VPWR _9128_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _9435_/Q _4906_/A2 _7408_/A _9291_/Q _4749_/X VGND VGND VPWR VPWR _4751_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4681_ hold60/X _7126_/B VGND VGND VPWR VPWR _5540_/A sky130_fd_sc_hd__nor2_8
X_6420_ _6440_/A _6420_/B VGND VGND VPWR VPWR _6421_/A sky130_fd_sc_hd__nor2_1
XFILLER_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6351_ _6779_/A _6666_/B _6603_/A VGND VGND VPWR VPWR _6352_/D sky130_fd_sc_hd__a21oi_1
XFILLER_115_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5302_ _5301_/X hold462/X _5316_/S VGND VGND VPWR VPWR _5302_/X sky130_fd_sc_hd__mux2_1
X_9070_ _9161_/CLK _9070_/D fanout441/X VGND VGND VPWR VPWR _9070_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_6_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6282_ _6311_/B _6800_/A _6591_/A _6278_/X _6281_/Y VGND VGND VPWR VPWR _6282_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_170_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8021_ _9337_/Q _7933_/A _7990_/A _9273_/Q VGND VGND VPWR VPWR _8021_/X sky130_fd_sc_hd__a22o_1
X_5233_ _5233_/A VGND VGND VPWR VPWR _5233_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5164_ _5040_/C _5127_/Y _5016_/B _5040_/B VGND VGND VPWR VPWR _8829_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5095_ _9339_/Q VGND VGND VPWR VPWR _5095_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8923_ _9467_/CLK _8923_/D fanout475/X VGND VGND VPWR VPWR _8923_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_71_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8854_ _9084_/CLK _8854_/D fanout445/X VGND VGND VPWR VPWR _8854_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7805_ _7648_/X _9467_/Q _7813_/S VGND VGND VPWR VPWR _7805_/X sky130_fd_sc_hd__mux2_1
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8785_ _5207_/A1 _8785_/D _5335_/X VGND VGND VPWR VPWR hold14/A sky130_fd_sc_hd__dfrtp_1
X_5997_ hold901/X _5761_/X _6005_/S VGND VGND VPWR VPWR _5998_/A sky130_fd_sc_hd__mux2_1
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7736_ _7648_/X _9435_/Q hold86/X VGND VGND VPWR VPWR _7736_/X sky130_fd_sc_hd__mux2_1
X_4948_ _9256_/Q _7339_/A _7144_/A input61/X _4947_/X VGND VGND VPWR VPWR _4949_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_178_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7667_ _7667_/A VGND VGND VPWR VPWR _9402_/D sky130_fd_sc_hd__clkbuf_1
X_4879_ _9433_/Q _7729_/A _7027_/A _9120_/Q VGND VGND VPWR VPWR _4879_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9406_ _9461_/CLK _9406_/D fanout423/X VGND VGND VPWR VPWR _9406_/Q sky130_fd_sc_hd__dfrtp_4
X_6618_ _7002_/A _6618_/B _6618_/C _6618_/D VGND VGND VPWR VPWR _6619_/D sky130_fd_sc_hd__or4_1
X_7598_ _7598_/A VGND VGND VPWR VPWR _9372_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9337_ _9483_/CLK _9337_/D fanout473/X VGND VGND VPWR VPWR _9337_/Q sky130_fd_sc_hd__dfstp_2
X_6549_ _6891_/A _6635_/A VGND VGND VPWR VPWR _6894_/A sky130_fd_sc_hd__or2_1
XFILLER_152_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9268_ _9420_/CLK _9268_/D fanout463/X VGND VGND VPWR VPWR _9268_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8219_ hold978/X _8196_/S _8217_/X _8218_/X VGND VGND VPWR VPWR _8219_/X sky130_fd_sc_hd__o22a_1
XFILLER_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput270 _9119_/Q VGND VGND VPWR VPWR pll_ena sky130_fd_sc_hd__buf_12
X_9199_ _9437_/CLK _9199_/D fanout409/X VGND VGND VPWR VPWR _9199_/Q sky130_fd_sc_hd__dfrtp_2
Xoutput281 _9132_/Q VGND VGND VPWR VPWR pll_trim[16] sky130_fd_sc_hd__buf_12
Xoutput292 _8819_/Q VGND VGND VPWR VPWR pll_trim[2] sky130_fd_sc_hd__buf_12
XFILLER_160_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire375 _4457_/Y VGND VGND VPWR VPWR _7425_/A sky130_fd_sc_hd__buf_6
XFILLER_139_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5920_ _5920_/A VGND VGND VPWR VPWR _9035_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5851_ _5851_/A VGND VGND VPWR VPWR _5851_/X sky130_fd_sc_hd__clkbuf_1
X_4802_ _8945_/Q _5715_/A _6043_/A _9091_/Q VGND VGND VPWR VPWR _4802_/X sky130_fd_sc_hd__a22o_1
X_8570_ _9231_/Q _8388_/X _8379_/X _9207_/Q _8569_/X VGND VGND VPWR VPWR _8575_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5782_ _5653_/X hold129/X _5782_/S VGND VGND VPWR VPWR _5782_/X sky130_fd_sc_hd__mux2_1
X_7521_ _7521_/A VGND VGND VPWR VPWR _9336_/D sky130_fd_sc_hd__clkbuf_1
X_4733_ _9082_/Q _6021_/A _5727_/A _8951_/Q _4732_/X VGND VGND VPWR VPWR _4741_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_187_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7452_ _7452_/A VGND VGND VPWR VPWR _9306_/D sky130_fd_sc_hd__clkbuf_1
X_4664_ _4667_/A _4794_/B VGND VGND VPWR VPWR _5918_/A sky130_fd_sc_hd__nor2_4
XFILLER_174_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6403_ _6781_/B _6887_/A _6967_/B _6482_/A _6227_/Y VGND VGND VPWR VPWR _6403_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_190_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7383_ _7239_/X hold318/X _7389_/S VGND VGND VPWR VPWR _7383_/X sky130_fd_sc_hd__mux2_1
Xhold901 hold901/A VGND VGND VPWR VPWR hold901/X sky130_fd_sc_hd__dlygate4sd3_1
X_4595_ _4635_/A _4956_/A VGND VGND VPWR VPWR _5727_/A sky130_fd_sc_hd__nor2_8
Xhold912 _9224_/Q VGND VGND VPWR VPWR hold912/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold923 hold923/A VGND VGND VPWR VPWR hold923/X sky130_fd_sc_hd__dlygate4sd3_1
X_9122_ _9485_/CLK _9122_/D fanout404/X VGND VGND VPWR VPWR _9122_/Q sky130_fd_sc_hd__dfrtp_4
Xhold934 _7146_/X VGND VGND VPWR VPWR _9170_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6334_ _6802_/A _6334_/B VGND VGND VPWR VPWR _7002_/B sky130_fd_sc_hd__nor2_1
Xhold945 _7917_/X VGND VGND VPWR VPWR _9505_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold956 _9114_/Q VGND VGND VPWR VPWR hold956/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 _9028_/Q VGND VGND VPWR VPWR _5870_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold978 _9516_/Q VGND VGND VPWR VPWR hold978/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9053_ _9110_/CLK _9053_/D VGND VGND VPWR VPWR _9053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold989 _9511_/Q VGND VGND VPWR VPWR hold989/X sky130_fd_sc_hd__dlygate4sd3_1
X_6265_ _6802_/A _6279_/A VGND VGND VPWR VPWR _6993_/A sky130_fd_sc_hd__nor2_1
X_8004_ _9264_/Q _8001_/X _8003_/X _9296_/Q VGND VGND VPWR VPWR _8004_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5216_ _5216_/A VGND VGND VPWR VPWR _5216_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6196_ _6399_/A _6232_/C VGND VGND VPWR VPWR _6197_/B sky130_fd_sc_hd__nor2_1
XFILLER_97_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5147_ _5287_/A _5115_/X _5870_/C VGND VGND VPWR VPWR _9034_/D sky130_fd_sc_hd__a21o_1
XFILLER_29_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5078_ _5067_/B _5026_/S _5077_/X hold994/X VGND VGND VPWR VPWR _8778_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8906_ _9442_/CLK _8906_/D fanout436/X VGND VGND VPWR VPWR _8906_/Q sky130_fd_sc_hd__dfrtp_4
X_8837_ _9370_/CLK _8837_/D fanout477/X VGND VGND VPWR VPWR _8837_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_80_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8768_ _5287_/A _8731_/A _8732_/B _5271_/A VGND VGND VPWR VPWR _8768_/X sky130_fd_sc_hd__a22o_1
X_7719_ _7648_/X _9427_/Q hold95/X VGND VGND VPWR VPWR _7719_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8699_ _9052_/Q _8289_/X _8341_/X _8892_/Q _8698_/X VGND VGND VPWR VPWR _8700_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_100_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold208 _7337_/X VGND VGND VPWR VPWR _7338_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold219 _7295_/X VGND VGND VPWR VPWR _7296_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4380_ hold58/X _4432_/B VGND VGND VPWR VPWR _4381_/A sky130_fd_sc_hd__or2_1
XFILLER_125_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _6050_/A VGND VGND VPWR VPWR _9091_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _5001_/A VGND VGND VPWR VPWR _8801_/D sky130_fd_sc_hd__clkbuf_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6952_ _6964_/A _6964_/C _6965_/A _6951_/X VGND VGND VPWR VPWR _6952_/X sky130_fd_sc_hd__or4b_1
X_5903_ _5903_/A VGND VGND VPWR VPWR _9017_/D sky130_fd_sc_hd__clkbuf_1
X_6883_ _6715_/B _6507_/A _6343_/C _6314_/C VGND VGND VPWR VPWR _6939_/B sky130_fd_sc_hd__o211ai_2
XFILLER_179_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5834_ _9574_/A hold25/X hold43/X VGND VGND VPWR VPWR _5834_/X sky130_fd_sc_hd__mux2_1
X_8622_ _8773_/Q _8304_/A _8354_/C _9080_/Q VGND VGND VPWR VPWR _8622_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5765_ hold553/X _5587_/X _5771_/S VGND VGND VPWR VPWR _5766_/A sky130_fd_sc_hd__mux2_1
X_8553_ _8553_/A0 _8552_/X _8653_/S VGND VGND VPWR VPWR _8554_/A sky130_fd_sc_hd__mux2_1
X_7504_ _7430_/X hold719/X _7515_/S VGND VGND VPWR VPWR _7505_/A sky130_fd_sc_hd__mux2_1
X_4716_ _8886_/Q _5573_/A _7032_/A _9124_/Q _4715_/X VGND VGND VPWR VPWR _4723_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8484_ _9332_/Q _8298_/X _8370_/X _9252_/Q _8483_/X VGND VGND VPWR VPWR _8487_/C
+ sky130_fd_sc_hd__a221o_1
X_5696_ _5633_/X hold466/X _5702_/S VGND VGND VPWR VPWR _5697_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7435_ _7435_/A VGND VGND VPWR VPWR _9299_/D sky130_fd_sc_hd__clkbuf_1
X_4647_ _9404_/Q _7661_/A _7144_/A _9554_/A VGND VGND VPWR VPWR _4647_/X sky130_fd_sc_hd__a22o_1
XFILLER_135_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold720 _9250_/Q VGND VGND VPWR VPWR hold720/X sky130_fd_sc_hd__dlygate4sd3_1
X_7366_ _7239_/X hold277/X _7372_/S VGND VGND VPWR VPWR _7366_/X sky130_fd_sc_hd__mux2_1
X_4578_ input17/X _4500_/Y _4575_/X _4577_/X VGND VGND VPWR VPWR _4578_/X sky130_fd_sc_hd__a211o_1
Xhold731 _7532_/X VGND VGND VPWR VPWR _7533_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 hold742/A VGND VGND VPWR VPWR hold742/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold753 _9091_/Q VGND VGND VPWR VPWR hold753/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9105_ _9551_/CLK _9105_/D _5929_/B VGND VGND VPWR VPWR hold98/A sky130_fd_sc_hd__dfrtp_4
X_6317_ _6317_/A _6317_/B VGND VGND VPWR VPWR _6672_/B sky130_fd_sc_hd__and2_1
Xhold764 hold764/A VGND VGND VPWR VPWR hold764/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold775 _4363_/X VGND VGND VPWR VPWR _4364_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7297_ _7279_/X hold798/X _7300_/S VGND VGND VPWR VPWR _7297_/X sky130_fd_sc_hd__mux2_1
Xhold786 _7245_/X VGND VGND VPWR VPWR _7246_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold797 _5438_/X VGND VGND VPWR VPWR _5439_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9036_ _9219_/CLK _9036_/D fanout467/X VGND VGND VPWR VPWR _9036_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_130_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6248_ _6248_/A _6794_/A _6248_/C VGND VGND VPWR VPWR _6250_/C sky130_fd_sc_hd__or3_1
XFILLER_130_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6179_ _6795_/A _6547_/A VGND VGND VPWR VPWR _6556_/B sky130_fd_sc_hd__nand2_2
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold80 hold80/A VGND VGND VPWR VPWR hold80/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold91 hold91/A VGND VGND VPWR VPWR hold91/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_90_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5550_ _5550_/A VGND VGND VPWR VPWR _8872_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4501_ hold60/X _4878_/A VGND VGND VPWR VPWR _4501_/Y sky130_fd_sc_hd__nor2_1
XFILLER_157_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5481_ _5481_/A VGND VGND VPWR VPWR _8842_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7220_ _6018_/X hold214/X _7226_/S VGND VGND VPWR VPWR _7220_/X sky130_fd_sc_hd__mux2_1
X_4432_ hold31/X _4432_/B VGND VGND VPWR VPWR hold32/A sky130_fd_sc_hd__or2_1
XFILLER_104_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7151_ _7151_/A VGND VGND VPWR VPWR _7151_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_160_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4363_ hold58/X hold82/X hold51/X VGND VGND VPWR VPWR _4363_/X sky130_fd_sc_hd__or3b_1
X_6102_ _6167_/C VGND VGND VPWR VPWR _6402_/A sky130_fd_sc_hd__buf_4
X_7082_ _9143_/Q _6048_/X hold65/X VGND VGND VPWR VPWR _7082_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6033_ hold898/X _5761_/X _6041_/S VGND VGND VPWR VPWR _6034_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7984_ _8206_/B _7991_/B _7984_/C VGND VGND VPWR VPWR _7984_/X sky130_fd_sc_hd__and3_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6935_ _6935_/A _6935_/B _6935_/C _6934_/X VGND VGND VPWR VPWR _7000_/B sky130_fd_sc_hd__or4b_2
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6866_ _6854_/X _6864_/X _6965_/A VGND VGND VPWR VPWR _6911_/B sky130_fd_sc_hd__o21ba_1
X_8605_ _8899_/Q _8312_/X _8376_/X _8949_/Q VGND VGND VPWR VPWR _8605_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5817_ _5817_/A VGND VGND VPWR VPWR _8987_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9585_ _9585_/A _5083_/Y VGND VGND VPWR VPWR mgmt_gpio_out[31] sky130_fd_sc_hd__ebufn_8
X_6797_ _6715_/B _6197_/B _6547_/B _6976_/B _6828_/A VGND VGND VPWR VPWR _6798_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_167_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5748_ _5748_/A VGND VGND VPWR VPWR _8957_/D sky130_fd_sc_hd__clkbuf_1
X_8536_ _9318_/Q _8372_/A _8369_/A _9326_/Q _8535_/X VGND VGND VPWR VPWR _8537_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_108_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5679_ hold918/X _5505_/X _5691_/S VGND VGND VPWR VPWR _5680_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8467_ _9211_/Q _8356_/A _8304_/X _9395_/Q VGND VGND VPWR VPWR _8473_/A sky130_fd_sc_hd__a22o_1
XFILLER_136_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7418_ _7418_/A VGND VGND VPWR VPWR _9292_/D sky130_fd_sc_hd__clkbuf_1
X_8398_ _8398_/A _8398_/B _8398_/C _8398_/D VGND VGND VPWR VPWR _8399_/A sky130_fd_sc_hd__or4_4
XFILLER_190_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold550 hold550/A VGND VGND VPWR VPWR _7125_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7349_ _7349_/A VGND VGND VPWR VPWR _9260_/D sky130_fd_sc_hd__clkbuf_1
Xhold561 _7309_/X VGND VGND VPWR VPWR _7310_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 _8915_/Q VGND VGND VPWR VPWR hold572/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold583 hold583/A VGND VGND VPWR VPWR hold583/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 hold594/A VGND VGND VPWR VPWR hold594/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9019_ _9475_/CLK _9019_/D fanout481/X VGND VGND VPWR VPWR _9580_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_131_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1250 _8898_/Q VGND VGND VPWR VPWR hold845/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1261 _8984_/Q VGND VGND VPWR VPWR hold526/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1272 _7124_/X VGND VGND VPWR VPWR hold550/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1283 _8886_/Q VGND VGND VPWR VPWR hold423/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_401 _7989_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput170 wb_dat_i[15] VGND VGND VPWR VPWR _8763_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput181 wb_dat_i[25] VGND VGND VPWR VPWR _8739_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput192 wb_dat_i[6] VGND VGND VPWR VPWR _8760_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4981_ _8801_/Q _5002_/B VGND VGND VPWR VPWR _4997_/B sky130_fd_sc_hd__and2_1
XFILLER_51_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6720_ _6719_/Y _6128_/X _6717_/Y _6619_/A VGND VGND VPWR VPWR _6944_/B sky130_fd_sc_hd__a31o_1
X_6651_ _6651_/A _6772_/A VGND VGND VPWR VPWR _6653_/A sky130_fd_sc_hd__nor2_1
XFILLER_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5602_ _5602_/A VGND VGND VPWR VPWR _8895_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6582_ _6987_/B _6956_/A _6582_/C _6582_/D VGND VGND VPWR VPWR _6583_/D sky130_fd_sc_hd__or4_1
X_9370_ _9370_/CLK _9370_/D fanout477/X VGND VGND VPWR VPWR _9370_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_118_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8321_ _8380_/A _8363_/A VGND VGND VPWR VPWR _8356_/B sky130_fd_sc_hd__nor2_2
X_5533_ _5533_/A VGND VGND VPWR VPWR _8864_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8252_ _8926_/Q _7933_/X _8020_/X _8946_/Q _8251_/X VGND VGND VPWR VPWR _8260_/A
+ sky130_fd_sc_hd__a221o_1
X_5464_ _5464_/A VGND VGND VPWR VPWR _8836_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_60_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _9161_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_133_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7203_ _6018_/X hold352/X _7209_/S VGND VGND VPWR VPWR _7203_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4415_ _4674_/A _4748_/B VGND VGND VPWR VPWR _7605_/A sky130_fd_sc_hd__nor2_8
X_8183_ _8858_/Q _7927_/A _7956_/A _8888_/Q _8182_/X VGND VGND VPWR VPWR _8184_/D
+ sky130_fd_sc_hd__a221o_1
X_5395_ _7645_/A VGND VGND VPWR VPWR _5395_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_99_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7134_ _7134_/A VGND VGND VPWR VPWR _9165_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7065_ hold79/X VGND VGND VPWR VPWR _9135_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_75_csclk _9359_/CLK VGND VGND VPWR VPWR _9288_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_86_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6016_ _6015_/X hold445/X _6019_/S VGND VGND VPWR VPWR _6016_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7967_ _7967_/A VGND VGND VPWR VPWR _7967_/X sky130_fd_sc_hd__buf_6
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6918_ _6918_/A _6918_/B _6918_/C VGND VGND VPWR VPWR _6918_/X sky130_fd_sc_hd__and3_1
X_7898_ _7904_/B _8389_/A VGND VGND VPWR VPWR _7898_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_13_csclk _9210_/CLK VGND VGND VPWR VPWR _9413_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_168_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6849_ _6715_/B _6673_/A _6195_/B _6597_/A _6733_/X VGND VGND VPWR VPWR _6950_/C
+ sky130_fd_sc_hd__a221o_1
X_9568_ _9568_/A _5100_/Y VGND VGND VPWR VPWR mgmt_gpio_out[14] sky130_fd_sc_hd__ebufn_8
XFILLER_167_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8519_ _9213_/Q _8289_/X _8341_/X _9309_/Q _8518_/X VGND VGND VPWR VPWR _8524_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_136_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9499_ _9501_/CLK _9499_/D fanout470/X VGND VGND VPWR VPWR _9499_/Q sky130_fd_sc_hd__dfrtp_2
Xclkbuf_leaf_28_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _9467_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_182_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold380 _7760_/X VGND VGND VPWR VPWR _7761_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 _5908_/X VGND VGND VPWR VPWR _5909_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1080 _5835_/X VGND VGND VPWR VPWR _8992_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1091 _7719_/X VGND VGND VPWR VPWR _7720_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_93_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_220 _9165_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_231 _9433_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_242 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_253 _5174_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_264 _5174_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_275 _5285_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_286 _4834_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_297 _5901_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer3 rebuffer3/A VGND VGND VPWR VPWR rebuffer3/X sky130_fd_sc_hd__buf_6
XFILLER_127_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5180_ _5180_/A VGND VGND VPWR VPWR _5180_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_142_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8870_ _9181_/CLK _8870_/D fanout486/X VGND VGND VPWR VPWR _8870_/Q sky130_fd_sc_hd__dfstp_2
X_7821_ _7821_/A VGND VGND VPWR VPWR _9474_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7752_ hold503/X _6048_/X _7762_/S VGND VGND VPWR VPWR _7752_/X sky130_fd_sc_hd__mux2_1
X_4964_ _4964_/A _4964_/B VGND VGND VPWR VPWR _4964_/Y sky130_fd_sc_hd__nor2_1
X_6703_ _6703_/A _6703_/B _6703_/C _6703_/D VGND VGND VPWR VPWR _6704_/D sky130_fd_sc_hd__or4_1
XFILLER_189_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4895_ _9192_/Q _7194_/A _7571_/A _9360_/Q VGND VGND VPWR VPWR _4896_/D sky130_fd_sc_hd__a22o_1
X_7683_ _7645_/X hold426/X _7693_/S VGND VGND VPWR VPWR _7683_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9422_ _9464_/CLK _9422_/D fanout421/X VGND VGND VPWR VPWR _9422_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6634_ _6818_/A _6632_/Y _6794_/B VGND VGND VPWR VPWR _6634_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_22_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9353_ _9427_/CLK _9353_/D fanout479/X VGND VGND VPWR VPWR _9353_/Q sky130_fd_sc_hd__dfstp_4
X_6565_ _6589_/C _6790_/C VGND VGND VPWR VPWR _6566_/B sky130_fd_sc_hd__nor2_2
X_8304_ _8304_/A VGND VGND VPWR VPWR _8304_/X sky130_fd_sc_hd__buf_6
X_5516_ _5516_/A VGND VGND VPWR VPWR _8857_/D sky130_fd_sc_hd__clkbuf_1
X_6496_ _6925_/A _6618_/B _6955_/C _6496_/D VGND VGND VPWR VPWR _6502_/B sky130_fd_sc_hd__or4_1
X_9284_ _9328_/CLK _9284_/D fanout463/X VGND VGND VPWR VPWR _9284_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_173_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5447_ _5447_/A VGND VGND VPWR VPWR _5447_/X sky130_fd_sc_hd__clkbuf_1
X_8235_ _8905_/Q _7962_/X _8077_/X _8935_/Q _8234_/X VGND VGND VPWR VPWR _8238_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_160_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5378_ _7011_/A _5378_/B VGND VGND VPWR VPWR _5379_/A sky130_fd_sc_hd__and2_1
X_8166_ _9263_/Q _7958_/A _7971_/A _9423_/Q VGND VGND VPWR VPWR _8166_/X sky130_fd_sc_hd__a22o_1
XFILLER_120_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7117_ _7117_/A VGND VGND VPWR VPWR _9158_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8097_ _8097_/A _8097_/B _8097_/C _8097_/D VGND VGND VPWR VPWR _8104_/B sky130_fd_sc_hd__or4_1
XFILLER_101_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7048_ _6012_/X _9128_/Q _7054_/S VGND VGND VPWR VPWR _7048_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8999_ _9532_/CLK _8999_/D fanout446/X VGND VGND VPWR VPWR _8999_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4680_ _9260_/Q _7339_/A _4906_/A2 _9436_/Q _4679_/X VGND VGND VPWR VPWR _4688_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_186_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6350_ _6345_/X _6230_/X _6346_/X _6347_/X _6349_/X VGND VGND VPWR VPWR _6352_/C
+ sky130_fd_sc_hd__a221o_1
X_5301_ _5951_/A VGND VGND VPWR VPWR _5301_/X sky130_fd_sc_hd__buf_6
XFILLER_115_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6281_ _6281_/A _6673_/A VGND VGND VPWR VPWR _6281_/Y sky130_fd_sc_hd__nand2_1
X_5232_ _9505_/Q _9158_/Q _9162_/Q VGND VGND VPWR VPWR _5233_/A sky130_fd_sc_hd__mux2_1
X_8020_ _8020_/A VGND VGND VPWR VPWR _8020_/X sky130_fd_sc_hd__buf_6
XFILLER_142_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5163_ hold994/X _8780_/Q _5017_/S _5016_/B _5021_/B VGND VGND VPWR VPWR _5163_/Y
+ sky130_fd_sc_hd__o32ai_1
XFILLER_111_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5094_ _9347_/Q VGND VGND VPWR VPWR _5094_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8922_ _9089_/CLK _8922_/D fanout433/X VGND VGND VPWR VPWR _8922_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_84_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8853_ _9184_/CLK _8853_/D fanout443/X VGND VGND VPWR VPWR _8853_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_25_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7804_ _7804_/A VGND VGND VPWR VPWR _9466_/D sky130_fd_sc_hd__clkbuf_1
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8784_ _5207_/A1 _8784_/D _5331_/X VGND VGND VPWR VPWR _8784_/Q sky130_fd_sc_hd__dfrtp_1
X_5996_ _5996_/A _7132_/B VGND VGND VPWR VPWR _6005_/S sky130_fd_sc_hd__and2_2
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7735_ _7735_/A VGND VGND VPWR VPWR _9434_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4947_ input52/X _5901_/A _5642_/A _8913_/Q VGND VGND VPWR VPWR _4947_/X sky130_fd_sc_hd__a22o_1
X_7666_ _7645_/X hold414/X _7676_/S VGND VGND VPWR VPWR _7666_/X sky130_fd_sc_hd__mux2_1
X_4878_ _4878_/A _7111_/B VGND VGND VPWR VPWR _7027_/A sky130_fd_sc_hd__nor2_2
X_9405_ _9469_/CLK _9405_/D fanout458/X VGND VGND VPWR VPWR _9405_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6617_ _6850_/B _6428_/B _6597_/Y _6266_/X VGND VGND VPWR VPWR _6618_/D sky130_fd_sc_hd__o31ai_1
X_7597_ _7436_/X hold270/X hold75/X VGND VGND VPWR VPWR _7598_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9336_ _9398_/CLK _9336_/D _5070_/A VGND VGND VPWR VPWR _9336_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_165_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6548_ _6790_/A _6793_/B VGND VGND VPWR VPWR _6956_/A sky130_fd_sc_hd__nor2_1
XFILLER_106_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9267_ _9283_/CLK _9267_/D fanout484/X VGND VGND VPWR VPWR _9267_/Q sky130_fd_sc_hd__dfrtp_4
X_6479_ _6479_/A _6736_/B VGND VGND VPWR VPWR _6859_/B sky130_fd_sc_hd__nor2_1
XFILLER_161_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8218_ _5139_/A _9515_/Q _8013_/X VGND VGND VPWR VPWR _8218_/X sky130_fd_sc_hd__a21o_1
XFILLER_121_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput260 _9129_/Q VGND VGND VPWR VPWR pll90_sel[0] sky130_fd_sc_hd__buf_12
Xoutput271 _9126_/Q VGND VGND VPWR VPWR pll_sel[0] sky130_fd_sc_hd__buf_12
X_9198_ _9437_/CLK _9198_/D fanout409/X VGND VGND VPWR VPWR _9198_/Q sky130_fd_sc_hd__dfrtp_2
Xoutput282 _9133_/Q VGND VGND VPWR VPWR pll_trim[17] sky130_fd_sc_hd__buf_12
Xoutput293 _8820_/Q VGND VGND VPWR VPWR pll_trim[3] sky130_fd_sc_hd__buf_12
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8149_ _8149_/A _8149_/B _8149_/C _8149_/D VGND VGND VPWR VPWR _8149_/X sky130_fd_sc_hd__or4_4
XFILLER_87_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5850_ _9001_/Q hold38/X _5868_/S VGND VGND VPWR VPWR _5850_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4801_ _9434_/Q _4906_/A2 _5493_/A _8850_/Q _4800_/X VGND VGND VPWR VPWR _4806_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5781_ _5781_/A VGND VGND VPWR VPWR _8971_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7520_ _7517_/X hold925/X _7534_/S VGND VGND VPWR VPWR _7521_/A sky130_fd_sc_hd__mux2_1
X_4732_ _9451_/Q _4836_/A2 _7056_/A _9135_/Q VGND VGND VPWR VPWR _4732_/X sky130_fd_sc_hd__a22o_1
XFILLER_187_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4663_ _8902_/Q _5607_/A _5493_/A _8852_/Q _4662_/X VGND VGND VPWR VPWR _4673_/B
+ sky130_fd_sc_hd__a221o_1
X_7451_ _7430_/X hold706/X _7461_/S VGND VGND VPWR VPWR _7452_/A sky130_fd_sc_hd__mux2_1
X_6402_ _6402_/A _6440_/A VGND VGND VPWR VPWR _6482_/A sky130_fd_sc_hd__or2_1
X_4594_ _4594_/A VGND VGND VPWR VPWR _9116_/D sky130_fd_sc_hd__clkbuf_1
X_7382_ _7382_/A VGND VGND VPWR VPWR _9275_/D sky130_fd_sc_hd__clkbuf_1
Xhold902 _9416_/Q VGND VGND VPWR VPWR hold902/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 hold913/A VGND VGND VPWR VPWR hold913/X sky130_fd_sc_hd__dlygate4sd3_1
X_9121_ _9485_/CLK _9121_/D fanout404/X VGND VGND VPWR VPWR _9121_/Q sky130_fd_sc_hd__dfrtp_2
Xhold924 _9392_/Q VGND VGND VPWR VPWR hold924/X sky130_fd_sc_hd__dlygate4sd3_1
X_6333_ _6334_/B _6871_/B VGND VGND VPWR VPWR _6872_/B sky130_fd_sc_hd__nor2_1
XFILLER_115_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold935 _9400_/Q VGND VGND VPWR VPWR hold935/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 _9520_/Q VGND VGND VPWR VPWR hold946/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 _4754_/X VGND VGND VPWR VPWR _4755_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 _9522_/Q VGND VGND VPWR VPWR hold968/X sky130_fd_sc_hd__dlygate4sd3_1
X_9052_ _9187_/CLK _9052_/D fanout450/X VGND VGND VPWR VPWR _9052_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_103_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6264_ _6802_/A _6610_/A VGND VGND VPWR VPWR _7002_/A sky130_fd_sc_hd__nor2_1
Xhold979 _8219_/X VGND VGND VPWR VPWR _9516_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5215_ _5214_/X _5181_/B _8794_/Q VGND VGND VPWR VPWR _5216_/A sky130_fd_sc_hd__mux2_4
X_8003_ _8003_/A VGND VGND VPWR VPWR _8003_/X sky130_fd_sc_hd__buf_6
XFILLER_69_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6195_ _6609_/A _6195_/B VGND VGND VPWR VPWR _6195_/Y sky130_fd_sc_hd__nand2_1
XFILLER_130_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5146_ _9034_/Q VGND VGND VPWR VPWR _5287_/A sky130_fd_sc_hd__buf_2
XFILLER_69_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5077_ _5068_/B _8780_/Q _5025_/B VGND VGND VPWR VPWR _5077_/X sky130_fd_sc_hd__a21o_1
XFILLER_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8905_ _9442_/CLK _8905_/D fanout436/X VGND VGND VPWR VPWR _8905_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_84_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8836_ _9427_/CLK _8836_/D fanout477/X VGND VGND VPWR VPWR _8836_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_44_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8767_ _8767_/A1 _5870_/X _8735_/A _5149_/Y VGND VGND VPWR VPWR _9550_/D sky130_fd_sc_hd__o211a_2
X_5979_ _5979_/A VGND VGND VPWR VPWR _5994_/S sky130_fd_sc_hd__buf_2
XFILLER_12_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7718_ _7718_/A VGND VGND VPWR VPWR _9426_/D sky130_fd_sc_hd__clkbuf_1
X_8698_ _8776_/Q _8304_/X _8324_/X _9083_/Q VGND VGND VPWR VPWR _8698_/X sky130_fd_sc_hd__a22o_1
XFILLER_60_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7649_ _7648_/X _9395_/Q hold84/X VGND VGND VPWR VPWR _7649_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9319_ _9376_/CLK _9319_/D fanout425/X VGND VGND VPWR VPWR _9319_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_153_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold209 _9447_/Q VGND VGND VPWR VPWR hold209/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_125_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _4999_/X _5000_/A1 _5014_/S VGND VGND VPWR VPWR _5001_/A sky130_fd_sc_hd__mux2_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6951_ _6994_/B _6951_/B _6964_/D _6965_/B VGND VGND VPWR VPWR _6951_/X sky130_fd_sc_hd__or4_1
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5902_ _5629_/X _9578_/A _5916_/S VGND VGND VPWR VPWR _5902_/X sky130_fd_sc_hd__mux2_1
XFILLER_81_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6882_ _6882_/A _6882_/B _6882_/C _6882_/D VGND VGND VPWR VPWR _7003_/A sky130_fd_sc_hd__or4_1
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8621_ _8974_/Q _8337_/A _8384_/A _8854_/Q _8620_/X VGND VGND VPWR VPWR _8624_/C
+ sky130_fd_sc_hd__a221o_1
X_5833_ _8836_/Q hold24/X _5842_/S VGND VGND VPWR VPWR hold25/A sky130_fd_sc_hd__mux2_1
XFILLER_34_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8552_ _8997_/Q _9525_/Q _8550_/X _8551_/X VGND VGND VPWR VPWR _8552_/X sky130_fd_sc_hd__a22o_1
X_5764_ _5764_/A VGND VGND VPWR VPWR _8963_/D sky130_fd_sc_hd__clkbuf_1
X_7503_ _7503_/A VGND VGND VPWR VPWR _9329_/D sky130_fd_sc_hd__clkbuf_1
X_4715_ input55/X _5901_/A _7588_/A _9371_/Q VGND VGND VPWR VPWR _4715_/X sky130_fd_sc_hd__a22o_2
X_8483_ _9452_/Q _8310_/X _8381_/X _9364_/Q VGND VGND VPWR VPWR _8483_/X sky130_fd_sc_hd__a22o_1
X_5695_ _5695_/A VGND VGND VPWR VPWR _8933_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7434_ _7433_/X _9299_/Q _7444_/S VGND VGND VPWR VPWR _7434_/X sky130_fd_sc_hd__mux2_1
X_4646_ _4667_/A _7158_/B VGND VGND VPWR VPWR _6032_/A sky130_fd_sc_hd__nor2_4
XFILLER_107_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold710 hold710/A VGND VGND VPWR VPWR hold710/X sky130_fd_sc_hd__dlygate4sd3_1
X_4577_ input57/X _5901_/A _7266_/A _9229_/Q _4576_/X VGND VGND VPWR VPWR _4577_/X
+ sky130_fd_sc_hd__a221o_2
Xhold721 _7327_/X VGND VGND VPWR VPWR _7328_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7365_ _7365_/A VGND VGND VPWR VPWR _9267_/D sky130_fd_sc_hd__clkbuf_1
Xhold732 hold732/A VGND VGND VPWR VPWR hold732/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9104_ _9551_/CLK _9104_/D _5929_/B VGND VGND VPWR VPWR hold85/A sky130_fd_sc_hd__dfrtp_4
Xhold743 _9186_/Q VGND VGND VPWR VPWR hold743/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold754 _9326_/Q VGND VGND VPWR VPWR hold754/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6316_ _6324_/A _6828_/A VGND VGND VPWR VPWR _6839_/B sky130_fd_sc_hd__nor2_4
Xhold765 _9230_/Q VGND VGND VPWR VPWR hold765/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold776 _7037_/X VGND VGND VPWR VPWR _7038_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7296_ _7296_/A VGND VGND VPWR VPWR _9237_/D sky130_fd_sc_hd__clkbuf_1
Xhold787 hold787/A VGND VGND VPWR VPWR hold787/X sky130_fd_sc_hd__dlygate4sd3_1
X_9035_ _9434_/CLK _9035_/D fanout450/X VGND VGND VPWR VPWR _9035_/Q sky130_fd_sc_hd__dfrtp_2
Xhold798 _9238_/Q VGND VGND VPWR VPWR hold798/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6247_ _6244_/X _6610_/B _6628_/A _6249_/A VGND VGND VPWR VPWR _6248_/C sky130_fd_sc_hd__a211o_1
XFILLER_103_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6178_ _6178_/A _6178_/B _6232_/C VGND VGND VPWR VPWR _6547_/A sky130_fd_sc_hd__and3_1
XFILLER_29_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5129_ _8997_/Q VGND VGND VPWR VPWR _5130_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_84_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8819_ _9476_/CLK _8819_/D fanout414/X VGND VGND VPWR VPWR _8819_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_13_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold70 hold70/A VGND VGND VPWR VPWR hold70/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 hold81/A VGND VGND VPWR VPWR hold81/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold92 hold92/A VGND VGND VPWR VPWR hold92/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4500_ _7111_/B _4685_/B VGND VGND VPWR VPWR _4500_/Y sky130_fd_sc_hd__nor2_8
XFILLER_129_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5480_ _5306_/X hold506/X _5490_/S VGND VGND VPWR VPWR _5480_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1 _5826_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4431_ _4431_/A _4431_/B _4431_/C _4431_/D VGND VGND VPWR VPWR _4507_/A sky130_fd_sc_hd__or4_1
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7150_ _6012_/X _9588_/A _7156_/S VGND VGND VPWR VPWR _7150_/X sky130_fd_sc_hd__mux2_1
X_4362_ hold50/X hold857/X hold73/X VGND VGND VPWR VPWR hold51/A sky130_fd_sc_hd__mux2_1
XFILLER_172_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6101_ _6101_/A VGND VGND VPWR VPWR _6479_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_112_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7081_ _7081_/A VGND VGND VPWR VPWR _7081_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_59_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6032_ _6032_/A _7132_/B VGND VGND VPWR VPWR _6041_/S sky130_fd_sc_hd__and2_2
XFILLER_113_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7983_ _7983_/A VGND VGND VPWR VPWR _8008_/B sky130_fd_sc_hd__buf_8
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6934_ _6873_/B _6799_/A _6871_/B _7001_/B VGND VGND VPWR VPWR _6934_/X sky130_fd_sc_hd__o22a_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6865_ _6865_/A _6865_/B VGND VGND VPWR VPWR _6965_/A sky130_fd_sc_hd__or2_1
XFILLER_179_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8604_ hold959/X _8017_/X _8603_/X VGND VGND VPWR VPWR _8604_/X sky130_fd_sc_hd__o21a_1
X_5816_ hold648/X _5690_/X _5816_/S VGND VGND VPWR VPWR _5817_/A sky130_fd_sc_hd__mux2_1
X_9584_ _9584_/A _5084_/Y VGND VGND VPWR VPWR mgmt_gpio_out[30] sky130_fd_sc_hd__ebufn_8
X_6796_ _6794_/Y _6343_/C _6560_/B _6960_/B VGND VGND VPWR VPWR _6880_/A sky130_fd_sc_hd__a211o_1
XFILLER_179_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8535_ _9302_/Q _8354_/B _8331_/A _9406_/Q VGND VGND VPWR VPWR _8535_/X sky130_fd_sc_hd__a22o_1
X_5747_ _5653_/X hold336/X _5747_/S VGND VGND VPWR VPWR _5747_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8466_ _9235_/Q _8322_/X _8333_/X _9267_/Q _8465_/X VGND VGND VPWR VPWR _8474_/C
+ sky130_fd_sc_hd__a221o_1
X_5678_ _5678_/A _5715_/B VGND VGND VPWR VPWR _5691_/S sky130_fd_sc_hd__and2_2
XFILLER_175_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7417_ _7239_/X hold259/X _7423_/S VGND VGND VPWR VPWR _7417_/X sky130_fd_sc_hd__mux2_1
X_4629_ _4635_/A _4667_/B VGND VGND VPWR VPWR _5750_/A sky130_fd_sc_hd__nor2_8
XFILLER_190_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8397_ _8397_/A _8397_/B _8397_/C VGND VGND VPWR VPWR _8397_/X sky130_fd_sc_hd__or3_2
XFILLER_123_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold540 _8875_/Q VGND VGND VPWR VPWR hold540/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 _9086_/Q VGND VGND VPWR VPWR hold551/X sky130_fd_sc_hd__dlygate4sd3_1
X_7348_ _7239_/X hold314/X _7354_/S VGND VGND VPWR VPWR _7348_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold562 _9239_/Q VGND VGND VPWR VPWR hold562/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 hold573/A VGND VGND VPWR VPWR hold573/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold584 _9375_/Q VGND VGND VPWR VPWR hold584/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 _9351_/Q VGND VGND VPWR VPWR hold595/X sky130_fd_sc_hd__dlygate4sd3_1
X_7279_ _7494_/A VGND VGND VPWR VPWR _7279_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_77_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9018_ _9475_/CLK _9018_/D fanout481/X VGND VGND VPWR VPWR _9579_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1240 _7434_/X VGND VGND VPWR VPWR hold355/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1251 _8873_/Q VGND VGND VPWR VPWR hold899/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1262 _8939_/Q VGND VGND VPWR VPWR hold583/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1273 _8933_/Q VGND VGND VPWR VPWR hold872/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1284 _7184_/X VGND VGND VPWR VPWR hold203/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_402 _8002_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput160 wb_adr_i[7] VGND VGND VPWR VPWR _6182_/A sky130_fd_sc_hd__buf_2
XFILLER_49_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput171 wb_dat_i[16] VGND VGND VPWR VPWR _8728_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput182 wb_dat_i[26] VGND VGND VPWR VPWR _8743_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput193 wb_dat_i[7] VGND VGND VPWR VPWR _8764_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4980_ hold39/A hold8/A hold76/A VGND VGND VPWR VPWR _5002_/B sky130_fd_sc_hd__and3_1
XFILLER_51_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6650_ _6748_/B _6658_/A VGND VGND VPWR VPWR _6738_/A sky130_fd_sc_hd__nor2_1
XFILLER_176_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5601_ hold638/X _5395_/X _5605_/S VGND VGND VPWR VPWR _5602_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6581_ _6673_/A _6551_/Y _6959_/C _6579_/X _6580_/X VGND VGND VPWR VPWR _6582_/D
+ sky130_fd_sc_hd__a2111o_1
X_8320_ _8320_/A VGND VGND VPWR VPWR _8363_/A sky130_fd_sc_hd__buf_2
X_5532_ _5301_/X hold495/X _5538_/S VGND VGND VPWR VPWR _5533_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8251_ _8876_/Q _7953_/B _7973_/X _8856_/Q VGND VGND VPWR VPWR _8251_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_9_csclk _9359_/CLK VGND VGND VPWR VPWR _9416_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_145_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5463_ _5315_/X hold110/X _5472_/S VGND VGND VPWR VPWR _5463_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7202_ _7202_/A VGND VGND VPWR VPWR _9195_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4414_ _4674_/A _4858_/B VGND VGND VPWR VPWR _4414_/Y sky130_fd_sc_hd__nor2_8
X_8182_ _8772_/Q _7977_/A _8181_/X _7983_/A VGND VGND VPWR VPWR _8182_/X sky130_fd_sc_hd__a22o_1
X_5394_ _5394_/A VGND VGND VPWR VPWR _8810_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7133_ _9165_/Q _6048_/X _7137_/S VGND VGND VPWR VPWR _7133_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7064_ _9135_/Q hold46/X _7072_/S VGND VGND VPWR VPWR hold79/A sky130_fd_sc_hd__mux2_1
XFILLER_113_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6015_ _7648_/A VGND VGND VPWR VPWR _6015_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7966_ _7998_/A _7991_/B _8002_/C VGND VGND VPWR VPWR _7967_/A sky130_fd_sc_hd__and3_2
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6917_ _6976_/C _6917_/B _6917_/C _6917_/D VGND VGND VPWR VPWR _6918_/C sky130_fd_sc_hd__and4b_1
X_7897_ _9500_/Q _9499_/Q VGND VGND VPWR VPWR _8389_/A sky130_fd_sc_hd__and2_2
XFILLER_52_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6848_ _6897_/A _6609_/A _6195_/B VGND VGND VPWR VPWR _6950_/B sky130_fd_sc_hd__o21a_1
XFILLER_167_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_494 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9567_ _9567_/A _5101_/Y VGND VGND VPWR VPWR mgmt_gpio_out[13] sky130_fd_sc_hd__ebufn_8
X_6779_ _6779_/A _6781_/C _6779_/C VGND VGND VPWR VPWR _6779_/X sky130_fd_sc_hd__or3_1
XFILLER_183_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8518_ _9397_/Q _8304_/X _8324_/X _9245_/Q VGND VGND VPWR VPWR _8518_/X sky130_fd_sc_hd__a22o_1
XFILLER_182_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9498_ _9501_/CLK _9498_/D fanout488/X VGND VGND VPWR VPWR _9498_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_136_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8449_ _8449_/A _8449_/B _8449_/C _8449_/D VGND VGND VPWR VPWR _8450_/C sky130_fd_sc_hd__or4_1
XFILLER_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold370 hold370/A VGND VGND VPWR VPWR hold370/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold381 hold381/A VGND VGND VPWR VPWR hold381/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 _5909_/X VGND VGND VPWR VPWR _9020_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1070 _5863_/X VGND VGND VPWR VPWR _9005_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_93_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1081 _5831_/X VGND VGND VPWR VPWR _5832_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1092 _8932_/Q VGND VGND VPWR VPWR hold516/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_210 _8682_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_221 _9187_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_232 _9467_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_243 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_254 _5174_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_265 _5174_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_276 _5285_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_287 _4951_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_298 _5901_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7820_ _7645_/X hold496/X _7830_/S VGND VGND VPWR VPWR _7820_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7751_ _7751_/A VGND VGND VPWR VPWR _9441_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4963_ _8808_/Q _8807_/Q _5068_/B VGND VGND VPWR VPWR _4964_/A sky130_fd_sc_hd__or3_1
X_6702_ _6419_/A _6503_/A _6441_/B _7002_/B VGND VGND VPWR VPWR _6703_/D sky130_fd_sc_hd__a31o_1
XFILLER_177_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7682_ hold97/X VGND VGND VPWR VPWR _9409_/D sky130_fd_sc_hd__clkbuf_1
X_4894_ _9264_/Q _7356_/A _5562_/A _8878_/Q VGND VGND VPWR VPWR _4896_/C sky130_fd_sc_hd__a22o_1
XFILLER_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9421_ _9421_/CLK _9421_/D fanout461/X VGND VGND VPWR VPWR _9421_/Q sky130_fd_sc_hd__dfrtp_1
X_6633_ _6633_/A _6811_/B VGND VGND VPWR VPWR _6794_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9352_ _9416_/CLK _9352_/D fanout425/X VGND VGND VPWR VPWR _9352_/Q sky130_fd_sc_hd__dfstp_2
X_6564_ _6839_/A VGND VGND VPWR VPWR _6790_/C sky130_fd_sc_hd__inv_2
XFILLER_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8303_ _8375_/A _8398_/A _8357_/B VGND VGND VPWR VPWR _8304_/A sky130_fd_sc_hd__and3_2
X_5515_ hold607/X _5402_/X _5515_/S VGND VGND VPWR VPWR _5515_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9283_ _9283_/CLK _9283_/D fanout473/X VGND VGND VPWR VPWR _9283_/Q sky130_fd_sc_hd__dfrtp_4
X_6495_ _6651_/A _6495_/B VGND VGND VPWR VPWR _6496_/D sky130_fd_sc_hd__nor2_1
XFILLER_106_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8234_ _8875_/Q _7953_/B _8003_/X _8885_/Q VGND VGND VPWR VPWR _8234_/X sky130_fd_sc_hd__a22o_1
XFILLER_172_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5446_ _7011_/A _7013_/B VGND VGND VPWR VPWR _5447_/A sky130_fd_sc_hd__and2_1
XFILLER_172_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8165_ _9231_/Q _7979_/X _7993_/A _9391_/Q VGND VGND VPWR VPWR _8165_/X sky130_fd_sc_hd__a22o_1
X_5377_ _7025_/A VGND VGND VPWR VPWR _7011_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_154_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7116_ _6015_/X _9158_/Q _7124_/S VGND VGND VPWR VPWR _7116_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8096_ _9220_/Q _7927_/X _8023_/B _9308_/Q _8095_/X VGND VGND VPWR VPWR _8097_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_141_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7047_ _7047_/A VGND VGND VPWR VPWR _9127_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8998_ _9531_/CLK _8998_/D fanout446/X VGND VGND VPWR VPWR _8998_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7949_ _7949_/A VGND VGND VPWR VPWR _7949_/X sky130_fd_sc_hd__buf_6
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_74_csclk _9359_/CLK VGND VGND VPWR VPWR _9392_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_147_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5300_ hold37/X VGND VGND VPWR VPWR _5951_/A sky130_fd_sc_hd__buf_6
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6280_ _6556_/B _6558_/C VGND VGND VPWR VPWR _6673_/A sky130_fd_sc_hd__nor2_2
XFILLER_154_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5231_ _5231_/A VGND VGND VPWR VPWR _5231_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5162_ _5162_/A VGND VGND VPWR VPWR _8997_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_csclk _9210_/CLK VGND VGND VPWR VPWR _9469_/CLK sky130_fd_sc_hd__clkbuf_16
X_5093_ _9355_/Q VGND VGND VPWR VPWR _5093_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8921_ _9084_/CLK _8921_/D fanout444/X VGND VGND VPWR VPWR _8921_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_37_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8852_ _8852_/CLK _8852_/D fanout444/X VGND VGND VPWR VPWR _8852_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_27_csclk _9303_/CLK VGND VGND VPWR VPWR _9466_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7803_ _7645_/X hold725/X _7813_/S VGND VGND VPWR VPWR _7804_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8783_ _5207_/A1 _8783_/D _5329_/X VGND VGND VPWR VPWR hold44/A sky130_fd_sc_hd__dfrtp_1
X_5995_ _5995_/A VGND VGND VPWR VPWR _9068_/D sky130_fd_sc_hd__clkbuf_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7734_ _7645_/X hold737/X hold86/X VGND VGND VPWR VPWR _7735_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4946_ input11/X _4500_/Y _7113_/A _9506_/Q _4945_/X VGND VGND VPWR VPWR _4949_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7665_ hold93/X VGND VGND VPWR VPWR _9401_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4877_ _9329_/Q _7499_/A _5551_/A _8874_/Q _4876_/X VGND VGND VPWR VPWR _4883_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_165_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9404_ _9420_/CLK _9404_/D fanout465/X VGND VGND VPWR VPWR _9404_/Q sky130_fd_sc_hd__dfrtp_4
X_6616_ _6851_/C _6616_/B _6616_/C _6616_/D VGND VGND VPWR VPWR _6618_/C sky130_fd_sc_hd__or4_1
X_7596_ _7596_/A VGND VGND VPWR VPWR _9371_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9335_ _9367_/CLK _9335_/D fanout422/X VGND VGND VPWR VPWR _9335_/Q sky130_fd_sc_hd__dfrtp_1
X_6547_ _6547_/A _6547_/B VGND VGND VPWR VPWR _6793_/B sky130_fd_sc_hd__nand2_1
XFILLER_192_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9266_ _9466_/CLK _9266_/D fanout472/X VGND VGND VPWR VPWR _9266_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_145_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6478_ _6839_/B _6672_/C _6478_/C VGND VGND VPWR VPWR _6483_/B sky130_fd_sc_hd__and3_1
XFILLER_161_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8217_ _8849_/Q _8010_/B _8216_/X _8105_/X VGND VGND VPWR VPWR _8217_/X sky130_fd_sc_hd__o211a_1
X_5429_ _5429_/A VGND VGND VPWR VPWR _8821_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput250 _5169_/X VGND VGND VPWR VPWR pad_flash_clk sky130_fd_sc_hd__clkbuf_1
X_9197_ _9469_/CLK _9197_/D fanout458/X VGND VGND VPWR VPWR _9197_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput261 _9130_/Q VGND VGND VPWR VPWR pll90_sel[1] sky130_fd_sc_hd__buf_12
Xoutput272 _9127_/Q VGND VGND VPWR VPWR pll_sel[1] sky130_fd_sc_hd__buf_12
Xoutput283 _9134_/Q VGND VGND VPWR VPWR pll_trim[18] sky130_fd_sc_hd__buf_12
Xoutput294 _8821_/Q VGND VGND VPWR VPWR pll_trim[4] sky130_fd_sc_hd__buf_12
XFILLER_58_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8148_ _9358_/Q _8020_/X _7990_/X _9278_/Q _8147_/X VGND VGND VPWR VPWR _8149_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_102_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8079_ _9259_/Q _7958_/X _8077_/X _9347_/Q _8078_/X VGND VGND VPWR VPWR _8082_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_1_wb_clk_i clkbuf_1_1_1_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__buf_8
XFILLER_124_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4800_ _9134_/Q _7056_/A _5630_/A _8910_/Q VGND VGND VPWR VPWR _4800_/X sky130_fd_sc_hd__a22o_1
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5780_ _5650_/X hold404/X _5782_/S VGND VGND VPWR VPWR _5781_/A sky130_fd_sc_hd__mux2_1
XFILLER_187_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4731_ _4731_/A _4731_/B _4731_/C _4731_/D VGND VGND VPWR VPWR _4752_/B sky130_fd_sc_hd__or4_1
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7450_ _7450_/A VGND VGND VPWR VPWR _9305_/D sky130_fd_sc_hd__clkbuf_1
X_4662_ _8813_/Q _5388_/A _5596_/A _8897_/Q VGND VGND VPWR VPWR _4662_/X sky130_fd_sc_hd__a22o_1
XFILLER_135_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6401_ _6401_/A VGND VGND VPWR VPWR _6967_/B sky130_fd_sc_hd__buf_4
X_7381_ _7236_/X _9275_/Q _7389_/S VGND VGND VPWR VPWR _7381_/X sky130_fd_sc_hd__mux2_1
X_4593_ _4592_/X hold972/X _4964_/B VGND VGND VPWR VPWR _4593_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold903 hold903/A VGND VGND VPWR VPWR hold903/X sky130_fd_sc_hd__dlygate4sd3_1
X_9120_ _9456_/CLK _9120_/D fanout404/X VGND VGND VPWR VPWR _9120_/Q sky130_fd_sc_hd__dfstp_1
X_6332_ _6802_/A _6874_/A VGND VGND VPWR VPWR _6758_/A sky130_fd_sc_hd__nor2_1
Xhold914 _9296_/Q VGND VGND VPWR VPWR hold914/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 _9336_/Q VGND VGND VPWR VPWR hold925/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 _9456_/Q VGND VGND VPWR VPWR hold936/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold947 _9508_/Q VGND VGND VPWR VPWR hold947/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 _9029_/Q VGND VGND VPWR VPWR _5870_/C sky130_fd_sc_hd__dlygate4sd3_1
X_9051_ _9051_/CLK _9051_/D fanout453/X VGND VGND VPWR VPWR _9051_/Q sky130_fd_sc_hd__dfrtp_1
Xhold969 _8453_/X VGND VGND VPWR VPWR _9522_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6263_ _6263_/A VGND VGND VPWR VPWR _6802_/A sky130_fd_sc_hd__buf_2
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8002_ _8181_/B _8002_/B _8002_/C VGND VGND VPWR VPWR _8003_/A sky130_fd_sc_hd__and3_1
X_5214_ _5213_/X input38/X _8796_/Q VGND VGND VPWR VPWR _5214_/X sky130_fd_sc_hd__mux2_1
X_6194_ _6228_/A _6194_/B VGND VGND VPWR VPWR _6195_/B sky130_fd_sc_hd__nor2_2
XFILLER_69_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5145_ _5275_/A _5115_/X _5870_/D VGND VGND VPWR VPWR _9033_/D sky130_fd_sc_hd__a21o_1
XFILLER_84_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5076_ _5076_/A VGND VGND VPWR VPWR _5076_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8904_ _9184_/CLK _8904_/D fanout438/X VGND VGND VPWR VPWR _8904_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8835_ _9172_/CLK _8835_/D fanout494/X VGND VGND VPWR VPWR _8835_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8766_ _8766_/A VGND VGND VPWR VPWR _9549_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5978_ _9028_/Q _8709_/B VGND VGND VPWR VPWR _5979_/A sky130_fd_sc_hd__and2_2
XFILLER_12_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7717_ _7645_/X hold418/X hold95/X VGND VGND VPWR VPWR _7718_/A sky130_fd_sc_hd__mux2_1
X_4929_ _9376_/Q _7605_/A _5518_/A _8858_/Q VGND VGND VPWR VPWR _4929_/X sky130_fd_sc_hd__a22o_1
X_8697_ _8977_/Q _8337_/X _8384_/X _8857_/Q _8696_/X VGND VGND VPWR VPWR _8700_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_166_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7648_ _7648_/A VGND VGND VPWR VPWR _7648_/X sky130_fd_sc_hd__buf_2
XFILLER_165_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7579_ _7579_/A VGND VGND VPWR VPWR _9363_/D sky130_fd_sc_hd__clkbuf_1
X_9318_ _9486_/CLK _9318_/D fanout413/X VGND VGND VPWR VPWR _9318_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_4_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9249_ _9449_/CLK _9249_/D fanout474/X VGND VGND VPWR VPWR _9249_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_69_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6950_ _6950_/A _6950_/B _6950_/C _6950_/D VGND VGND VPWR VPWR _6965_/B sky130_fd_sc_hd__or4_1
XFILLER_66_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5901_ _5901_/A _7284_/B VGND VGND VPWR VPWR _5916_/S sky130_fd_sc_hd__nand2_4
X_6881_ _6881_/A _7001_/B VGND VGND VPWR VPWR _6882_/D sky130_fd_sc_hd__nor2_1
XFILLER_62_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8620_ _8939_/Q _7908_/A _8358_/C _8869_/Q VGND VGND VPWR VPWR _8620_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5832_ _5832_/A VGND VGND VPWR VPWR _5832_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8551_ _9190_/Q _8400_/B _8652_/S VGND VGND VPWR VPWR _8551_/X sky130_fd_sc_hd__o21a_1
X_5763_ hold892/X _5761_/X _5771_/S VGND VGND VPWR VPWR _5764_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7502_ _7359_/X hold127/X _7515_/S VGND VGND VPWR VPWR _7502_/X sky130_fd_sc_hd__mux2_1
X_4714_ _8921_/Q _5656_/A _5529_/A _8866_/Q _4713_/X VGND VGND VPWR VPWR _4724_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_147_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8482_ _9372_/Q _8346_/X _8386_/X _9348_/Q _8481_/X VGND VGND VPWR VPWR _8487_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_175_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5694_ _5629_/X hold872/X _5702_/S VGND VGND VPWR VPWR _5695_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7433_ _7648_/A VGND VGND VPWR VPWR _7433_/X sky130_fd_sc_hd__clkbuf_2
X_4645_ _4665_/A _4956_/A VGND VGND VPWR VPWR _5738_/A sky130_fd_sc_hd__nor2_8
XFILLER_147_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold700 _9195_/Q VGND VGND VPWR VPWR hold700/X sky130_fd_sc_hd__dlygate4sd3_1
X_7364_ _7236_/X _9267_/Q _7372_/S VGND VGND VPWR VPWR _7364_/X sky130_fd_sc_hd__mux2_1
Xhold711 hold711/A VGND VGND VPWR VPWR hold711/X sky130_fd_sc_hd__dlygate4sd3_1
X_4576_ _9197_/Q _7194_/A _7356_/A _9269_/Q VGND VGND VPWR VPWR _4576_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold722 hold722/A VGND VGND VPWR VPWR hold722/X sky130_fd_sc_hd__dlygate4sd3_1
X_9103_ _9473_/CLK _9103_/D fanout431/X VGND VGND VPWR VPWR _9103_/Q sky130_fd_sc_hd__dfrtp_4
Xhold733 _9294_/Q VGND VGND VPWR VPWR hold733/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 _7182_/X VGND VGND VPWR VPWR _7183_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6315_ _6800_/A VGND VGND VPWR VPWR _6315_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold755 _7495_/X VGND VGND VPWR VPWR _7496_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7295_ _7242_/X hold218/X _7300_/S VGND VGND VPWR VPWR _7295_/X sky130_fd_sc_hd__mux2_1
Xhold766 _7280_/X VGND VGND VPWR VPWR _7281_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 hold777/A VGND VGND VPWR VPWR hold777/X sky130_fd_sc_hd__dlygate4sd3_1
X_9034_ _9551_/CLK _9034_/D fanout499/X VGND VGND VPWR VPWR _9034_/Q sky130_fd_sc_hd__dfrtp_4
Xhold788 _8880_/Q VGND VGND VPWR VPWR hold788/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold799 _7297_/X VGND VGND VPWR VPWR _7298_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6246_ _6744_/A _6744_/B VGND VGND VPWR VPWR _6610_/B sky130_fd_sc_hd__or2_1
XFILLER_76_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6177_ _6181_/A _6633_/A VGND VGND VPWR VPWR _6232_/C sky130_fd_sc_hd__xnor2_1
XFILLER_57_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5128_ _5068_/C _5127_/A _5127_/Y _5128_/B2 VGND VGND VPWR VPWR _5128_/X sky130_fd_sc_hd__a22o_1
XFILLER_57_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5059_ hold44/X _5059_/A1 _5065_/S VGND VGND VPWR VPWR _5060_/A sky130_fd_sc_hd__mux2_1
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8818_ _9484_/CLK _8818_/D fanout430/X VGND VGND VPWR VPWR _8818_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_111_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8749_ _8748_/X _8749_/A1 _8765_/S VGND VGND VPWR VPWR _8750_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold60 hold60/A VGND VGND VPWR VPWR hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A VGND VGND VPWR VPWR hold71/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 hold82/A VGND VGND VPWR VPWR hold82/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold93 hold93/A VGND VGND VPWR VPWR hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4430_ _9447_/Q _7746_/A _4424_/Y _9199_/Q _4429_/X VGND VGND VPWR VPWR _4431_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA_2 _5851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4361_ hold49/X hold22/X _4360_/Y VGND VGND VPWR VPWR hold50/A sky130_fd_sc_hd__a21bo_1
XFILLER_172_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6100_ _6141_/A _6228_/A VGND VGND VPWR VPWR _6101_/A sky130_fd_sc_hd__or2_1
XFILLER_98_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7080_ _9142_/Q _5809_/X hold65/X VGND VGND VPWR VPWR _7080_/X sky130_fd_sc_hd__mux2_1
X_6031_ _6031_/A VGND VGND VPWR VPWR _9083_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7982_ _7991_/B _7984_/C VGND VGND VPWR VPWR _7983_/A sky130_fd_sc_hd__and2_4
XFILLER_82_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6933_ _6923_/Y _6925_/X _6929_/Y _6932_/Y VGND VGND VPWR VPWR _6953_/B sky130_fd_sc_hd__o31a_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6864_ _6969_/C _6864_/B _6994_/A VGND VGND VPWR VPWR _6864_/X sky130_fd_sc_hd__or3_1
XFILLER_35_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5815_ _5815_/A VGND VGND VPWR VPWR _8986_/D sky130_fd_sc_hd__clkbuf_1
X_8603_ _5130_/A _9527_/Q _8013_/A _8602_/X VGND VGND VPWR VPWR _8603_/X sky130_fd_sc_hd__a211o_1
X_9583_ _9583_/A _5085_/Y VGND VGND VPWR VPWR mgmt_gpio_out[29] sky130_fd_sc_hd__ebufn_8
XFILLER_179_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6795_ _6795_/A _6811_/A _6811_/B VGND VGND VPWR VPWR _6960_/B sky130_fd_sc_hd__and3_1
XFILLER_179_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8534_ _9334_/Q _8298_/X _8370_/X _9254_/Q _8533_/X VGND VGND VPWR VPWR _8537_/C
+ sky130_fd_sc_hd__a221o_1
X_5746_ _5746_/A VGND VGND VPWR VPWR _8956_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8465_ _9283_/Q _8316_/X _8327_/X _9259_/Q VGND VGND VPWR VPWR _8465_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5677_ _5677_/A VGND VGND VPWR VPWR _8927_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7416_ _7416_/A VGND VGND VPWR VPWR _9291_/D sky130_fd_sc_hd__clkbuf_1
X_4628_ _9204_/Q _4416_/Y _5656_/A _8922_/Q _4627_/X VGND VGND VPWR VPWR _4633_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_190_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8396_ _8701_/A _8396_/B _8396_/C _8396_/D VGND VGND VPWR VPWR _8397_/C sky130_fd_sc_hd__or4_1
XFILLER_163_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold530 _9295_/Q VGND VGND VPWR VPWR hold530/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7347_ _7347_/A VGND VGND VPWR VPWR _9259_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4559_ input25/X _4460_/Y _4419_/Y _9365_/Q VGND VGND VPWR VPWR _4559_/X sky130_fd_sc_hd__a22o_1
Xhold541 _5556_/X VGND VGND VPWR VPWR _5557_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold552 _6037_/X VGND VGND VPWR VPWR _6038_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold563 _7300_/X VGND VGND VPWR VPWR _7301_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold574 _9185_/Q VGND VGND VPWR VPWR hold574/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold585 _7603_/X VGND VGND VPWR VPWR _7604_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7278_ _7278_/A VGND VGND VPWR VPWR _9229_/D sky130_fd_sc_hd__clkbuf_1
Xhold596 _7551_/X VGND VGND VPWR VPWR _7552_/A sky130_fd_sc_hd__dlygate4sd3_1
X_9017_ _9475_/CLK _9017_/D fanout481/X VGND VGND VPWR VPWR _9578_/A sky130_fd_sc_hd__dfrtp_1
X_6229_ _6891_/A _6794_/A VGND VGND VPWR VPWR _6230_/C sky130_fd_sc_hd__and2_1
XFILLER_77_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1230 _8863_/Q VGND VGND VPWR VPWR hold881/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1241 _7078_/X VGND VGND VPWR VPWR hold875/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 _7273_/X VGND VGND VPWR VPWR hold687/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1263 _9099_/Q VGND VGND VPWR VPWR hold894/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1274 _7398_/X VGND VGND VPWR VPWR hold430/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1285 _9338_/Q VGND VGND VPWR VPWR hold713/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_403 _8796_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput150 wb_adr_i[27] VGND VGND VPWR VPWR input150/X sky130_fd_sc_hd__clkbuf_1
Xinput161 wb_adr_i[8] VGND VGND VPWR VPWR _6080_/B sky130_fd_sc_hd__clkbuf_1
Xinput172 wb_dat_i[17] VGND VGND VPWR VPWR _8740_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput183 wb_dat_i[27] VGND VGND VPWR VPWR _8747_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput194 wb_dat_i[8] VGND VGND VPWR VPWR _8729_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5600_ _5600_/A VGND VGND VPWR VPWR _8894_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6580_ _6507_/A _6343_/C _6314_/C _6362_/C _6314_/X VGND VGND VPWR VPWR _6580_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_176_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5531_ _5531_/A VGND VGND VPWR VPWR _8863_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8250_ _8250_/A _8250_/B _8250_/C VGND VGND VPWR VPWR _8250_/X sky130_fd_sc_hd__or3_1
XFILLER_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5462_ _5462_/A VGND VGND VPWR VPWR _8835_/D sky130_fd_sc_hd__clkbuf_1
X_7201_ _6015_/X hold700/X _7209_/S VGND VGND VPWR VPWR _7201_/X sky130_fd_sc_hd__mux2_1
X_4413_ hold53/X VGND VGND VPWR VPWR _4674_/A sky130_fd_sc_hd__buf_8
XFILLER_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8181_ _9099_/Q _8181_/B VGND VGND VPWR VPWR _8181_/X sky130_fd_sc_hd__or2_1
X_5393_ _8810_/Q _5392_/X _5416_/S VGND VGND VPWR VPWR _5393_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7132_ _7132_/A _7132_/B VGND VGND VPWR VPWR _7137_/S sky130_fd_sc_hd__and2_1
XFILLER_160_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7063_ _7063_/A VGND VGND VPWR VPWR _9134_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6014_ _6014_/A VGND VGND VPWR VPWR _9076_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_702 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7965_ _7965_/A _7965_/B _7965_/C _7965_/D VGND VGND VPWR VPWR _8007_/A sky130_fd_sc_hd__or4_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6916_ _6894_/A _6815_/B _6894_/B VGND VGND VPWR VPWR _6917_/D sky130_fd_sc_hd__a21o_1
X_7896_ hold993/X _7904_/B _7895_/Y VGND VGND VPWR VPWR _9499_/D sky130_fd_sc_hd__a21oi_1
X_6847_ _6982_/B _6846_/X _6931_/A VGND VGND VPWR VPWR _6911_/A sky130_fd_sc_hd__a21oi_1
XFILLER_50_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9566_ _9566_/A _5102_/Y VGND VGND VPWR VPWR mgmt_gpio_out[12] sky130_fd_sc_hd__ebufn_8
XFILLER_167_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6778_ _6778_/A _6824_/A VGND VGND VPWR VPWR _6867_/B sky130_fd_sc_hd__or2_2
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8517_ _9381_/Q _8337_/X _8384_/X _9197_/Q _8516_/X VGND VGND VPWR VPWR _8524_/A
+ sky130_fd_sc_hd__a221o_1
X_5729_ _5729_/A VGND VGND VPWR VPWR _8948_/D sky130_fd_sc_hd__clkbuf_1
X_9497_ _9501_/CLK _9497_/D fanout488/X VGND VGND VPWR VPWR _9497_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_163_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8448_ _9210_/Q _8289_/X _8341_/X _9306_/Q _8447_/X VGND VGND VPWR VPWR _8449_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_184_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8379_ _8379_/A VGND VGND VPWR VPWR _8379_/X sky130_fd_sc_hd__buf_8
XFILLER_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold360 _9039_/Q VGND VGND VPWR VPWR hold360/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 _7685_/X VGND VGND VPWR VPWR _7686_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 _7668_/X VGND VGND VPWR VPWR _7669_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold393 _9273_/Q VGND VGND VPWR VPWR hold393/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1060 _5829_/X VGND VGND VPWR VPWR _8990_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1071 _5865_/X VGND VGND VPWR VPWR _5866_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1082 _5832_/X VGND VGND VPWR VPWR _8991_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_200 _8034_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1093 _9292_/Q VGND VGND VPWR VPWR hold259/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_211 _8682_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_222 _8883_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_233 _9467_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_244 wb_clk_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_255 _5174_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_266 _5174_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_277 _5285_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_288 _4601_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_299 _5901_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7750_ hold175/X _5951_/A _7762_/S VGND VGND VPWR VPWR _7751_/A sky130_fd_sc_hd__mux2_1
X_4962_ _8806_/Q VGND VGND VPWR VPWR _5068_/B sky130_fd_sc_hd__buf_2
XFILLER_51_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6701_ _6518_/Y _6441_/B _6759_/C _6700_/X _6882_/B VGND VGND VPWR VPWR _6703_/C
+ sky130_fd_sc_hd__a2111o_1
X_7681_ _7556_/X hold96/X _7693_/S VGND VGND VPWR VPWR hold97/A sky130_fd_sc_hd__mux2_1
X_4893_ _9296_/Q _7425_/A _5750_/A _8958_/Q VGND VGND VPWR VPWR _4896_/B sky130_fd_sc_hd__a22o_1
X_9420_ _9420_/CLK _9420_/D fanout465/X VGND VGND VPWR VPWR _9420_/Q sky130_fd_sc_hd__dfrtp_2
X_6632_ _6399_/A _6973_/B _6660_/B VGND VGND VPWR VPWR _6632_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_149_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9351_ _9461_/CLK _9351_/D fanout422/X VGND VGND VPWR VPWR _9351_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6563_ _6563_/A _6563_/B VGND VGND VPWR VPWR _6792_/A sky130_fd_sc_hd__nor2_1
XFILLER_177_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5514_ _5514_/A VGND VGND VPWR VPWR _8856_/D sky130_fd_sc_hd__clkbuf_1
X_8302_ _8336_/A VGND VGND VPWR VPWR _8398_/A sky130_fd_sc_hd__buf_2
XFILLER_118_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9282_ _9466_/CLK _9282_/D fanout472/X VGND VGND VPWR VPWR _9282_/Q sky130_fd_sc_hd__dfrtp_1
X_6494_ _6906_/C _6788_/C VGND VGND VPWR VPWR _6955_/C sky130_fd_sc_hd__nor2_1
XFILLER_106_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8233_ _9086_/Q _7940_/X _7993_/X _8985_/Q _8232_/X VGND VGND VPWR VPWR _8238_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_145_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5445_ _5445_/A VGND VGND VPWR VPWR _5445_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8164_ _9359_/Q _8020_/X _7990_/X _9279_/Q VGND VGND VPWR VPWR _8171_/B sky130_fd_sc_hd__a22o_1
XFILLER_133_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5376_ _5376_/A VGND VGND VPWR VPWR _5376_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_154_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7115_ _7115_/A VGND VGND VPWR VPWR _9157_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8095_ _9396_/Q _7977_/X _8094_/X _8008_/B VGND VGND VPWR VPWR _8095_/X sky130_fd_sc_hd__a22o_1
XFILLER_86_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7046_ _5951_/X _9127_/Q _7054_/S VGND VGND VPWR VPWR _7046_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8997_ _9532_/CLK _8997_/D fanout446/X VGND VGND VPWR VPWR _8997_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7948_ _8206_/B _7989_/B _7996_/B VGND VGND VPWR VPWR _7949_/A sky130_fd_sc_hd__and3_2
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7879_ _8996_/Q _7920_/B VGND VGND VPWR VPWR _7887_/B sky130_fd_sc_hd__nand2_2
XFILLER_23_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9549_ _9550_/CLK _9549_/D fanout500/X VGND VGND VPWR VPWR _9549_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold190 _9476_/Q VGND VGND VPWR VPWR hold190/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5230_ _9503_/Q _9159_/Q _9162_/Q VGND VGND VPWR VPWR _5231_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5161_ _7902_/B _7850_/B VGND VGND VPWR VPWR _5162_/A sky130_fd_sc_hd__or2_1
XFILLER_123_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5092_ _9363_/Q VGND VGND VPWR VPWR _5092_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8920_ _9084_/CLK _8920_/D fanout444/X VGND VGND VPWR VPWR _8920_/Q sky130_fd_sc_hd__dfstp_2
X_8851_ _9084_/CLK _8851_/D fanout447/X VGND VGND VPWR VPWR _8851_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_64_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7802_ _7802_/A VGND VGND VPWR VPWR _9465_/D sky130_fd_sc_hd__clkbuf_1
X_5994_ _9068_/Q _4507_/X _5994_/S VGND VGND VPWR VPWR _5995_/A sky130_fd_sc_hd__mux2_1
X_8782_ _5207_/A1 _8782_/D _5327_/X VGND VGND VPWR VPWR hold11/A sky130_fd_sc_hd__dfrtp_1
XFILLER_52_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7733_ hold87/X VGND VGND VPWR VPWR _9433_/D sky130_fd_sc_hd__clkbuf_1
X_4945_ input20/X _4460_/Y _4944_/Y _9156_/Q VGND VGND VPWR VPWR _4945_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4876_ input62/X _7144_/A _5596_/A _8894_/Q VGND VGND VPWR VPWR _4876_/X sky130_fd_sc_hd__a22o_1
X_7664_ _7556_/X hold92/X _7676_/S VGND VGND VPWR VPWR hold93/A sky130_fd_sc_hd__mux2_1
XFILLER_20_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9403_ _9419_/CLK _9403_/D fanout482/X VGND VGND VPWR VPWR _9403_/Q sky130_fd_sc_hd__dfrtp_4
X_6615_ _6732_/B _6449_/B _6255_/X VGND VGND VPWR VPWR _6616_/D sky130_fd_sc_hd__o21ai_1
XFILLER_137_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7595_ _7433_/X _9371_/Q hold75/X VGND VGND VPWR VPWR _7595_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9334_ _9367_/CLK _9334_/D fanout423/X VGND VGND VPWR VPWR _9334_/Q sky130_fd_sc_hd__dfrtp_1
X_6546_ _6546_/A _6948_/B VGND VGND VPWR VPWR _6987_/B sky130_fd_sc_hd__or2_1
XFILLER_180_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6477_ _6477_/A VGND VGND VPWR VPWR _6478_/C sky130_fd_sc_hd__clkinv_2
X_9265_ _9483_/CLK _9265_/D fanout473/X VGND VGND VPWR VPWR _9265_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_133_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5428_ _8821_/Q _5402_/X _5435_/S VGND VGND VPWR VPWR _5428_/X sky130_fd_sc_hd__mux2_1
X_8216_ _8216_/A _8216_/B _8216_/C _8216_/D VGND VGND VPWR VPWR _8216_/X sky130_fd_sc_hd__or4_1
XFILLER_133_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput240 _5241_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[5] sky130_fd_sc_hd__buf_12
X_9196_ _9276_/CLK _9196_/D fanout461/X VGND VGND VPWR VPWR _9196_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput251 _5170_/Y VGND VGND VPWR VPWR pad_flash_clk_oeb sky130_fd_sc_hd__buf_12
XFILLER_133_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput262 _9131_/Q VGND VGND VPWR VPWR pll90_sel[2] sky130_fd_sc_hd__buf_12
XFILLER_160_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput273 _9128_/Q VGND VGND VPWR VPWR pll_sel[2] sky130_fd_sc_hd__buf_12
XFILLER_161_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput284 _9135_/Q VGND VGND VPWR VPWR pll_trim[19] sky130_fd_sc_hd__buf_12
X_5359_ _5375_/A _5378_/B VGND VGND VPWR VPWR _5360_/A sky130_fd_sc_hd__and2_1
X_8147_ _9406_/Q _7931_/X _7933_/X _9342_/Q VGND VGND VPWR VPWR _8147_/X sky130_fd_sc_hd__a22o_1
Xoutput295 _8822_/Q VGND VGND VPWR VPWR pll_trim[5] sky130_fd_sc_hd__buf_12
XFILLER_99_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8078_ _9355_/Q _8020_/A _7973_/X _9195_/Q VGND VGND VPWR VPWR _8078_/X sky130_fd_sc_hd__a22o_1
XFILLER_114_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7029_ _7029_/A VGND VGND VPWR VPWR _9119_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire367 wire368/X VGND VGND VPWR VPWR wire367/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4730_ _9158_/Q _7113_/A _4585_/Y input64/X VGND VGND VPWR VPWR _4731_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4661_ hold33/X _4667_/B VGND VGND VPWR VPWR _5596_/A sky130_fd_sc_hd__nor2_8
XFILLER_147_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6400_ _6428_/B _6818_/A VGND VGND VPWR VPWR _6401_/A sky130_fd_sc_hd__or2_1
X_7380_ _7380_/A VGND VGND VPWR VPWR _9274_/D sky130_fd_sc_hd__clkbuf_1
X_4592_ _9115_/Q _4591_/X _4886_/S VGND VGND VPWR VPWR _4592_/X sky130_fd_sc_hd__mux2_1
XFILLER_162_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold904 _9360_/Q VGND VGND VPWR VPWR hold904/X sky130_fd_sc_hd__dlygate4sd3_1
X_6331_ _6802_/A VGND VGND VPWR VPWR _6331_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold915 hold915/A VGND VGND VPWR VPWR hold915/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold926 _9256_/Q VGND VGND VPWR VPWR hold926/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold937 _5390_/X VGND VGND VPWR VPWR _5391_/A sky130_fd_sc_hd__dlygate4sd3_1
X_9050_ _9184_/CLK _9050_/D fanout443/X VGND VGND VPWR VPWR _9050_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_6_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold948 _8041_/X VGND VGND VPWR VPWR _9508_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold959 _9528_/Q VGND VGND VPWR VPWR hold959/X sky130_fd_sc_hd__dlygate4sd3_1
X_6262_ _6262_/A _6556_/B VGND VGND VPWR VPWR _6263_/A sky130_fd_sc_hd__or2_1
XFILLER_88_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5213_ _9010_/Q _9118_/Q _5453_/C VGND VGND VPWR VPWR _5213_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8001_ _8001_/A VGND VGND VPWR VPWR _8001_/X sky130_fd_sc_hd__buf_8
X_6193_ _6312_/A _6312_/B _6739_/B VGND VGND VPWR VPWR _6194_/B sky130_fd_sc_hd__or3b_2
XFILLER_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5144_ _9033_/Q VGND VGND VPWR VPWR _5275_/A sky130_fd_sc_hd__buf_2
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5075_ _5330_/A _5334_/B VGND VGND VPWR VPWR _5076_/A sky130_fd_sc_hd__and2_1
XFILLER_84_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8903_ _9442_/CLK _8903_/D fanout436/X VGND VGND VPWR VPWR _8903_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_25_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8834_ _9172_/CLK _8834_/D fanout494/X VGND VGND VPWR VPWR _8834_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_64_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8765_ _8764_/X _9549_/Q _8765_/S VGND VGND VPWR VPWR _8765_/X sky130_fd_sc_hd__mux2_1
X_5977_ _5977_/A VGND VGND VPWR VPWR _9060_/D sky130_fd_sc_hd__clkbuf_1
X_7716_ _7716_/A VGND VGND VPWR VPWR _9425_/D sky130_fd_sc_hd__clkbuf_1
X_4928_ _8968_/Q _5773_/A _7077_/A _9141_/Q _4927_/X VGND VGND VPWR VPWR _4931_/C
+ sky130_fd_sc_hd__a221o_1
X_8696_ _8942_/Q _7908_/X _8335_/X _8872_/Q VGND VGND VPWR VPWR _8696_/X sky130_fd_sc_hd__a22o_1
X_7647_ _7647_/A VGND VGND VPWR VPWR _9394_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4859_ _9393_/Q _7640_/A _7623_/A hold90/A VGND VGND VPWR VPWR _4859_/X sky130_fd_sc_hd__a22o_2
XFILLER_166_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7578_ _7433_/X _9363_/Q hold78/X VGND VGND VPWR VPWR _7578_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9317_ _9480_/CLK _9317_/D fanout413/X VGND VGND VPWR VPWR _9317_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6529_ _6732_/B _6898_/A VGND VGND VPWR VPWR _6530_/D sky130_fd_sc_hd__or2_2
XFILLER_134_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9248_ _9476_/CLK _9248_/D fanout415/X VGND VGND VPWR VPWR _9248_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9179_ _9181_/CLK _9179_/D fanout488/X VGND VGND VPWR VPWR _9179_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_73_csclk _9090_/CLK VGND VGND VPWR VPWR _9194_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_87_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_11_csclk _9210_/CLK VGND VGND VPWR VPWR _9421_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_26_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _9465_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_98_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5900_ hold20/A VGND VGND VPWR VPWR _7284_/B sky130_fd_sc_hd__buf_12
XFILLER_81_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6880_ _6880_/A _6937_/C _6880_/C _6879_/X VGND VGND VPWR VPWR _6886_/C sky130_fd_sc_hd__or4b_1
X_5831_ _9573_/A _5830_/X hold43/X VGND VGND VPWR VPWR _5831_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5762_ _5762_/A _7132_/B VGND VGND VPWR VPWR _5771_/S sky130_fd_sc_hd__and2_2
XFILLER_22_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8550_ _8701_/A _8550_/B _8550_/C _8550_/D VGND VGND VPWR VPWR _8550_/X sky130_fd_sc_hd__or4_4
X_7501_ _7501_/A VGND VGND VPWR VPWR _9328_/D sky130_fd_sc_hd__clkbuf_1
X_4713_ _8891_/Q _5584_/A _6043_/A _9092_/Q _4712_/X VGND VGND VPWR VPWR _4713_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_175_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5693_ _5693_/A _5693_/B VGND VGND VPWR VPWR _5702_/S sky130_fd_sc_hd__nand2_4
X_8481_ _9412_/Q _8506_/B VGND VGND VPWR VPWR _8481_/X sky130_fd_sc_hd__and2_1
XFILLER_148_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4644_ _8862_/Q _5518_/A _5948_/A _9052_/Q _4643_/X VGND VGND VPWR VPWR _4649_/C
+ sky130_fd_sc_hd__a221o_1
X_7432_ _7432_/A VGND VGND VPWR VPWR _9298_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4575_ _9253_/Q _7321_/A _4483_/Y _4575_/B2 _4574_/X VGND VGND VPWR VPWR _4575_/X
+ sky130_fd_sc_hd__a221o_1
Xhold701 _7201_/X VGND VGND VPWR VPWR _7202_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7363_ _7363_/A VGND VGND VPWR VPWR _9266_/D sky130_fd_sc_hd__clkbuf_1
Xhold712 hold712/A VGND VGND VPWR VPWR hold712/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold723 _9354_/Q VGND VGND VPWR VPWR hold723/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9102_ _9442_/CLK _9102_/D fanout436/X VGND VGND VPWR VPWR hold71/A sky130_fd_sc_hd__dfrtp_4
Xhold734 _7421_/X VGND VGND VPWR VPWR _7422_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6314_ _6715_/B _6343_/C _6314_/C VGND VGND VPWR VPWR _6314_/X sky130_fd_sc_hd__and3_1
Xhold745 _7048_/X VGND VGND VPWR VPWR _7049_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7294_ _7294_/A VGND VGND VPWR VPWR _9236_/D sky130_fd_sc_hd__clkbuf_1
Xhold756 _9358_/Q VGND VGND VPWR VPWR hold756/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold767 _7102_/X VGND VGND VPWR VPWR _7103_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold778 hold778/A VGND VGND VPWR VPWR hold778/X sky130_fd_sc_hd__dlygate4sd3_1
X_9033_ _9551_/CLK _9033_/D fanout499/X VGND VGND VPWR VPWR _9033_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_170_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6245_ _6721_/A _6724_/A VGND VGND VPWR VPWR _6744_/B sky130_fd_sc_hd__nand2_1
Xhold789 _7311_/X VGND VGND VPWR VPWR _7312_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6176_ _6181_/A _6633_/A _6181_/B VGND VGND VPWR VPWR _6178_/B sky130_fd_sc_hd__a21o_1
XFILLER_162_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5127_ _5127_/A _5127_/B VGND VGND VPWR VPWR _5127_/Y sky130_fd_sc_hd__nor2_1
XFILLER_84_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5058_ _5058_/A VGND VGND VPWR VPWR _8785_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8817_ _9476_/CLK _8817_/D fanout414/X VGND VGND VPWR VPWR _8817_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8748_ _5271_/A _8748_/A2 _8748_/B1 _8727_/Y _8747_/X VGND VGND VPWR VPWR _8748_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8679_ hold970/X _8017_/X _8678_/X VGND VGND VPWR VPWR _8679_/X sky130_fd_sc_hd__o21a_1
XFILLER_166_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold50 hold50/A VGND VGND VPWR VPWR hold50/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold61 hold61/A VGND VGND VPWR VPWR hold61/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_36_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold72 hold72/A VGND VGND VPWR VPWR hold72/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A VGND VGND VPWR VPWR hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 hold94/A VGND VGND VPWR VPWR hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_2_0_mgmt_gpio_in[4] clkbuf_2_3_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _5235__1/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_16_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_3 _9008_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4360_ hold80/A _5021_/B VGND VGND VPWR VPWR _4360_/Y sky130_fd_sc_hd__nand2_1
XFILLER_140_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6030_ hold547/X _5690_/X _6030_/S VGND VGND VPWR VPWR _6030_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7981_ _7981_/A VGND VGND VPWR VPWR _7981_/X sky130_fd_sc_hd__buf_6
XFILLER_26_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6932_ _6989_/A _6989_/B VGND VGND VPWR VPWR _6932_/Y sky130_fd_sc_hd__nor2_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6863_ _6869_/A _6863_/B _6863_/C _6863_/D VGND VGND VPWR VPWR _6994_/A sky130_fd_sc_hd__or4_1
X_8602_ _8848_/Q _8400_/B _8588_/X _8601_/X _8627_/S VGND VGND VPWR VPWR _8602_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_179_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5814_ hold436/X _5687_/X _5816_/S VGND VGND VPWR VPWR _5815_/A sky130_fd_sc_hd__mux2_1
X_9582_ _9582_/A _5086_/Y VGND VGND VPWR VPWR mgmt_gpio_out[28] sky130_fd_sc_hd__ebufn_8
X_6794_ _6794_/A _6794_/B VGND VGND VPWR VPWR _6794_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8533_ _9454_/Q _8360_/A _8381_/A _9366_/Q VGND VGND VPWR VPWR _8533_/X sky130_fd_sc_hd__a22o_1
X_5745_ _5650_/X hold710/X _5747_/S VGND VGND VPWR VPWR _5746_/A sky130_fd_sc_hd__mux2_1
X_8464_ _9459_/Q _8360_/C _8411_/A _9339_/Q _8463_/X VGND VGND VPWR VPWR _8474_/B
+ sky130_fd_sc_hd__a221o_1
X_5676_ _5653_/X hold121/X _5676_/S VGND VGND VPWR VPWR _5676_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7415_ _7236_/X _9291_/Q _7423_/S VGND VGND VPWR VPWR _7415_/X sky130_fd_sc_hd__mux2_1
X_4627_ input7/X _4406_/Y _6007_/A _9078_/Q VGND VGND VPWR VPWR _4627_/X sky130_fd_sc_hd__a22o_1
X_8395_ _9432_/Q _7908_/X _8387_/X _8394_/X VGND VGND VPWR VPWR _8396_/D sky130_fd_sc_hd__a211o_1
Xhold520 _9311_/Q VGND VGND VPWR VPWR hold520/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold531 _7423_/X VGND VGND VPWR VPWR _7424_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4558_ _9277_/Q _7374_/A _7678_/A _9413_/Q _4557_/X VGND VGND VPWR VPWR _4573_/B
+ sky130_fd_sc_hd__a221o_2
X_7346_ _7236_/X _9259_/Q _7354_/S VGND VGND VPWR VPWR _7346_/X sky130_fd_sc_hd__mux2_1
Xhold542 _8885_/Q VGND VGND VPWR VPWR hold542/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold553 hold553/A VGND VGND VPWR VPWR hold553/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold564 _9327_/Q VGND VGND VPWR VPWR hold564/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 _5440_/X VGND VGND VPWR VPWR _5441_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4489_ _4489_/A _4536_/B VGND VGND VPWR VPWR _5453_/B sky130_fd_sc_hd__nand2_8
Xhold586 _9415_/Q VGND VGND VPWR VPWR hold586/X sky130_fd_sc_hd__dlygate4sd3_1
X_7277_ _7242_/X hold222/X _7282_/S VGND VGND VPWR VPWR _7277_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold597 _8950_/Q VGND VGND VPWR VPWR hold597/X sky130_fd_sc_hd__dlygate4sd3_1
X_9016_ _9181_/CLK _9016_/D fanout487/X VGND VGND VPWR VPWR _9561_/A sky130_fd_sc_hd__dfrtp_2
X_6228_ _6228_/A _6967_/A VGND VGND VPWR VPWR _6228_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6159_ _6181_/A VGND VGND VPWR VPWR _6973_/A sky130_fd_sc_hd__buf_4
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1220 _8906_/Q VGND VGND VPWR VPWR hold435/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1231 _8866_/Q VGND VGND VPWR VPWR hold422/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1242 _8958_/Q VGND VGND VPWR VPWR hold870/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1253 _9070_/Q VGND VGND VPWR VPWR hold546/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1264 _8871_/Q VGND VGND VPWR VPWR hold387/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1275 _7082_/X VGND VGND VPWR VPWR hold465/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_404 _5279_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput140 wb_adr_i[18] VGND VGND VPWR VPWR _6078_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput151 wb_adr_i[28] VGND VGND VPWR VPWR input151/X sky130_fd_sc_hd__clkbuf_1
Xinput162 wb_adr_i[9] VGND VGND VPWR VPWR _6080_/A sky130_fd_sc_hd__clkbuf_1
Xinput173 wb_dat_i[18] VGND VGND VPWR VPWR _8744_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput184 wb_dat_i[28] VGND VGND VPWR VPWR _8751_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput195 wb_dat_i[9] VGND VGND VPWR VPWR _8739_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5530_ _5291_/X hold881/X _5538_/S VGND VGND VPWR VPWR _5531_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5461_ _5311_/X hold383/X _5472_/S VGND VGND VPWR VPWR _5461_/X sky130_fd_sc_hd__mux2_1
X_4412_ hold31/X hold52/X VGND VGND VPWR VPWR hold53/A sky130_fd_sc_hd__or2_1
X_7200_ _7200_/A VGND VGND VPWR VPWR _9194_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5392_ _5951_/A VGND VGND VPWR VPWR _5392_/X sky130_fd_sc_hd__buf_6
X_8180_ _9048_/Q _7923_/A _7997_/A _8953_/Q _8179_/X VGND VGND VPWR VPWR _8184_/C
+ sky130_fd_sc_hd__a221o_1
X_7131_ _7131_/A VGND VGND VPWR VPWR _9164_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7062_ _9134_/Q _6048_/X _7072_/S VGND VGND VPWR VPWR _7062_/X sky130_fd_sc_hd__mux2_1
X_6013_ _6012_/X _9076_/Q _6019_/S VGND VGND VPWR VPWR _6013_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7964_ _9304_/Q _8023_/B _7958_/X _9256_/Q _7963_/X VGND VGND VPWR VPWR _7965_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_82_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6915_ _6915_/A _6915_/B _6915_/C VGND VGND VPWR VPWR _6972_/B sky130_fd_sc_hd__or3_1
XFILLER_82_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7895_ _9499_/Q _7887_/B _7904_/B VGND VGND VPWR VPWR _7895_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_22_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6846_ _6925_/C _6846_/B _7006_/C _6929_/B VGND VGND VPWR VPWR _6846_/X sky130_fd_sc_hd__and4b_1
XFILLER_23_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9565_ _9565_/A _5103_/Y VGND VGND VPWR VPWR mgmt_gpio_out[11] sky130_fd_sc_hd__ebufn_8
X_6777_ _6835_/B _6983_/A _6987_/D _6924_/D VGND VGND VPWR VPWR _6784_/C sky130_fd_sc_hd__or4_1
XFILLER_167_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8516_ _9437_/Q _7908_/X _8335_/X _9277_/Q VGND VGND VPWR VPWR _8516_/X sky130_fd_sc_hd__a22o_1
X_5728_ _5629_/X hold831/X _5736_/S VGND VGND VPWR VPWR _5729_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9496_ _9520_/CLK _9496_/D fanout470/X VGND VGND VPWR VPWR _9496_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8447_ _9394_/Q _8304_/X _8324_/X _9242_/Q VGND VGND VPWR VPWR _8447_/X sky130_fd_sc_hd__a22o_1
XFILLER_175_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5659_ hold742/X _5587_/X _5665_/S VGND VGND VPWR VPWR _5660_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8378_ _8378_/A VGND VGND VPWR VPWR _8378_/X sky130_fd_sc_hd__buf_6
XFILLER_117_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold350 hold350/A VGND VGND VPWR VPWR hold350/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 _5927_/X VGND VGND VPWR VPWR _5928_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7329_ _9251_/Q hold46/X _7337_/S VGND VGND VPWR VPWR hold67/A sky130_fd_sc_hd__mux2_1
XFILLER_104_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold372 _9412_/Q VGND VGND VPWR VPWR hold372/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 _8835_/Q VGND VGND VPWR VPWR hold383/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold394 _9305_/Q VGND VGND VPWR VPWR hold394/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1050 hold14/A VGND VGND VPWR VPWR _5057_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1061 _5825_/X VGND VGND VPWR VPWR _5826_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1072 _5866_/X VGND VGND VPWR VPWR _9006_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1083 _5843_/X VGND VGND VPWR VPWR _5844_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1094 _7417_/X VGND VGND VPWR VPWR _7418_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_201 _8105_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_212 _8682_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_223 _9318_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_234 _8898_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_245 wb_dat_i[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_256 _5174_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_267 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_278 _5285_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_289 _4904_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4961_ _4961_/A _4961_/B _4961_/C VGND VGND VPWR VPWR _4961_/X sky130_fd_sc_hd__or3_4
X_6700_ _6700_/A _6700_/B _6700_/C _6700_/D VGND VGND VPWR VPWR _6700_/X sky130_fd_sc_hd__or4_1
XFILLER_189_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7680_ _7680_/A VGND VGND VPWR VPWR _9408_/D sky130_fd_sc_hd__clkbuf_1
X_4892_ _5228_/A1 _4889_/Y _4890_/Y _7129_/A _9164_/Q VGND VGND VPWR VPWR _4896_/A
+ sky130_fd_sc_hd__a32o_1
X_6631_ _6736_/B _6781_/B VGND VGND VPWR VPWR _6660_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9350_ _9461_/CLK _9350_/D fanout422/X VGND VGND VPWR VPWR _9350_/Q sky130_fd_sc_hd__dfrtp_4
X_6562_ _6562_/A _6562_/B VGND VGND VPWR VPWR _6563_/B sky130_fd_sc_hd__nor2_1
XFILLER_118_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8301_ _8301_/A VGND VGND VPWR VPWR _8398_/B sky130_fd_sc_hd__buf_6
X_5513_ hold437/X _5398_/X _5515_/S VGND VGND VPWR VPWR _5513_/X sky130_fd_sc_hd__mux2_1
X_9281_ _9483_/CLK _9281_/D fanout474/X VGND VGND VPWR VPWR _9281_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_157_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6493_ _6906_/B _6736_/A VGND VGND VPWR VPWR _6788_/C sky130_fd_sc_hd__or2_1
X_8232_ _8975_/Q _7947_/X _8008_/B _8231_/X VGND VGND VPWR VPWR _8232_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5444_ _7011_/A _7013_/B VGND VGND VPWR VPWR _5445_/A sky130_fd_sc_hd__and2_1
XFILLER_145_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8163_ _9407_/Q _7931_/X _7933_/X _9343_/Q VGND VGND VPWR VPWR _8171_/A sky130_fd_sc_hd__a22o_1
X_5375_ _5375_/A _5378_/B VGND VGND VPWR VPWR _5376_/A sky130_fd_sc_hd__and2_1
X_7114_ _6018_/X hold151/X _7124_/S VGND VGND VPWR VPWR _7114_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8094_ _9316_/Q _8206_/B VGND VGND VPWR VPWR _8094_/X sky130_fd_sc_hd__or2_1
X_7045_ _7045_/A VGND VGND VPWR VPWR _9126_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8996_ _9532_/CLK _8996_/D fanout441/X VGND VGND VPWR VPWR _8996_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_15_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7947_ _7947_/A VGND VGND VPWR VPWR _7947_/X sky130_fd_sc_hd__buf_6
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7878_ _7902_/B _7991_/B VGND VGND VPWR VPWR _7881_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6829_ _6800_/A _6828_/X _6457_/X _6463_/B VGND VGND VPWR VPWR _6834_/B sky130_fd_sc_hd__o211a_1
XFILLER_11_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9548_ _9551_/CLK _9548_/D fanout500/X VGND VGND VPWR VPWR _9548_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_10_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9479_ _9485_/CLK _9479_/D fanout405/X VGND VGND VPWR VPWR _9479_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold180 _9213_/Q VGND VGND VPWR VPWR hold180/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 _7824_/X VGND VGND VPWR VPWR _7825_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5160_ _8652_/S _5160_/B VGND VGND VPWR VPWR _7850_/B sky130_fd_sc_hd__nor2_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5091_ _9371_/Q VGND VGND VPWR VPWR _5091_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8850_ _9084_/CLK _8850_/D fanout447/X VGND VGND VPWR VPWR _8850_/Q sky130_fd_sc_hd__dfrtp_4
X_7801_ _5392_/X hold517/X _7813_/S VGND VGND VPWR VPWR _7802_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8781_ _5207_/A1 _8781_/D _5325_/X VGND VGND VPWR VPWR hold36/A sky130_fd_sc_hd__dfrtp_1
X_5993_ _5993_/A VGND VGND VPWR VPWR _9067_/D sky130_fd_sc_hd__clkbuf_1
X_7732_ _7556_/X _9433_/Q hold86/X VGND VGND VPWR VPWR hold87/A sky130_fd_sc_hd__mux2_1
X_4944_ _7111_/A _7111_/B VGND VGND VPWR VPWR _4944_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7663_ _7663_/A VGND VGND VPWR VPWR _9400_/D sky130_fd_sc_hd__clkbuf_1
X_4875_ _9345_/Q _7536_/A _7571_/A _9361_/Q _4874_/X VGND VGND VPWR VPWR _4883_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9402_ _9467_/CLK _9402_/D fanout475/X VGND VGND VPWR VPWR _9402_/Q sky130_fd_sc_hd__dfrtp_4
X_6614_ _6857_/B _6946_/A _6614_/C _6613_/X VGND VGND VPWR VPWR _6616_/C sky130_fd_sc_hd__or4b_1
X_7594_ _7594_/A VGND VGND VPWR VPWR _9370_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9333_ _9436_/CLK _9333_/D fanout460/X VGND VGND VPWR VPWR _9333_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_165_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6545_ _6293_/X _6378_/X _6544_/X _6908_/A hold85/X VGND VGND VPWR VPWR _9104_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_146_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9264_ _9436_/CLK _9264_/D fanout462/X VGND VGND VPWR VPWR _9264_/Q sky130_fd_sc_hd__dfstp_1
X_6476_ _6778_/A _6754_/A _6754_/B VGND VGND VPWR VPWR _6483_/A sky130_fd_sc_hd__or3_1
XFILLER_109_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8215_ _9036_/Q _7938_/X _8077_/X _8934_/Q _8214_/X VGND VGND VPWR VPWR _8216_/D
+ sky130_fd_sc_hd__a221o_1
Xoutput230 _5265_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[30] sky130_fd_sc_hd__buf_12
X_5427_ _5427_/A VGND VGND VPWR VPWR _8820_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9195_ _9195_/CLK _9195_/D fanout467/X VGND VGND VPWR VPWR _9195_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput241 _5242_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[6] sky130_fd_sc_hd__buf_12
Xoutput252 _5166_/X VGND VGND VPWR VPWR pad_flash_csb sky130_fd_sc_hd__buf_12
Xoutput263 _9140_/Q VGND VGND VPWR VPWR pll_bypass sky130_fd_sc_hd__buf_12
XFILLER_133_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput274 _8817_/Q VGND VGND VPWR VPWR pll_trim[0] sky130_fd_sc_hd__buf_12
X_8146_ _9206_/Q _7938_/X _8077_/X _9350_/Q _8145_/X VGND VGND VPWR VPWR _8149_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_160_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput285 _8818_/Q VGND VGND VPWR VPWR pll_trim[1] sky130_fd_sc_hd__buf_12
X_5358_ _5453_/C VGND VGND VPWR VPWR _5378_/B sky130_fd_sc_hd__buf_2
XFILLER_114_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput296 _8823_/Q VGND VGND VPWR VPWR pll_trim[6] sky130_fd_sc_hd__buf_12
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8077_ _8077_/A VGND VGND VPWR VPWR _8077_/X sky130_fd_sc_hd__buf_6
X_5289_ _5067_/B hold431/X _5413_/S VGND VGND VPWR VPWR _5289_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7028_ _5947_/X _9119_/Q _7030_/S VGND VGND VPWR VPWR _7028_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8979_ _9283_/CLK _8979_/D fanout485/X VGND VGND VPWR VPWR _8979_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_70_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire368 wire369/X VGND VGND VPWR VPWR wire368/X sky130_fd_sc_hd__clkbuf_1
XFILLER_171_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout490 fanout495/X VGND VGND VPWR VPWR fanout490/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4660_ _7126_/A _7158_/B VGND VGND VPWR VPWR _5493_/A sky130_fd_sc_hd__nor2_4
XFILLER_30_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4591_ _4591_/A _4591_/B _4591_/C VGND VGND VPWR VPWR _4591_/X sky130_fd_sc_hd__or3_4
XFILLER_190_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6330_ _6871_/B _6874_/A VGND VGND VPWR VPWR _6330_/Y sky130_fd_sc_hd__nor2_1
XFILLER_127_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold905 _9288_/Q VGND VGND VPWR VPWR hold905/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold916 hold916/A VGND VGND VPWR VPWR hold916/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold927 _9320_/Q VGND VGND VPWR VPWR hold927/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold938 _9280_/Q VGND VGND VPWR VPWR hold938/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold949 _8828_/Q VGND VGND VPWR VPWR hold949/X sky130_fd_sc_hd__dlygate4sd3_1
X_6261_ _6311_/B _7001_/A VGND VGND VPWR VPWR _6268_/C sky130_fd_sc_hd__nor2_1
X_8000_ _8206_/B _8000_/B _8002_/B VGND VGND VPWR VPWR _8001_/A sky130_fd_sc_hd__and3_2
X_5212_ _5212_/A VGND VGND VPWR VPWR _9560_/A sky130_fd_sc_hd__buf_2
XFILLER_88_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6192_ _6192_/A _6504_/A VGND VGND VPWR VPWR _6312_/B sky130_fd_sc_hd__nor2_1
XFILLER_97_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5143_ _5271_/A _5115_/X _5870_/B VGND VGND VPWR VPWR _9032_/D sky130_fd_sc_hd__a21o_1
XFILLER_97_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5074_ _7025_/B VGND VGND VPWR VPWR _5334_/B sky130_fd_sc_hd__buf_4
XFILLER_57_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8902_ _9442_/CLK _8902_/D fanout436/X VGND VGND VPWR VPWR _8902_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8833_ _9172_/CLK _8833_/D fanout493/X VGND VGND VPWR VPWR _8833_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8764_ _5271_/A _8764_/A2 _8764_/B1 _8727_/Y _8764_/C1 VGND VGND VPWR VPWR _8764_/X
+ sky130_fd_sc_hd__a221o_1
X_5976_ _9060_/Q _4507_/X _5976_/S VGND VGND VPWR VPWR _5977_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7715_ _7556_/X _7715_/A1 hold95/X VGND VGND VPWR VPWR _7716_/A sky130_fd_sc_hd__mux2_1
X_4927_ _9224_/Q _4454_/Y _7481_/A _9320_/Q VGND VGND VPWR VPWR _4927_/X sky130_fd_sc_hd__a22o_1
X_8695_ _9073_/Q _8388_/X _8379_/X _9039_/Q _8694_/X VGND VGND VPWR VPWR _8700_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_33_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7646_ _7645_/X hold621/X hold84/X VGND VGND VPWR VPWR _7647_/A sky130_fd_sc_hd__mux2_1
X_4858_ _7126_/A _4858_/B VGND VGND VPWR VPWR _7086_/A sky130_fd_sc_hd__nor2_2
XFILLER_21_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7577_ _7577_/A VGND VGND VPWR VPWR _9362_/D sky130_fd_sc_hd__clkbuf_1
X_4789_ _8875_/Q _5551_/A _5727_/A _8950_/Q VGND VGND VPWR VPWR _4789_/X sky130_fd_sc_hd__a22o_2
X_9316_ _9420_/CLK _9316_/D fanout464/X VGND VGND VPWR VPWR _9316_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_4_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6528_ _6862_/A _6528_/B VGND VGND VPWR VPWR _6729_/B sky130_fd_sc_hd__or2_1
XFILLER_181_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_7_csclk _9359_/CLK VGND VGND VPWR VPWR _9272_/CLK sky130_fd_sc_hd__clkbuf_16
X_9247_ _9398_/CLK _9247_/D _5332_/A VGND VGND VPWR VPWR _9247_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6459_ _6850_/B _6596_/B VGND VGND VPWR VPWR _6460_/B sky130_fd_sc_hd__nor2_2
XFILLER_106_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9178_ _9178_/CLK _9178_/D fanout487/X VGND VGND VPWR VPWR _9178_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8129_ _5139_/A hold989/X _8013_/X VGND VGND VPWR VPWR _8129_/X sky130_fd_sc_hd__a21o_1
XFILLER_114_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5830_ hold383/X _7648_/A _5842_/S VGND VGND VPWR VPWR _5830_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5761_ _5761_/A VGND VGND VPWR VPWR _5761_/X sky130_fd_sc_hd__buf_4
X_7500_ _7302_/X hold928/X _7515_/S VGND VGND VPWR VPWR _7501_/A sky130_fd_sc_hd__mux2_1
X_4712_ _9251_/Q _7321_/A _5506_/A _8856_/Q VGND VGND VPWR VPWR _4712_/X sky130_fd_sc_hd__a22o_1
XFILLER_30_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8480_ _9420_/Q _8402_/X _8378_/X _9356_/Q _8479_/X VGND VGND VPWR VPWR _8487_/A
+ sky130_fd_sc_hd__a221o_1
X_5692_ _5692_/A VGND VGND VPWR VPWR _8932_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7431_ _7430_/X hold402/X _7444_/S VGND VGND VPWR VPWR _7431_/X sky130_fd_sc_hd__mux2_1
X_4643_ _9220_/Q _7249_/A _5784_/A _8977_/Q VGND VGND VPWR VPWR _4643_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7362_ _7233_/X hold778/X _7372_/S VGND VGND VPWR VPWR _7363_/A sky130_fd_sc_hd__mux2_1
X_4574_ input97/X _4488_/Y _7729_/A _9437_/Q VGND VGND VPWR VPWR _4574_/X sky130_fd_sc_hd__a22o_1
Xhold702 _7098_/X VGND VGND VPWR VPWR _7099_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 hold713/A VGND VGND VPWR VPWR hold713/X sky130_fd_sc_hd__dlygate4sd3_1
X_9101_ _9442_/CLK _9101_/D fanout437/X VGND VGND VPWR VPWR _9101_/Q sky130_fd_sc_hd__dfstp_2
X_6313_ _6788_/A _6788_/B VGND VGND VPWR VPWR _6343_/C sky130_fd_sc_hd__nor2_2
Xhold724 hold724/A VGND VGND VPWR VPWR hold724/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 _9390_/Q VGND VGND VPWR VPWR hold735/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 _9350_/Q VGND VGND VPWR VPWR hold746/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7293_ _7239_/X hold289/X _7300_/S VGND VGND VPWR VPWR _7293_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold757 _7567_/X VGND VGND VPWR VPWR _7568_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_9032_ _9551_/CLK _9032_/D fanout499/X VGND VGND VPWR VPWR _9032_/Q sky130_fd_sc_hd__dfrtp_4
Xhold768 hold768/A VGND VGND VPWR VPWR hold768/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold779 _9202_/Q VGND VGND VPWR VPWR hold779/X sky130_fd_sc_hd__dlygate4sd3_1
X_6244_ _6744_/A _6623_/A VGND VGND VPWR VPWR _6244_/X sky130_fd_sc_hd__or2_1
XFILLER_130_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6175_ _6175_/A _6633_/A VGND VGND VPWR VPWR _6178_/A sky130_fd_sc_hd__nand2_1
XFILLER_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5126_ _5126_/A1 _5115_/X _8705_/B _8705_/A VGND VGND VPWR VPWR _9030_/D sky130_fd_sc_hd__a22o_1
XFILLER_111_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5057_ _5059_/A1 _5057_/A1 _5065_/S VGND VGND VPWR VPWR _5058_/A sky130_fd_sc_hd__mux2_1
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8816_ _9487_/CLK _8816_/D fanout411/X VGND VGND VPWR VPWR _8816_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8747_ _5287_/A _8747_/A2 _8747_/B1 _5275_/A VGND VGND VPWR VPWR _8747_/X sky130_fd_sc_hd__a22o_1
XFILLER_71_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5959_ _5959_/A VGND VGND VPWR VPWR _9052_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8678_ _5130_/A _9530_/Q _8013_/A _8677_/X VGND VGND VPWR VPWR _8678_/X sky130_fd_sc_hd__a211o_1
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7629_ _7629_/A VGND VGND VPWR VPWR _9386_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold40 hold40/A VGND VGND VPWR VPWR hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A VGND VGND VPWR VPWR hold51/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold62 hold62/A VGND VGND VPWR VPWR hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A VGND VGND VPWR VPWR hold73/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold84 hold84/A VGND VGND VPWR VPWR hold84/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A VGND VGND VPWR VPWR hold95/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_4 _9008_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7980_ _7998_/A _7984_/C _8002_/B VGND VGND VPWR VPWR _7981_/A sky130_fd_sc_hd__and3_2
XFILLER_66_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6931_ _6931_/A _6931_/B _6907_/C VGND VGND VPWR VPWR _6989_/B sky130_fd_sc_hd__or3b_1
XFILLER_81_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6862_ _6862_/A _6862_/B VGND VGND VPWR VPWR _6863_/B sky130_fd_sc_hd__nor2_1
XFILLER_50_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_8601_ _8701_/A _8601_/B _8601_/C _8601_/D VGND VGND VPWR VPWR _8601_/X sky130_fd_sc_hd__or4_1
XFILLER_34_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5813_ _5813_/A VGND VGND VPWR VPWR _8985_/D sky130_fd_sc_hd__clkbuf_1
X_9581_ _9581_/A _5087_/Y VGND VGND VPWR VPWR mgmt_gpio_out[27] sky130_fd_sc_hd__ebufn_8
XFILLER_50_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6793_ _6873_/B _6793_/B VGND VGND VPWR VPWR _6955_/D sky130_fd_sc_hd__nor2_1
XFILLER_167_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8532_ _9350_/Q _8386_/A _8657_/B _9414_/Q _8531_/X VGND VGND VPWR VPWR _8537_/B
+ sky130_fd_sc_hd__a221o_1
X_5744_ _5744_/A VGND VGND VPWR VPWR _8955_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8463_ _9219_/Q _8391_/A _8367_/A _9475_/Q _8462_/X VGND VGND VPWR VPWR _8463_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5675_ _5675_/A VGND VGND VPWR VPWR _8926_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_72_csclk _9090_/CLK VGND VGND VPWR VPWR _9434_/CLK sky130_fd_sc_hd__clkbuf_16
X_7414_ _7414_/A VGND VGND VPWR VPWR _9290_/D sky130_fd_sc_hd__clkbuf_1
X_4626_ _4667_/A _4956_/A VGND VGND VPWR VPWR _6007_/A sky130_fd_sc_hd__nor2_8
XFILLER_135_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8394_ _9224_/Q _8388_/X _8506_/B _9408_/Q _8393_/X VGND VGND VPWR VPWR _8394_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold510 _9458_/Q VGND VGND VPWR VPWR hold510/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7345_ _7345_/A VGND VGND VPWR VPWR _9258_/D sky130_fd_sc_hd__clkbuf_1
X_4557_ _9445_/Q _7746_/A _7043_/A _9131_/Q VGND VGND VPWR VPWR _4557_/X sky130_fd_sc_hd__a22o_2
Xhold521 _7461_/X VGND VGND VPWR VPWR _7462_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 hold532/A VGND VGND VPWR VPWR hold532/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 _5578_/X VGND VGND VPWR VPWR _5579_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold554 _9075_/Q VGND VGND VPWR VPWR hold554/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 _7497_/X VGND VGND VPWR VPWR _7498_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7276_ _7276_/A VGND VGND VPWR VPWR _9228_/D sky130_fd_sc_hd__clkbuf_1
X_4488_ _4878_/A _7126_/A VGND VGND VPWR VPWR _4488_/Y sky130_fd_sc_hd__nor2_4
Xhold576 hold576/A VGND VGND VPWR VPWR _5404_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold587 _7693_/X VGND VGND VPWR VPWR _7694_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 _9343_/Q VGND VGND VPWR VPWR hold598/X sky130_fd_sc_hd__dlygate4sd3_1
X_9015_ _9464_/CLK _9015_/D fanout420/X VGND VGND VPWR VPWR _9015_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6227_ _6897_/A _6510_/A VGND VGND VPWR VPWR _6227_/Y sky130_fd_sc_hd__nand2_2
XFILLER_106_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _6895_/A _6158_/B VGND VGND VPWR VPWR _6950_/A sky130_fd_sc_hd__nor2_2
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1210 _9438_/Q VGND VGND VPWR VPWR hold335/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_10_csclk _9210_/CLK VGND VGND VPWR VPWR _9453_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1221 _7415_/X VGND VGND VPWR VPWR hold699/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1232 _8883_/Q VGND VGND VPWR VPWR hold846/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1243 _8801_/Q VGND VGND VPWR VPWR hold49/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5109_ _9227_/Q VGND VGND VPWR VPWR _5109_/Y sky130_fd_sc_hd__inv_2
X_6089_ _6504_/A _6089_/B VGND VGND VPWR VPWR _6739_/B sky130_fd_sc_hd__xnor2_1
Xhold1254 _7839_/X VGND VGND VPWR VPWR hold378/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1265 _8981_/Q VGND VGND VPWR VPWR hold406/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1276 _8961_/Q VGND VGND VPWR VPWR hold413/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_405 _5281_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _9483_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_41_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput130 usr2_vdd_pwrgood VGND VGND VPWR VPWR _4941_/B2 sky130_fd_sc_hd__clkbuf_4
Xinput141 wb_adr_i[19] VGND VGND VPWR VPWR _6078_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput152 wb_adr_i[29] VGND VGND VPWR VPWR _5124_/C sky130_fd_sc_hd__clkbuf_1
Xinput163 wb_cyc_i VGND VGND VPWR VPWR _5123_/C sky130_fd_sc_hd__clkbuf_1
Xinput174 wb_dat_i[19] VGND VGND VPWR VPWR _8748_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput185 wb_dat_i[29] VGND VGND VPWR VPWR _8755_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput196 wb_rstn_i VGND VGND VPWR VPWR input196/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5460_ _5460_/A VGND VGND VPWR VPWR _8834_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4411_ _9311_/Q _7446_/A _4406_/Y input10/X _4410_/X VGND VGND VPWR VPWR _4431_/B
+ sky130_fd_sc_hd__a221o_1
X_5391_ _5391_/A VGND VGND VPWR VPWR _8809_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7130_ _7128_/X hold916/X _7130_/S VGND VGND VPWR VPWR _7131_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7061_ _7061_/A VGND VGND VPWR VPWR _9133_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6012_ _7645_/A VGND VGND VPWR VPWR _6012_/X sky130_fd_sc_hd__buf_8
XFILLER_39_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
.ends

